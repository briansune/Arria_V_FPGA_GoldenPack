��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t��PlͲa(֤�aI��ԓ�/F�O��1%Uic+j�� '>_h�����u0L܌�>��5���ěd���?��"�z�Z���ݏ�zc|�	�;*�vA�4R����	���A�︭�d�ʀ�I�չ^Ա4Q��5y��Z:�]6>��06��a�����;d����{�ˈW_J6,�x�$���1|駆��1�t�
�@�!��Xju\��k߇�M+H���/H�8�ƌUM!}��D&W���G�;�����Vo2�2���d�o�2��lEb��9PjJ�]���d�/��)ps��}���Ul�ǄH�S��l��q�Y�/�b��D:�L�8�Jz=HAR�hW�A�i8i�ܢs�� �5s9���P��'��쎇nB�����0h<��ګc������W���Bu��=��!K�����eK�.��}�u" l����M�7�"ɼ�~O863נ.̹�%𵷉�D����xg�^l�qn/�֕�Z�gh��%�����a��t$o�5��ޢa�C�س%�\9��u�A�~�1%��+���
M�<����}%�[#ZKu�������#���x)�1抛�VUF��o)���}4+�>G�5T��!ì�8��ӷ���r<Im��GG����R��pV/E	�x��z����M�T�f�oI[��s��h�'���Z�FVY���e4�7�
��l_UH�T�A��c�~Ȍ��iFo o^���/e����$0�I7��F�+Z����ݿ93��qM/��H䥐�?ѳ[��� ���i��(��t�f���є����O;�1�Q{3q���/��lyfb���lP��f*o��s�u�'�(a�q��/�-��~R���K���v�M�R(��}��?���i������=e�a��*���~�܏�Q�3Yـ���{��Y�Љ�!�5�����`
��2T�$�p3S07�D�仌[M(�H=L��jܝ�a����$�q"%��Ѕ���֚��Q;��}��z�ᔥ|�6\c�|V)-����3���b�"���
���"aE/4r�v=�l���I73/�ʸ-Y��%<7U>�}�s��l����hN7��u;y�b�h�A߆χ���t-3Y�2��j���b|=<�V�;��1�A�e���
jX�s
�y���%I\qS��I8]��p�ȟ�u�*��\��gqZ/A���l���,7�rWG���0'�����:kS}R~,���V�:���Æ�����_lG��nK��@ÊOu}0vDϑ	�3���K�C��ҝw��FmX���W,q@3�J:���=\?�h{���-}�z4���
�sw��e�����~[���bn!�1�+���7��M���PMFlXI���?ӗ��ߒfں�Գ�!>?������*dWx����&D��b�FUæ�� �
Xj��#��ʗ��=ԡq���i��׾)���u�H8�YU�Ҭ~�u�S�$�s��3�˪:@v���S].��!D��so�Ԋ/�$�U�zˬQb	 ����D�ց���y|�`d��9U;����\`��an��`{K���p8
��ȁ [���y��i��̯p'r?�N�-]�fzf|��{vz#5^t�я���D��E�ǚ�
��,��qh�<���ӡs�li����ղ�%n�M)g��'-Ŭ�C��6���S���	�����*
es�}n%��'2�VjI��(4�����mS.��8$f��E�u�qZK:9��J"��P��1s3�NwT�4f�}�L)�W����+o��`��NY��Z?� ��j�j*���4Y�����CU�� ��sO���	�h*��T\y��n8�׀�(;�.�/"&�	��I�Jb�x����f-����bD 㹺LB�4.��x�`47Gw���:�R�-e�/�hHi�=S����R��J޹���=�%jН�A�K2��G���8������,Ta�&}W=��_�� �?��%�p���bG��VA�NL%�Qb�O���_���+؍\5>�dki��-wz?}6^a��=��g5_uP��ή-���<��Gn����%gm��{|i�p���q��4j�?d�,/6{U�-[���΢U��8p���6-�W�S��2ܒ^�&��]7��@�@46�d�[��~�������ǥ�Ѱ{��Z��sr�Rb�܀׻��	B��{�z��
`���AX��Tr&x�~�j�{'~'�X����p�0�9s.��/d?��G��d�YB�D�gx��:�ClЌ�9��o������G�M'�;Xx�p��Ezծf��O�a��4vs���G���@�z��Mj��;������G7��ZhY?�L?�h��ذs2�{��Dj�t��ܤݸo���'6ż�6J�t�G1�H�_O�V��Q�O&�#�q�����4Jd�(�f��K랭�����U���[K@Q��S;�:S�&�U�{Qo,�����ΛJ�:�M�"�F�G �9�K��>�� �5��j�91Tݑ�.בefo���9�͂�tQk���
���+���[�.��P ���w	�g�-r�d���� ���b�	"?ɰ�Q�o�^B�[���+�����t~�EU����W1\�R�!�#�j���Է�f�U��P|�Td��n�w���k���id���l��	9��$_�v�JH�eb9���i�����B�-й*�S��V^�Ufp�?��:����T-Ea��}B�H�lR��2��T�=R�>�p$�s���-��vq���� ~�(O3�L���ñH�O0����P����|��1�|�>�� ��|��P{�ᦊjAw�����T4[������n��A-US*F�G�<��t�g��I3#��H�xPSG�(G�Kf�^dG�̳;o��h��eF9Z,v�?��"�(�(�0�m�ul|qaV*����������Ʀ:
�A��ޑ^�k�qb�i$�O�07p� �<����ܰ�5�[��SD >�֚S�zצ�L�HI�E�(����1Q.N�Uy�A��jk`�4-6�5O������X�&9l��o�nzJ0\�~�
8�h��:=������_����@X�~�8t�4]�'���#�^M��Dj�=
]Z�h�:�1�hȇ	�"��ų�D¨���r8h�@s]��zݧ,�`ъ�ҏ����h7�>��Nc��P��r(j!|bCӛ���?R��/F�y0�m"�/>O��!���.v�����m��r6z�h|@q�~��1��#�9���[�'G� �%Amg&ْ�ĉ�՘z:@]�i�\� V��JH��$-��#i Ls�m�(�*��GUxNM8�^JE��Տ�<�V�P@��F�Hg**/��ty��j�k�P�������l�����yM2��YgG�wvfX������do:(�k]uX谬�r�@%��~�ς�_�h���3MRB4L����Ȧ�($G'#��sn�Ȟ���F���sꑛ�.��El _�(�P����?�0�oĦŘ��K�U�QC �$@�aV%"�RFr��k�yw�ӕo��s���V��i�9ZZ���N/$͈�X��S�t������w�}����P�F�����Doe� �JMqgn��cUR�?N ��&3���CqE�u��c�����G{�B3A��P:$<��-^̐�3.	B˭q��D�+�>1�v��T<��M~�����
�������+T�.	;�v�İOC��.�����t���-��7���&}Qf�ˇ����6��th�1�A�?O	͆���v���� ��|���1|c�<�ɻN��v�(ʦ(�'z;�'�ഫ?�hתf�>����@7o��+B�����7���	�2�AI���~�0����s%���烧&�b^�$�*�T�
����F#� �l���gZҡ�X���yw^�cab�E���36`g��ݝ�Y�����(ޘ@���s��(����D*��Y��[����?�=��U�ӑ|k�gȊ��'�S�
�4xڰ85h=�d��1� P��L��(�����Z���h����1.��5�_t�VW�ss��O����Y�}�����T�˾����d��]�ܓ6�>xA�H�*�oh��UҔl��x0�eT/�N�B�n^��--��i�~	�2&�rK�2,#�8Rewr���\�v�Φ���¼��dMT��q���Klg�G���Fmv�+ѷk��G`tB�م,jpH�D�ʢ�yxFTn7��^�5$����ml{[FR�M��'�R�Ά�B\�h�yK%D���jEnpg~�-";B�'$Hz@Av1�@ߋt؎~�z����Y�0/ږ��f�?r�<��H<=�6��r^�pǔtQ�aG�v�(��fb��ʳ��}�f�6�g%J��'�܎ߠ����6W���m�|�%%����iby���0^ 0��|��F���h2��9Y~�%�9�o�n��]���a�n���nK��Ǧ����V����Az)���jT�Dv��L�?~�ypc���Ϸ�
`�]�d:�vl=n;�f�;�j�#��Eϰ5�� �[3�G'�Z٢ŗ`��{y�f�ؘzў�j�'Фq��%��2h���"��)�|����KꌍVB>�M(�'��iYC�l�ɔ+� _D���e�R�D��D����pjf8����C��keA���0�1�h�,������^�_o������K�V�KDEZ���&� �B�LՎ�y��QY<�z��r�ٌ��~�F�5V޳�/���?ꆳ�!�ZπP�H��)��,U6B����;�]$�N�T���:=�ɡ`@��oQD̛���eq��{B�t�Vft����*H�v��g��O��|�7�,�ڔŖ|��LP��p$*6��?ؤΣ���dn��Yn@
(��xmx��èE��q��V�<"7�ojm���>I'�F��"����Q�M��3u��q�3�M��ez��g��'d�zڎ�M6 X�I6]M31bo��=T��3;\cʹpi�C- *G)fs�L��׈�qN�:Β)Wnd��HUSc���ue;4 0������a��['����K�	N����+(�G���HP�iX����4�H�>��.غ��	뇜��_�1�F��TG����2 xC4�p2�/�~�M�@�����Zۚ�+x�
��bu�&���U�Wʑq1s�P@���⓽�`5�g�qJ����XЈ��k��$�H���z�JC�Uy6��BZH�&cH@k��*��j<?�7���XdA;l4��Ƙeü*iҖp�(ї��wT���.���{w��E}�Z�vOHU�~�.`";�ݪ��ո��V�5�ѕ���(@���MZ�y�6�z�c�*��k_���:y���ͨ�A6���rj��"��fԇ�J�X����(-������$H*�0ʈ7�W�AX��/n/��O2V�_�]gc�:ۻDc����Jd+�
B5�ƒV5��ΏR�Ai<�B��3v��I�n�,���l՛T�t�-R�VKT&��3���kM�h�q���*6嚵Z��)�iY�[�@���&����'q�Y�T�T7,�B�:�]��Rh;Bp�M