// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tKNZ4cLqZl8plEk8SCrUkapd/cStBo5iS3z3Gn+Y3I+2va+RRWO/znILgmVGEkJiBolYg4IXuL23
kzlJX5c4YstBNswXqmHP1i5zAljKP1I8/7fl1++8xfnqJ1YkgIrH+8/Yx1X1zQzGtWSVQ3YjBC8S
+CqidQ6Ta3BDLoJvE50NasTIddkwlkiBjkeibKDxYRUXdLz5vxoJo28+OazgHQ8325WE+Mu7/jTd
1rqQ09GEDNU7gEsD3JpELg5SEMiNWKBxOD/HbY/ykQSPH/qgP8jVEbTfR4PLNKiTSN884BjEdfmq
H/GBtf+bnaIWD9R5ZLhkASsHUizYIaT7aKODeQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 93792)
j9d+Fp5uJDWHL/kjyyZSvybqxjlTscS9lcu1m7rw9SIElAiuh4xvfsPBewyDRuBlye95ZGPT9zst
7mhm+0PyPDW1gGMWRiFbO7ZJ18reZDdd9wcVbezVwwiIF5j8ZiImKSoukVF7Qzn3V44Ttp0jXo2d
5HAgkBUpZvPaTXOW7USxkk104QO/WpZ+4nxRuBWfSup0IzQtxdg3A3lPlGp+RRv2x4xMspJH+4Qj
4jg417AhC5AfxFf0OsSG1sciorCryExBZkudlK0+D1twPdhYqr5TYv4O0VUsSYcpulxB5EfYmlBF
jdhBE1qetmLlq/foCg0P7zl3RDtwNr7VGbOxwaFj2TgL93G+pFxTu6BzgO7afQgZ1nBbFhBM14vq
6UZbqwaJTknfzYjF//dofFbVBnvGUJBPiA82YZyBT4fId5OTFFQjS/S/vTVApkL/VUYdv57ZhKz8
KmNbDt7x+4Bb3+tdTsVgsYjcez3bJNIMFTle3VnjCP9wa7anK09F0SjzYqqURkdXcPUNFSbxhtRP
S6s65dTavYbFptG+VMFFjvPmtVQoU8j1LY9bMrBPcvNo5mmTgPuocqBFra/u43oF6mf0jFAoBUWp
M6DrHFLtSSxOIJRzlH6+JPWXvhwyH7QgeqbxUYSxeljKcJ2bmJ+TDitWruAMa9OXZNz2Z+F2JOsm
ijjRPvz7Pt1uJ/Xc3t6ES/x0JWIVI8pudWYnIhcqi5Wh3rRKpHlVKBGnOs6Uk1/f58W22mMhaLRz
LG6JaLy7XOtgRwtj3qPFg+P+//VFaoSxDpWZIPBzuKheXMbtu3/h7TNwDoRMQ6yOlc4zR2m/9L4y
fYQfFR0s1zDA0kgG5wTvc+RPtzKfdtvdLw9F8Ffc8u4rR39Y4vKj9C6WzX5B9D0QFNnldbx0pQQy
1yrLPS6di+T+s56b+lXzV+zoJ9NSO9NFWtn7KEu/Sx1SFCND1PLLmwI6kLotK/ibttkfz8FfJaqK
mv3tNm1hE8+egwId88+2dcrcowVEU8j1m/cbr207SVc2bAbdrViCp9Q9ps8SyfmZd4H6jPb3Qdos
n9TY6m+c+bWmYJLV0iHQyFlYIbILIQsAMp4GcVYYjucegMZNwfTOiPZmZO2QH4Iw4ifvAqKwIV4l
X58WYtQYaC5QWJlo2d1DDYKMqGrCezWTeQKbvHyGjyU+2lGEb5Z0iKqG0WDDdgNG+yHcVyeHt1lN
HzxxpP96nXWC8Ly4WyoSFdJxMUl1kRg2c6pOgjlTT5LxQkHRFkEtQkySQtIf9nDNGRj0VwMFyVZh
b9ErwJTGqoOJ/wibGx5XjOle+UrmLO7TpcfP3+6ANgMJ8GKF/aLiZ22I1UNfzTuarj0ngmX7U/Yw
tJq8oHNOGymhJl6uAZM6QopsZn8si8c+m4up82kH6c8hIiCyquRs4ZbC3piFRRI6PeD5mpbYSD4D
YZVLn0N64+yW9B7mkY8SAI9kds6ekTbWZnN2cdmlguUeGAOh6CQU5+Nwps4k3sJlSeMvn9PZU7Tj
Xn9I6it5AsfgasTm2bwvqu8G5AnTelaNiBT979b3EG3A2TRVqMmPrapr/cgo5GuqAw2mJIN5fPw1
0Gv3oqzUjqjgJM0v3p/hy/uwyVm2jIgEXDf3nOvxbq+ADWJlipwpPZ2GjrIF0T5tqKerFBM1PTDt
doCysMyS6jEFNWyAccmyZr4gzyXgCTShD6y/nMSzt4E5/P7gC5CaFkn828IvyFvAZN8Di+G0LAJQ
gCRG+Lq2KL1AdZtlw6ufcx1JH5TtI5KXO25WcYoE7sD1Mw7P+CKDEjlCVydCZnERRMi4EWhFztH+
lC7CCjwUQkmoXfpUuJ69oERrf5UisNwoDJEQqhqskN3tszNSoPt8VpfjrUQNdWOR6Vi+Bj107ORg
ud4+afCYY6+34KRQe8yuMvezi2Z8vB4yaVtKEErQGLxHinYx2jjsLf6O/PjmRT4morFDyI+jiAJn
UoKTL8bsAGApAoFu4ZgcfmsC6WN30PCKeIjNVeuC8lSAX0TeZfirW3MPF7z4b9uMFzzPdCxkD4X+
u6MpSdYeIcwMkyW+d8slHPE7NBisglCCpXXkfWNYTbQkPFZfXzOBpTdIMKxd7gYu97oY7PwOZv04
GODmkhTKy0dk5hHGQ+dn3xQ+YcCeZAbu83omKUWoqG4FrxOBalfGMY6ev33nN6U0xy8JdDbVS2tb
z3NKeuXfUd5eAepgS6k/QJcPhwn9D7bxLjIo+PGjpw76mXcNBgVD4Tlo96xNhJMA+oLl0YLWOcg+
8HNtArTSovoFBw63VBE791ECps+SAhcfl/qpS7l9YnPf2BnYouycH3Mj/jaLR8fbNGot2lYCsf9U
pmVWhhNXrEd+N68IlYLTGFuzPHaSjeqjHQe2pKQELXa0PSIZaLLO7qeNlayKBU5VzZFh/20w7HpW
egOpGeRRP6PzbzCt4cI+exzOy9Q6aZtECpz5/XisjKtLzmFtXq0edi7CuVZcbfcJKs8EWxJ9uObe
AUzIUNiUzuyc9NxI1gvFSUJOdm+w6/ZADLjgi96Y0Sn1MgSBZYJ5btHZoyjWHh7gAVXQm+XctCPP
KDPeTiSBZsZX85WAMT2RgcB7stWmLzQCKEgfxpAtR6P0UwAUqkrqBQipdqMBVPe/kdWaVXpGEKiy
XMdWRKPnbJehzUIBH4tgft8Mo7B/eI8JT40sJqSm6hTxwitGSotWikID53PobUfpIgGEZXijtM1V
MB3UTIEbjQDo7mju54HGp3UBBDuo2GYpMoXx7Y/vsuQBagrhGouT3rEbLFybjoXOQer2FEVV/IIy
Wk94dWLshXfgdVLCqgIVkf957sVWIo+9uOMWHgJcWVoYGyBDN3y7jADOiIcuDN/Q+u2TfnFTWb+o
O/UmkONlRfQiGedGbh/Rrbd/pHr5HIuDcy0uqTeKYJHZlwxdxb35GOQBpznkQ59oHJfZUbPIY8BD
RU+ZVJD1njuhEEGVUsjyX4233eqHbC2zKzq2TD2Doyo2Dfi94gSIG2/BXoYVwHGwoAWIs8hE+VcZ
Qia4+/hO3QBfi2p6g1a4+wSemAvuHx8SR+1zzu07hA+VqQNK7y1baYkG2oczDWs22M/UAMtcQYv9
BktGPHn88BJZueoi0aoTmqSAgpJmBdhOPWVNkxgWa9LcVoiex5r3IpV+u3Tdk0vx3N/BQ8ByifFM
j+naNBoH8q0wkFfmKtOr6zHV/TPsTrbmgunTWj8oBNxzr4vYV6EiCLZRBrcoGA7/BWXpiHtqKjLt
QXOvVAT7LkoghCmXSrODlAezNX4sE3oFAkGi2tesIb6qeAIdb5mHS47SdUvJjrTL3aiFq/InCLhj
Lkx9rEgS+x3N2lgu4AIiPOERc7iwiKcq5jZPoYUjpGJ5cK1MAqbYMPGpj2rMWy9y7n1+poMaEiU5
HSpk1I5Bf+GLKMVkvXMrVesaEb1uALrA9Rff+WEk+fJjBu7EbHrx59ZhyrHaKR45ad9Ul0x/1piJ
PEhNq19+1YFVIlYAq0NPSWZ93dkJR5ecDdC0gpznwKRwdEo/8NDvo4piFoarqagzeAhmX7r/xrHu
O3P7mXzHfUHS9bF0X6Zsq0IyBzGMbYi5JAfg2TRLUFzTyDIl70alXbsdLnA772l3WojUg4AI7ZUK
YP86yD9Hi3WgNBmqqbPFl0o/JMRAtpvnobrXYETADOkTEaweXtj34QGxP5e0wn97ozFaDoiJ9NJd
BFE5R4YVhycJxD8Rhll36c7vKLVwyH6HmewblpiGVeJsJMVJftKQ9xxosQs/ZSArwk3keCinkibZ
iumjcsTIE5hCuXgJfPCBaeu8XGr9phelwT5yd1gkaJJwsLCxaQezxSPeFQUD0e3+V0gP8aGbLiEO
WMELIrkSS6DfSOFglTRSoYc5nKHX7L3Y3qmY/JHkDKhrQcSl4fjV9yYo9oOck/BEOBeUqrFdhxal
ULOKaRfEcJwDbhNIjr1AziGaLVsN8QXy0qD5AP33Bnb7mK9ShYirJpw71oK0w44mJOivgDSVY2Dy
PrXByrwg9uNWmbORfpPbDdPLIZOjexC8wTwxqKA0tay04SfApE9o1/yfDkyvb2czAiKNpud3Tj+j
8z1EG5chKs5tO8xLGjKEKPTqQQx6E2OcU9dLPNgpa0pGfHNUQ9epYYqLSzKqQqFCFAigDEhjzsAo
Nsuu0vtLIa/z6IU5bnUesD7MjkVgQi3nbGX9DbZj1ADG7liayw36OOxO6nJEU0wfUdhIyvhIWVh6
iIqVHyMdVz3K/BNWPaoiTHm+qjHJBcMfI/p6X0NsPGB5PN8ny/iqsYu0HVPD5jXp6uUahqdWM8dX
bQMvJ0EcBz2oY44XmU5MoO7PSdsEAU0n718YpFrzRS/LK4zbcC3GvBN2jgKo2ed6hLgJY/2Gw3r0
CErmQlBY9ns2bnAJrMaVHec8Wqc6O9DeST67PsZk855Wo8W+gUKa4tUu5ZYK/rTrR68aT+/iOq/9
V9P5wWbSdMAr2xQuF18dAx4HkC/jkyYj5C8KycL8jIqfnqE8429owt+CZorxcu/xo3lQ4/mEOj+S
81s/yHt09NRVEtRr5B3+nbE1lJZ/uRQ4UQfuk8SmI6kO1+9xPaZzi5nYVAKYG+Q5JJIyTidR8qSk
3MQDkh8JUGcLofopGhHLttH96ZOZJ8Ny42+K8x/Vr6XdsQwnwp9KJ8Ll7a40adfgoEF2MstHYEX5
xWOYdF/Yw2zUcpSbedgTab8gmzSoqFjpogPeMpJzqS508x2jQQMux5BUaiAWs0QJi4AmNkJeTo0D
ZNydVbb78hoRVRCjCWxzirwyQOC4FQHcrZX4R7UDIFrsfGYWglDMFfL7+JYthXzUncwt2co6lqlf
L8SScHn+hoO4uIneJEGpYqUsVTU45/Ev9BwevoOD8kx7qUqwEEHPXzyx1MPrsdezqx+rc8nXKeO/
P9DkzzywlFk/c0ocvcvZ2vhoRYlH4nfDmWPo10GLmOthChD+dvnYpFgD6schEnDwM+1+KjZCFJGq
cMqXTLYYZL+0lYelpaG6SGNxquErxZgKsu3k8d0ll8iYTTDqkONIgQwc/RHtzAEy8X/k1AypkTxT
bkIaH8NQ51rR01tcWRazzbzQgbJ9sOO0z9MkkmVGe0SZGFxj9AR7YK1PdEiujUvipO1HclcsaZmf
sJg2RiCRPTBnG+gJnzMaZ47Vni+IiRvQz79QTQfSGPugz+N1idCCR1DFRVCF8ZX5k3bBo/V6HoUo
GerKVkfcWzmnxJdvMmC9IETLXY611gZ7UK23x4qYcOqYHLan9TcwLYZ87QwWJXexeY2KbQaKndmc
XAItwzQktDozxFjaoCUNOOpiI0LTLQ86zMDb8lH8+T4RRmDz9vdaxQiYh63HtAw6/LQ9p6bR6ZXM
JI38LgBz7JDqBW+W0Yw+zuBDUdtXv/g1B1Co+w4Qha+gwnIZxyr+gY1lNX97hpeuWiSTB7EtL3AY
8PZW3O/YmRbpp8WXWRKJbIUQ5mupApwgl3Ca/xur5ygDe5jY5+UVHHJWkf8gw6giZcgYieQyDqmC
hmmhRHsEMknVfzMp6NNksCmQmMXNTaxRaKrr8y6Lfrlk6HhDo6GcS0CLvkux2gxOgH24NUWmCBl5
da13LuPk6c9BQVK9SdhVFi9SmVQCsUIZ0HhWRfghf2Vxg0uC74nQAigWKqczu0NWeYph+zGxC+Ds
myUgGnHjDTnhXaTR7o6LF9fkavu7ZeQL56I/MwIOci/wNrTfq69Rq6Fo6t4B+J6ICUK1N3dbnVVh
vgLukDOj0J+8rmQexuMV4n6d0U94zNA4akPXhqMkWWHCRymAcqjZivHTDbpxm5DLRH3DeQLVPDrn
V4vnGSxXWSXAzFfogCbpNbRTOIYmbIUH/tfDho+svqHBD6hpUgo1Ls8ZF71325KsdTfINx1eRtH4
AaUY8d5kBMtQuVU09pMPbVauH6wvmFCial/4wMjiYRGw6IucFj795bHDUZ7UqGPGM2BeW0KAASPE
wCQUZZHwh7L8g6jHFHN/WohBkMnSMZXbX/HyujaZAKxjYMbNzV8vgmD4bWKYEbyQvCFRXNqWnAQH
WOfrLS7jPbRUpVyVrSehtpLur+QVeVemlt3NShrQRRvtJssGvew3osrBW9jLz6HeCBgB4A7qzJyQ
bH98NuSpscQPPTsx8Gt4OzoB4PuogStedAknJHGb4BAp/FhF8o7AdyMPhptSmjd7Blp1TK7O8n13
zEREhxMLwKrIw5YM3rJKgqe9S7AKnZjZ0HDkYdPDe5edAk1kDlEUxTuxYTk2jhI5Ip5LG+iwJVWl
3v+ONzwc0fUIqoUYsiwdmkCToVXQ0WDKA4OrvjzomOw1bQ778NLgBHYtGIVjfH96RPnexSF05o6y
7Vu0UmMIwNxV+u/ZEIl9xSw7C195cRtPYHlucx1UvqVahI0qB9qoAoI2ndRoY+u6F0qm6sMW9uwh
RdxejXidvdojd9SoQ79we86yAQeX2/lQqu+7702bACBGJnowDgobHoZVtLaezLBXW74C8R2O1BLk
AgLOcLSU0SQRrsMazjkKv2xzJ4NYWqjAsodWLIzbGuL1MWQmNXnLttjiLM5oU7GecdZGqQzOYvAi
mZH81Cw5r4MCg7hSGgQuIc1U3m2ddci4Mwf6+atGXaBmwIwnmkW1YUHbtiIwD3vOtdG7De7qySyy
HigJa/mUZMTigxtwzVPmH3THla5OPC3yJXxCaNuM4I2uFugqNheS/mFelFdSDRZkezuAfCQ7t32O
VMMdVOkUFhOQovxWpDJUwC//pM2OC/xIxIs/1XPTnQMCPIdnOOS/HPQ43iKN9igDlPOz5lqpzMm+
yho4dGAAEqMKM3aykNd/JmsodZAO4GJWarSJKUDbLqie/cImXN/gLcc3j3YX+npunJiJ1rpGfm04
RsLahkpeddwBte7YUMfAzpTmxt9UoYAlK/GmvE9LS0VTS88p5IsdEgI9MkzyJBm5d3/ndXLt3gjy
GIMaGBTeieCVIMl2p+50ieLXSR+dDMyjSF9uptCN4zn/LjQUuKxKI1jtWtHZXxIx+RD+bRI82gk0
Bux7F5blzLDWYi2s9+Q5SF5ci6rKcnlYouAwn5kwjFJZFS/ITNFbJXMtPNtNkHVPE9n2eJ4Ta2Lq
tOfsMHLt6kNlHcSV06fAwqyPnckihkhbNGZYPkZi8MAbpvitEk9jyRaAVjezDMTnCx8KWrCehZUo
nzK3ipacqtMKpI39Pq9gTCT5HkJ0BVek8JroGfmOshSZB9yawitA6rtEmd8SGjewTnQqwsrQPg5q
nrxiNtZKXV1IhUmMlAU4NzjGLURQqo+fKIbNnoYYWZov5zAZ6u3gAYEczftXiEkIpCs++340uxyM
RSyj3VsrGvTt/5YRzp3u79aWyBmqPZ4l/sg5s+MN2uetuSMrKc1IOeGPSSLgVmvtcCKgg9cjD32Q
nFRerD50tI0+hTc+HGqhhVY6tmJiqS9ymputBKdY6otyg8VT+hrXg9FGwDezPukL/NCpERmBQ6CI
EOtBN2qw8aqt1zGzhi/p3N1CL5bFfaNBySri5LMG72YSPLr+gcxUngVuyQIWWSEke8NTNq0B6YUX
Qq+VnIM6TN70ywO0BgDxyfefeAHiclSu92wUEvrNJWs3YpOm/Fg6LgcP24IYTyUKkCQ26oxgeti6
Us19ATEGnzU8T3ZWE9phmHP0paSAN9EbYRqv0VfW4X7ijfwqHRerfbq3LcPr/1akuvIzU7m6UPxq
ZcxI5Fh8iknoG4mx3ORRzTzCNjQ19QU/s6NVuK0ouDaOwOLFkCrGV3/DCgTcZzRpY1qUVOHXZPCF
Ahltv9whilzhgsaX6Y/TqOikvXEFsrs2kBDrIgFsRWUvijto3kQVajfDBGk8TOWnmnZ67m2c2oE1
1bqhSRWZzgRYUt7dAXI8FA3AFJ1AWKHaTI1J8eMPdnR0mRSJS4d0LtVKi5Iuc7mQkN/tXj0V+Jq2
Wt8a1hX/JQQxHI20B2+r/WERsKAN1XQXeL77Y08stlbNvxwcjkWn7TfWs7rb9WCQA+L5TeMFbFja
fk+GHGnqLVKTxStl7bdBIUDrnOAs2p3qGlbYERqwgIiwNUjmCzYt6uOtebnFqE6tnhw1zAQpmJQ5
R3ZJFwt+NOqLIBZYQl0izJmSL0PGOathCyUWxDQbyUW+ECyO2PjP00J73RfGrCLJ4CYfBBxfstY+
rbhuqYij7vUG+tSzWmscWwwuVNvUTAZjoUP+/CrCm3hWLi5BDHssz7W0fXx4gOZGHG1zoK7JTMzc
g6NdWQlvswIQ4fBRLga9LrzEEi+XPbpd25m7KCQBrRQZK51LoHwQIJJVoLLls25LX9X1CEPQ22Rt
7aO11YdK2ouv2k/lIPkfSh+UB4SB+Fd1bekUPGQm00H1G34Bd7h7lKpmSmyZRtNhu1zJXLZXh0O7
mEIM7w6C+kHun3KY8CwM9TQNlCheerdNkeSspGqx4WxSgSvdndUuJ8FhU9PCeKkShG/gVJahEZLg
DxoSmhJ3QKunqmh/11QX7zV1zGNHpM3EGKoyTXjyvRO/folu9TJG8vbFh+gO8ac1k8D8PshOX09H
CaAu6sf7vv8zUMfQ7BMmJjWMsl1Y+M2IN/S7nd4lTVBvLTVXq8yncvBqdqA/jsR0biy0t97YeWa1
/+aSXd2i/qEYplXQJTHrPbUjbefIX+eXOGwnaL3sECjIgasKJdJ7w9wpsaCCY4cd5aN1gAjB0erX
30Jwn/Q4KsdyI6+fqBS/oGHVyYB1kgV97mLK0KKUL9cVqxo1nyj2BOTB7kdxLU7pRhc3OhKCB1Vk
6SuFQ7oTENTPmO5FtT+inyZYqyji/fOR15SAN+lO4vW4aB2S8B80uiPXtYaVVzJIn1RQcEX80efs
1b9hFny0i06AA1Gw0TCj59CHhm5uaZtR8DIELEo61J4PodN/aEIM/s/MLC58UQeQQ4D/qBdNIvZK
kdylSNo165nH57pbGKjRtOQZjadhHc+4pezxTTlJLXfCQ5zX7RV/r/EFDMiu8nZWja+2fy7NDNvV
e3GDUTC4tuDO38JU2hcXXN9EEL/+so9v/O/48rg5sH7x44Va8vZi7PBD/Oq+WtrzB3rqgHDfEiIn
vlFFfkgTjef84d0mfYBJEz3RbiSi2E9WDFQo0cwXT4nX3zzgkKpNqLR2u1zABnS8FhVX6RfjDtz0
6lfVBvm3k/ikBqYxOMz9lJLc4+UYQptuew31Cgtu6OD2tegd8XVeQ9PERMj1iRObJvFBGDjBDUfD
43T53amadDKlm26HGIrTfcOT4htDl5yFdR1luqlt4QwNnHkcTCjMuxC2sWUfQ9+cbQD8YWR0ifm3
fi14uIO01GCVrwcbSAYT22+3j5DWr2U8NxwSdwICdJRye8+qtNsoiEQIIkBTQIKLDp1nbKjSqOdg
ztxIZLIDb9Uq++gvNeH1CU91FOYq+PG8/ZhenmSCbNuhEOsd7PKmdQg5sMLx504ndtp7NIUvuBdR
3G5o4QC02bZh5UvjJEleb/16X8QrjyXUn9p+DgPpkynfsTh/ZiBghLUxckgDudqMex0/M3mW31/N
1cgxyuE6mLVS1nSLPxy3nLFmjwwpPJwsaxuhaHb7zPPqn5+IXGlw1hRf0LnPPRsqn20p2BbeZhRT
d8TshKgezDTIHwoiHExMtkS/pzETKeKQQyJcj51NLe5r0675Mcx8D++nAHzCCJQGSVUedsRY9/+H
uipScD3vxTaBRUCc9yGU7GGoa6D0Fga2N0uDLOvnyguENBS5zB+fdShFlRBqfmKbY2fn1w6nZAP1
yug/ljJaj5ZxeegEyz8io1fl4ddiN+2Sprkh7gZKvMY8uaU6ZyFuUqT/q1zOsLSrMBMf04WybHfP
Hvr+p7Xvobiyi90116z1uPdWAwLU2j9emhHlgqinhxdanBBYNDsrO3aC+s9hcHMYGreClCnEcNOp
fL3opSPisghJ5QZj0ptp99WEZufa7LHmg5Ih6ZI2CvxunRv1uAlC59pGps6VBgpyWS+jZfDcBNen
+/AWS2GXXKNBBSusF+Z8h2yTfic7a6ORt4Evn2xja7SN9IbvclwqdXSbBzgMDoz53RcIwnCIAZCx
rvPiHet1iy8NwF0+HDkVZrAIQecQCV0dX4khNjX/kq6XJLbfpADcF5IcBy2s8uGejXZ/q/dfq8ab
T7UzZZV6wnITNEC5hTEhkLSI3KRwS4X3wUJ6pMC/Ok/4UcunFlcyEAxbVtxdBvrEy0AOvmFXan3k
mgnIB84EamgUnMEY2pPxytT1jTWFxh1SXUdW6DxJjDok5ZWwh57AeW2F0ZvYdKVpz7awF98NxyMe
Q6XAiPoecAayLgi/5JkHeD3a+EKy8D0MUC0DwvHkQVZUcOt1svF2XsYxuEUfVGd+2o5vXNSFgDjK
NC62o63fnqQv0CZgjxrgpd18xmfFSvdgscFViS2CTjP+0qcUmtG0E6Q3vQYGC6Qu/iVOYPVKsN+j
J5boxlfTDEZgGIOjTtA9XQZkgAmfyvZ4zgtyKOKtCo7CFl097pwu8F25KzZY33B1OZ+JAFHVJVXA
2qWjIkOMUv6lKP6ulyk69ItcIsBxD8DJELJFr4qBE8BnRiLXEVJBOnWzAW4JqKwU4339gWhd1wzK
RB/3Plm7OJN+/0xciXzYMTOQOaSiyi5T6mmAAsqCCOfi/R59X2alaijmQG/hobvThldmyEaeDy1n
5++DKUCj4sTSllk2VnItDbO5r5d29tfQNHtXvoiXZvbPkV9T1jfSMDxunRM4vSvywDI+M1Ps3AyJ
SoJqxljipzqINtBwIyhmrwtwom/IA816pWZ630SD/vMaE+3Uq/daVjno0eU8l5kq2RekO2ps6rbl
IcCqflcSZb63MYHSgd/psRRgv4K2pnvBDaSmR1YyJfPvSGCEbPfmnay770jUuNjbtF9oGDAYndKq
f19Q4Fr8LGSlpRlqoarNKKCH/gusfPwg1lyO3cZpPZUaykOfX2q3zB7IP3c213MX9hjbHutA+JlP
VukQOgaiWzwSjJTdeuN7K8rzPHhW06GV6EKRref/00uDVNOlNAVHsW+SZtjVg6lgC0XnFsPJu959
SgaYIq5/xL/PeZ0YDkHRxE0dZXkecJJ+Y7blfJQ+ojEssYy1/ZbXeqyw6jo5l3sizseuQOkjUxWS
W/6vLM4mSU+N6jBYOBnJOAlU/Wr6x0UeTJPDvKzQoC50u7GdeZpOdgEl/gkZ0GIds+XLKMQUH96K
q0XIMkllXtSz5PXEgbjUP4/JgxLR8d6nJkSdnnLnke9dL0zcWeK6fJsYvzvRQ6Mr7cwIiG9oWD2H
JCNnC0xoS5OMbzq4GM7oGxJPm2LXzo/6ptBcmhW3QDGnQErm6wBqV0DNkYX3q2y+Hm/Ppr3b6M1a
PvJqURw7OvJjykBxgbCrV1GJvOU8Oeh8n7g2jGMsb4Q3cX02Txxtc4EexUnAu7tI9sY6Dw3Zeckw
unR25NbeSUvBU2r/sLQVWBrrJwRqlEr6eXWeT4DVEZzenZXGvcJL3shxyM4pgpGlxVrUbmvBLJ3E
XIdqN8r0eJNf3hehWQBX5TnVH9sq5ew5hJqmobjiobX38mr7CEUyl4DuffH05v8YuPP+Rz9Xt6x1
3vjDfbrRyK+lG1+2owSjEXJ0NLDBd8PrJDdfeCDh3p3kZd/p0SrPM8aDjaAXHF+G5vATMHXd6Df8
ZrJ/gbmvn2VS1hodOqaqQ7mq/j3O0QDIgPgzsA/JThCQ4H7Tw8w0OF7U3EcG2KityY/GBkMPxsyx
OroaL4o0KF0j5vA7sLJTJmgdis3Qwm8ckIoFL7+LbEfxczfxvTZWhM396gsIanBq/P53n623Mk1E
ktGESB1FX8lAMbjhNoQGdyJRezLuZz3QD0GmoVgtytJCsMTUnftjnTboUWf+JTKtVHOt0XBtDVJA
hQUwHFiypHei+9JRgNueQclMOiq+q5Ld4FJHaMxmEPD3Sy1rUrPavq/NxbxphxwikC2JDLNmU49i
G/j4QUkxmCbwSuZ+Dlh5/vgRqkSlE4+YrWCDR23IcwBU1Teg+PXi5TZ5F0kk/XXmDvdMocsH7/SE
3lyJ8Gd3DqTnFwFHK+93KAB0mNi1fdQ/7ya6vWfSXWqNOdohRM/TWCFusDaDOmHqqi4QexClr5kU
abV7CLD/YhJKfrF/4vY9Pnk4q0EF2js/MjPr5MGfOY/UNjPH468YSw0/pe46MWLy7TEuEou2T89G
LiQiR7XJH7RxIasFoHP2M8DBaqn44n6Tz5qTXVUZpzlt1H2CVYZC9PESfX290NuNCNL0/L7EFRku
r47VS74ICgvs7bi4cgFxYSOXhNKH1ZXEKwK58x9M0eqSXrkdwOILUBUcze9vCsUnslHp/WFpELol
8U3sbeDN1vT58VWXqk8nOUtjEfmOMpmgcvPrz3JblAVn3FN1Rkh2n36Yf+8mGTRMbLeNUUgPppBJ
+pFG3YcQF+UuNVBHviGm/tHb75HT7egNH6KyTwQTCDbua1MjBsomCD03S/2zEcWmG44NkjUIsOTM
yom8RYqjQOvIu8grDZTPjerRJ08JG1ErFzwfiIUPkiEq1yHkTeWmpnM84n7/k5MPjGHFkohwhNhY
YH7/mWYilpl+amE4Eot9y+Ae1v7ENHRYO0Tw+gN15Zv6XuLeLiS2/ks8BRSOL9oVC2hsacssR94U
V1Jd/laZ3nGThUKjiPRCpDASf8SroWpkseJz+ks2qI3tiyCaq8TwmLU4Az0LezP84XEDiYNNlLRa
aOnZkaTdA76cb7xXaZ1ozHr0DUF5xWbP7YXHbRt7J5Jq2pG0+ZI/UIPJngsde+kMDUG39xUULbwS
7P2x4H/qXjH5vjcq74xkxKvcfiyUKNjKSZo7TmIvRiaYzUDk4zY04iHem4h1e4AaEBZACcxoUccv
M1a/s7FgLdYx6Q63y4Vg/m7p+dijMYDbi1rIhwJujNMH+tSBB2rnVM/kp14rpN8j0Jx6BpJ/huit
tnJ8ra0aTWJiTWjpkPHpKnfLqC8tMMwuoblMNVTID0gOgWNEYx+PGYnvT18GwDbwg1YMztK6Yl+N
i0UzBlBQEmisfGvqx/GUG36cLoLdslhN0AasjXSROzkTdNm4ARzs35moYePsQzBjocmp0vAQS7Kw
HssHzd4PY9VuTOBGnr1cXBNabZXMLu1bpWJuTBcapj+VpWOkEsTyRB2fG6VVDNpWhaKzNTkZhthD
+52V3DlEub4t8rc4y1QzD0vS4TCKZh3bGzhgE1pjZWYvCuDmTZp2MLIAxju2sLmcjT9LzqRvKT+A
xdFfhjI9rYID8GQCozldjDx60rZ5yNE41dkj5n2jtSU70dB99vJg6sBX5SfU7VYwDjM5ApxxBkTh
oBH7/93P0V7Cjgh982+Se3VLMtUY6Gxh31tWunwJnE/61ZaXnEbmzEdvn26aGeLO3r0Zs/wohkBY
FkjVRYgKyIHZDC4OpazKP2wZva9U82xgzS9C0+X1p427MxOD6CEXD8TaMyUgIld4BHfSxXhJBakR
YpMomqaHc87Y/1UoE+mtvUL66X98C2wES/dIaY3HVfyKx3k8x64Ga/sHiq44k5ypou0kKpnMiGYm
wgqCsU0kSVgMFhX/5CFnP1Eca7P5l8jfkKOsk+pynFmySg+VfHSLFK44LzfleTjX2k22fX1wqLQE
Qx5aIoQrouPbo74fFJ3TXr0z9OuZXJWck/8GLiR3bD/IFnM3luqtUuJfo/4JmfJs6DJXAChZf7bj
H18ZZgxHmQVeRi0F3MKIr8UzgFzNI6K66mPq8X3m17Jml1zQszqoSagwACpP1hdYiO8n/kg1DHLU
h/FQDqeQj9ihGEyS1kdhCobYD5174Qi2IEBLFIjMj+CUcQU3LE2xN0ZyIRJu0QqpVUBJpizjOBJc
l6JVNEw4xMAqSR40aeQ/NiCa/UB0EkZJUCbpk+4FwWICSBXpYez1azPkngmgkJGeFHgtddxbBXML
GG8gZPB3P/nebwdWMnWP6Dxz4l0f2PgNTsZVKBYS8SlodmWeVW2BDcYrx0nMWlwC6Dx/j1EjPRi+
Z2dCVFYu7tITNBHaIpNARtXLxCeIKiOmHyE+HV0QLeflB3deAJq6co1zlVv1WlRQ2FIBU4lBD6HJ
KsY48f5earUVZ3Nkd6neESpfKSQqULqqLmIVaUpmQkhSoiCS4gerqCzkhZumek4LV1u0FS0hBY92
LdYnz5/DqRPyE2vnIVKysh/+BwDDrjspsmDtMV4hm8xaTJ7GdddkrBb4mb1g/viy/4bTKM8RwaRa
VBGh0ho2odCIiHQl2oDqJc7pt5JNerCP42y7q1Upg6XjdkLtI0zqi+vtVSrqTNtQ8Nes1an5PuDe
mWPSb/9fFMIBzUyAP08FFwNoUw0eQ+pEbxzfcvGinsEDe/pjvrf3AazZeJtMK2kBBab5oqsfMKHU
emA2QO+qPCOqONXwBGUjj/MPylXlwPbGUusPPz6ZcYNYl13Id1eju5tCapggcCuRCeOhaxd1TLZI
GH0c72kjLX2sP0+l1dMXsQRnB41h0BwSx36JgZiVL0vKFKz8LKf21DVcrB7QOW/NNkEXIYfRRA/O
70OxhDs6jp4GO7f/dL8/9y6YSZBV0OOPiwf6GdBwWC5CcaKz29tRDy0q+7zR+tfD6CEpSgymRhpz
+PJp1PGRqtc3RR3N1H8mmYneV/eHuN9m10G5MoI/w3nvg3T60fGpiMCTKW+VPJZ51NuK6q59PC8H
/t96UPzjnzk74Wm1GKGLVQsa+oKjnTK3Mgz7mMcNS82cBh2xG3UcIMD3Ngtbcw2IL0ipVNBxhl3T
kNWOfsZpbzL7ZB0KOxzAO5TsR/vDdCsvlAN1TOmaFXUytWQo+yzt1rV2P89t7e8d9LxtrbJEb8Lq
GRppoHwha/501NXdR3XKqI2QxxXUltTD8W8jQN0ZeADcBIlbmb6O6NExzx1FG0Y18osp+ynXvnxJ
OJB/hG1Drq6GvAO/PHgfBtC7wT4McEuvbJcWKL5JYsQ71RvgEkeQrPEuYHbgti08629NS7gIi9RI
Ms1i8KhKRWq2TV6O50SYj5jmwaYakGxgBVZYK37w/uVaW5QSpyZVLARTrp83ltdJ4Y+Wf8bkbd/6
/yxwtJgFtbLvl7HSjCZeV0L2kjWTRdwto8eILktfR8eFZpj87fMUaM1RyA+2O5RYGDUUT9Zuc1De
l3NqPlMkHQLKZ/CZbP3qM7MzjZB51xbIv4NnhDKARDAp2Mx/CuIwp1oi6juE5byqGit7cuM5qMeH
XWzNJqCblCvzbICBZSENILMR0kv+tsEho2BlTZVIKB+BiUf+ADGTsANRAZ/9yzid28m4HzOecPUn
Gr2K+8jrYZBizpFFvAsM7VKXfJ5H/PRN3GMCk8YScxfrXrju+zMaCA16qoVHi8E+zBbcNbizF8/r
uMyfT0LiAUqlU3xtPijYmmEMcXDkLplOwDw99YEGH6SmP0q71tVJhwAFo9K0pVneud6DIHQtUUp+
0B6Ml1YRhw7GsLV1GjOAnkovpJXti/GgrRYfakBBQRzqBVAtZLYoVv2Ih6rhr0ge2wl5jMJCGE9k
usGHvxEKoBWRq8t0IpGrPQmHRzh+/TSPsnZfg1uWTvfNZjoD33x4DlaR4sNiH9a28HcnrL8lMe81
/fXYo+xFbwH6qQ1ZOivxgcNzGTRpuzlguTU1nCX/089xGh3A0/577CfAfo2O/L9lsp4XIhi48pye
EdnHGv6knJab4eAJQoJ3t4MIui12TYofjEAH6j7pJ9vSp4T8/ZZdiNLEvDFpHjBHpQAtXARkBp1W
MYnIrnDM76TpVty5UwnL+Gv96FuBg1i8Omsk1d3Wb5RSOFnVocT5zczuwKAoUvsnf9qEhEvARDZl
rsWD90idKsQbRoEr38UumpP0Yyv2P8f/2AU72PmDb7wuDiRNsZNHf2/eKvmIsmmMQAG3WTF/hx+D
wOSEt5gbBXZBzaTHHmA9VzshIdnzT5/YV7vAWdjiuFX/zoSfp4gYfAUEgmYU9HtxfOTr3nIFZErx
z/t6uDXyttcbswvQZDDcf0byO/jorfUmbGDIB873c+QL5LkKUUGeKyXimWVkVmGiaxbae4kRzEQ7
8mUamgEqDXzIiUwqOjLpy8oZ66T3AqYwZU1IQaOovDZHGwXMBmvZ4+pt7LGdKAJYuMY/q//3L8KI
2Xu7wDJ67YK/VGHcsQn9RUo/xyIzbBuO/ozsvSV3vtruvZAEvFjO8sAkEEn7+9oljNfWQxpR9XCC
/St9bKAJJ9SIGOcZRdm/hJmOdD3Fqc3vt9Zfk57YczLZPsNGE/mazawO8XR28R93gS1Axq54tFd2
jK9abxR2gOhfmNjmK1Zm0SDs+j3BB4AAATNm5pHC4rA69yOAjsaoHPB62fjILurFmHvX24CL+YWt
GrTTQC316RG2kozcatF11Hj5MekDZJk2qQvu2vtDqzuqLeoCtGEZwDgaXcbW7NDI8Y69RLCsBRJS
wTv22Mfz+iO232CijkTWfWRgjGZZ5jaieFrEm/YQ46BfaCUyZy63y2BlAqLo7+UzQdLc5KqtZZUU
RwPGUwkYdzQM3ilZoFQSdjeeu0UkcTEI022HKSZdKKAEWl/d8+zpLi7rsf4Q1Vmr7dhaHY6dh10g
7mbIWzoP/hFtKGYZeY2BjMSH/Je03XgQlCebQTjOzl4DAITghUsmHW42zcwV4hyMC6am3l0vQk+S
rPzrxajVs9pIovT7VJnb2gCIh77h3KNXS5V44JZNGK/cZpl/gHdLSUZRuLFx6d1P+Da3b/OmLcYX
1NmjdcZ3eiXIb0YXwVPoZzodqgVkS/5xUDm2HJxlAZreNvuP5X0J1nE90UZYsRUVj8vHuP6SPV29
o78gjVoY2TV/LFK6SQPCkTqq1yPrDvq7StxkBs9WfL+vRYBE4/tXFm81tcTSgTu2DujBG4v0nJHB
7GLtdsJ9qPSGrebQr8PmfHygVR0y2PWBaBxJ5c+kmGaQxw/M2PCfyIG6wC60g4/Cvw8yaxmY53ZV
G2AEImke6XJ6kIZpIhL3gnLDqtvpcUwMpT8vrbspPPnZmyLFMRpauckTHU8M6qCslLSAEjVy7Bni
jxNTdbIWTcdYgxwAqh+27llI5pZRV9VCpw63CspuzRPUg2/c0K7aoxOvUkNTfcQmsNoDNIPHjRjo
p18NCweo8j5pdHCAUqj6V9k9+z7LVykg2KRvakJmx1ELYKzjgOs0eht+zTT4QmPVEX69iEl56nry
U85E0s/iLI0KWVvv1YM6fHA0K7/2TeG0sbXo9yNNEQjN30jVB/yVIcVGiBLD8E8vsD91T+1xepDk
T8EjNg/ddpTIFrzOgQlOPDI5w9UFSkkwf5wXYk9wAfXy7YvTnUYYlycBl4nkZkbeI7EbCpD6hpJw
nsQzXBq7ovVZjZWXl2QfPNQXsLdAAeoR+C33ovmXuol9Bz4yNN22SoWbeqhQJlDpcTQ3dKYrRdEx
IrBO9MJT5TpFatoVDiU+VgEdj3oe6tmwe7VdbcN7/wn380GWL9WT90H0cxRyK/CaJn1Ko3Il4CSq
2ns/Opv8NdNF9ePG8L0Z7peI4+umD1uBI6SVaPirp2HUGpjCqYeONmeq7kBQ3VTv+rbIrPe28bxN
mMA7Lalr5gagZAdrCH9ocnXuT+KugP/htMkhQRfbp++IAWA+BSha9ESGYW5v9RmyjTfhRJLa3UDC
hlYLm0yK545Fj+Oeff2XBco/yDUt06+pEg9ooWJxIpJR6L9SheLL8d2ZHkX0zjF/vBgFfx+zQ9+i
/rv2H3ek2PrDTL6ONmmaX4hqPeuaMfm4JAtyB3A8iPFs4BkQE2rfPPihmklF2IIWgdwDAXiT3vLu
im1oJSKQDEQhsRAdxN0+7CIDzjLrUEK/XcZ8O/ZhgLatdYj4VfgJOFNry78NM0RBMLcVm1khbSFZ
GDNOQHnp2faJWUjBKFoX1vzvHp2QbwiBwZG31vYTsFC7N4xFuRfDv2BEJACKgKd+doTjqjZqEihx
L15fgBYHsvRTeurtic5edjzr4M3dU/L8LAlZbQvL5WZciCYdtm01W5XDWxYfL7QzoqmcFXK4kaUJ
VB+MoGrhqyzzXQ3X6ZGFZZkJCzjxw8PSYyMFSSsMxmndxcOKg4RUkGCEsduRah7n4Sw0n9GDRACO
Ey3OI7nopBDcJoiQmXYrg0NeOa586wj/hBUCu9iZugJUI+iaJENiMGy6FgoUBiZYp73vLPNCJFDg
eoYXU5FhhWL8DcMPqkbZuUGMjeVGNqhZnq8InM8ouUJ3CYIcrPSl7gVU0/4sGuttEZaQ0MWH0AUj
Z/n5FeeIHY2qLRJMQVaP0PeNS2OneGF4BE0Fu3JyaxynxLVjf1reH2ufek7Pq+BgcbmfKkbU3j7O
7MJnxHpSW9cq0jWlTtcqbt7cgSnHvq98fFzz5ykJ11wExWcALVpe+BbnP2UgK61KY4R0+lGsqXBG
lySNDvubDu5Uiwm/+3c8I9kaBOPZAxwWUw7pGuAvUpD5WqTYmiHK7d8CUTiuAvXM591bj/BG/SFQ
h+19J1YC+Lqwyr9kaJuqgRU1N910sVkdsIQfgYJG+XFJNShZ3Um98VUYK8zqWHkpKXiX7IAWSoeS
Nf9fxNmVAn6Sbev5ZsuCL2bNh5GtNIHVCXO+Fyx239BDZ5Y/jONFbQpGnBaQEksOURAyQLe/pMhC
us5bitQEPRtaCkPqzsBuhKj5Nk7ZyJkZRKE4EKELjzf3mV3T53FK4WEnaDFjODvethllSRswSgUd
bONG7leIK208I6Swbe+j9baPT28wlzgOhQJx70LRJGt4pDthqooXQJhwf/DghswC76uQ5cTpAjOL
jfBRFW62Dh6psdE2lilr1wMEaM8BEKz907vYHcnMSwdxVl4HySaCbCBRpZMDdr24JsC4aJWidBK5
fAwXjHKVSZ/YQyBCkAcXV5DRvjjoueimihXAKbB8YaT1hjX/N8iRIxcJeUgSo1YAOJJ+1waq2J7U
u8jFBV7ns5NIVM3TeM1V0GkpCpSF5g9JDEmv+kmztEa29GhIYmv0q6KR+LJEVKP5WFOrouhPia5L
+84t1usmF7Iqlst8ev4tpKDRmCcdiX7Y79jG3svJBzcy6rbmyGvtMlGZI6We4HqGUQngqm/6BgMY
SSKMe3laLLF+cYksIPGExFu6FJjiDhejhoajrLQVsuM5lj+ir43tMa7ITNI2FCtInomBuyqahu6g
J2RvdmeeuSoWDW1EcaRxVQDmpeEOClxMNm1/LWa04xAfReE6tid7aVeiLRMYJDXDkgmiFwyLp3S0
lKviCeNEIMnSBgDGxzGwOs9No2uTMusBkvaMiBJdtI6ceX6GMbPgQ1HbBaGs6s53ypp/GNWKlt2+
761LIJw2LUBfr/vGGwy4+PEL7N0Aa4hbUrVe8dn7l8tyjmIajPw+T5GhHsow6yu/AOs/a+igqLGD
XO3JxcXSTgFPBy0pAxDAO1yaOF47e/b2tZKH1LBFS4p/cQ3dn/KG4BnOF7VA5ayTdOvF/AGAO2W2
3C+5Cx1GyHQes9nYaDEt2aDHBMXV4yldKVb6hwFnhxvvNCrWZ00ko2uiDdUeW2+5cWtRb5/tOqY4
KnTBp7xb6clh2EORtXcS10q72WzhpdFYJI6nTJA4zoF2vgFi+Zal+UmrhTExNE6HdSzD70q6bLzu
bUKAzc/BvAiHkKeVS+PwiRRSVngEBHFyX1cXOqGvKKprNu3jMTVuufl4/sam2UArV3abYTcgFEiU
AkhU9Y7ILs08yTL3xUUyG5K6i5mtmpeS0Zy40voVdvbpM8Lu8uoU8Auooywcm92FA7gXnyrvUrZI
vEnhY83wvpOhgzsu1gCXvYf5MhqbOsmCUrs9iSFH9G+3N9Qb8yT4FVbVrrdBpxvljXT5ao0hdkvx
3kN82VJFSxVHqzx9oeGMu6Z1VnqG/vC5y7jVkGfH3e1V1RA1few0W0F8p90TnAYAGoG+iDPQkKY9
SwrBCwILf7sAo/Jy8Rx5LB77oGN8r/CZUlH3IPV1p02bm0YWvEuArjz7ElF/4ZNZQhGcYLKTdL2I
Hp3VdLseqevY0HDDP24a8xs6+unaSw9SCEGaioJ9mk6yEGt9KCM61+Nyr4+DyWi4rmy0Y170Y0/u
WAb3NNWjjSGj+hHhQQhIXRUS8GF+zQZ+++kXvhSIX+Mj7xcEWIpxdRROFRK1ru/EftGk+/jl35ip
PmutWnL1Sv7niPistUZ8EjOtE8pyrV/H2lx5zfv73MryaXNlVZH99jxjfZ2X/5Dv4W7yK1hrj9ai
QW/l/5r1h23f8dqWhKAd9zT3uU8QpgDvzHqVrqqJ8GiH/asC0JtAqXIR/4TcBGFc88WUua0XcUgG
p2w6f1302CbQ0VpARLUigI+1Sr8o1JGA+iL9nPzZtwNMWDv0A0/uSit5TZe9utSGGysepiDxFULb
sTwTFyG8UgTTh874Zhmf9law8VqpXOjklA+133Po/1aMMFom9n9JnSB5Q49JMdluO1HihAnKeVBM
b3tUy+AxJ6wn4+Kv/uhheqFRQGHDWhC2lW45p5sMpw+OXxOE4WcLTTkIYrPE/67xcBEzUimxHGJW
JvFlEKZ+coaaRL/FAqNBMvWNmln8jzNIbPXYhtu5hkEWKMJsE8f43tU8YzP2iORQS8fkjmIDbtd7
fxQ8pnvkOPRsu9j0NNf8MRzY3uNbgIZIR+KvUYtW+QTq0fKVdaDAK4+KA/C5AJ5gK/w1mMlIOgEd
cq7b8iZ/zyzzVdxcYTCGn10FWFHaJmEnAjZoMK6UMZgURI7QqxaMDJ6jTw1MYk48zLQ2lqp8BPmZ
tJ856To3BpHOfxRq6/YP6l+yYNDJ2MjmYFV2M+uFn48jPSWRe8fD3/l1Iz25vVH/PXOTFXHC5nMy
SKLvJ8mJTmhB8mjfEm2OHvtZfW1Nwmk/tdIY2aqQPxw6eVUTR7nDj8LM39evLMtLbr6+nAg7sR1+
+5g5dZsvfuiMMUXps6Db9C4L3NYTHUE6jEQterATmWVMtRkawgKU/Er0wWLxcbjmiroGiKhmPZpI
uFpYPUXg2fIybDE1AO65NxjtjoKSgOfalj0xtm8dHeeaiY61bErTcctmkRsX0fOV0qJKBmc6sM1C
9c3KEn467XZLTsTsPB7CSiJkoXb8rUnnjMp8NU8P0XI4oe7Y9fWH8rHmhCLnW/QFJgvl9vWYOEVh
w/gO0SNjP3MTM8yyQ2pJZSnsRLYvoigBikw0WtkkHXxSvKwAseKN6Dsu7zkh4iVUVpI2dj+RRFE/
07iXTvEBhje7MFwNvt2GWeImhEVZaUGKLzEOnBJPTf+vVuDgQ0CwTmxH4sOe6PW+nk5ZVhomxZ9u
OzrBTiz3zeK1RLho534dL4CPhuC8HCuqvUd3zoVVOiarBna35+GTppr0kVVSijF36arvAmMCa6zN
kDWhxbcBBLg44iO++8P4licLynxyncsv0lStIri6cWgvo1Yjc9Rfl+nroo7xJZ5jXae0Z/D6yZHp
ME+/M+yicQpF3w8RPEfR5Qq38oGVOuRDeWxLJevm14wTcHVXNLeaJQZY7moGy1JKz0MYFnSw+gtT
2KM6CDrHGCMTfBEvILXUA9N72Q8ubcUcXBFdOZ923y9dvmDhdgiu7erZ9OyeFodn0UQ2vI97nAgj
0AX5ca79Qh8e9OMKmCm7GXU3NZil4z2B8ArYTybHGs15a2ckRR38PRJBUHKBUagCGp9cd6P8P5F0
2sOeATtkOg/9yMCKSQufTpU9vb7ZQgHnuJb2jmRVgMScRGCpEWzkl75JvFUjpKORtQFa5dvTGwbr
fFgydLNWhX4MjLC0z6vTno87aCgYr6b+H1ngfw9AG8KEe6+td4UnULaXgk4DjUcnJFWYNHhkHaXT
M4ZLbTQFCU/cizrev2OJqJWiZfpnF1Tw77HG3GSngbHbyBrWDgaT6/4Py3/OYRJxp7WyScnSLlJU
BddWmWq6+YOsv8L6LPtnzzG7xdoDEaxPofwZkcdV5BevLeJRon8W06JytlyeX0tztRz4uGUrS/8t
5LIn1tmrt2O18PVf0GBOnjdU4L69DmFSyTM3bBy15293zNh2cqkgl//5OIT+c+JBW/kGNfwdXmDT
IRZM+r6gB0hErMmP1c0LdK8r+zfgUoifAHBldXpKMTPDsFGEOlq8BQktkp1+LmOZIbBToE72Y6L1
nZZuQMxUmJKXE3NBAhOpSppxmeUqHKq+mq6psIQbs0FbcvXy4LLbZ72Km89jx2fLENJpFRmNAfxy
7BAVSE6oHqNBO8ygFVTOjFW28i1rA4Nn9tftfsg6vUbcepxl9JIcLOncWj8YwANDXLuC0DsOOHnh
s32liVjDq3p864oQKLhkUj5m48LD7Ip++KX06F0+kh5xxuR7kO/9cmCPYHf2kCMLqe8E7YlD0MDC
frmlASlv54cm62qiozI9VF02gPQxWJuCn9f1GQE7iWY1x4t2lMkJUFKiBJhjzlSZzfM7+Qh2MYdf
SMm04hfCnJL07ZGBXE8NzptRKIIKeN7mFST9TgaVp//zyggrnlIXDVUdkGj9q3otxa5sX8X4WcVn
6kLSBnPtgAi81YZBZG3a/8NnupIXpG8sI7RddsDz2GhHF2vMux4MahaCrlvhWM0Md6FnsceqhIkM
fKxdjI5I8jVA1yyxgp3lMvkalPnMME08JCLB+W5tph5EFR0hXtXA05joAAb22QNBXTQk3noYyrnD
pOx1I5Ge+zoaa4a/QHSN6nQbD1l+kPJIViH2m1VMtVh96PksE5vCxuYaNM7rAp4CxEytsB0eEWbX
iJ7WMBVs1dilrtqiXna05KELO14OC1FCPHf1oKGoS24J6zRp2nuC/3aUD/d6FJ6aUGrHdjFQja+A
kqRqP07Jgtuq9Xi+2DX73sdTQ68Xc3dOErPHFtBVJwVTa2pRM/LPstXojURoI/dVlMQk2va4x8J/
5vGjbtGKM3dIq0evrxqsgHYnv+fT1uvH3ymUJPmsqz2VUjJCam1STe1Mw2RedSssAmSxlohlb0ux
BdDpR2bGQ6G0cIkB00/MLQHrw5nNjW/48psbL/82pIzSNkcOccKsQitoJQ5qgCRbLipj0h4M5uxO
F6/CeB0rPpoM6Q9mIq1OjpTBjssjip3vO5IY8tca3xt+gIfrAuX21Jpg+Pl3WbQXqBilYB0a/fQM
xDOCnKzdjqNkJEpSLi7BDczmvvOD1rcX7uBlYT/Z4zXBTNk12r4E2fXtDvCgV+YxaTyoh6zyxfXT
gSo21dnsybGBiFvrLKwywAgMdHM+T4QHOI9B2jO5R6k3r1bpjNz/eOzSUwfZWLD48H2Zpmd6fRw0
ciSuKwTnA3Qq8jYr9IXZ35Hh73ewbwu9dxZM429rTy7/+BCcHoPxU4r8D2avQfpLthtrkBS1DGK7
se1SLmxYlFp2Dj+d9crfyFsFEiES0a1t3mPKek1DPI/zLERUvEwZ0c0e9EaFkvX4MvoBvjC2crbX
QgBEm3oSimy5yVQeChW5LfqC1tivzY5hdCs24s10yCAhJ/puO/M3XIFzVwb8H7NLN4VLih0MREGF
a4RV8Rs6yBwW5aOUuCN3mKqLaaCjWiKWXFZ2NPTKQaK/Y4npQoYIOPJ4fNQfARF6i/tqrAiBa/iD
1ksYmCE+DGz4IBiMmBfANKA2OllGMghQBrhVVKFuYjDVLgBmVVtCGoDAA9LCavu5bPvBdyEGpJRQ
fYKnOLhk3wlSJneMm6dZt+yNROYn3LPjdd3455i1+Mq7GpTwczpl94h5aQrpzzfocI+dFokil9ey
jRoifwRbXVqT2EO5Gn831zn518JWpVp6Mlqgw08+6KxcnMNPFT2HGuA51mfL1hEHa+PGBdXzMwTu
ZtzxDaDUdlVJwKChxXrYOIGjEPDBfl2TWLhwYZNzQI5HvcN4bvVJZaaGFc/6oeVHVn9ovURwbXT0
rQ8q3xVg4usglGajutftar2vpkXk7CmWAP3yhbUa1+TTTgCu81qcu9EPDrUKLcw4XvMRndTGlSGv
AFaZae7OwcvPoBqCnJI6+FfL78KCSdUF+j2qQfx2z6MYX6cB6+4te2UAk2z5m9Gqbk40MuEM8tiI
NQykcyweYUJH/hNLc6y00AoOu9+F4XJYH/nwvDEu8cdvHHEORG8JmptcEQA6xgNUMKovUOGPMj7G
4e0xcbSAbBMGGa7rHN7FPBYAD6I8BmWnjzWgylXMlh70rl4CpzU5LvJWY24z6srljzjQWB0xifQW
NE581xGXQGxlfyv3/T4nXNrCn5lcoNgH7hlYAk0GVD5vqVSJQFYovh6zAdHK9pvbVZwFn2WEw1UI
B5jl46Bq6+gNFD2/1GYRNIoSqLBmJYYCvfLKkDBpjQgKEKqINZ/eAtlZiZCIkf3F3PJsjXU1QrvV
0VGR3oVOwykMsRscfitupsZw/vE5aeFfAzWb2NUN1BJ4kZ+YVAYZMMDrG2mniIPvj6JB/8QfIhQd
Kz7fikdtjL9CGwcyyVUV0k+WMSAQExnvQrobKjEZBbY/kzfHBLNpn9mORoRvKuZufYkWJt/Qgg+E
K3gnK8dQgiFuGbnW+lufl6UU8ytqvFlkpUiF+CPFepvx/G5WhUNGNr/+O1CQHieVluMNaSw6kEmV
42SxyiT6bxYIeBiNMI2zjec7A7pTubID2+UIi8NL9U88s3zRjCobkyVskBcFCCiXXKvB+RJJp7wo
sP6nFOrq+KaNHYCZJER3stiRSv7dbvnLxbMfjo+ExrY4Qz6kDS+zbOqfCb950aQeEBXbTmxibmsv
hcTTnFz9byTquyxpE5/6+fkqjMgVF/mASvdCoO7zas41LU53UfPG9k9LzRjHGalwO8tAbLsxIKYd
vnyLWnRnYLea4N3G+MAt1jRUxLdpqJHXCqn8G36WVt/agl4XNgyIhXDvlupTYhbqdbkh6LZmGE67
AnZplquBu9oJLkFar2cVVoXzVDCQqscrjPD8N5oHb9/1gt4RD5XfQP6+6sM7Lwtsp4qgYCuzu6ts
p6UIT+Zo3kPq0fc/kJYtTn48fFKSKT5+zbZunMw14q9Oi9/69NxOnPm2QYXpykiOJfUXmh7rEEHB
geLEfT8XzYIK3Z1f8ZBInAZ7E0yiL/7cXe3smubiblbdqN0pdeTvLs9LMOb8L+PWctRCZQxFxbp2
xXr/7PwLabWZ/AxfIxtgCLzrEk8aGzc9qQ9tFHPK0ebHXkdvGo7rHqgZ6GKmUVKN7B0ctJ38nJfr
+iQVKxfkBKKlWB/ON5Ej06n1gH5oi3+G5t38Ho17zpBZvWVzDHCpcfo8HcUWluP7SCo1KBRdzhny
YanUfIHPN+fweOtSzUDwzeo0aziV+yZ/oAbJnY69rTx420auutFNdp6ga9gNumA1qNr4LP+7Ky2N
W1dBWyZ6CFfwY41AuHR2MTBbQhRuJiEoIfmuSCT7h7gmu8tEp4kER00jD9vbpwsag9FcUWWKdgPg
fr865CAZgX8GPXzmCkke9T1Agp2CpPyHtO4TWf8nCasTkjqrUwEHKmVyzXyBQ6FVr+BwgwLV+RoF
k4XYAdubWJHpE8QESGanN1vwUSSXXPU/Pzp72ZijhBgxQVym6dUKFo65j2Pfl/lQaDAgeuMZ7m+s
JS9rK+d1YhaWkgnwcgHCUSFULF+WVeHJlz8CRoz6EmBaivYC9fDR1h+riZspvAfUcLlxsfjF1kcq
iU2pqb5NHJdh03ECEbX0w2aTSDkHyriZH6xtnHIO9l7rX4NFjRGS0XjKbyp/0rPWRmoqHPAzhW/q
ivbmqBwiRfVQQ8rJoSVqbJpboJBEZiQAalH3/U8CVUT/J5TCwNTb4QVHXrBCB5042VgPB6lLvxey
D3qkw+tKdFyvTKD0lnyb1clWCWNs/WPejXMIKyGZGvybRb5Bc5dRKJsLLwAlKDm52Zlmq8/MBVKp
RB7zvvwiueFTCQfBR48AFIdeW2FqgUZ8iEVbOaU9pbjt20lBfuZiM6l4xulwQbzV/oFb27udjKed
7wt6JXDKExjFoLM/yT3LUyl4LJQGpUVbpUm5LdXl7GpeqGZVEb/kxlom2EgCBLjPT+0SaIUQEz8j
Sowtt8EnSWT6s8cg1RniNzQYiCCgq3VOPquTU+EfpkX8UQv7pqZhJ371mECKORUuINjcFbNpply2
vp7HsvvKqs0A1uBc3Ygj7nkulKDFNY6pAtvLM+38cNESI+0a0Sa+aGLBqigeybih+BJY7eac2Cei
LBc9fEZn2RiQch+OCYoj5W4jq2tNjrWCMdJwK61sR48SRePH3KJ2xQ+YJcpsP4i9DNMEEb7qmGXR
ELQui9cYI12KNFRbH4HbKPwM+eZtDhNFYJGLEqagjkXCyEptGbiAoYEkTHNGTtZoYyIxvePUH0NT
Afl3Gt7Z9mNunAmJhFoQ78EqgM1A/rL0+gnBkpSqU3C1jnw3Vi8gYlu5114JugbpjIwTjVRfqZlI
s0CLP8UtVuILx1+8Q0vH2c/hDcyLetccGXnS6HZRqdXwjD+kaa54U8KgzU0ciE/Rts5pFGyfPlX2
zk5Is8040wBXz85agKl63+mYyL3CXZ2Ez2nfQSjw7gaejjnhAlTWbsYdh7DemoS9UzuM3JuDWs5j
XnDfde+7PFg2zxtVWQvdmsh9SnRCDq1AFqM+CF+R2VC/MpuaCmwhrY3MY79w0Uwu2o4GIRuqlWDF
lhKT7Is2+Q56oHCNxgPwpbO0RFgvnLgMogTfbx3jenJNnzDtcuEvl8t05BN0+L1Kpo5gp3QL4Uq5
fesx0vmAguoPWIQNNb2finpNzL6un6uOAdtlWX/B5Ln67upyuBBok/55tPRYisvbkNif/ubqjcDO
cVJv5k1pGppZ8V6n5YuSAVzpHOSnxdjtapDgo2QwcCuLMqSNebrqYTCfrMyiEGvysPXQf3rhvZtW
c9An5RbjvjNnDIrscVniyUJS/wBYE5Kt3eZHZ5MbVPSa+e6DhA9ywE6Ci7xXMJlY7L+oyuR+kpkK
A/EiUnOHZTj/sXlPaCYw0qp9GdmQsd157C2hQzzJDScCzcwaOMY+oBnXm1KsasEjFsw5/LnhhJQN
rR4UvllEsqXR8dtivbpr5vjlFg7lNZtNuSYQOn2Qiob+b+SpmmLE4Wfn5XnxBOBigrrBm6sRJcTN
2vHgtXoWlKBO2TVfA9ZATu72AmIUDz7l+pMzmOxfgDZmO0ZQQX5EivR8HSy2qh8V8giKceEQxH1L
Y9fkIVrLopo+5HSG3+7vL1PSnmsb5kCDXIeE3+wqQbOAdH5V5AUDJRa0GpKXZj55ID2UwFcR8ZDD
Rntdntd8utahA3cqdqMlpoUno7RI7jUQmFeOAfk/vBntuvf+ZlIzj9rKgUBj6rd/GN+eUDwROLDj
lYkuFmtXGw3KhY04B1yO84pAu68bnqFtYfrNCy0I8QzeyLGC97Z40KtQr5EcSPCD/rDWzmFf/iRs
azMd2RTdsMK1M1hkqwxrz+e39uIdsQZWprE6RaUiFUyo2CdzniSWYfLwCHU819ub3kmFmgOGevjs
PdfsByZVM3wEXZWCFAoI5DRfbRuzQ4080J1rUwuE102AH/oC5c+oMSU26qQ0hyrnU8e0TnttFD3e
R5PtYsY7V4y8oMgGkobEjJS9pNVteN8ot9cqQ61uTy3h3UrWLvEg7+m6RWrs/PJdIDu26RbhbOgn
JqDusMo8NmlooD88qpwCFQuhgVkEvF3waERSxXezZiMZkOIS1ZRRQvd2DW+W0nx7AlvknO9378LT
pO+GE43ivEeBcCERVj5SBj4Ozj0INiN97z2EMs2fOVLsSSwSUBc5Kz55M7ulRxRUKgDA+hmQ6BmD
8zMR/kp1j1EB4OKvuR440W35vNLQ1YRhwBqy2L1Npv4vfYVa7krYixhrGu9eKJVDOvdTGpTn0kRX
rUYpxXcu68qlUgzJtctxnwZ0056/pRszlYW1PYbm/luY0UH+IjGpzjzY12fooS0/b+ycoPUhEfqf
0Ns5/c0mSiWO6w5qHOLfIU3nrLE+B/jbFwQ89DYWTpEivenilMb8g3jGvKMGIidNGkQ8zg14ginT
hC9mNenWC0jSKw16im+xmoyJP70w8Bo6LrObut/FK2ZyPDR7R03qlFxl8XzmBLd4znS3fTkiWluG
u/g3n7S6+C4wjQEGKs6KcNePpVe0LGdbBa1Ah/Et6Uu/VW68YRHwMJOW789kKjD/n85FxkUT3pAq
LL0HWM62XJl/tvuD1YnyVHnltg7DscbvlitP4Ok84KPA5IV5kq13X/gaPKGErXzcEqtH6TBQdRQb
KX9z95S0uZFzAlEDods6LjnuvpHrQhd2WhGI5aEv6TtymeiQ/oEayo0nCkVKnpwTC8TkZ2qFJv/e
u+AvXuJ7DHbCMGb/nL/pC3XpcvGYQjWZjOjWHpZu7qlubejvpXNUYUTp5Huks0EFC6hNeDEx0jDc
wuUCsIWxzAVM/5G3QFRGHKdmhmSj6CIfHODAu3tmr6IjHACC0Ob+ITixdg+uhXB+bNGSflfIKWG0
Kug5VtG76g6DVOxpGeWmYhR6omE7XOnyZMz4Ub15OhCuhKZP9umVzfMSu1FRlU3cFKriXP/+zHIE
rbCQvsTRgj2aMd+NfVpqIwrwlVD7FrWxv2KOmz7+gtMq5HRCXvxJY01x0dnjNg89EcmlwRfuYxsj
ghCASBmgfDgbL5u0yzrRvF+Bvv6lNdKZNuclgaY/0D3x/z7ujqA4KzKJcVXXSapStgZA//LmlXlR
nzUls0TyHQCQSCY0bKSPwKmlOgUTcM95iMu5InuJoIS52Y7x8XzbjD84J/ldeMyK9M+q1TyAHBiI
IuYbivVftQhNi0ACHoveKy05Ekjf/Jg7fOtzCq80sWV9SQ8ACxydoi+ncJmrzAo9dr6PtylMtba+
atX5750F4ZQ24R9h3NI4EBjtVV3V4q2IRPhjd0e3OX7+lxROSBGARs57mxjXRSPCcfUuloZWS2Gz
H6ld31+yrlzyHrp3tqw4UKstoYRxddB5mV+KjukGHqEqCnh7ywINUSBz3LiCOecr0D2qR6fmRZ+0
2yL0fnyIlZtZqJCyhV17twWpRhzGewCzFQvmqE0hvDPkO0PXfF9YE80XXDrRuwnuChf0tLISEyT+
F3lL+2rEP7JU1czRnJFNKdXIYWCxIbCi8eqKmInzSmt5IgParonr2LzWuy9Lo7FXvoxr8+Yv5PMw
RmO4y0QDyUVCa0bnffwbWMiN4gRO8oMyDG31bW0cnVPCC6X+Ds8iaTg8w5sfAy/gltAtceoISarN
Jg20b6SgBU0fqN16ezRytpREevFkYDG1j0EIZNwruXffFgwqSmbAIdEyJWuIj6HVGetmLMw5v2C1
waLCMHmiTC40ILU4wKUOaKwPSY4sifClMYV1IOvhRk/2BmmrWdsisDwfY8uxH9qEHyOe07YAdwLM
bdBEgRQxhRWzdaOT+tXk54mwm5YfVBH2nZkf4qIfcTAjs4O5GRm0D3De29msGyrohP614GPnt+s7
WKtJnoGhfTxQtb7q/7wQ6Hfw/83Ey5Kkdn4hP5XkMVnVKRCx0MaUocANMRXgykfo4WH1hUCPhIA0
2sCCBqPLujIAvwlxjdkRtw+UCamIvXt7GyM/JHD4Swid+kH3INby1Y8ZQkFt4HI2vdAANgVeNlih
lHuuLL8yBJr/Mou7gKv6Iu9fc9QRIFX6oSd8NxSGzILQKwI/VKHcuVzqnqN+Z8dc+IE3D3tqFn+V
vAq8U4iHV18SapcwTFsX55a1A0o0ioKVVD00ycoBJ+nq4QAaHWzjauSOYp7hJc1ZpMuXZAesGE7D
bnwAm3ufuNN7+Kg0gQt0rY0BZwNGwrjOSvIOJKht4/q6lAWLiWOllidWQ+kPrbsi3C38Wvil/s1A
EyFF3SY+5bhDyZclYPFE69gmxWDAzwFAkkSwsDB1v+tSfQYZ1uRwzXp32KNBGXG8lliF5q9Q2Qq1
SJ/9bR6LFVk49BthlNpy0ge30lqZOUwNQuki8Ksg82M7+trsh50u45kE/HYqfAF13GvWDnRFwrsJ
hvrQOAIXWS6QX1Eq4ISu3LSmp66bn82iSrFPbEWWQSh3ulgBPOAJog/qOBBJnjAXTc/gkhsK/MyM
c6AL8BN2vTXcpT4PFh+hR+0CwqJX3rhd2/KXSyjUhf9z7DjYCKYvDd94nQVpHXlXwIGPWRjfU9Rt
JpD3GAv9+d3OxQbmeXY+4SeA5eykZP8r8Rt7ag/oOekL8lCP2NEGs7TIYeELky/uwcfmvyyJp4/J
jb37roQJQ104tW+BAIPgBlafKkTY5XKliYqL/kk+MPQSX/FN6FPkPOD9t6pky0w4SnabZDUs3dzS
jqSBC56tP82834qZACXv7a1Hg8RZt1FmM55ljh4ihGqU4J+nnlAVmGl27x9y9FBFgf9eGTS2dzl7
H452GnzwVWYgRrviJw6nKkBwT0PAW7xYpgQ3qbt7mFq1TtZKhf0TvKqNK9hRqZ8cd2pSvo9Y8exG
GNQe0wTsHACr1PGgSjBTVymOqUaMvRqX+Di/B7P1MZMOWPt3G8MKZCzjGZuFlnk4nN1YvxC88xGr
rCB/DpOSaEpqeG05DIO3E4rR7gy+MX3KFrQaADHBoae9O3szI6cVFksplvZpsVroD+djF7Jjd3NE
DjhI2TXvWgTaFOLCPw1HwfL2ZT7BtigUdD/YWJWCGFOFvOSBx+HIAeZX1C8PEhixJ78wnAg1lAAk
wP5Le470tk3XZrCHMfpUgXYye4RDkzYviODAwRMUTm7DzT4Df1oKo79dD+lWfNtblNTaxQM8Tcrl
w0CfzZhIpa/eUEhMYk1rILWtymBAXV6RB3hbiujLuUtUXoPE9C9YI+0mRoLyL8qiMDAzrCCGdu0a
t8yGBfeL4LRiFR/EjnUGj3gDn2glXzj8bllZLW8XkCY4POOiKk1vw6ur/uwL51Jldwc6fRtR4L6b
RKYl8qc44xKTdfrr4u09WTHVlUwBxAdQhTYLXok89k/pSW+7aa+y+PGpZy0fdDZCquYzQMVqoFyP
7FyGNK3Z+2E4ChOQpyiM6/Ms0duSQxLmNWwL2baAx1kuoxVnw3Bo28Mpa3sEibPv0IJQzKwLvQZH
r9jLrpGR2fCmd7YGlIUJ0jozeXOHav7G27/iLEvGTP5JY9Q+v28r9SEVpasqwwSk7QubdX6IgEGh
4mP8pa1BIukIRQWvtCMiwflFDMtexbfZWdSR7WLqDEwNJg80KUHgIsVK/Jsk+SFPBeHYBdeHb3mF
J11dqsgOm2l73XQvQwk7jI7dadNEdFLZmPGQMSbawHKTAAk+vHHIF2629aUy6FodWorTQ/R7jbkr
OOtRX5vJTIEw382jwFJXLzOqaRQTZmnlUt4zVHau2IlbOHwMYod6t2dblyx2ESlY2/HcVMph7Hak
HiHkyIwwMDZGBYp91os9mOwy1kHOcV3+5QXGdfD6VrEf6APxe1jGXvuKm8A6wzqSvKI0b9NXaf5D
p3vRYGxQuyRFiiI06+GqddI60yok819i2EPUOZCf7hQoE6RPK8OVZpXwEqLF+50FLzh/BefGEwSr
jxB4hv0oC+KW4GPS4wEOL0syO2RYXF5KOsjWPGiQyzXOdipynIv+5umM7CwucIAlkGT1N0+1jw+H
S0wzEbsAVTbNoEFud6QzAsHp+YFHKCI0496aS0s7v4YFBRgbg6lX0zr4ckHdrzdWQaP57qVw5x8i
w5MzcrOZBTPx/6cC3wWS7WcE0eAFXbPQHpp+l0tGaBEu79S5cF3LIA1UnQvx3R5+EVO8uXMR7p29
6yVo8mvaiRZvSPzOdQS+xQvmy9thi0pcqBGVfoFzXIA+IBQicuZf9NYvwEX8iWfg53K7ey0m/Q0B
t7npUlErsD/8M82aas0FHg4Lzcu7DsKYP3j/XFxYHLJMZCdPMn5wTKsUiStzi3dUcUOjzw3BMClj
A5lOvevX6mCSVDKrbfQKh/fwsO6U1K7WkiLp8rQz2rctmGoE/8eqEucsEpxHteOO57LmzN02mncq
a08nu2KqSER7y/Dqa5EJdW7b++rI3yQDU/eMJTo7AjPM8LGJp3Cs14Gjn+zkhIV/ulRewbOrqFTK
z/fpJQYUKNpN6oiMp5BiGMYrITnAu5bi1s/WcW85fQBrTH3GJC8PIOgldxnpoMZaKoSPHhNVgar3
uzprHGcx2U14QXhqKRbKi5Sf1boawwEfVH8J/d8t266NbJV81tEZeXoNJJEAXFnbqVWOdV0scRfT
Ar7jx1Tn71nU0/bv+DgjmzsakQLMCc/XW63mmnlrw71X3DvQOOgDhY3Hg73gw/N5Sml1JqFlN2Mz
p6+x/yVRio629fmrIvo4rvTvhDinL38neoSXKcDVNvQabmymeNATKj98yIryq2Uhib3uk8DAby5s
5l7M97q0pVOAaru6Hm87Xsp03xVr3J+gPmcEpq8SZqHWfYiWBCAdsaUqkl8ghtGIcWJJQyy30q3Y
oGO/U1z9sN6Knx1owwoOhQez8UkbFiou+1J93/047EnXUDC6sWhUNAI2tBuEVHPfD1pIvQEjnpOG
GsIz/uzpNKtzhCLNS9hikk6o+uAbLYYEhCKvTuqCAFIPBToNzFfqvPmw2GAoLi93kMYFsBQRqjSG
nS8kU6h11sGbG0gqSl0IKuPHMVL8j0/19csjhpIhC68VUBHytEvCdUw/tzdKIjJCFsO+F2Y8B3tI
/2CENVQe01JwMsujPHAQIwDM6h4megvIj5KzIvNQY6nl1uBlHFURZJakoOpjARzwhSCizwSlTqmb
tNGgDPtMFiKXm6jvbexIgEOWI4QeNy2gqux0eIHaxtc/FphkdiMT6A+BAGUV4y6XR2Vqf0DLPWRR
Jay2KWpWBegsDmBSdmAVxSPIyuYkxjyGwnIz0K7ebdlg07Ru7+lPz4t5mSKIOEW1+Is2NA4M5GfN
w3Nj++HOCSbR88lae3Lb5LDt1hRKfA9QAE1Ot22HFNFlQ1XJiYzPqxEwdXc0Y6mVoeI1tWqMt4Rv
cGIAf2yh5M3XicRfXH9v+ic8z5ZOUHwGkxDoxCeFNyt73TlPhGKbMBT0WDS00Id66JCw1/L0c7wY
5MXeCrFI7bZOOaZNPCNscP6AlIJWy43U4LhiwJ46xcUdlE4KvHN2tmDZhCuZMuRgcnJc3h6/EiZN
mVUj7Aycqzs93TTiBZs3GXMKLkyXaYUIfIMHw6ky4iM4uAzqYjXS5XeQ7puDqcjmj5LZyveOFQIu
XqtsTwzrmHzf2epJHoFEK2EWJAeDPSMQ9AlUjOWNsQXMG2DaAuR5sqkF3uiX+XYFWw1PSU2yHP+N
Bn58UcUlqUYLNSCJ3Kf3zJHymzaBCpTj2w7DlCD6HXnUSyoEx4Le94ETV16QDsCA5Ga4ytQl+gYu
LlPdfAcmyHXTCo78fb28jZeUo/2UYf7tDylT5jfV9HKd1Queortgprha8Llbg5hnOJLcnG0IxkeX
ogLjvYFOc0JLWtscVL5pibVMklyErNyNKxXaiA2z+v/LriW7g//nEOZ9Y7Js4Fzyq+J0hR0D5mwy
ON9xpgdesGkX2xz+ra2FgjLZQcNgZ4RFcAKs8vU4ASe1kiHv/ga4qv9Jbh/qAxvxZrXLdXC82jiM
rWVgVtArnw1V8gYVKl7E7Zr/UObsOEdvHNDpR4UIwVyosteSTP/gCSl0x0AWB+8odD/IdaoAx3mT
/Rf0L+u54UIcv1DB9SIHhWSP+mC9NAZ30D+5a/NQ36SLBjOOInVqiw2lp7yXLUJX0hMvBQxL+CAO
5mrahbeIEwCAIR79NXSJRizs9wHQrRoUWvILzp8c9h9/9xknY1a3WXVaEIFdw/yv59hes2SK+XfM
ZOkkJPxGdyA8cwqGYkq9V2X4DFLL9Y3wbLgZ7tC9AuiAz5aTM0NBURH9k6PZx8ZVYSVQWsmkaYXX
eZ0n3Py7yKfJWiiJSqouPs1uRA2mwEAlsCyOqfnNbSR6yxAPYHYKNr/iX7tm5t/fhyAj/VZBkhgR
6833qA39PRM5he3PEuxdlGicZmCG1GgoVdXoTtvQ9l3iWnGcsn1Is+p4irdvaDr6WrfZZUcSTahU
zIna0JD7v/f1RnLjpb75iamBhi+LJ69ApP7rPIpw0pAq7mx9xfb1yT3/ddT0fbTTBCjFCh9sK6ie
+qU62nV9V8JTMCQ1tYEgcI1b3i7hi5+8riKKJDazLpVbtm9o+d7eiXMMbZeuk83xreyo1g42B8U0
THksz+tndKiOVxZjtsFckWb8o1kvfB3GCgVR0JokUJ785VB2JYuioY98B4ix5IuutRkHFsahrEpY
k3sMB+d/tYQdSQD9SJ0c3Wvsj5nO2dGBzJ50p2ytcWR0D4EWoCyTGN42sP20hnwEB+fKxfxXu1ov
7crdLNNPC3wR1KJOPJXC0H7PHzrHelsMz0v6cMr9jUUXsXK7W9wMQyuyFPZBMbF4Conts9eUJGt7
eN5NHn+/grDDnbJ6wmVSC8lN8hDlRJ/ZWRQibI7ZDXhbSC4XcYES+iaaPPxBwVn5b1dKcpP045Rk
4GUNCBHquQ0swUXpHHnOnLHvVM0J4Tu7/C+bDiS9zDU/jMZMvROM5vz3UKCCIHxAD8eDZ0BeG896
Ly5ev9WMUajfVthCzYH4W0B5dhCYfx4KltTfiYaOYOvWbjRURKh6aIM5aifXQ5oiEF476iG7/cc2
j2W+dBg577PWdMobwCTVw6ILwNfUBDkoV03yYgodZpTEsqPt+8nimxoetS1ZiyItURSZChNybLWt
Xc0QayDD8+6HECqrt9u9Jy5+6H78Bf7ev32Y+JuQpY3jChY/vDH8AWdNqOK2D8+dKr9N+XmpX5Q1
FA5tv/9ZADwmsh5LmU3+4FQIAm6ZCG+IuB09anbKZFx01S4slzY69Mf2w7hSI5mizXhsxb5c6zKi
wEQkH66/zhRWLAHx0plfUmWbKrFviXDtp+sd74ETXHxQQk5UwZD+YKZBwcA/f0nSgkhfjbTmhKfo
GUKhXcbchr5Nv87d7okDD/NhTyoutsbaGCBBPC/ZgM/HrgHaqnFx7z7M3I9c6+uAqexOPhfRmWwB
ariBPu8bKdnKPgdlzz1cXmIJaHg5bHCeSzxcS1oabKauA1E4288UsIKfvMMDi3jI6y7qd2iZiTv3
OI2B/kkcyplp6yBc7FBv9qAQ0H0eOaAQCZ06O0qm0FJPhkhm7PDlXu3IgTqeHLRc6qM4+1+2bpAF
WP9XGtsNXeENN3w0/OKZAs7BPypQ4V9ry/u5Q3indr69bfpQOjkzxCoWDmoW/PrFhKSbdLSlhHEX
HVYRYM2MESynhyYAAljsRZC+fLIWnpeolMRXTRxDDzPUjhYyJV8L3IeEJXh/VhjXYSZcZLhZUwjG
22edDzTt87D6jRkDF4L44S/xpRuQCPVIY+kSf0xUp0e87RDWmUe6MsBODPXrxRAipDcsBW1MuOw8
c/y7QoYyUYoxMkqIo9TzBZ8cMTvFHRO6V1lpZhZVMMWo80rp7JnfrjF6EbvNkWa4m9Fs+gkbSwI9
Szat3NSn5n0aEXUNjFRYuKvvn8T99Dn0GQwYWHPvIO51u3uJYN5/aU0dfgXNxjjTcg/FYsLFB+CK
0K4JMqL/VzKa4M7fsei5MH82y94JRUld629YsFepfENxHcl0c7SVuGO6yd4InX51ozMOLIQvDV9R
TVmOjWZuzautLyIG0ICp+hiZS/6QQZYtZaU0T4xCE6jZhxnBrLG3VsF45YhmpN02vWOGZSSqhDoH
6juWjDrxCAH0vkn6H+DaCxpiGePGgD9kxdWMf99D5Mmj/EPWkEmNaAsRc29OrQ//33f7QQA2Su5Z
RT0uUN8bFVfiw8+YUI2m2Q0YynIAlIfFcj7Vf5395LG9fyMvyzXJ+13/FXut7IfNZ/CkcFnXLdn7
tSoYv9xBDkADhxWuoP9X9xZcXKLgKdYw1k/qjPjAC8zXl4Buj7JsE7z1a/a9Du/SsDQc1qx4D9FM
cw2ZSLvzSefnhhZuzWNkzWsotozbdtXg6jQ97ZeB5fVj3xCBYcNPFLWEFi+QxyY42lXWm9gmBU/A
d+bSZ4rU29vWa/TZbsmCKYWPpxOXeB3FgCkNxUAIa7qaHtUqyeRF5WljBGRbLAjkvxOHhILkHayw
mO08wOQli8shgHKNuhFKAtPpMtO+wMCsqHzbplfBjRg40yY7/M0iR0Ke5aXtRdfW3XKAnSIa+047
/TcqT4lflvrCgBRo9RzlminIpbvOxz/3x6Hz4eUxeSINIw2ibimPUU1XvFP0oGz7JTlmN+uGf/NN
mhNQ5se1tM5XdClv4Tk+WkUHdBFxm4J3/Jo669yzFCxY8/e+NiZkwPzywd9SubteGZ2CL5Zie0XE
qDEO/TkeYYwH2pQ08CMJkac5q0DmaT2ee9g3ZUpjSertoLpBuxZu+Q2tt5wolnvUKXoj4J1CEzl1
z4h5VtQwFDEZVxXU7wpJFhwKo6zib3/04jznvjy+C4571+P/IFXwHpbBMXC0v3YZHXQgi5lg/1/q
VoOao+fHXcpfzn4o8n/0Bi32A5VbGkW7nUDgH4NeQCqTPCsmlKED6gpZbzhU3lBAoE5YBVAX/S/M
HL0Tl1zqW2Tz2tc2f9v7U1z4YSZ9FW3xklQ97c+8BEFsbDN0ZmE2CTkLx8fk+XMI96p6+tGGih5d
gDh/EvCavnNrdE3cpT5knLRumwEeh8IyW6rYLDg6jBHTCgaRQOJMZWk2la1EWyBHvdjlKqO43g5z
1Fy98EZgYjP9oaiBdjz8VDJOX1f5NBbR5p9V6rLFZm+rxkSQ6ac2nx3faxD64QfI0eetqD1FOSjl
1/S/MihSIE9cDolYO48pS9M0ayfQcsSJS4NlATettdpuF2D26oHItRUb0qlgGUtaqGZvgbCkrhR0
j3GMKyT6wsxmXmmGKKO8ZlX4tRB2iTYGGKsLrjdnWkVeQTpYeGpkSVJDoCD5xF1JTpznulwX8QK0
eQjJ/1/d4C7pfhez8hdoaZXpMuZPyKdYBn6HD+TOif6usYFsrRkNwfg/2Xk9gE9GUX+kD8rdVGdC
YuPaS8zlXt0ee9JXhYDC4Xg1gHo4ucaHGRUJbSxu0I8oZTZJIfLw2xXvLthTG2S5WYCFMPbH9lgs
JuF4d3ifxPD2sBwC0jgFcRNC4wWu+WFYCcug1LNpAkxK6RV2f+5TtgFroVp1nx2SCDVLb0wAXVJF
9X29uyEX6aHLTjb3KMx+5Wi1Ey3nwu7p0BEZwXdvJzFwz9u1eLvoe9wa3m/Omshxj+gtCzyde161
IXcNfpFHnmLmHZaBp20ar2XBZhgShi3oUXbRhO5rwzAb77zV8ZcnF6wxjd0Gw60fPsi4BU7HdRnB
KFLvG8CLUqRtSlclMHKoPRfGsYhR2eGGuxM0hmgHStJMA2iSIKKHavv1RUrHnh/+SYn8X5FcshfH
kvov8f4mFHd3HLzkIYEgnabQi/qr4YmaLFesm9/phfQ2DRKf6pv60dtFJ5c6rgRwFr6Nvc6jMCgY
03RLJsUxc3z4RgM+6QfEPDmbTsD2NhLoLp8tpdd5gS9NvcWMIG+jj4nUJPomXJW9+PS+903tyoV2
0ZETTwD6FZb08s48Qom2GsfqfDwyFjOevsUJliPVAjhp0x11dQQ39O5xARit2p718wPmkMwJYbmJ
83V1WhPeQEADrEFp+x6QWFi7MrwpPlLSqHiHH5xr17NIQzZUfSDX3x8zqcjyzS20RqhZ5iC1mdG6
q2ERYaKQZ6mQi4eh8oWFzjEezAZHNUO+4YROm4pNvzZXfmvlkPai3yvKYlU7U+ShX+wH3hX1Luqt
4n4ikhDVDHMNJHydKHif5e85C/hZtXSJJo7IinwkZ6LqSxoT0uHmSgGUPVBqFT8ntnZ6vt6R726c
gsY9Bcsc5Jlb3izNBT2yFQQqJ+5+a+IhVaym3SQNacA2zoyHueum1VqpqIslyz4wdWclgieA5nRU
z0n0Rlso9h3JGZU9j5snLDeJHAp69IKAZy8XkQDnYksfkWPHF5MDifeXdltF9HYgjRUAsBB7SNI6
uuvWWoUJyAbNt5J8vTCs+GmphTMH4fMmjZUk6176M7X3JgAKh+UKj1tnMjU7u3kKJddBDFsi5lY8
cAFcPScoRrjU9EfM4q3zMNSdj3AdLOUGKmY54IBaVGrHAlkcIuiLuK4k9Fx6XhftK01qVDdRfUM7
jGGkPc0LHUZMBGGkSmYdAhleImnKp/xrbEvrR9kcgGbHW8/Asshf/uYBs2IOpsiJfcM2KKI+aviV
a2Zy9a9KOiKT94T2NUrs9VaWWgefUKtGHeto617F7aLQMd7uAxkmwyDSJodxPrvQRSXtVgz1T1+p
VRxrJzX9vKCm+VVZujY2kh7e64c1Pxwsc5IGVQ/bg07O0adPsU0MLkBhX4jwOJxn/HQ83SHhv1mz
vhIt9rYWpgGG3nVt7vUUXoadbn/MD0Fekoxz0c/WhohKIGZfqOFkgGvVfuOk4XtWVTg2ITf28z06
oU2AbT6OWF5FyLrOFmK6er0nlyYgKp+CtsZEiuv64+5SjXitwu0jz6DBXYjEvkm5XMwvNrYwpz1C
Y22NYxmlhxz1fBsHkqLs3kqGo5Z0KFDduvlW8HaJ82fglmCo87sWAASQgNmOhaiuiLmV0RzLGqKE
vGMF4Ky5Hc8v8BrORdl7szzazEbdFbWIjq+sRo2dOCo3tbC9e1p22Lv96e6vJXS7FRnCs/0RCIwK
GP/uQB5ZU0MHSXxJgx7GMdyg+NvZugdfxHEH8QbgcZITm2/9Pq7E0OirATyTUs8tijZwbda0nze6
209P8Ue93fudpy670+35wykri5TvDcvYQ/hez1sbBnj0SaLoG1IB7o6UzTbI372IVpu+lO7DCt3r
GNZ6zrD/7CVEiamAtMJSwFv4Ixe8aLzQrqOYidLQw9jdAD17U4fNUl6tFoqZPQLZ+NZYoyzxWHmY
9v5FUX+SLm4plyl+M3As7N/iHxPyugdicHYlQkpg9XMDEN6pyEXXdMs90u2/5f6x9yr7OIeFLmyK
dHSzvo/+fuxZ3dqcQS80oCnRdqjiNX4SHk2Cot3euH2nX2OdOdpGwdzaQhcz7L3sqGy1jCeqWV8D
q6D6XiIW7Cj3w0u7s0zxgjyKfL1hZNnsjpHpzRyBM+r1IExtDMSmngqKeiHvbjXV16LJi4CPMQQt
ZooDQv8RViJ9gMQSS01qxMJw/KbA6jajvVdPQ0JBmwIw/VyDFAFN72HK82CZvcCk9ZJIMYmwQWiL
P8jhQBIg50igu1AIDCOdCq/BPP4iEcyy09v44b9LqLHDBPT3BoDvRlvC8SfkV4g6mDPe0td6F1Eo
KCB1jgK1QnKHlm0FFJ8noH1EHJpSYcexST/3EkuQ1t7KITGuMRDBytyqygFsQmmMsUHVLDDqkz45
agUbTBTzTLZuUYlchdFO1Hw+BI66zHSHOAFWBgeJfIIKtOD4iawKgpBrNPfuI4ODRqLXTdoXDYAC
WKlQf/sS44uEP+K0Xd6rlaK8X54jTAqhQ7ndxLE52NlIG6GildYEIqdmB+qZK8TZ5C/nrGL/W8KG
Q3XdlfdKAgTJb/0YVPPQXQJ9BPsx/oiv18jQ13Tr0DFKNEnakZk5MJQEewLUfBvBO1BoCDb24+c2
cECF8HZkI7D/M5sk1gjDKtpSQ6mZgit+POEjQhGDA55H3tiSx8bYd58tqBCnbC8rnhFCP5JaSFpj
Xb3eaknGOvcprpbsHOCkrzhSj2aCV7mBFGXV6eF3DnhLd/V1SeACwknK6k+5NUt6iFgTBRvk2Nqw
V4Vixidao6BGw7NFOuikO6v/dYMqsb1VDKNm/lx/UdLV1eu+pU+VZQtTMTSWg/Wnd8BUjaoX9kGm
vGMcSrDo4SYamlu408fH2H9nwXpnhQUEWGLtOEApdNegNIYVBXR/2ksvgTeWFxPGb57fcYf3+LiS
oHhEx0q2ble2MvWNxdCZgIxdBYwrgsRVm4vdfdViyOH5szkLAcUQfLLdbPfX0/HC6iCu4Ngw3n3O
Srwg16nLjHbW8mKM72jvcG8t6xVZQGCxBEz8n1cYeK/SKuZ2689YetW+rmW8EK2HQlUV7mh1FsMQ
+I+I1NZvI4Fd1MtaWke4P37dGnXKzlZlly//gLDALs6toiUdT5zrO0Nlz52JMKmqOFaRsvvTulRQ
KTqSFkmbp6EiZ0zIaHfSOo+VxQ3FaX1PARNHze4nR3CkhW3OTNGYWfY5SvIya8pTk/R4udWrTFBT
+EmT3VkRijoeKI+rgq+mKKeqB/nRb/fuVHeY9hdHqgPlGUW8wQtagiIksu+z7oOjCf5dtF3FK3IH
BisRYBDDApwTLodQnTfNSFOOqG8A6s1IXrKO1xtxUp26TlcJp6z+6sDm2c3RpMhL1DVr92e+mLKH
vkuKD0dNYLWTUaAeFKb0yasWhuPGX0dWB3YKqHpk1NXgzBtAOuaLHXrQqsX11kd+mVueZ4zGXJEw
Joc1kwpagUDBfcwwPs8fx9MDe33Jt/QShCOGKOUUGHcwr9tRxjbS9ZK1ZFXIcVnAiRjdtVsx0EHv
oXzsxn0+dhdHxMeoCNJiBzia6FZZq7CpF3VWI7aBlpCvGD8rG4P3KexfDmw/lEPfIWvwXj/7ZyDM
8vW/v0vffiz+qdDwvjOpTJl7VNTKlzpmtTyAiJR6C/VhKTeyg3BWrI9Z+netFB/kdWNyHO06ujCH
nT3J/6AN5RLYeGewxl4+P0FkihBF++tCtDGyWlJP7fGt733x12IXjSBcd72NTXEi/rNtNZ24ZVYe
L2iXA0n7RvaAh1QzEciz3zEAcOy33IWA/np6YfT4Y3N64MI76Yn4/c6tVS11FVAu3cFPOoWa93K0
fzZhuBx3bx8+bp5HIl+PQkKOEbQPSJME/VSDsykaJoGr3WFye5deQYMi2/m1EhtkHZmUhexEC8hI
JQlzyW21ZuSYKUDPR4C1ZyRKQlYfHy13xfOKLyKd38qSRyITR8U0psHM6jqSXHF7FqOOe/imNxxW
KgxW/GwtptHvcKjC46Ned4roqNg3eP4pDPYESOZl9dBnMtb+o7EDU+AIdSHTdcFsrT6YzZLc8lKz
4L8yxxrsCcK5fNzhDrBXcomb9R5FjPTsOB4stkzAhi4UMR19v63h4yZoUBB5/RiFQV18PJ03kXsR
cq5AP72LT8oJF5XkDCEcEKGSSHhbzCvIEqmRu28DliS4xGq4LQ00N+0PNifLXUx1pp/6RW0JFV7m
O2lmZzqE2nrxZkMRnYqaew4DrqRL6vrkpS7Hr+s0riFjrHg07t77l5kzshwOLNSeWpwiObhdm62U
qZvFBbfRv/1f6QDoXjSScCOTtyo03VoVCEl6knrn0gkG9ODQi1Y1nF+nUcmh4DNCUx5e7YvQjaLW
NUfsBxS0FeUq26N25/PPy0LsYvSD4wn+u3oMWTmLKSJvsmMACFZglW0vM7lQYUgletmodtzN0lp3
aN333wAx5u2J7xFCIeHZUoWEWRjpRzE5b0CzwT6EmGbHqsu6Vp+fYyRZIBND6YSGhen2uBwS2UcF
pTsjRjGoQyt7f2s7FUwXcOJA5Xc35eK9/cLcxD1q14fSr2hahjNF7zQVg0iHNuW3JPOXT2gL3FUT
LXTBZjqTpyu2qIksRrvNASVmuF0iPn2EBd5QFlKeqcRkCdhbodEBo9LrQHlA8OSseQEyzAat2O5L
2M7M3gmRKzMepvk8W343luNgEiI5VgXPBi4nPWEg6GjqVTL/vCMhR6M+WQ6eEp3JLK9AeRBIlYXd
QL/OnFon4CKCCi7Jz8YZpfyGJadGtTTK7WT0bBvfO70Hm04dio8YQTwXsLnN0TIz58Kc0TSMpXT4
yRR02lLxTwhY65HN+iL97f+GxWeWAR+zm6MRA8jBRx0Oh+x2ZVD04MQHCmgoEHeT8p6f1cw4dRNH
pS0D8j0ifDUubxae99wjFNi1+VjD2laWbP14JhO26TkBZ9Nb6kdXx9YF548/faaYLyBUfBbdDbir
nHEEo4fP3iES93u6+cNootf8ekME4ihKGqvKJ91oIKpdLVeYnVvbl8YWUJ+gfW4yj17DlmR+ARc6
uU9d/OVvS0+OPKJk0UwfwyN+84OYbh1tT4pbgQO2HHq89PfZT7pDAsvBpkLqL6FF2P1yKTGpvaC0
jOjadPg5lbjSTsgQDMtzOHFMHB5OPUFX0BdlXd3D5xZ/E6iOOrLWEg2PMg2MnUH8SdV5ewqacA3S
slx/euVUT3hnFsXzT2v/8DY/o7EnVn/L3vWr03LmSp7siQfgVvwOL8PRApiHIKwnryQ8bPky29nS
zNWTxdI0PhRSZBHmXE0LgtmC5+4nzOdc879kIMrhWMlbV/xgzTQHKy3mJdOKo35/K0uW784D3rME
bd9vm878BladsPGY7SbIpNoz9zMrYYDFmsh7ODvTPrlq5McGS5gnXZ4INxNxY8+z54npVPbyI2sW
obSKCgiovyWn0gxu3PpLcPXWohOul8ywuemBfvNkoVl/NW1HVhaIo9w9RZGXjpqUkvEBXoH/WK55
sZuKdQUzHNeCLVA9GC0XZtbdgHVi2Fjt0lfWIgucVocTM41QODsi0+m+ULe2BHaL7Am3KT82ESe3
BL9Deb+1MBEFlaBsyLmFObViQG/VhuUeo5hMhq1hS7mNkesEXX5xJoWFTX/rZG8yJswSY+re18N1
pGS47n1/y5KJM0/lVljPy0VLi+VbU+0iKeqS1ictFzTgZceFhWNwSe3ElOnic1/5RSfC8yrNGl56
WLqRGGIDr/ltmT+1Lfh/1O3edLlCWyJnoo5m9hBMtB9/2DjXSYmcOI6X9PDqAtI/JJApNQFDfi9a
hG3tlNi5jKfo94Z5PLVCNiyQNoBROfLbuyY9tSppA8h0UCLQ8SMd4hyIkxGpmgXVCAIdGTE6EpkG
c/NJxF8BGdspsapb6HG61VZ93TDfTnP4vrIEj3ODRGkN9f5LUP87l0VsqGBoaR3ix6yzMDrfR0cM
wgbQ5pARKzzDnUrqyyPIFYTw7aH/xTTnWpgOCL+yeQz9r6zM9AzyQnubGU42hhlSJGi5avG9T9Mz
ZJOpzqXi0G/jZtCxkmhuDba7/KPFD+Y1fijKR35YoaF0AQVrFB7htYV6vE1nd17CQdDRglKApwrf
eBNjVFKGOLQsBbGEqbONh2eTA7/9mwDTT5x6wV5vjCXauzK0ny1bPTzaZ3GyQMUaDCLHDqDC0Nj6
JFP7ttQmoYT3poW/jpFJN4hsVZBOxl+eDpORqkAckl4EO0MJTue8I9nXsv2I6WE3KiSrGdoe47tU
94Wvm225eqxOpIhGw3GLeMiHRa6pivsCynPyq1yOYy8k9cFe7m4mQi5dqIJzGrTAZcf5E/Y1Hbyt
bqhuN1AzvA5s0fxE/765yF7m6JfFP47vm7GuhXQog2An8s255d6Jb0YjKBxaOeyVL0AKv0y9GZwG
6vISpzCO8ipLrRN78h1YZzpUdB7zVCrrqwQMCPVQtrymlCQJDfyZ7gFqac2g3SDo1LErAzxGK+7u
ID1gCshwKsIQzcFg/o6j38ULvQa+eFLXE/jD6yR1dz3UCODhyWTXuLcWIXQp2y6OaIN3KKQ/V8kx
xSZND8gNmDUFFm7+pjbD8hSf4vTQScvtEv5yC5qaIH2aO7Y/IQ9BT542mtSt/OzoYQTg7IyA6Gez
bSvTaATelfRbNM5UF/pPU8W6fkqaT41DvskD/Ivr+oHzhcitRrjW3ju3OeDTiuAWxmwTTToCsKL3
LQB3CnTqqXSpqsLuOxstBms3TtVzUpHlU2n4vpCnCb2Gik4RMCv06gKPzcFEOcceCOS7Fmqr++xJ
oRuOhNvpuLNq75/evHe0VZ+8eipG9lH6ds20KuIG9RXcwKExrAasRFJIUMP/qiLE8MWgGG3PRvKN
2+6Y3IWc+e729D/1sXlfTiiHrrfdGHd8ttjlUL3wFBDSC+xCIpJa4jrB8PM3zSOAUGtFGfYLihd0
QiIcVU1dZmYvY+XjBpwyRp17oepRb9w/TYvsEYnQ1pAJGO9GM+tvn3wcY2n6lXIisr+DpVrDS6O9
lajoxBsUJre5mBf+bduI6ZGiWxjexKv9kj4ojt+y/BUgEnq73tAgHyfjiU3A7UezDg3UJtIzV5bm
a5qefJdeqCRuSpQRkDMxuRfxMga236GxW10s3OEX87xey0LZoYEmWieiMJJb4gF6svhAS2TaUl9+
XNvsdIMptYFb625opUuItYSYcibpASQxt1uf+M/P/zgPeB1cHQPoykdqztu2OoPtaONc0syLmwQq
9dhBw6Gr/X183Ppbo2IqKA9J1akpxVh3gWg7x6PDQWOM/EsAs3ZmsLQtSt1whjPBMGCQ6OGtBFob
hTb1E+Soe9j9sqwmg9w/IojQEnygbJB3fOJwzZxCX1ntFXS/178Wq7wmd8xxfW0pm0gZ9YcRfd2S
1dGwhuuqRPBTMWhGLeUFB+y6LdWJgVjmQ6qfstN39ZlfGHqUaWYgRhdDfZhgXR+TuLBlgc8BBe+N
X8MOUpgIEgbOhcLytw9gCEtwO/w1IjweXN2rm1KGba+x9x7VpG2jDJWCXgMaP2q7yF0mT8dBUKok
paka9l4BQs+Jl/xBkaZ740i+2BMtF2cnZ0Tj58NKZ/lKzep4h7i/av1RIemC63YySfk5TBGIA+7J
e8/Ql+ATLiYsz+DH/vK7JDKyDCwdBC1bcSHQLjJHe26qUA9gwx4WOtGWRrWmSEphmuQ86FiPufDf
agEqd2QxlGUWRLb6OAo28CxyLPgm/ZZ0+eOIBSIIUk+mRe5nK7jMCDjgUSkC6dCWEAVPLv5rfxeE
31Tz/g3Krx20OHVcoeGJor+4WVEUArLuf2s4vJTV6MBP/xQOntxKmTEDfZtLGLuCdcdQiK8yXq6L
mUGibnuuMQkF+FPW18ZCLRFyecblBTMJ4hRbXoNVsiOAY7fOIwkEcZNzaxpiu2hrwpnS5l/5yvCB
cs1/DlGMbnKAg23irx646rhzDPi+3srh3zqjbJtjK4HLM7yTTr8D9G1lhs1ZMPhwWuv5+JzyCe4N
tMTgO+yIhLt+3zeYIKc4Zy/yJQPoOWgD99+O8U6vx0CxZ2Zun3LLIoztzNzJmTgDQz/6442IEG7L
xeDVo4s1fMwWvVfvmGUlkjgRyii1W7x2B7WrgCztWKB56rWcFkcDp3CZVj0IE+A4uggihApwA66t
Cw9HplyfeawS6IhFtVWtttNHpvaaR3iV1dff3lB5QWvvIGOIx+Py1eubrwTPa2Y9GkEA/IW7tR32
1MK5lfW6KoBs9Zz0b7UjbjgvEQ2SDhooj/HmJCJAaReOOIdORm9O+F9j1osfbIO5u+WcyA8gtVd5
EHSwn3YhRqAEsOx4ZDkkysaveExJnGkWSSjb6ZBDKTF0bSxHmLUI5m5pVimdzLbKrxgkAdPV1EdN
c6h7YAb7orkXCGTCH51jT+AzUetaV2ShGeYyJ1OKFxc6Y8cTRwwE/t1qGZwAzg+SlfFjXvPkNdpB
AR1G7TTNvQarNogwh892u9Xq7sTRIVJSofWN/1AzVYA2igFkFZY6v9hjMckgk5FC/aoflNcL+QRw
k+gLTEUb2Stv2jJxV+LtA6ra7K3boe2MUkIvE2GJAgUOyLDO+SSA+Ur1Nv8hCHH9B5489wwResEV
Z3P6H4+Xw1CJD1BL7HRiaGH+DobxR5wAnuY3T4hJ9fhZ98U4uiqqY1LaEWWEABB5nPNocUlt0MjD
ca5fFy254SRWuqErUX3aLT/qPlCe1BFYysBq2EWCqrv7eyBY29w1+9Fx6Ov+mnHoYYzSviLYkj9L
SGhHiaKPKDImrGxZLP5J0Zbq1JGRx3OjTOamoFcR90ZiXFH6r2NkWNqnw/5HSUy6foEkqiriSp1M
sXeaEL+jXUZUH+fLMW/iULixeoEZQi6x5R0ZuRs/F5Xw8wJgppFJi3MXpUVUaWch2h/yyzoggral
9wS8/1XT+sJj9yPgcOeTPW6+F2vdu7iE6bz8hj8Qjf+RxY8ZDk3CXmlAmfbY16CQjEuqkKUuBllp
gzZSO2NaDbO1dNPhA/jPU2B1+6HOK/Zupzubt4evqffldEd71fNUdXTYOEAetJV3CXzHiVZNSXUb
pWnOpCgdgEUfog68DnMphqWtXWpvCmX4FdcUM7wE0AvkHjyi4+uQ17bWBCUG/pAEUKLhNFYoLyja
5P2b/lfZJt5gonIMKyNYu0/jURcKyvE6aYhRlmzfowJjFgtgzKTQJtIs4hSW/MizwRPdWonOOGA/
fiJcurHQYdpfNuDswTTRbG4K0AxaPWocanGBFjwXRYEOk2mk0t2/MYGkWYFsV7xgx0gJyXaSIpyf
uknoOA4a2BspqLEdpbpXMjJQdw/XfEmStaxa2axKC41SutWgc06uUA5TqG6D+wB+JocpnAGTkRqt
TtiP6rOFJsfrzgpT3PXyJbC9W25fJRwG1tbOUSIkT43QbCuFSG4xHh5irL9Tz6jAK3q4hJuw0E7G
poOuLHocU+jGmjx6nuZal7N3l9AIhSafJMI7frJIIGCxuNYfaNL8t7vI/R56/rRaLxbD6hnlhR6x
ejlaPvcng+r3r/z1c+penoPtapGQFqWOZc6p0f0cwGsxCbP1gKZoTPut5JsfmpKDwy2Jtk6Fw6SG
MXxH1WnAyiunXIgGcVo7qO/WV9oE8C5ejNdj6XfQpi0sBPVc10YsCwlxTTuwdftwmqAQmQ/wQ58Z
rhu42vfQdhLzIoEdnmQZJ1aEA0JUQJtijXq97gNloDFJWlS8CrbWZB/hLlEs989aLDU4/oSGsd6k
suehPgFz8z027D7e1ZFZFcyyaS8w/QWD5n6QOZJUN+mC0m6vGH8jpElMtPR3yLNiL4g+S5EgBVj8
dfZIEx8EF9OJhPw9fuRKG0aIbPmaHH4C7U+bX/bXGGSW5qw/IPf+rPRnsE2LfiCc6h9epS/5opfB
UQfLr5ahre16I0hWUPL21GlzuC8Mlw/S5qYt4nJm0f0Rup8ulHaimUqiR5OEa2V38WjyboMe1VB4
/VJP6yKvFleWB+7BTe4UdHH+p5GB4fYeSRQDyCA8uJo7E/h4lXtMDUH+FvhHQzLOxXVi8/6HO9vt
QmA8chgfBRbGhD5FfX4EB8QoawIajum6vMjTvDCZajPFrxtPu/HZhb2tHnK/UXzqoaF87qXcLVB+
X2J1t32QxtyYx1HeDEMnvdp+0UvGGMIl9IOVkJUU3Th3CIZihGu9uo7o81IEw/CpUWWjQ2iTMvTJ
QlB8kOk/UssP0BSsWdQneFEvIw5Bqe63juYNUBdwwkRt4kqEaapqOTHZMPyKTcVhOH6Oa6zBem6C
fXke0CCUbzFAQ4IzWu1uz2frwffEk+L3jXDK+Dj/5zJm7k4iRyAxxV50QdyFM9dbVnmAvqi9avf/
D5ygsuYUMqzUbEE+PU5u6DpqdapPFg4frrYVso1dTy7dpQDth4fhHVZQjfE3M6DQ+sz3wEr0Kg24
MDUsNk2jt1A+VcLgoulK4ecjvYyRZ1YZ3HDO6cUselZNWyX/CLUHlqr8u/ZohptonUdn7n62HCc7
mwpTjri6lk86sxYEylJDpIt29FqeTXhDnuIvZjEg9L5fQ70Et34T2sDWqUOr6JJq9+dUQTbPP3rt
ZjVJcsOlUzeLw6kT0ofmESQ874/ezoswUiVsh18qeZZVqWQOs/VzVppGGC4gHur8AV4K8xa17cuG
iAxE6eRSz8CnvjnW6+ArSy5LlJSNa8o+u/RSqsJ6EuiMpBH61wnk3GLxO7PIwDHuGpe7i1uJ0be6
pTqPxBvn4tANi2FEnbOp+24lW/EanEJLfuOatfKb0AyR4KMqaJ7caf2Qkeg0VIvutKrTUXQZ9lR6
DGt9dRWnTth95llIx8V5CP0VcbATjNJ/5zilN9yc14jUhVQCeOEGeVYmOtAebWhKzXZXnUE4rCbc
M3Li6GXN4m8VplrZlKSHAJHGssvDywFoQ+k4zXRgxzI9lo2s1ihmbU0zILzGz+nPBOd/UzJJuGrH
W1Hx1N7x8YHjIZSgMXPKmG9fAvnSVEuAc6C0rGkFnHgPjtVC+qhJ/3HIJ8uBDGRUKSOLAAJi+DKy
LheMU2BTacuCXb6jwZtaBzfXXlFjlBw6WKbvvq24EtPi2vETBh6NZF48L4st16u52DdMUkVA59HP
VzAOdxbkJDlnU73cZEirIFxyFNU2GQ5G1lrA/YIn+EXWqCZ/GYlo2/2NuZ1vSWygUJ+AUigPy0DL
+CEFSm672iD2V+QD/6wzrtFT44mso5UloGYs7EFtelMpcqrk38XlpxFCS53vvXorO71oSiLUpVLF
d1F9oZEAd8I2W6iu8u9vLC8H8rgmASEMHFQma+YXD7E91P3fpJFY1uF6dMtL2Pp/hE9OIPVEK4oq
RAo+Pe9lX1518Ng5gqR4zt8nO9uXZfcg2gX4is51C4zhudXsEc4z6XAGEfxFfxupRaZNLmJC30I6
6QfjeZu/n63ACyqd5tSawa76JigsGSlxU9muUW/8t0tz4bnFUXPYKz7C2W27OzAqe1yFPtMlyyD1
77pG/nVLLQ67IEaSt2b6rZRXPQ26XZHN6OtCW8+Y5KNokSfjmCp60402VUDXbLB0i8ehdkKlZ+NG
LkV7QElCMiMFcHAtPm08QS2K+pRab2yrIlKiQGpQnjb+Pha68y6zIPc9TTjGHrXuK5JgQ0NUJuga
l7d5iIeWapaTJ86gbgLP1OJcqbO6tlVyLF/0Hk8XZvJqq3mYVZWQMdu4HerCitGILAbyBh6Dztns
ORlyicM5dZyl3c4Q7ONt3yZjUxPq8TlFoi8Mp5Y8W2TbB/jRukMFMBPMF22rbhLtrJRuTOssoWHA
W3Kdzwu/9jSS4X+BBRthuWeuCkFS+GTk7SMcLAkK20hNNhwCTvjmIlV72yE1YFVv9EOif7se37b2
ShvLINFLKCXgwO1KaDflJd4IT9ymSGxB5s8y9a0DrKnXdd7IgpaetIUMl0DEXKSYgjs2EzK0UPsO
PI5RedHs3RgzSXZNxQ0r84OgqYuzHQODLo/stvbpRh1oku0UzNUyRuyPAqGBwGY3AGuAkytbjiGw
ua9nXQGqL0yQMW0vaf3dhBUyDewuAv11NYbZBjM12wJKgR2P+Cm3mGXrB7uy3xCjRGXMBJDE+5DV
JUE4jC1HjdpHRQfZEwrDcLKQdTsm5DQauVkapDfQoj1gNvfK+TRbGY6e5CzZG8v+/P0OoNxc7qSD
JKaDm1n7Mhvb8JQuI3B303iiJTMPwNzvfZu0X0duG5RhMXr8hL0WbctQFapirJ/kVE8ND4Yta4dY
pDgo06oKNmM8w1+dVjlx00Ww3h1J3PQy4NZMQ3Y9VYjV3hzhpSnmWLcfoyQo5Tt5FgKBT0u8Vpw+
ZTo0wVv+eDFvPZVTepaucjjfQj1QgayOV+ALlInDP7aQpx6ul8SO6rOXQ65mypGpJCA3YzIhcM5l
guRndpILnZMVZITwa/idrseTMAF5EkfAoOrHOkkJ0gaLFKDs5AAEFgWd21oNaZ23t2/3FYpiSO1t
4mJsyEJ6YfjlRwxwpIz2KPXf7MhfjKiIu5tCZT41boR22Ae82S9P4N/wCPby+O9osc6sQys7+DUr
VfXWTwpj9+I3KErU+uLR+r5AT10rc/X8awW9F4ieuVQRwHMcMIjFzURUnnF8mS3HpitPToO2PC+D
9U/RCSWYSZVpaYnPo+25floAdnZ46CuW/J5OGHvC7pW604HCgmNrER3C6+ECuVHsOFM5dIRJsgQq
l+9d4CnnwQv9jErdzYKzvI4KbaVFROrIhjyLEUDM4TOKmSRt5OsjM4rJg+Fb2B51XEdgKS7aD+PH
PTSmtJFeQ9yo0siOB2a2l0Zf0evIofNjxWsTzEzSNSZ3tiJDaUo/LhhLlSlqqa1hj2IOvZLJyPmQ
o04O1oPsbA8o2Mf1eDBLWZniRr9AtGmG6oFZGamvIFoqXdJsomjKXMNV4KM7UQGm+S5vXIxwtuZU
4svuUycNyAps3lGzaeVF4G0nifB/KltgFx+8ubJMHMwIW9ox0hRYxyJTZ0puMcXgLXvQWyXzE4l4
J/xe94wLoMXm26bSkfNhSgw0YqfwojBTukh0YMSPjWrI1RtuIQtaraMqThCzuvEsKO50Z4TuxmQG
b+KsML2wasxYD4Avf5g2XL4xApy/Mx5RvHUQGY1BNOG2K+ZWLw8wp+9KqKQEBTDTZObXNp24BK60
UEuHzYkm+0aQcLj8UEg9xq6fkeDKkM4sJa3xUqS0J1Fclq0Crgw4oXusGDMwlOlw6HD9jGy2yTUA
6tmbaUY0ruCsL8hyj0Oj58R+nr3p7T5h0xEzi0Zq8c152pM0X1nk3C9vcgm9zlCnkoUeqNj8GKWB
sWB7NfSPgGOXSUFIKYbpMeh3nBf+b8/JIn8tgwkRyKhbDTcstGtIYc3NVbAQE5emcp7jBZLWLt0W
2sypW5asC1bPCH0bqjmItxy72K/K6fR8QchPTD7wgyBBVHmyovBSFcI8s2gRq8lWZLwPEISKM7KU
I2/qRbaesGUsSSnHNDBpnU5Cb8ulaUi8VMklZusaTwl4NHAYi4beml1Dkx5FC/KLGQCOjtUqRK3H
5T7UIEFuynk2gHnwkW3I7W4HJcPkhmjoIgKyN5d5Xen/o7VunFYJPlJbIPjlw/91A5CkPVH7AA2D
XqIBbmcKEgMycF8lFZIeuhx5fqVzVWI2nk0aKQWkmc5NHwnpK81uSxXSbvt3QtyOUx9pVjxAfQ7o
I5loEpZ0j2hGBlg7aNDet83omyK4mo9OivHZpQYexzApRuddQ4gEokAy43552DlFiZuoMliL9QgG
GEdSSemvf1XbchQqIyb95e5/BRdoxa3P3+1cMvsETDSmr73mDMPmMcFVAliLSQFniXKXFdhxnHsG
+pYAup5Pz4aClHmHaX17HDqcfRtzVSEOf+cATV4VoMt/D4c+I7U+Af0sHwxb6NMZFJA8yRhZxUS0
LGchr8aCZO68Vc9b7IM2Z0l1nydpV/y0LY08d222ep8ALu9TGMinuDLmaygAaYveAxdGPX3kBBGL
Oq57ilB7gyoMghmbE+3xi99JBtTDxPE7bVgDxvjklwV/QhyWLyjz27aXbfTPDpRrvKvi0BGsTkxh
dARvlsiB48Ttpvy9biFOWdqieYpAvCrDFvlnBjWjc/1ztpelYayK7awOYOWX4wjL4baACnKHILTe
fYCMhGhDcFo5oziav2MT8Ui4xW9JYuMvnS7v9BjsnPyBqzonHWK3UgFjZdWFwmErSd02eip2BGuo
1vvyGMNQf3Ap2oyb7wLCBanPfP9Wj3JS/26Ms5IoTATK/bk3ihAsOwFU9m0ne8WrxZnroyWGpE96
8Mt6hmh3jxVte0NxrTpBlhmRjjinA+JbCSTnaJ+QJvXDu38CAsshJaXsRRjFcrRQjD8xYfJcKF9c
7DxBxrasiiT7iVusnyzTgkd7tHGi58ZFmlo8cdKgi8kYhv4e6YSLSnjnbdZUwwbmXx9ECqapqLkE
nRoVR4V5d+jtgdfKHJd/Cgq9dUt6pxdYQ+M6KjiHHLNNk1GD82RW+e1ic5HOpxBj2vK+TC41OCkQ
hG5WxJbMiL/iGYq26fySZLBKhBb/zVnbUnV9E1Mj9fQJ9kfYeoquB8+u5dJVBXxoJixIdwdCRjux
0nnJT7knKVTUlLrq+39pWAKMtNhIbPc2ccx9r5VwuaszA4Cf++5BlW1lKN/ouoRVqpIYSW1KmcS8
HJE872PlRCrxdfMXYGeJaKz+SluPilknpSMNgOtVc7mzvBGYMwVmBcKjP+HxLMpD67YexNMl4FzZ
6x1AyrdCFXbIDEAf8A4Xvj9BXCWJdNDExuL5Obt1MSItn+HYkL7QHexLXzSCKsrVpD2ww540kire
6bR6Uc6tnASvejL5zPw8Ar0YwglFiX1KylcyJt7Py7MtEPbpRZnbPsQNTzDkow6DGpTJtYZyIe8g
KtvbfqkSO0zG/OW82ym3yqHMXULsTDOo7JnvPPB4dlzSdM7pTkEBAFS1P7gGRXGa/npRmOZlnQIp
LgA8d7zI5dNv90zDEoiUuxn7jtQzWbCO99G8u5CbhcuQ382xO+Hy4HeS9u+THJrxnYx58i5KFW5K
MAXLF0iCX2HkHEbJu74970HQFmKHJvDFXDuGqXWp0Aarx4D6i0QI3Cwl6ZnoQ1twW1+Bs19+Z0Hd
rQIYdJVmZUOi6sIgal8TptjpsSZggqX4syPhn8mTu1MLmWGWjJPHstcHVlWpTt4I071aisX4xFZ8
8dFVA7MNO+bWfz7oae+SBZuhiDk5cCPMsNsLaLxBTKy66Af1w17ltEhszLByQHRic6/ey8sDKqGZ
4eWhqSW3zMwsFrOWxhUqvnukXbViHU3KphuBPfdIL3wfUp9S7mkagGMkolQXdfJkbwBoa57LrqJI
clxWwVqYUrqQhVs5oNlmk1WzRxHny/PhUCwsK3OyYnnXbvDR8+DZDY/yFOrp6HBB3A32btuzH3dD
d6x8iR0JSOM3R7nwgr7UvCc6Z4WBH8njht0SeHr0HJWh4HZllOMvV6SuPj19xYrYUYusLDRmJ4kv
Gp12aN/Lrxil/TMvPuBM6qYbclmTXNYLS4e+xUZgB2d4g/r2wfHX+XEpOeASVqPDFk9eEya31Ot+
4JwGLpYvQSNAZkEgCjx59NNeaGGHZMOTPFfM1mg7Z10DkqM+Q0v/1DxU1GW9BSecR/A08UpfUJzD
o+eYJID5QP/1dYJ9n9Uz1vi6mBWs6MbBsYo03znxOFzHjr5OAHA+rHBqh/9vXYEp2h4Xjyo+IGkp
RIOW1EIM/SFWlH3Q/Y1AABiUPplDE7mtvLGZNHzblHTDFZhv4aHJHKQeJO907DNn3G/e13qydpo6
ZcL6wG+zeYnGgPl9ijIEEvxq5Ua1i4f45Elw8+pLw6k2jVl46kk36gFtxxtyuXs+3JKGR29CsTF4
iUYePnOXYA0hXOwLhiU1WDFyo36fe1mtFm01a3pb1qm/I8EhBR2jQ4MIEA0EbXEicIfkoXw4sphZ
q32Y+rw+5jaOpTT11T0mlBzuXvWB4apyhmi4qwdNhwzQ6g+u62AVct1BR3CASS+6Xx8EdKNCVLNO
G8us6geoLWXXEuoOqxJIgIQYO9ld6mL+Jp+BCGsgoUzUldmmhQMQLPWv19zrFYoSC1LpeAl/LpQg
x3mTW1j9FGFF11xWCkZH2vIEhLNemRjF58d/P2oasLXDt2AWLcw0oE2NMlc3dU1dgS4pmGlGYhBg
faI5ldA3hDCKJ2JqBuWv7zPOVQw5yP8lXx42Yl5UGu0adr2a42y+MkaJAavFUxFLaWH82xsnV+qH
1cQhcBEPf6lX37FCc0QqvdX1moVrDhc0Th4HM6SPSE9Msf3rFUo+NqE7zbdRsuOA9qVQ2arFyKvm
kUplAJhiNZULqHExHuZL48lh1suFRTNKJAg62t1JkDq0ll8KY/gLlii2Z7Q5dycSmV4wldGLB5qm
1zHgOiq3xt2q7yqy3pwErxxNCb1sN7PL02qdTD8kUqkHGCcV91/VV47jo8DblJHxrirIFw9H+YSU
rcBGAwuuwy7IDqu4p9aHRBu3DIcNFjfy4yu3J63c+c/qzMwoYqYId67NIZ3gsR02P7qmrylx6+nG
mojunD3TxTorEKcGZ9rm8WcYeAa063ETKbYom9e6K6r8h2FsX7D3aheTOxwpyMOxixCE/OaQxdhh
027QP7q2lJd8/BxflbVgH5envDzkt1n3BlFk8TStNZI1h4sQnH4HSlpevVDCGaU5XBhagh/J9x0d
UGSBPbWuYX6ATLRYEqKCBlCp61ExeVJaaTOvO4CD7z3M52l/f9CF+g8ohmaVujXSgwqNUqteZ1lT
hjtlySWzCEB7T7tXPHJIIdjF6KWx+f77sHbkH5giE7syIuWVUlSJkQ9oIZwLVHSSTnvXKe0PTLP8
MvRWBVSXTS9jiB9KDXnfQj6p+OExVrxAaQJ76JxprA6A3oIoNn1znRgCdd6n9yzy/ZBzrG3ZIue8
9ip+4HnbRdu4d1roqzLdZ/ai6j+WE4tG8PqPLCGa9m85SN4j0YZrcZcHUnkRJIQR61nuLr73/jEh
kNf4KNEv+CaWiB8xd5mym7h8UIfreK4xM8IQOt84efdFJt1hnz6Et1w3T3Pd49kxVAWVWLJ09mBz
RSp4cXZmMXC0i4C6q70JiJiWtZnBWIPQYMmiNzUOEbSCK8eFmMIKyTHx/hzc9g8l38DZYRGY2eAz
DRD+5gSCOf92NH6an2fPZytWoA+bdyqvTvdWS1Wgyz1gnxoiqKoC9BHkZctya1gf92e9u8awHYNH
X1sT8biBxh1F77Wjv///1wloetz7UuQKtt5mFf55AnOmMsI5wUztvjfa93ecl+uUlRtn88/o4ah2
fpDQlGTDqjx+8u+A45XzQu+RYpvSFHr45yPFXRr3qRMubQZOlnvpa5R80iL8/odv/JTtb/56o95T
zSZz8fy59fzW0b0D0I537I1JeUohTV0Y5ABGQVQLuY4lHx0uTS0sj5SHWdaVHjsYgC/Ow4wPvA67
5ZqSJNpFwHCR2Wr6WgwrXTCx+6dlSR6nY9NiXgT1rzohe6QZhKRw9XlqB45eDn/wnDhq41HcCxXt
FORe5bxXPJF/She6LPJU4FfMMTRQsveX7wbnFT9J109wu9ih2sMvVuB2ZIPH9PBsbUaHrQbRaKlJ
iGG9/WlHxVWQdimSxbM38LGGKZmtkPtGhbvigW+nyUrMYp/QD9qu/Y8sZH+V01bdWg8qMfkuYAX1
CdNdPuAWT/NYZaXgx53XTfA3lcr6hrtpCH3cc/7bSQ8j9SbNo6ZAH6q7+s9xpUDiVVYsE+HtR/nS
raGCmbVRj4+ZwdEa3FkgP1roBmPH+Yq5kPFYJ6L5qOTcoWYQb8FUA6QauzrjZaMrYqQWGwLxnkO2
YFLo7GxNvHIPfnBFhjhyf1K3cLMuzIlj8u6U8fdLrNbn//xd6aIWx/CAnwSySr+JfP/pFez6RdQs
gfdOBxHmbRTuMOYUhS+bomDhm/0tfY1goygtc/GIzERa4EqkoRzNncdMVWpgIohlj+v4cz0g5yUL
4oCXLqi/1JapCp9km/AGqvhecUufqY7DneKjIB6VDLZosP9ppKp+QQ5LLqlQq4wlAPx870iGSEVw
zkuA3VHKzhjfwwlqgqotVXh8eHVlhr3fT43EcOteeE5j9d+6IuDLjz59950m/7N2GMOlzlWY6qBl
j0afiqRi0Sh4Ju0JrR/q+u7w6rnbdTirvrUZXC9Bt9Pv34yXqITKEruoXe9NzbevzNq4/1F8W9rd
O9LkLix0NREh9HpSlbvtoJLbpaumBe2AQxGzghHTR5H2ndUEuILW7G0HfyUJq7aWrC7+6GZ2oyFG
m1r5sw14K1zF6IhnefiRbfRylcRMUhfkqa//WmiYprPjbi4v6k7nKFCLmdN69QuzVo2qqe6/OjEB
bqJjXY4TzBaCMJetT9L/Pr5t3Lxrbk4vFqKXjXUjQBxwbVNLlg1PwrcXHVJQwQj0Xe2kaIweDA0T
+IWTd2SRYY7qSOs5TnAJelIYu4TW47EqkOQ8W4xgytnYuc08mqdJ8DUu3Ic/wv1+CgrOAN5pzTls
z0YZaNWvz0XcpezdBn2lLqIAf0HjvFDmEacercuyQ09uXJdUY8jkIdccKWAX1HnOMrimrgVdgIg3
Yx7qpv8YV1OW5AFcIS/yAM18m/ui5K75lFtrz6dBm7nWckIqgTVmmZo0lBGfq1Zh4uMfoSvjAVya
4M3+7Dwl7nkiYIjt5TBxRUDMXg4fJUDZxl6SzZoBKYtqf/knlTTgmg2XvENxGP3gsuH1T0b8hEP2
VfccAhFCPbxOTNB3KvDCt16R4I3rOABZ/Ld/ByXPIcXKCFXex/C14PbCykn2VGBeboPXruXAGORN
sZDsArX3ft4OkV+uLqmdulJ2i3zYWy3PjSRZ007Qpq4e0DsI+9Db9Rz7jJ4zyeG11Dl0vFFymNr7
//5rFrUHNU4i5SYwfB7RFpKnRPrsPEWbU4nC9gRFigtSk9p5Zz8z/7FxnE5m2Xby+AuOg80OT2Tu
73aD0hZb8cqbKx4wepao9ZQOaX8hSESTNf9VH3BJ/b8bsZDfusRPzQTvdE6RLxpDJQQM78kpVO31
nzej6l+8UaYvmBYhZFsHlvlnJ973cBQkad57kaapE6z60bfFE5UvTKHRz+VVTsDZVO/uHswSWH63
kRy5JjOfsdOdKO+OvB8ySJlKkuJNPZ5aVuX8MS8KeD/3Nye6RmAWI6wMIgXsCpygdSlxIaoSH2ro
JBsLuuMEXXVdSE9RYuPDIU6HvL/YCEsb2sv2mXeNhf6F5SRkX37QKfp7vU7sTpOCfxprAsD0kL8Q
OzmyFEZv2Qv44EUPt6ga6m+92UEyQVeJuIzxE2lJAzHuECjkGFSwCCk9Mw4u3EHWwRovdd0QJ/wZ
l9uHnU+p2DkodWR3ihLMSBdj7B7XYDzWycEHVAy0siDLlXnH1NHwFdyaiuPnGlGx2mOlmQgN07je
9JSoJeSofNYg4iPBvmlHKWOCjiCfQpIlyGMjRu+5sLPc4hoa6KxXPQxf4vPD+6L7lb7z1tHmqONZ
xWQjxZjEv5E8LoCk6ncfuyyaBfJtU1fm8U83VvCxidibMa1QpoaSm9o2a1u2mNSZw6fDxruLmX5m
WY+rZHdZLfBa1DjkiDGai7Vfd/JKp5Wr2QmMvQS6aoe63SJ3MK+DIOpxmg1vJxohhjjIm4GAw+Kt
YWe0bQ/BXRnehL/8txZgAHijBv8ekeQk0WLuj46iRnY9QyT81XtQ3X/9ydSBzHLZoAmihd+LUfQ/
BSc9n9bV6ua2DCvsH941tTKFB86s1sNsrJRJ5C3eJXlWAIg2fjEzAci5WQfR4Z5m3j0d5yA8veVD
7HyZOpLPPRxnM8F3aBtq/M2dOSSXvBbCvW/3WNZ2aN9kj/tkGu9wDwoGCKkdKQDfoQn/iv5PHexD
TptHPkYrIV57nehEmRavPXekgbHkECxDbWpqNMJHK5ep3KUiFF5YS+md/p2O1BWru1AVIMXmsYjl
2ktJC7Y6g7ZhbbfCgfBhd2dK5LJ12HOlKTQT8Pzbby2eqr+WJrTPYhCVyx+Iyhej87edZKesbxiA
9EesC4DAJkYJ4+SXNlAEpH2SCYoyw5ekcUCb3FXcVPy5nPTivNqljGiG/l9Sp0OtzMw3Eq2Exr7E
mwtfckY2Qfy0d82OwuDATz6q5QkqFaY0Vq4g69BpDfrIRG6ic4w8Q7mvUTLy+esej70pWgmZMce2
GHf219sGsX9a61Av4zKNa+mDRuKkAFyJp/2m1YrQOOmClWz/GjMJ+hH+Cb7l2cylyT8YSrXIIC2H
ygBxxVxU7QxyZ4fYLVIaXwBECIHgyGrZz2bs741pCFf/T/nwDb8Ry6G3NTvW7iI9JzoJsKaPbC9Y
YcMyrRuhlIdcBFr7xcK/tg51I7omzC3WyHaeFww9nOQ7QVH+oaGeuZH5F9mGRc2fkC95nfxXkEDW
cb6D/wBSP9GdoNVq4eic4Vg4pGqkXEY/xa9/tKN12LQV9f5l67KBUHCuKE83EeLgoHs39H8Be9wn
EO1zwvLj+heNVVlN+Q1+2cE4CIKVLAWCbh1qarQjn/MYt9NK1khAHA6VsaLR3DTAC11YXze7N3Ae
8/uzHEXSvIud+rPZLzfYGBYFa7OFmKhlbNwW3YxtEq6oWLTz4vefTcvyXdhvpEPFx4MsZkcwmqtq
y6+FDjVWzW9WPgi9v0WGG0gMGzJQw77BcRpm8sOrLhkSjGmzlSu635NACuptC0fGgXtkDRog7Qt3
fyaNF6zNBAtg5Up2sIM3HKHry/PXv6KR75O4mcKONaAE7Cf1EkBIBb2ULAtU2UG1S3qi+edftNQ0
GhPdJkPiv7swkcU+M36GO3w+99Hxx6Bx8fdgHv86WuxEU+6CZzQ6lXMlBChPDaP+0j3Qa8sa0Ov1
V49hvPowHlMlVTuEBq9Ue4QVD2ao7x8WKFzpBhY40SMvE5vIhPdGsxPPTI/qhukCvjpWY37+1TxD
iCjiczcu8tXmzU2UekyQQMMi0RuBz/t6UvqF29zBjSNIGPV9hKKuzS720ceCZ+OtjuME8X6lPsih
mwFPa3Wf5i0M57C5hCyy+DUvjb4mOfP2H51Yx/Q7XLrAPHCzAzZ9nVXne2lssA5Qjr+Ws6uqy4H3
jn6J+SUy7CKXAjWkRoGOWkZoDZCl1IAyhaiwSO97B3U7A3LeIy8/Sc4Zg7r7guVWnrG4cn/4Na+8
9n21lL7wSoSftPimYntQtgevOlK3pJTJj7cjanqG4F8uwEZPBGeHvsNDXNOpuq4U7AkLZHhiQ2eK
usJL4rs1gVCLTMokGwRoCP0Z07GBaVLXs4gBQM+MRPlteUbr2RulH7C2/+Mz3eCzsSf7laAWfOgI
w2dtkFtQiF4wt1yVE35qc7JFfB6i938toBnsDceS2nS0Fu7ofWDI8rv39oeyJ+3zJrgnkyBC8RGu
zIV3o53kl0S49LVtmhYDU0cKhsbvq7XNJz33VblkkvYXLcXMQI1TE3dytwWM3k+zU0joe2ANp/LT
gkExCNLGNy5youYP8lhdjdxV6H4DYxsbm6mnWb2K5IqoS1z6OqaOqyiQoB+hOXDeKwKMoe68FxVm
JeIEDwB4FBK4lfkM1KlA287xRTxbQ6Lb8DJoPyKPWuI6v4A1PiPwSYluGg4kFpBH7NbdokiPJcap
Z8/Spt5MPU6We9o9FWRSRsXLwU+/TXasGfEzgE2f+seGjto92rspPYvnUDpyPXN5SYkByJ4pZwlF
XWPq/YAlx0tLY9xt5ljDyHri8VUpOqf1mNvhNzFoKy/dvHH56qcSLl7nFFLe+HALDenvfnPEFOAR
sBqVQ7xE6zf4VWQLUKEdOtfmIthkspIDii30zaE2/CjebhQXakBDLQyIwnztUv+DyEUg1y5E2yGR
JbYSC8y7m/wzxjENsRe5vzqMG0LOQeqr277seYVXj2kYrqS5kbb2SxHefyhy6sZFyyUljlws10q+
rCAlTvZ4Ia9wbaL3VBlHVpJyaW9urJWJyMMdMRRFPpyIf9G5vUC/xiNZy2Eroj4mv2/Ut6LOwi2i
YCrY+ssazPYu3XL4mISRru4ELAyDkDVc+m0BoxljGbPEqJk/AAnqc6j5KgDGJr7z01TKWkLOIJvz
Z9ziWrFUtoLk0uA+vxSpEm4zz5mqOP0xYej245K7lsy4G0mFMGSZmnPzx3ooQePWTxBEfFNJFQ5H
xxCWj02QIK0q4uuF9iGEEn3WtiCWtKojMvxG+PKmP/Rixg+nDWAqfOgXTFiia/D2/A22KpQwZwAI
UGb1Uq/SWwhC1Z/RnpSuA0FiKwmJt4PXVs54RAex5WR6noAgt1mgDwsVnd6mGWOkV8h19dZvYRtI
jvAXngm3DpYz440GYVtmMVnUF11ifwsQXbYtuW57lM/1T44BFPNVvAJRWQ/aB1g2rV6jy4DGezjY
fa/Q3s1CKf7RHoCAdtdTNuMEwq2vfovnelK6wrDdGGmqcibQWIXXxefNXX/J+m16i05adJMxVyqL
3Tn24DzPztcGDLS0+z6EiduLOcj3d1TfLoYFwwhVQEiscrJbx2jVYWV2Kx2mDRujSpwqigDbX2v0
MrfiF5OhlifASxIxGBPpVqILqZHsJ8aWwn+xeAWqk5UPvx0NW6Cf8shIruDdF2up0eOz94OpRYF3
SVJM+V+vB9p4WtKz8JWRYqqyX3CrJqkgrugfd18jGO/HxAIHKg2fpjZmpAAWMM2HhY3ptgkaxwSK
VyVy1vnOZrDdjk90RakARS7NnbrU0IlLL7SHyy8SY8xB6M1SXpVhvl6TWXAF7gkuQTay1iiusD/r
npNLCvceEdHJi8KqVxeluD1VvBBxwDFIgCJYT42+0clgaCfM2UpnZ8XWTRKb004oB8eoUAIR0TL9
iG6Nc8EW9snWT7Ud0GQ2AXZiW7barJhTNzugN/YBx48JThL9RZdT+HBhrOeGAwEDGTu9oxm1bjsW
eVHhbQJZOKbRCFlb18AuaZWQVTNSEE9KneTqCoTSzaKIk1nZzbG1Lq/BTEKKY5O+ibXh5du2TmAN
68cuBfl3OfySNO3efPEr9DhlmnGVAuilTXaGXaVmZO9LI5233+aVWXx+Hf15a6uU5hqLAAykXs/Y
ZYPHy5YiE+6rKYMrwi4pta62g7ScF9Y41EP2dygUCi78CZgLER9jUm8Gtqk2E3GPJ4VkUWO6AZbp
5Mj5rgMiBXuKZzUZl4ZbwWmCTp/xX6j87vld/IJ/0rOq0MbOqA+1scNlygT7g1SHPyHbLy6/A5Mf
DBKiXp2hgW7l0chPjazF6h9gx34i0IUGIF6fjm3GQmgvW3vO5QMb1TXnPVgsN4mfvCbi0hZcGGWR
Lk+c7+AnBt61UG6/TQSUgliXvEH5SUk0SlxIhE75rBMeta4cuZvJSkobxiesgNADB4FDV2HDdYov
MIGita1U7UF/PFzqdZTa/fa5IApg185F1G4s7JXBxaPccoyxUIJbCZjVn6SLiyZEGUARlruoNYvV
up95O5AzbqLgHte4TO3ifR0ZcEAH/5vcaCcCxk0zyy0lP1N0i+f3XiDp4uP3gHm8Sf7aX+iZY62y
JykYcIV8K9UPzkaEdl+9P4N5lrmEgbrExcO+lDVKzMqgKJ2H1HEM0gTvmsatNPoIOt7Z6q4WRAlv
fu6WMRiYwMAlJVS4j7wVBWF7etJw5XCx/2UeJoUgVkypRWYeKGJadhHXebWAPbwlzMDHmVAP0eBz
qY84U7rM9S8Q7u5Y3ieyXTwxgqkEV2U3GYPgj5Dl0cTIkBJBh8a58EOCrECHYiZiGJAoQ7H6eYrc
wJKlx0VRiuclWhUl1LXgACRlLr5kKR4ZYVC4SINgtbFy0qvEQDNv7cBuYDEu4ocZfklIzrMmaoPe
f6mgZwyWpqtoRIkiEcoLORbr4fqe3wvFP40iDGTjFx1k2BWYvp7IJC0MMFyG3GhYYDyRrWIFInDn
up1bs+izpCT/LLZtGbrmsyKC0liuDxJm5JthMGbmSDuedpicGRZEIlS20wOU3fY5qxDv2fMiGbGU
TJr3YaSTU8F7usijZD2+wfeBEqVt5Se91OUwWRJDRLtWQ5tKlYgPnefnSx7dExImUz0rERLvr8+f
W4qDbh068dr2z4Kbl1JUDo4d3kZM5gNVGv0/4gaa66nJYJnoN+CEO20fTbp3TpVoGzfdY8RExqkB
z/DQ9ohi4GkHZdbMtP4V4c7xg3bj5n1yg/z4vRcS+xvIoeFpWqOZMrJVdHImBhXb/WFTdSrNmltr
2rtxtuJnD2oqf4nPEypCzGLQ2fGOGUDnr6XaesZ9dPgOU5SyYWGQWABetRja2IC7h2/qsa+N/2dX
FW42oTnIX74ex8VPnZcdOQCTjfUv4Hzgqbfzg+I2u+Z6PfrfWzboJQysq59XAay4Ww8WBcQZuh9I
tJRc0G4ZyGlOZZUkTvBdqhUXSWURR8+WaeavPTZ+xedwFP0Dn3ER8h9HOeIjLM5WYSZuNTvQWLmD
JUFTo66g6n/AAjFtYiB4bkk681g+lOLzKDrqgv+Jz4WzGmU3I2GWn++WfLZtFt0IopSbXmflte4Q
T2HlVgRTJJSnZvlbZCGo8aST5eH8xCHy1l8YewMAcCXv3g+pdxogQ5QOiJ7qYyTziuXAVWnG9FB8
SPRqCqBXBvh/Xqs3AM/UqJalFsGtDb8vvVuJpeMIJ2jTNZYvcUOLoz4FvdWvW11/6bHjhHR8dATX
lv/vXMj28hG4r1VKV1WiBgJ+ORtjdC8LV/21cp9rgzZYoxvv2JqKalLBz4mjOqtJCJ5sL40FaJun
OB+O4TLb6Ur12LpmUVVIZJKMHhbh3CYolCGVzH8kW0NRqTege91EMuiGHD/F0acgW8bZG+5JPrHg
1zd2Gc/3THDRQ0FiciNxp+D0C5exlP7BBkuKLiiJ4drUPMgAqgGao013msUoRlveTvgOXMvVSDNa
m/IZrHRqJnM1keS5urJ754m9bERUJCHgPQ0x8MLcphITnc/xdSjAs4A7X/ZBFcH60hBgBffLCKlV
pyTxjftp6IBQvR/phPK1GfoLEw85sjxc1GkBGzOWTWpDSkJYdu9O0OZ1CCFUPR7i4AHe6dGhcheT
waCQKW2F6TSF+jfjhsce8ZLUDkR47oy27LIF8L+z4lZus5Yu9T3jLKLP/pRCXK2/slO0etz2wk1X
Flo0cqXg8VKlNlyhe8W7rOXbTyrQhXMfHNWoysP9klhvYQnG2Dy6BKWt587vrKGDUSogNFI+tj4y
Nx+tKdPgEByUSDMcJXsRL3vlrrcWErnpAUOWHozEIM+UhW7pI/SWAi5RVyAvcxNKDkyHFxS54dMR
Pqf3UVQ4s61Xr3FYH85JNSu5Rp217LR6P2DwT31bw0PDqHw9YVvOpmA18+PfqrbXQu72IQ4ewZyc
79LXJpivEXgN4UihMozm8AyXQzIAWkcj81qpaKzKAGgHH5ShtIY2ckk92syYvC70kDhPe0+2k7Mm
t1iZU5fItEbgCkj0ButqJf1XvuhazMFkqrK7/FxQD40gOr2n6t+0HJxUS6/U6VQrLR25T0DeTj5d
dR5Dzm2tr6dS8t8mFRnu7hNFVHjcSeDPXjjRQ/wjbhJ+V9qKAe/ojNLqUA+anrINlAy9HWeBpiag
crauZZelSdFKGDRHhQAM/86+Dd2uO1D7fkaWADv7RJtnhQ1MRHg3Kb2RreJqzGMmwDMktAtIgODq
ub59zpcii8DcbWX12BpoA4iSmhyRBx8h1yd0gpg8Q49PToNoOSD2xoP3OpDk0+kE2phLrQNG5AaI
AdwcSafIhfrWWCWUcRlL3yCPcyL4SuaKlAHDyd0Tiaruofi0ciBmL6je1AK5gn6txvzKZvMZV2ed
HwCwK6OmFh9KhMDmU1mVnX2F8Vk4OjcKbZ0PRD6pjGs7xhevGW5k54Shr3ET+2FRDUqmx0UvX5/h
uMd5RctMLPjl6uxC9PoSRwuMRThJQiP460xQ5N+PQYfBPi7I/RAls7d3LN0VubbVTv1FbSIS6Xhh
On4xrmqKXhZu3OclJWAgmLL7PU1VB/cMOSo+Tpe+JjgYfJKoqHTfZXrahylKiS6jm8B2FF4nZfPR
P57npkMjxeeU7K94KKXfuUINvandGuwxMoPUgUtt8SnUc+Ty2E4J+yTtvFNntxzXdWVTG2l8WM60
84AYJiaixY4UhUVJQJ2RAhkfWfIuWbQXDQTCGICh1Zjh0Gb80Z5ZOIKEY+zDUVEjrVI1iLJSYn/6
ioXAjG2fxy9tCtNI2UWhcDaNRc5cg7Ncs8ma3+d4iVhoE4benvgrdcz/32680KkhnrywhTw9a6K+
gokUkdZiwHVWpIyPGJsdewt6W8VtIz4vDlyJ7WS7/CbTl4sqmiSyLbl9BSrSW28usjilULozbLZf
1phuJ3X0crM8Ym4zG2abL0fK7QL8E19pTX0dWUoZ5JDRbjGAbFjd5KMTLTfvp+9TOT/y3msF9P0T
SawGs8Y8PGzC8CW1aDdq92YpeRIxSYzwnJy0eEt8wiKgrbMv/oz7Xf3OA+djjqwYFSd7mOPFPZrf
919wXTQFX9O9kIS5bG21U+K1lEzEFXIo26z1QBZrdLSBgeu51uwiWou1r2vUhJiFlTpkJJvn7QVv
Zb1mfMDcqDY7+8VKeZe2tOP5gGFX2tIG/FxdMKyzO6vW5FuazIukHBiv5mMRMdtqZFLh98EGKcXw
M0ctDZqhV2aFso56YtEfTaV9iiYCVRMMIgbst7zoS1d/sXaTpjjf7QBb2Yjb+HPMxuAS9d/fc/5W
IiNGgVWeK2Z3ra3+LnqRtln36xwFT8KkL7GNWi6DzgAbOtV/cM3P1mlaNU1Dsv8eQ6fk1LkzbcFj
o1MWQe85eqV4CpOAWAIz2LatE6D5ZM3Y85Wd7xQkapO8GpPdoEXh4PcvBVohTEbrFXO8+rlGKcBT
+qkqeUK4ITlqsjswY7ZEffxsJKZRA9o9bDxcugKUjTckhSOcUL9IsD2Q/uGM0UEiuQTm89tGE/b5
jzd+TCqoV/4CvjRO7w1+V42EvquwlL9QpSwsMISSWfjHyUmMn9JKvFEANCVXVPp8Res1OfBs/DZd
pt0FLFcgqTGdrRT9feYM3wYZfqct2itBdqAq4z04MWsuK0iDHYEi6xH70rExGAnzg8lK2a31lo3w
cekV3IKVkM3yVZCfrwYbSvDguMSYjE9s126D5XftY94eghSz3iucwIA4AHY+rUB94W9zLEQojPx1
hXORa/aj7QQyvfNAHuZP8ux5YYzrWRFlYbju+QbhPuMXGHpykL6H/zJh8KQFsyBiZDZZS50VrpM0
gMrBew82T3iixEMzCaZN6alQqHFTtFSSGJfb8RfNrsUwEK9oTVJU0EwBVcgx17CZAYOhYN3Joc4w
qom9g0yM2sDTNqHwrxu+KQ5YGczNKfC/aUvpYX4ra6Bfp9ntRnVV+rFe7ARuM8zyg9DH1NusNcyz
AJj8/e36nojGAQG9oKgmlterU6PNVf3rNkvfzDKYet+mgUtNIPiRKSaDT4nc6tPL5tH6VyMOULcj
w3S/0w7r3Jh068TtvJZWrJjSG2lC5+5RIV5fMVnJlmY7RtM4MgKBBKCc9BrC62eqzUpphV9LQ/+v
5XFsSP3+ZlHyCgFS+5iBU7FC4tNzxxlpFTMEEdz3Ow6UkrgXKuzaAdGn3WKgxD/l4gKVGK9Y9c6z
Oizi9BYeeKaPTREo9YW1Ge+pPkHwH41ST+kMuSjZwuFyXVk2uXGlg6zQH6B2k3eFwdAqKGLp57CV
7RZkdGTJx0cVyJIKUWP39IDpHmf6xaRTzk4HoEB4zfoYKrG3vqR2b866xx1nPU1kawRZBkvqfjJP
Rl+6DSx4o9hkaSHI6a893nuRTGglWv7h1fAqzM6Q/dUUngeS5d2m6PSjZrz9VMCWjT1GT50iApHu
VOo96pZJ4v+hbCe6FHfKEVr5LwRJuwjzbYdz+qGIN+BwkTsvfwrwmRwgu2fbIikVB+aB9/+pQXta
bSARs323jjTqjLewTb7/fEwDWtQMPdDM+/eRWWxeF0ogjo40EVMeeU+ZA6NAX3GAuk0pRewBJMQh
sCm2uZ91FCDUiZdvNDPm6/V4ZNVWL0qTsqHSIj1xxJ2vUqPmPg1WxFbcWngZcAnRwOFNYp96Qayw
6AiDdUvem59aPkSd62QtJSJnk0E+vcmTeApzxM1Dcg1vkSP3uYQKQGbsM3Zh4ICwzWrnNosQmBWA
r2DDvrN1115K8oS012TSNn3fPoWaHqwcA75LDkFMzqu4MfdkERU0PhacPknrwHpzQgQcy8otg9SF
UyYAn8okX8nT9fGGL7I4qHBbkZtKEwEWBvhpQqNA++odBIs8eBGVJ9n/pTe1OCaxowdMsktcc6w9
JEdHrO80ZFYVYjvOOZsvZ7eKl4Ii4L6+ylctvNFBMxaQzju37834GSvR0b1KoBLrbUCL8+xDYDv8
kkomqSZJEzJnmorIGXmum5jQnMLUam9cr/l5aZgAI4hS8VbdhebQUiuqGBkOH1XhnzI0hnXehMDr
i8J6wvDUHr0gNGF+QQXnSW/ML4ga9b32wgcIFRy7SSdC8QvlYlN+8NqcXb5UGjVNu1iuvTOjqbLT
2Zwz4/oxImhnSh0d3ksAgKaOIhww6ArBdFzJ7oKlIgNWMMn4CV4TFynSUu1Nq1jXcNtrsXbBRxyK
zyfuq+omVLvZ5SE96x7pp08T2R0DPClNJThSvEs1inG3iKwuz3WzwVPUwa4vmEWycLRwe3w4jBM+
vGySj3AhbnAuJfChu3pmBem0kdHdtduGgCoy8clBPFIy1trPGIUFZ1tNkMb0sM1G/VXYddI25A7I
r1pjo9vxgsEocKpmvXELyo3PH8ZPCljiJsgTblM8AbnE5MzMyBRNq/ISSCBkCh4CFyTOTGK7322B
ALbtQlKfbFH1kMUts8p7LzR89jzi4b1IsFroPrJF0mtEgzo8KyNrUH6urDuGT3Q6JOrEyF7LyD9M
nnp8/B4ZIxImfkdd5a4wnaRZot7Ujh5qkcXEEFcIswsTlvjHulWixObo2pwUJ2LY51zwoLw3cMzK
jo5ltO+4tpblWdttDILF3cmwVyNgN6C4zQ5B2ekX41TMWyH1GMUAah3fQjzw7BMDLzNvYASUitOM
xGqctQ3Vj/7RiMIuE9LbD+sJZH5TQuyR5aDszUdfocb9fSEpNBlPmL6WawAXcfEEXYAn71V/mY4u
ifzHAQ57cc3I884G77X66CiXzFU0vB4E4BwQKzFRyglwHGYeMAkoA/dkWfhE2Wtvmetp/lEgvV7K
bjzjBCmAo62MCkTZbFezH4Ho5/lciFU6nk6uhbJQmcKZviwGTmThxHfTqBM4t9O4akdIGDuYkHvd
kr6O6sxVtMHgGvNvKvQH2lhlHSfhT2jUlkzbuA6XrE3rkjUI0/LzdmoUgkTEEuKgbE6pSc1i+jhk
5kRySWLaOaLkEe35NR5nvY8bees0hIJiZpxER+IUysDa8X/keOUqypFQODqUI3f3qQxqK2dYJqo5
+oZrUWDdEb7cL669nE9qnLcR+R4qP+U2ele9r4Q06wHHind0HifGJK2mag6aw3O80TYaDfND9rEh
uuIvg+shJ6Qac0hv4OwkpS233UwqVsM3C+YsRz2FTaCsUwkfWcygeDxlbhOaKpf1ZqNAqhefm/5Q
C+ubprh2iraZPY6zpqdzNQslHRQ9qW6Ldi6DajUHNB/J1oslbkPlaQ1Ch0PFlsBYHt2RBH8BIR8f
KuKdEsArc3fPGDqJQ1jtIOejihCWetHYTViSTjy1oNzECWcEF77InGt7eQQk/bXHI8CsqDf4qX0A
esKdsxRptJhFoc8j0ySF7bxadZiEgFQp+jb1/6LLshKgx6z7P54fN6v2MJAhVufJNtpKMHESLHLU
KCVf3+U4qB2hxbxNeN3mP5wB7LRNUhFusK+1CYqwqEi3i7xKGdIy/6ol/hZnqMcfcUFDjiDpEdGl
bmhzhZK4cmxNqyMlxDXUcaMfUIxeNjRVM1QAqmzKvtz16nyYKGKTNK6xkJw4tkQWY2ZOQcUCHlEU
TJcgDIcJqimAKVgzgt4qL3na1426e12Wn/sCxPOLfGJl0HJ8H6P4UP3q+mpwgbkhqUWFXXjp2Jyv
XzlYWKWpL4Xu3AUQEkZ5B5dQ4u8W7KDok1GamVqlJLqQ1cQ6hmZa2kGG2m2hKDq3b6KkTwtRABwY
px5ZwH/lM85++ZvxWNXglsRymseZHGGwJR29I5BesomK3x7lIyk0CO0MtGBHtgFGVnBagxraTPPO
2QD6Q+ES3cxHXJAGTLSfcQu7ESGX5R1a1uc50VbIh9TlcGefISL2b8fo1alLb6LAeE2HetyGovSN
C3GnLYXvpv0BLKk/FDSx0e3WB5kWhOCt02eGc1bU/VZa0305+V8qIiu8QABOri7/aABVvnz4SyS2
WssbR0ZQ/ekwNer8d5lua52p4w+BHMqGudeavEuCM/F41dmPzPAG3ICEB/itiDK+x0f4K+HPf/c7
6uq9v9uA56w77XZ/uiSFaoCkVJPSgh0i2YtdIqk38vrpZPFGi+QO2UhUJR1mlVZnIB0DUbiuCIHa
W47X28i0BvMsX/kOhtS32UqTpLCVu2/kBiNxzETiegcTWiJyKer0WbRERl7zZGcXKAZIbm9THfyI
zyshuh9cdfLQcGmDfNCULsKEOSa4L4uwCwQMwyCDt0q0cm8sa66/nbOrYifMH7SP13IHAowHU8k6
8Jj6EdgtousqBTA9idrmZgdxeccRfAUiqee1EwdEo0Cmc0+9t8ac/tUOCE724ncqJHWbiuZ0I6Qw
tmfEUrEBjC8e4IXVk9/oABzwr3eGw3U1EkJ5V7VITqkA1kbT0B2CSceEYBogrZHwKyx1jKvoXqX/
PMZ9D8N1c1hX2VUsppzCeWJQDDccDiJW3DZz1Px6lIwX8g1d0yHrWvmj8l6JLsYGLd5cSk71/F1A
7DLOJD38mcYqfRYaylzpPbzJITz5q9aczqKK8qxQsFtg0RqPE8lV07ZdKmr3Iz88jmsj5U8h8nsq
GJ4f0RmmcjBJu0ud08QH7W3zy97F4nntLnRIz5bAV/KIwPm+BUcQw9iUh/k9DDTr/uVhIlR4TJ9o
4FeL3js37BGrvp9Kq2/MMAaCXpuhaN6f7l8uqJ3NR1Qtq+688t1KnSa7RgacVRGQXgH06d4LQeP0
Qo6p9DHaS8S2ek0fOiwm8vMJyOH7tG1JSm5tNCUWoltqczuMgpmqeP2t5SS/gWxtxfeb/cXeS7jw
kekfyqC0Mt8urgetpDk5g0uafhS9Xb5BiET9Ylxvg61WwabIuQMFkF6Fpr36AUFK8BZKvfoRslxl
DcQo0Hnko3C7ODMOcD0wgY10bua0IleLkDA69Cm6SFgebCIE1770AW/W6LD1H/UAwPG8kj8yzovU
gCZlZcXu18Ch1tsJfDKMjgbaiEzPHWk/Wh7LxEMyHl9yyjyzyhLE5s4kjDPgZ9vR6tqlR8UNbX2D
9HW3Gg8YIQM/rAWC1itOWQkDqKBF4T7G5U0qFF5jS4sltrFgHJixxSc3/syZuJmTxlq45QTtl5A4
fqadG7BnuHWcPesO3YB8bCMkHoBNChcJcHBQGqoHFO9POzmyDoPuOuLMGMLiQBLx8wdTcfm6D3iJ
ukKl+TOPBTy66lFAgauox1/OoMbWpebOlmZyrauOhl7fJR5/l2202txCM9y2Jyjnj53QmE/tBgk6
5hewkqKAb4eE6vQtf0jpmTssfLfu93+Q2NwedVkW58dpCXR4GXaBS+J8pAyERYRjPncc/0ysGDt7
Q7S6Q126Xq4wTrIgjwpmRSnlbEB15JtyJ3LoDWsfjlxwJX89dXMV6p6QQF6UENvcfQF77iNvgrcL
8YCtO9kgdDYLMR6Xf9LerRUj3TsnJOKflU/CxG9JLNlnJNot4lwyYLrcUbdf39YWNrVmtearqru6
adPAfNN5IAr20SACQFynjFbCS4AjsVcgXkLgIEdypWpWQgxRnfmWuX8O246a7udSELZmycQcp3+g
uHuKeuJTnbvFIS+6MY3sMVBmEHmcgzs5lCrVyeToW/DOITmn+/7qoBs36wAFyOKCZ8IFp8HHbaJk
4HjbeoyF7vTZJG4enG+1hMdCtO2RjDMnc2GoGEgMmgrism9Oe0sBxRgHdYa7oc2OVQ0CSw80swUR
wAGEcCpSLXe6B5nmPGwTE+b901fOCB+qNsnmLccBdqNVzOOoft2e3epkFsfQ7TvGku1TM2aVTZX8
aTx7WKAlsArtYMFY15pTOCgmlDd6jdi5j379WW06tOX/ur7zcrOrkqx6RzHmxfZuk8y5aplLYaON
FVUjtmDi2BJuQvRZlMvn9nOcfwQjSpFqtzRdQRvnhy7EXzjXMUW+piaVWimMqjmDsr9CFvwTwaxQ
RA6Az3igcZawTPP8Jx3QpaOfLYKW3is/ccnppoIwDltoYZkZdFdwMHyxTZqiU7r143J4SI20DzQt
jUaviAcL3cYZrVklJEjJoveq289XthTagc/7A4Ab7nF/jRSjjDwRhBV06PiVol1XjjgoHHM7Uj7q
7nLrzguO+0b1JFeRkvxCrlfnkZvnagjiE2d5fBE56iTZGgE/Mvar542LHBe9xHnO3INuP4/L7QnJ
TA42rbe3wWyRQv2PS5vfdaLRQYrfXDf1cvCm55swkP28mDULlbXFW4ybQ3fdtPLGVIY2rSSqq9ms
S2QCAk3PHp8UrOyQchy8fUw5TouwjQIRMcxCf2HZZbZ3dr32uGm83kDSigJiiJmCAm27abCJtcZT
4d6GRw422mdnR+uk5gavEehllkVxcf2a1rmQQiaCYXMPGhaMcvCpAzDPpChUNf1cuIRwJT9+uNpu
1o3klUMqxTt7gzwEkeFCbRG7ZBUvpxdM/22DjoKZErf222x5Ofw1e1x3VWhy8CwYEZy4Tlq+F1J3
RpyQy3tnvVI6C9kDRY0eoXp9jW4HfNqeFbXryGWEaudjUcb7LDxbfg6Pqao8Eu2r4pKCGlFz1XuH
tPH0uJL1UL9lMDHW1PjIcW8Rdoh2EwIQX/FIpJALGph7Zl+30fShvT0cGKauDrucE/qw49mT083A
q/orLZ70h08dxO5y8BAhbXnT18UnzXPpwlZkNqhMa7xe05zp+pHmH8dJLJWT49OwenVYDXYigreS
YBKe9oJ2MIZgOy+0gK2u2mS9weXJjwCQZZw7S9wWdQc6kk96Dc0aWlBwXpuu51fHr2zP++iE/ztw
1hxkiI2tqRr8mYrB9LGNJC+1e6PfDf2asd+t3VZ2Nc8ut8QHK6iZ+Zrdp7bZGy1+GmZog2gzV8Oc
MEt+lGq4kyXA+hTP9Stxl2kMA8RGXE9v5naGfQJPa6arRlJ5Y97WeH3FR+3J+KgNwHX1yv/RpC3c
bxOQ1vyHdhVf14HwKtlPVq5ZHqklnfD7bbM5fgU+TouDGx+0ucm6GjA1bH3WwJwZKHfHn8b/VPUY
OOmQ6SAD44dpoXZEa3mbRponMRK9HgbhoH81Vhxp9vsF2C2j4D8U6HUKL0+4/TGr4ty63FdvGDOT
GsBPuxE4Fgk6Q6ctx4uWHVM7FawqSgozm775sDYVV945FCjxvF+Cbvi0dbcNSDiuwCaO/ljC/ZQ4
gikp48SKHR4mkXIlCF3BKF5Ixm0sjbpLziTvK8mLSBpNarwPIEBZ28Et1cSeGz3uAJqf49uKaXaG
7VjVC5nPjDN4Kh7C1QF5aNOZ5dJGGqdTQB4TpqqpeGdJzztGUblnJb25eQwA5qEmz16ZqU6EW8l1
2KaGLerNO4d2UBxLR+125sslLy93Uvf1cW2JT/EhkIMoJRjCA4Ak0Qb6UeYlz6XOGIIlnw+2KwCQ
hWcPvd4n1sC8ONJxxpQvqhsqEKIGeUMHWV9auoTVSYP60zciw3HOzayDi6mjcUp4W7XzJycjIxpX
o3PpjJXybn/Dca35tDydrIktadCvh7wTH02FmrtXyxTc/O9dNPFut+gGkIgrAE/i2Ofy+A0WVujT
Z5VsrIn3YgP+Ig9Ng09jP2pAbSJmi+QJHN9KgGsfH+WNEXLQ5TYyclq9Q3TcFh5V6ezOdQxMYVJA
e5Xr5GA9rVVNQRXDZxFKTfoemQrbNIfnbdvrMhN5mZkB4Zz+m6LH2R13wii/JUYjjqmoY+MW+wZM
0PZT/s3UllrAdOfrPP31N9Zk6fRVvcxX4uCf0xaS64yUS8UfSOy6tRYcyPFZRlU4Y4QyBrAyPAKm
rrbUJgk+j9lniAOGdpIyRypZqC4fjXZzkBg1n3yDjqawU+kVIIKH9BEB63CEsttDoMpB7u+NmVZN
pG8VwjhwzC0KrRnvLRjVFHvJLin0iYYtn92jGqsi72zC8FtLJ5Yn/NYZmj3Fbe6SDXn3DdLaw5PI
QQ4BOXqALNUivcwF8i5hoP9bFXMM9DRKTjgdDVtbS3wsfx/tDt6XpzLMjPkG128esisGtwauRoY7
Orl+lGY3s4QEaEi9x1M7+QOa5OLR/MAyDVX3Fe7yApfTEgd4nSTKJrDMZbn/ZCgcdjbKKhyqsdjg
GiIzxCudiPP0w/9CZUzeUY1DZXYDuQ06dOc51LIUqYbJDZ8oTjcZywRCUvJcdgjV20HQ0Rk9/UEz
DvV1LauM+zSuynjashxKdlst/M0DUR+imG9LI3yCtzVy9bCxVXVkafipfeHkLtBEDXrDe3OAp01G
xKTA8P4eoG96taJddfYGLgMLFMdJ59Ie2/ysPmk/d5KYJMIMUJoS+wG/eOzRZR89Uet0ndB4WRK1
O0WmJn+FVSBEJU/0pGK/K69ZIqrfxypQnw1fvw83lQtZW0udpzk2SwSgxfh6GGDUc4/oeRNiSGAg
s4WWuhTj2LYyl00gv8Iq0DMA4v3ZyH4pNyT6HdD/LfHv7C9Ykhrc5dfn1DNx56dsTCb2pucowHsu
jIslw57CwTaIaWj3pzLjSqPAR+5g05r7hTDBgizCF/cuoQsYcOjuWkwcXwI3r8aFjGjeGfVvy23+
z5+2faYhsHO2NYbKz0RSjcrp/Nzr7VDbFgLY4OybRWorwaJeYxQUOaa6b1bkJ5hV0Hp77q0aCKLT
Imc7aZYTzXfcqDcloExvxHyGBNCRcr6jYfadwh69Gz2dxv6ddWMWogHsWPmJGoaG/55yYiT/Yxmf
lUmBjOd00ijxJDvn2wdzc4ggVBKDs3ha5YlnhHPE8dhC7h175AbM0IXduq8DqAdCQs8mt0KWILsy
W7+XhpSiqfY1FmmJXAplO3UrmROWLHr1+ej14VTxTk5tmCInipOz2ToYI9GVjhhlzecJqM8WoLhV
Reepm7yvj/0Ak2d2FTWQqRMq62IF1kX8VOhcGGravuFA7I5Vi8kZxXawMilBicDP/H4MEWVOGs8Z
qJAM/PEoMtzSrIjtqtEPQXBP5eyuyMGQfMqXAk8p1eQDkKvtDZySnIvUBCX3roc22Zd3FC1k8YOs
E1Cgpv9ZWm83/a47sA4tOi0UDLHlovLzVZdRt2FgF9UmBmIDLPvl9SADh13GDQ5jLTBFxrXZg6ui
HDlizzRn0jk3IS/DEasESSqnKllx78j/vKxG74MLX1jD7rIOv7hlgkyeftcEi09hQGamtkxny2Zq
s5mfMVK7h3CWFyWZwSDrN+N3Nf+Arrun/07LF2XfGt4QEeZtvVCGogrhbOjND2zzTMF7LdWzCYFx
kz52y+UDX+XYwSFOPlcSlZIE4yNk2gWt6g2qlt94OuuD4LO+/lDD2zX+PUGYMmrNtS23Om2x9zkw
3CZhawUd44W7dhIxzchoH0JyOtRGB+uN5y3/jmmuOuKtggGX/OT2usuJCZ7cj8YM49Uk8Hx2nJao
211qFw2PVNV3WAd/IHuqg7KsIs2ELHDoU7MZljtjcx1ioPiCdmL5GbGry/8uhvWUcwrpIWcq/nQJ
R/U94L9G/ZaO1mmL/mYgYSPQ1aG/0GI10XBVtqNfchuZte1ecIZ3i9XMWvpxaYv6UOqcf+X2P1Pr
r6v1zkDDm4BnNl6vhadHpN249USkujNdLXlC4HSe726aFwLMOiQL63GZz5GJRJRg9XqqOQ5iFgz9
gsxSZkxl7WMjPBCaqYkjYd8+Jv0thpEvYkFObd2zODoFKyzWAqJH00L+WdJwmH3JaYZsmYDIMyPU
uFXrvE6W4WWEq6TSe9PzklOuv2G115VMYIYtrDt7K6MuX2Ly3ZAELuasb0SyoR0QGPGhyDh4vj1W
a46ycZxbfN5KFfIRxtczH+aNY2UQXLUvT6//hI0J2CjNkBzwlt+HxJ7U09k12rGYPEP6TBxDxKyq
sv/OOPJpmChlXsFV7YifdSu5jPZT5m44GvPi/uZy5JHHyKR72QSJIIabEuguxrFd7lOMoQ2SQ6P+
hGtvm2JEYMM0f92d4GuHfGygZBvsD98urpOwGW/Ny3zZ0Uxs2TShuxzZ5VDfevLNDLv/iPNmCG3C
DDo571yGLfhZYR5zHNjPIJwQttWD+smKmEZDDVe5dWDtstbO0bsfjEm2cBSEt6CauAOVyUmpp+ip
vaU2nky2pOte9wFs2rWhvcsN/SbDUFgNjE0SSjSsf6ZHdsL20SQli943ma08zqnnzqdpIKniMC5F
vTIyYEjvInZ6hNzit0HccejX+y/zC+pWAQRAQjWiBmMgqZDb+bpbZUPadFRctNhYLJs0la+QBBpV
RR1Z8xR9nJfb9RSbNgCgAHTt7kYrv9m/At1596DXcCEtpqt4vb5ooZZshX1bXbDRJhhSlcwb+IQV
DQcllq6sL4IL6wBr/Mm0KMhdFN/tllDw2JE4qHH6fUEmZqeVMXorn0RiwRYT5cIXulDD9fW+98Yo
auPJDUEAYFmsFpnZ0bKTrImsLX287N13SM/vGNBCeNYyGYQglrihhird/+2v52378V7tq3PI33Yc
FZ+4iG04NLt4avopL2t+9gRKc89WT8h1Alu6SC+uQOZGyYGpwLYBQ287WtQvK3Iu0GqDcpq9UiDV
5QDu2/uC0MF9td6DXgMllPSiTQV4ySPRIHKaZ+jnh97eCOO6st8QQcZz6+F3OfUKMhuN1ONI/w/8
Aapyvf6Yy64IeZ3Lk3hk+fFkRfHtr8042l55fbp7aC8NdCO3guByJyaG6b/kKhWETx/vHTAG5ApL
WJP6dlziShwuZxusgfcPxHv43vL/qSbzFv30QNiH+STNdt0Ejkei7p+VQ1xPpXi8bhu3c6CJhWW+
1ZNoxHJaDsitD1FMrkhIcY3E/7RNS9Jk1Bb2j6r8BZwSfuqrLdNfV99CzjFxoOsuangNwA7zf0SQ
aM90daDksqJwxfxMwpv9swuMDGTlSm6rO8hcWmOZ1vFSsOKZsQsJXKqWuxGSEBuo1Ch3vwA/Qpu+
RCf/jdQAvAOsHj12st1NHO/Hihu8nXCA4WUN9woxbn7y+bKJqswZQAPLSLq+yNz6SimyvpPzAftn
dkkIRtVIZ54sqwwL4AenWIxublHmiZb9CAAngTsAM/pNbsOyQrZeb6jI1Q6qhzCjScOuahX+tpBx
ual8fT0l3hb8bQuafJ0eMUa/wqGp/CE3RSe9/VbCUt6CRk/Rw229jwYeQ2lGw6AKPtfgQTDvV0jK
j9gq4loqc14Blu+js9HBZ4PLJRZ/9scwPURRM2plkNEw2EUBWxFSifDpO6J0RFy7hXVl0kaOHi+5
XT/yGPnjrO57EB2cZ2wr9YJ87v0NQPdYi/C+gqOvfVBmI/dm59H1WuDsg8Fu4Haw03TGDHnohEXA
BXy/KpT2nQ1/yWDMBBtCNcjRDX+3REfZLkxAILJM1kBICCusPW7P80A0xd1eJ4+RzP1HmyYwP1mP
yn4P9BCqBelHWG4qMQTvY2FnBB4LLp5BCeRxr5fTIqmS9yIJfwfFS2a6Janp1ZQFEBWtJ9Y7uoKY
3lQ6BiSkXR5HlN5UZ3Z0aohc3ycz9Hzvd0GZkBbPAS13u8NHKdxJisLk+AKTa7RBtVYnS7kW5vbK
jOndYMuAZLxF/LYrfCPQm9udQB6qOVLiLlVXEKVFWq7WOWt6ZbWmdISqGpKM+EwyI7gKz12TUy5j
5LbmqSIhbuFEOGVoFpcEWhnK8mCfSecvY5pe72WoZcpgPLoG4WDPzseWGR3hiF7ypz6GmCYaOoXJ
ISkXN8st3cQzXZ+L7zH6iLAUr07uJ0t9mAsYJB/6VBWJ5uDIMCE8vV/P2DN+15OyjjJfs1VJojiS
UxYAYbkzepLmafL5QfDGa67l7Y5PlF2or8T0H3xFLA0t3Zrvm3+AV9RT7MyzK8YjNZaJ2DPyEN0U
UUsb1q6mFUDS4a72P2189hcLDirBKkvwAh77EJcNEz9AhTCqMFhdt45+eMQMSAXjcoIpEPXWUcu/
/DhC0oER88jkCVATvi+Zh2fNbN1XmgGL+ldqDwqfREyBCZAWRRscXE+X+/zfksg1r2f4iWYXrHpl
jby6shfRq6KuW4EwLl4MVPylEaFOGQCt9rt5R0xzWBOpo3QnwbNnpSdC0UhqqCcBa1wIgDyMx4vX
QXdPG3KVKeoic5TIgPh6lVWlY7jBxpq2ljxTzLU7/2JpMlXz3ZsBwSq6GknIn45ngzAbTCPiDqBS
Htl4EkhcQ778usQgKav/8IOXGyqgXf5JFbW74+tvhvpgCCONT/60+kUTYN+np3fl15xPFuNw9Zuf
wJ8a1UNqugOlD9TIf1yRbVh6P812LzZ54GuqFjnLVrosD0O4BMlYCyCAdaRoXh0yDk5fmKkBBNjB
UU9xgykIhDoRnHpoION3DTyKdj9FRrbaDCvEvgctrzbNVHgPniGB8DAsPylY+O6Xilp8yG18LvKj
tgo+1HXpivuxWxY5kW4F3Tcbu58/nfR5WG8b5X8XPH895sQdZP8+lkPBSFy3uvMoK/z4JkFFIzu0
1CcYjHdO3vaOpWUU/ltok/m/foP81nxbmcIo27HAPtKd0XTD2UbngJGZPvlNdU1NrpMcafrYlPag
ZKuNhwemelOzgpupeQ9hozaQVANQz+Q6RFmsiv/VP6RH/jAxgqmNgfXEwzX6MhHecNgH6VHMrKPC
pGnism8729KwrC9PMuTXL1khJL3BVabhqnmEArLWKuc1EM+Zwn9QpcZVoKQ87mZcXwxAqtNTvD1w
/hjvKmsQR+pZEWRUf5pF/jLxCVVk0rCY+fbomQlWrH6C1YUeYVUpUH4FWFLAdjJDxTNR2o9H8nxa
62HYGduPZFKuAnmlbGPiNTCFMQmxlvelI+V/J5dWHz00FSD3QjzzW5ZMEoFXsgW0Ra+a3MEt//bd
5aMiO0+n/jhfNgPIcpF5X3npfDf8pNdFv7OJtqgXEJXifJn/iKh7125jh3g1Gf8TLwXrklklnvHU
ldprpz5pMpsRiApXdQjNKQ+UNasX1ToZVdX+bHOzoe7vzSSOyf1C2eVTv+Hh+uYeOhxtiL3mqXFP
fuNtOhx3TpSFNC/CdJyyypmekrakpC0LZw+QncZlfbv1eFRxG3TiZuMDnDnNkmLS178cYPVkHXLJ
Gshb/Fi4WxhpiIwg27m0DPLVMoy+i7s6AS30TqfzJo+24qjxqmV9NZs86ZdHEdbh8kj/QYpMc1pM
8l+q6VGDxwq8798q01UmSZ8dMcoVPqhQSxKNrXmQhvybsa1XFoH8uSyytbTABYuXeLHty2w7ZEsY
yIujq217SNlm8VoXJEDnisQdSk2+icamSqIW5mSjsr6J8nnDLP5RapGxvhNZovEgcwI4atsELpHW
NSiecAWKcS7OLJsb6vxDalUD61xffKiZieSupxmNd1wW7hAM5gOoaid5nOggWa+ii4CxmJa3LcZl
4l0leg8MaU8mYqj/rnqF5oLW1PKvcXPScUE5/yaJc7KoLrfUhx1v31V8HS0RgbMQ3jfjrXEUmFXz
kqESugq3uzH5cwZHETNVLKStb69PAf0E+z/x1W6sqSWY/S48F3SXGKisAf5mT7m8wIpN1oXpuy5G
Og1pXGc2NCfHz+8hPU1LRBT8GU4G/cg+/y7etXu8n1ZWANKLtaaLh/1u6c5IFkfNbH/JBJnjbN+H
PazJxgbW/3808IDuhnMm+eLLrNTI+k3XD+QUwChVoBqVLPfj0yzMdF13ars+WITK/icn17uK/kYj
evazU5bbOvtqyhGPzF/lUY16A8I9zazBQgs3P3Cel5jJ3RujYDdnZ2SgVe33WuduBfx59t0DBZbc
4StkceIMm5l0y5nSr7xxRFdgU9U7ga9OzEa0+eCFDEmcBcuP4ZOXXl7WwAnAKmhW5gn7nXA2sh9r
5x4m0YaM0nJIsESLOqeDDEEpVAjmgUHygSb6TFusLFR1ujbfe+wrAWYaR0NfZZolJsCgO6VB4j75
oNRDVIVuGYDiUuY2zx4xjclRYIDTk9lqcnkF2jj0uSlZeAMeooqCwPMJn6b/MypZUaS8GG+YLGm9
LGSuuj3l5NwAf/Vw5inBJBOihzbaemxaly+ANvUWHluidXVevz1mExXBBGtXvD9gu6c6M+TEp1wk
LJCHQ+2SF76jyPKajNfYOEmz+jBCFIS2FUZ75q2nEDFwofutBCbpEO7lVwRaP4008SQdIww5zItq
0FuxeABdcE0X5CVLrkJGF9u+iIg27JtLGND5Vq30dc3xYxZWJY8Lt4sjDVKmamEjiatliNI2aspA
wPPwNK9j+tpeLD6p781NPT7xFZdxkhfPl+xBZSId6cPMWCGHlva9JsUv+HV9C4UGKWvmPJKfDd6A
Iq8ULh5E4JnaGoJH4I/GZovYliGQBJ1I22dp32N7C4iyG+CRlswNj6zlRHoi0ZcCn3lbpVALyZsf
WxYTQQgH6X3Y4uvVvZuPEed/gFtul0FPDCwq9C2E6GvujI26WU14tlptbiRsMlxIkn4gLvaScAUB
CErFttEHdSMNkl13VYVGFQlzQDEG13bw0xMqc9WSA4zIGT5XPDjFKZbaaHqRneUCtXrLRJOmkTMx
3fBE0oc8mCCjp+ZagLeXiPnhy9+mMtozZA4IrPpGJ1JeofLR96TB0O0Inl6QUjlMc9UzkompWp/q
BYmAFN0KLuIqRKZQl4JlS4q79FvjunFHH8ID/eCClklGctp780dpHy59khbcPW5sjzkK+y6x06co
P+30i5e5u1d4tsmYQJyOn4AWQ2ZhEoMHRW7WQKoKGJaJGggUD+iWCtZPdP6G7LdlPwYRiAKg958p
qDogKQGqyA6zyAPwG3+Sxb+XCC9yGb8bUKDhjNn5YHP/i+Avh6Dys25bvTr3WbBcmQrup3rYS9W0
y0+dpfKI7HIaAYCdtUdLx3Mo6GkL7I8R/2iFjJ6DqdSpV+HRooYe/KBpu8JhE8egQdoR7kG3ajZo
2FDD1ztMVURLNPTN+KiEVDuAJWtXc6LycM4RFOs6wfwCVIU9PgzcQf3Pu3qmjd7qi2qWcwxgSc3f
cBx0KYNmE9m93t1kopYTGrEJeXRRdc7nsWZShJgJ3j2p3F97Pwoz6hVcuiQp1BenIVXjyMc9vWtX
edJUav3Db0SRW9opJUeIBHK83ee2ZWdeDjzc0jmD+sS0II5SHY/51vVJDgUuFJrSjhklnfuB49uW
bbVbZwF93qIEdn8rq+1FBI4PN7iogQfTUsGBdnm3/+TWjbtxtOqEZPbaA5Fz3vYNhkDwSYutpRf9
fBTW4ByW0tnwJyzWMcWhiiXb+JjEkltx2Dbg/0s/alHAvwnKeNvh9q2d7C4HzLuiXNLbkNXH+GwP
bEy6CqThPceZ9+CvA6hTRaAisJbiBtvtSsznHUY9QkyDa/YsAlaFTQmWE03HKQk2we79eQDi5Ses
ccpqHRrOYXOGvnH/677CpMfT0W+jaEH/w2A+Tfd7ZX+Bi3I3/Cs54GpYg8SKklNUDTOW6j+mf8Me
1ANYMfCQhljb8YYO5KcVKmzMmO/eLe65ccIUzrL2/jeBDuGsDJr3IveYgp1JgKfxBANxv3Ny9Dni
zFMDtGE8mk+Uk6K5xN5p1jnLjOf9uDbY79Cl/+biZHrbFu55kd9BRPXTIbAOtxFQnbMFpz/CRL+U
s7/CBgGLH2f2sq9eJlJ3U8WIV1L/DSGuzjfVvbdQ27ICkHA7+GBW3ChnSJ+tHFp4iZBZIYoxjovo
fV0EwVZtLTHC+I4rttI2TqXoidhASPgxwi0XnrWjlJW6ubMdgEmsTVVOQUDuTqVS0BXryi8yBe9+
yTYV5dEeHrEOKU+uxUsZ5MLc0kqhbxMiAyzRgovOUvBWWVEaNy2TCt4MY1ueAlJ7Vp89MI7yRL9J
N/UFsTFc1nHnSMEwQ4mcmbSclTXAMeCJ5mitLvxhLjRDSJ0vokLKu0PgLTZLFIP1o7luZ5XYgTct
Jm3nq+YTtXMCzvS7JJTl8KpQvdKOP0ebe5+w3O7iynd6GmCP05sacItKHvmmOX4D6hMQOi1WvHTj
z1Zr7vht5PyG3s6GH6CJ5TRwurXsngNRUwE1kQMoENNECljbkXlFSPIBNHUS4Ghm51jqohvy6Stm
Ii0N9gjWrc3dS7P/a03I/SVKc2qMV0kdjXUVBbI++Pq9qMqNDc3lmVq7gPah92TZuEmGI3RRr+TP
VjuaAU/ovmhGRGYQIEJCWsEzqeZejgStXVqBtnwS28V92nEs4cnQG9svft3fthJmYawwrwUj9r4l
xE7Vz/iqLRbD3rzythLpx5StSi0M7J/1VJ+JeGtD/3qFeJOeSecGILlL7UxSxrsHB9RsswmtG3l7
Sf+8YmAJkmomMXmM3eJeUCpZHREFLcyGqlbIm7x8Me/PyTvxC3Xu7psIAwUCujPo/pLN4uMQBy9/
8P64MrcnZg5FvRceVmppgIBQY2cggRkJYoPyivvfXO2rYlR8/kseqgH1reC3AUMjGZvcWHqHKAjN
Rv2bmBS9ZFp0PBavnRsB53wTNm9DpXwoDB214QmfnmIfwuclLceffjODvxEqRQQTy4OH+QAUe0cD
k63E+KANpyObPcEYAW/E8k/2VY/ftUJMupwi1Bzn4UqtblqTtseIGX06MhpvmYuYkhCHH/nztDbe
7D7sDwB5jBH/Z3Q9UwP73vxyapFjsncT1dOHv8QAGFkLog59HpQ/3gFPBx+oe3+y+HiR/AGkFTNV
0lrRsqSQpzmaxKj80CvH8VCRsGehYirUZTZ1LqlHOoYox46B7Sbw06JQNzY+yzZvBjHZSjwt4ry8
2UXyecsg4JAu8rMoS961IJFsUpfBmIHKsAsyol512qdAc/OCBpZ9aRmXFiqmniyol9fLKRs3hFou
ULZyY9FKV26+omDmIAtocMrdTXBl8w12JMw6gYFhgccv9ueGkWSVlbHqd4sjRWphmHU3mOoYQt3E
6i/XOxzf4Vtno3pbixw3xXwlIQN2mDjcqgOtYf90biAvGGD+xjrstfyW5ebyMh5awYlgQNfG1u4Y
yXZgOYUNZAOufqONTk39I4zb1nNM2LcKl3MeDa7RcqEQ4DTTypuHSNRAHINABuWETOFIA0rOBPtB
QfI+bBUmBXSetLVKhm8ehHM6u6Gy7vuyCYlon8k3ovk1+iAxuqynomrOypep22MNPm19PicvHbIR
U5cnvStyy74vGtvIsRCAhOvz3Wi0ZxtIKWIljB8DU2OJ9r+tUHSR77jmmxx6UDOcCja9AiKfVY8d
FAp2hxkNHmrNKfPEKCG8rRej4ddI3+zHx/SoBlxgNIvJ2jSFrkmPy9zKkDbVs7putJ625gCxzYjP
b3dVVQ2K+yhp/1xj7e5a0cUhJrd/V0xJoW6zfleubd6/Jl3vi3DKg/Cs+69Vb8lzYRz+iek+MBDQ
yPpkcQQwAHHxACZ9IxZkBZJvyjtd8BB5YTqmEmhcqDJQogcZ3O7DJggv1LDH7yoZof1bdaXrdhqe
NYewRTymk4yvd70kHl3+RRMtYGK/TsY8EXJF67Ba5u92FidK3ieLkZac/zMKvvg+fn3t4CtJMlrj
1OuEHA/Dku+RrMKT7ht3c50mM/c48IUDtRc6qNf1v00crrTXrtkH7DzQJtzG+lBu8s3DN3YAEfHJ
vKaw6V2u75VVKwvcJGgVjtztiYdbQRPVyE7exqCZswwB/fOSWJ/H4FTTGbW4x7zLn8reFAcLS/cZ
zUmW2QPmHLrh9KQqGzkNtTmEdanRVkK9TgAaaUyjwUT4iB83imCXlbNFbE7b1TxwgsFP3ORtxHlC
lL69Jmr8cYejYl9sc9CzPktKmyYdbMInu04pJl6j2X4p4zX1llbe2ZkkeEXTS+pIcCviYe0WudIW
TlMY8vEb3Twk4yMgbXGMtsWr1wQWlpzjyP9GcHTw7UPiF/aPOXlYYi2FuCy3TSoF0qbw5TcmdIYl
DvA+zvP0ABFShhW3GCeJdAvft9HzrYZ8jSK5B8X+KUNWXnVzv2uT7I7ehVYIMso33WgbQ/L13B5f
yOLtmI3oQc7I3Yvja1vD3AxPVEHB+AwSUMfeqnE73Xu3ac/uVsO6eG+7WjiurpLLd2u85gL54P4o
ccN29poBq8jOTTwjbaSkB0w/X5ZuxKoVKi5rFaTkIx6Aq12eRg3gCxYTuN924RXRwVNu9qsIRhgP
atwa9xVVWWf28wSPKp9RDDigAsiZNhCHI7rD0Ps9YwqFwgGjO2/JTdNPzdmnIWDdSM0OjKMhFpSu
rwwjWb8TM/zWQ7DDjwElskW5KQl2Zvu9YK5nW85I+ZJp+ltN5ozCAbtu6V2mfTp4794fkT9ZdCH4
ILevq0ZD/sIEMwnHIyyT0qAszBW8POUW1BVQhTwBhtktsxzdVY2rNRNOSwK4uNSubxnEmb/iCy1k
f5FoEBwQdJB+DRWP8c1GXdRtIoJ1lgNXt7PpuB+Tnpe0GeGgtFxqmhhyEE3FKhdeyjOXmUIdOQLu
ukFze1l5iqah7fNS4m18yIK9ifR1ajMG9iLkF00ZJJ2aTbRuBUSDncnZfobuWqWAJ9oD7pL6W6pt
o5/Ul887m3mYPuYzHlreTZBq+azjTlMKQMkMulJljaBhh+IarFTVJ5/Xk4RALQRHTNiHXQJ+5ONC
Y0r5GyG6Ota9ezVDV3J7TzPlOf9iNOMEInN+WgFrIAM/sPL7ue696EBWJ7mXXJopwHjreadcKoqk
kpnf1Q3P8/EuYSUGnt1W5588G27NKIU7QYFKELB2f+r+R0dWegf4IRmNSxBl+0r/1DBapBRhWZEH
DOPUw/IEgPuLfpSobodhOOhERB94by626YuuZyCQolV6xg/29gsc/pilZMBuNryALNH12kStGAnX
dKRgLJSdJyOH0Fv17vDBgHilZHpKSG2z6+VSFYBvabDUXdIdXS505svijll/P7UkdRdPAFP3xO2B
pfpv5H6ZHJsKF8elh+d3kPgeHCc24SrTkQP/xPbdj9tqDVamx8yrH3hrevNC29iVCnl9jz6zU8o2
DrrcDbQCS+UAZFRJWP8wKNNTbfGRiNTidLhP3ZEloe3O/McByBgcWY+GDcymCYYe4RVYfFDV/spc
aWd6NudxPdRnMTkGHNd8bA6mWtlVH07LCybjfXXXwgDpblnr5LnV0Jj6UdkIBXyTKodpVRIV4wE1
kojJsWXLFdMro9ecg8ljiqTlMQhnFXHRBkAo7Ek1m9LIcambzC+nsVkNuoWQzlZRS1Y9jm9UFINf
zyg/BRF32K0eN13hrLkJU9gGw8x89h/DeS9PszcUjoy5Bd0fMGeWjjdArn8ehKEemh4md1E4IjYy
gOs5YCV6o+5CbJI5m+qvYRHN4ClFOI4jN5BzQvK56fX5ksSGYkp8fh4cbMYEThalqbbygOTUeXzC
dIBx9iTbo+Gt2jh2xGXHubMfPlSCar1lXF/ka6a3Qd0PEDttCRUYSjOGbSmaYgsam9GGQ/Y7Farj
Lvj/gFXVpDEA/0UzTNDIZhh8cIRj4OxizQ0V+I5lpUbkq16MCpXDU5AHhTMkCiXwEZh6kaqpfZC5
m6oNGbrLidJtYz5B92cvlbN6ANR/KxPqC5ZOoykeiK3PsQvVQNe1DQsHhBtiOb5aI1SiXosc1WXD
diT3ZBplahSwbR+UtO+kS/+z7vZII8lF5N/hw8nJbo+mtAGe6moIAjXVWcQRYujFhN0Jm7/qcYV0
kGme+sT3btQQe6Gm64f+8ieYh1h3BGvGHFpzHiBW1A8ow/PX/bc3XlPtJj0mGvyt1Vl9RgkIOP9b
7x6QmQ62VgdtPeRW/0+KsPk7YvVke0slOLAawIZlQcMhR3Ugf6pv0QUmWXU2zH9jV2SVv7VosesD
sUQa4kIeNubQp/VkXKNIHcuzWVxTCUQr+/a/Xyrlc73seHKGIw7aso2h+kYrU5FIDDvu1bn4TIW9
lK95GWlgYE5uKdYm91+H1iLFVdYIqe0UYC2Qa1yrHkZij0X2zlnFfrZODH5iCin7g2QnktRyqSZN
DmzeIn2011F3BcRJ0Mtr8PBdOTgkPDQH/Nu3YvOYZoCdL9Y+GgnAtGNiw+BZPPCUV2d8ucInfIfh
5ZqNG17gapFySGuuY4K3m8zJMZhc4fZ7aFhKBlyaykZrbRxQO0s3DnZb4UiBKzOZaOhqCtL0JdK8
CjeQzfQIt30E6ds7nKfIYY354ydo/GOPYoQTIIga9g7RY5DV4nnLGm5MB+DmHoeDamPG0D7mLgsa
euhKKD5ph8Y8tRPICX2Z9EqSpFS06UWF7zGOW2uSJuDqIUkPrj5qMOS7uSw9puMvFT6kYle9umKA
JrR97mUJoZQzBikF3drMRYLHeE0E91C3BFVvHw5nPId88nTH7alOyTh00SKpU52QmXD6mGuMQGkH
6nuz/OXLEbLpa9FbjLfm5xOI6NNYp14r30FeqeU0gzy2xwYZnrp9bgjZ6Gkzeouyj6gn6kHhpmCa
4sjVMO3uyLNUiJuoOoEklDfwfelMw3592m14d3N8BXknHxhGGkYEVoExyhO6pLXNkYf4koDuV3KX
osNwx4KTaGPX4a36+6cB/f6BkhyDcUD+y6p1sj+oVRNiG6lPqGZomPSTsQuJ9FXvaPXXSY3+GwaS
49nWU3oW4oy6GyXkxAXIHuThZEFsou/cpjPfqR/mfZKaAD/QD+54ofExnVHFAmcQtk4a3BPaVF3m
tbIXFcO+2CLsO5A1fbOXFO50fLwaTzZ+L5wQ7lk2yGIrzITorr+c2xQqyiG1g76GhrypEb7yh03W
+7ZHs+2DhebbszA4HnuKlrWLwXtKl1l2eM1m97VAQutLEwWgKvqGxnX52HunokTzMPheO6NUPbak
tixj5q0joeLRpNHMYmZ7ytSfCm/Vt+6RsEup3LiPknAnJtoDK73gd0f924OpPeky78UuuD2vagsn
mfX9vsrwv8sjC7VzNTi3E1JMLmnrSp81l4KzVK2utk0BKuPXx/Ub3o4mUXQA31ETCTX7giUBTOk9
mfsuScfvqDnLut1s7wuoG9LYtL3cSAejUiQmUbYEd1hj7nTkOPafZkmdGUL69Aw9n5lzGewXMMgh
aIUMZtTMDqsnOQNQm+yTxxfU8HaMNGfYpySu0gd97j9E7rwbnmytrUXR2nNpEafscyrYyym4BxYu
XeQT81Yazj2Z5oIk4zjWR2vQwXGU1tOxUg/Eet4I+ImxQ4lhBk5LSAgjVQY51MbZNjn6J/LiGpD6
2NlNQ5k4CTKuBK8zNmecokpCYTKmG99G05evR8q1USQeQSxGqMpvHiVgjAu+nucMwMtL7tjKJpCU
EygUdwb64qx3e6MbNhjdPNd6WbNysSe02rWf0qLx+Lmqqe+2JLCU/lrVzQrlGx4VYOKZZZuII6Ct
cWTreVD4thXjf1CdfGEhQFk3gbXNknkVfj78PKbkWQRd8e7aWiSZAJ7AYCqCCe+sTtMB6WVz2YQD
wbQLtwHe4hM7Ep/wKCcqaglf35bg0fhqapnxDpicq/zDAJKYkn23UrSu4KBsWIXgxzUGY50KEpGP
ycSktJwNVH48OafCadS3iweShI0DPTPJISnKLhe80f46cIW18UHADy8+zHelK2nONscz5j45KZMU
+NRXaKGvNDyULhdMMyUOINytqZK5CLA+8SAbiVSl6LlrVcR2xDE3kbn78kp35/YaouJeKSEnj3Af
xTc+oVF7x0bUgrHsjDEoIvxxYrijyMOjR1aKLDNL/tT7m0EmWIZtmzqEJBH86A7OQmqSsjXV1Y4C
xaEvHOj7rrTbZmTCi0RLBb+al4Sfdr5Eh2oq9rZrSZMpYpgNKpJCOE+8gnWP14t44HKkD6NSKLES
i7XCDvmEUHVkyJ7EZMIKvXnSatil9/OO9NdjQDWh9U+C3yjYjphrl5vxB3pBjDsv96gQk7cqlexR
NpUzcFeygM5r/7jpRjQyzPrC18jSydwSDr/Hs06LsjMYXU1SSvQm34fEbxQLo40WbpBt8qO/cHjz
goCQyqkLBgPCoGSjkjcW9YH/t84J/tsifhJoVpR4jQpEGI7ANoEiiTUg8tCIwHTrSKTzu4REztJl
NLby4ld76W6HbZ0WOvJweT+TQA+EmT04o7OJ6PtiFvz9pg+zvm9FP+r3KdzDHCw5/bEaKb95cvPC
8eM71iO5JWx/lV6XTisgBrxDIi5pJlpENPGcTeyfq5+UtoIDOVWhs4TA68bfG6Z2AYv5TdXN4/Hw
XmBy+fpiPNf1TGA9ufAniTMp2lfhUrnu36wI6aOc9Dn55fFGBcYOtxgYkHixANesqV/rRf1n2WKS
/ngpbat9RAaL6I+vrp3b+shtW8GDbIidJ7TJHTd+tsFwOEGZGWEELt+Hsr+EDUAhBeORljAV31Vq
rChEUHeHRaUdGAnCqtsvXtoaY4kR3YwyTShzLpkJv1gYXuWPeNUEbLu1u8afz8IaWISUxe+JKciO
Bwx1cmkPiMj2gC3XZs9R/OILhkHIWB8tcq7UuBqATVW6WTmifZPP6IA5zzTDPd29FAqbU6oFpkU8
pbndNbp9D5X/YQJESZ5uNL1KJo8wCq8ezSpyr/U1WhsOKv4jVLifCs21IOl+bc+si9Pdwg2bCI96
0Yi5HGigzMF4rROpgSPJ29Z9AMpqbk2XNe2YntgdQUOWr3IRx37pcp0NRYoj/KuxeaCo97CAVEI5
1obzP988ywbnoN1ffvTMZFpqQ0EsvUwTaFQoc8idf16pmi8OnZrCR/ifmD8WANlrB8/dCsEY+f7k
JVjOquHSILwFHRY9nwnPg9yUAR6eLGQBwnGjUxREJGbUF4UTQ5XyQaxzpL03cu2MRuqIHLTz7roF
ctYxJp7CwN2g1MUx+vf+RRqMyw/KCgo/Os4LQ37/ksggeb1UyArn8fPWd4GRU6o47Neb7dgCm48L
xBcQj7xGjfDBEkZ+cgx/orWD8YLZIkyrlrspJ8TxuUsu3l1LuH5pUwvDlaKR7RQeEHAE9g05PcYW
PnOeVoDkPVH3yx8r1YvUj41TJCAmeBL/5TMjuR4YGk+d8ovCrajqdU7VS4dN9OJfUToq1mLQwSZe
N8LJxNxyfNx5gQoye2s43gsRiyqMmgIZ7p1PBS0j+IUorJCv2PkLsv0PySiwfyPMcNH7mIq47rOx
9E4V57tUHqFbBijmr/C4spGyKXONeLF9RmUfrzkYhnxdeq/MrT6DLPVFH5Rs7676eiG0Z9Y8FFuh
74bGAhlQP9QB4t4MNEkVKqq03VdHArSm/LG2Ur+3jdPrYoGwX2ih+jGfzaHctOgFOD5YhEmJ+cRZ
fX70Ky/rxGMcX8zBCi61RDBEcTfgE90nGxzWtfllfwrG8Sv4AXn1RSAI4p1AF7IdZ/m7tjKLebNe
I3Q3WbTBMrHFTH8P/3mNeErByU1KmCXP7UhoUG7D74gySZdhPtPk6L10YXDzW6ykzJUdS7dEQwN0
S2O6LBdiZL1vfuJOrK0e1WlFG4gA9KXFMpHIJgbw+SUnapgGjj086EeMpsZu1vOtUGTbmxrfzvlo
Y+0VIP4tG2EQ3LE3hPHXbfQTlKLBTi2Lb6Ghue8y8W9QOuf4VO5vLkWKxhIuEpPE0+S0svKYpbY5
ayZspXt9PTvrodLlmi5vPAYimTOppBqBajACCaMiK+u4qVg1cxqmQfIpkzgS8ZkwGFgKI1iuW5dz
zjxZeD/hxWLL+ezdHAEzhk3bg6J0olrj2+kS4BwtMgUcDMdd86xn8Ibd2EcMCQk3/UKAYqj2zxWB
dlAcCBt6OCagboJ479CLOOM0GYigT46FlaOUBawbQ91VZpRwKNUOQ6QQCwQRIHowmlpKUTmpiLga
K/4b1SnqnRdn+N14qJ6775RFpUIYnFBI1LWIImaOnrVyv0NphudEMn6I0DWIBb0UZwdFME74oSQ3
1xQQzps5AMbva64//4rRGoyNSAgkVqTP9jYsNlcycYQ1wNtZvycFT2DQh0qyeq9CSj8Ckz6FjyTq
q9cF7y5t1N5FAOMyuR2P+SFbKo285eb8/G6HWwfJBsRIgjwa21lS3DPWvq3OD60O/6SM9OAVP9Z3
Mb03HaNlGLBdVYgMefYa7aPrqs1s6zI/8UBm2jB8tZHxxumE+rrj1SVIdZ6rOucd903XYorxNT38
RQ3SvdrssDriifziwcZ4btCt6+U+2VriXHo6ff6OZ1k96OXc0dYHxrRhkuEM8BYPS+H0tcmHSSPk
mazDTF3k2azjiKPUN6673YHKIVnj9cHDvb+R8MFLz0RxHwy8fJIN9nvnIxSCBF5frvJ8UjcZxc1n
QZuKX3JLyCjUq4TqLniag9MCtIws0UjlU6eJ8prHJnvyMneWtyod1R1A1+VO6FbS+/jfgM5+qif8
v1pDZH2F7iEBDUolfTCrolauhYQ0FGYRZRe7Xs2OO7rAE5PaFvD+jRWjeYA+zvVLGVIt0zOLba2n
s5X51E17yVVfgLHuHHp1ujocGomtyLc7iw3uptH2mcr9pYiQ036+OP2MVVVHPdQlRl2vU6t3uhT7
j4PVJEyDYQlRZ/zVsGkHeCkeCO1d+g/tMrYt5/JPZaa7VORA4ofbVqCxoIRmF2rgly6akoJst2gh
s7B06GL3kV28nhr1nzmFVyGCImtcjXT3iKRES30HkaYOX+6s/2J7l3sGXMYFe4JIxnqX0vUvCnU6
NJOV1dQ6DqVsnb9OwJd5aL5Vrxlhgyrq2bDUAmrYA1tPCVI/7pUTlenTM+DYersHNora/wwFWGmr
qUwq39k5rLWrJ3VII6VmnSNDVzL4Vu7vm9Ic5CWvidxP8czzqInMQMrdXnVKU3g9RTeQEfbOj0MW
yKhY+JLirx8uCr1fswakLxXie9NSYayMDZzKDtQvuqydz0uV1CeTv8rngQvpxwV+I9W2vk5mfQ4g
rdgpzh9acI56ch67sACh+g1w28Nm/+91GWgl/VktqsIzp5e5wW4VGKxbB198gm8GmPX/fXN4CXGG
6BvH6Vz8zWMLY8XwbqA5+hBmCs1HulRPI99gN55u+j5QdNW44iBcV6eIIswNBqYadPuOIOh98/Vp
4LSWTNDB7vqLrlG6wz962NBpT+p06OlRRAlz5n/X8mLJtfbeq3PY7RURVjsVL9iadjMoGa9IwYMi
z9d7Wo547RrDdXJx185Kq6N8BUeeoRujMD3lY9V/D91gaNobNnrXtv9oNrJMSHnaUUcoawQ0bT21
t9ztjX6KCmKV1PcSuR1bC4PIqgtubUdrNB0vH4WyQbsHoPePu0mR2obGES4HDs6xeiQl1OB0hIXG
4BfUYgj5wjSEYl9c0jLBExKvDSe/R9F6SWYdAZyMxdobApqMUuL9CXOBgWKlJA3hYRHO2SM5VZ9s
gNcWZ7cjqDpgAjohhSkTWfGMaUvGfV9aGLw871gZ/qsFkFMkFJhzE6sBOJvhR5IHK5HvG4CT5CtP
D8cX/EhMy1GBuz/KE8zj1X7AnWUdxJEI8BN5YqwPg8ULBA+xC/qeUY/wmVevnS4PJOB6Q//1v+H+
VIRN6se4pPA2LLwBmneWNDVMxj0zYMJBaLQMGi9g6z1fMZ8tejbtvADOOh3iGZJNqIHjNX3pWloB
w9cziGg7vnCnNCcV/pOuzBzwmFWxgafP6SpFKdT7TX7si4iDU8k1uSCM+K9HDQ6pM40h/wufrrcd
21XAPnv48cHSPqiNBPMDvYd2KLqRG0WlNivLZR7OwHroRwKsn7ERQkw2rnKuTf+buqS/pT+0a4+p
T1/YTq/G1LFVyzBMlEL+5XmkEkls7cpgXhTG6XFrZZD2Fw/N19qeUTBFt/6yMe/AkOto+yTVflia
mYAf6FOheOc71Nx7jg0ZcJHn9Hbo4ZZEavTWao6oq61SGgMkKCxkom9JtW7W3yzMHzHMA+EpXplT
sgmL1clMivpdaZjOi30PqPufyLHB2XbVAXoFNe9mMK0eki6sG15EDUxO581tbB3tZgij0e74zYqD
1juUvY4fuf+wvwvu4P5oEPodb+9EV6Li4XzzNhvRpR78u1+Qz6AY1RIdpdqlLYXCEhIlhspXTtap
MApMBDwhyfrAuUVOytnrGR9M7f0Xa4opfMXzBvl4yZKs9sNaMrGlv0Vw4k4dKTjQn7UdxR9Ke7fJ
YsthDFF9XnL6JOzpY6k0FWF05AxSExnVdqN85zAsJ51vdqp9HtQpZMhMc4kf2bDcds3xjHg9cSlg
1jYbt0qxq8kqS/bt4cnM4ZCwDy3avztuMQ1ad1ANTFDIHLO++BUHsjeQB+nvQVaVLYLbCx53dsps
KTUvMKR4ougRdUyZj8dC1JFrgoDsh0G9heBEnxjy1B/R8Ihh2eoPrGYGevon2cx128gITHDefA5M
J1c3TMKdbUtyI+ajkTcsZxpeG2Rx1dOqBCux6sAmcn/JkNb1VVhdtMUCtUDuj4qNvOAFACd5De2+
mgbut3UEzdK3lBGa3dHqmDsDpPmqI/2PLuYiGKO5wvOrpjC5xroSiy/3HzuwRS2SF0EM64+iaemx
e5gNAfG7DfuhuOML58eeVELX3LpmVouNAYtSeVbTfS0BTRDnOr9No4b/c7P6lsNW1YOHFkx8okKO
RuBR5pjtFa2gc01bQbDh27AB8e1HdP0uyTuswNV0ggQP1+4/rjrWExvgSY75RF2BBhzQ9xeelqAH
yFv4Yz/r+5LelV8C793008xL9PonFVHaWZOHNhh2vSZAtsfDTW4bH0znAxpOyp8BUYgoPFr00Wlf
68ty/UTx0Qq1XxYyBYOF50T2RY9j2OZuoxt5MSzxG7ZqkJtt9V1r/cVL1egE13ekDIopya4/9BCU
9DfQTheMIyyM+ViQHrI19OfwD8zPwOElc4M+f0F7ZBPttU4ZTiWrKq1CGmRI0f22ZissikLCp6A1
Bs9rcYPqF55MS3JcqsS7xAKx+2L3qehqh5zbQznylg0zr2W2zX4/CHUNHSNrN47leSaFIQth6UVP
zIt4pB9eJmAErbTikNrNDFaMF1KyjSzv3bGAUWRp4aUUEZ5E/HJ1Jw60mbEXmAVPcVw7pnm3QhtA
P876v4IxavWxngv0fOdqCKAwiX/LE3eHSyiYZL9KWH9YUivuI2Nx6TAgFNw8cfh7M5i7hqOGWJqG
6oIjJPNOdD+gCgI03pGT7KlxDZk2DxXEakHGwhlAwy9Pml9z2aGK+xCD8c8je/9tZYpV3F6YPYsM
aqjSWJ6wOLJ3GNZjyFTrquAhjPkjJEr6JgHY0O8/eL6pglWgXelsxK0t6nuiiu/hUDiyenBvvAG0
deOnM5gb+4GYnOuiuaRTer03Y0cTNuGAUeT9mpp+QP77AqbkRVIn30m2AiuBYZee2AXuyHmkAFnn
I434xAGTCIK6JpDg72GJHiXPTwdKf1P1x4zKe6mDXmL8BqjobnFUtnBdGm9ul5QKz4StSW+mNxyC
mgB54kQJo+nrZO7tvg+88bAabBf1f/w2wYGj77Cb4Cod6mSnnqly91cWeIzffkQI74JsTJKvxZKI
xs4WGSAtICvwv5Fp7aD5dzFX8uz6rectvvDhU1IgoFaKRB0vU47M+zsrfeCzSgqF1PADq9cAue4E
YqsWfO853W8H37M7Rcu+g/vIindGTqB+Jta3vBLklONJD7JhhnbpD1bzGpLD5oF+pecE+we4A2Gl
H7Jb2S+0v4r/IKwKZ+bzRVHi+Ko0pcXz+oOjnwM9Y5zzB0waAkYnwNZWwbE7pO6d+o5COT41WiA6
sARyU+d9hCeYkOK71gZbzBbqHkA4apsrkjm0FmFfYDbbPlq73ZvkUQuDzGA/sF2R3erMgXT56GK2
iTtWtKkREgaXjTkqCzIT0Ygn7o8338wbVhbD4522gSuuyAKubw4VWFjfOz/tQ8I+1MRSoHA2HeQZ
ehE70R9eYOET67aBv4aNN9uulhYlEPb8yGnESCRrSibpPxZ/E1w5pvZlAG400a6CApl9ZTvd0oJI
BSClI4Fq3FLLCFyDtZmznwla1nN53Ookt2R2/HsbFzJI5GqOMw/FSJGUSlhQHfYg6HUTK7EobHw5
c25ysn1szr/tURXBgI5xAGF2IOF6cN8mG6vTxbTP0fe04XGoA0Xsn6lAHb/PmoTh37dqsl23Be06
Qq/52GsCPCgdiAtOUxn//rMQBAZiZykwaIaChy+Ha734TxHwKvOPyuI+Jfs1LmN9+kdWCWiA0Rwy
PHlmvhMsr6UBVKrEGRwNjTn4s12wgylPJ6CltM/ZLIk4Sywl7Y8XCZKMwEzCtf0ieejdJbbZIt9+
5Ao2fGmE9Oiqk+DLfHbAFLReEMvwbM01PwknWwEjxxjGmtd3gyapcwA9dSKY9/gAZrTGohLg6fVf
z6g7QAl3HeI1ErLGs3bVyBQ0oknuaaqbj99FFwr7UqtdvKmS929eCd1Cu4Es/HV/uUiNtFvcHBIY
L09ooD76ohHH9fmTuEX5w7K6rAhjLNhNgwNmv5cSVmyjifDZdHN1Yw2RkBflce3/HDm/jyYt0Bw4
L/jRzWGS0BnuWR0XrZXjV8L+WbpcWzwFGPrI5c8M/JqGBFf8BkDEHrQv91O49bY9rgO8dD0DZsB0
cCoa8fjJ/TVbvwyikUjbfigSZDk4KbXSKuuB7q/3e8Yikp8UFpwQ2j9pQASgODa99XXwxJH/8Tou
+6L8gi5AcSlto4wotpAD5jx4ubYAP83ZBsFdCV9A8BW40ojhTDKskJKCRmtqUPkZao5WRTh3C9lE
ryWvWn+ynPIhAsO+Av1y6BZEqtKbObInRLuBCjWZ2NLo9FVhW1lpfBunaju7yUgtxTom2DjTpmTj
qw+vjv1vLHdKJPxVzfZxSl4h0CJzkhnbqhPykyG0gmXTDbRwOaIaMtY2AANB5N3isgno0jI9ttXa
RkJhkJS3xsxbJSL5a/xYuLv1i/lxDFbOoAl/bj4/pHYkP0YnKscsiMzK1o7wwwgz89ZuGlm5jUYG
HzsEYiyjhwt35sMtHLKWjR/zOsXTByGWLYMs/pyoJQRMlPjScJ8pUZ0FB4gF0prR6XN79QOPQ3DZ
5uQE2XTpYQhxjmsatmkoliMlbzER/hQcRPtdf3gcOaTlWK+avuiQ6xRBTopkt4hpGzEjAa51jWSD
uiYnG8WMHkm5gc0EMkOdBfiQII06W4seCxuZ+oTfmZHYD4Ucl3uNdHDU3evl5P/BQ94dmAJHN7GK
PS4WOMgwE85VWZ8oDr8m0Bufk/DUkT2IZn/fDJwEtoPs2iHh2k0eM56pigxcaJKJPz1Gf+vz7FGj
pxFzFFlaTF+NXTV3RDFxcZgOsru8KflH9f8nSrOtdy6me+5izO+hBfM7TH2HyRkngX0kGvkPMgMx
IEsanw4OqKDT0Ti8N/pOAXQbRrBWKDhtiZkkp5/JQy6xW5BSnTqVqPaNXkUTyzQpDso178azXzXG
HXuvzjJv9SpAVdcmqnUWRPWowEpJoAeUnH6bhDL/o66GU6UOGrbtHcigeO3OSdazg9/9xwHOvBbm
O8UG/Vo73Skw+r56vI7lOiHMtpvJ1pJYo+hZXvMhu7u4Ol9yVEcX4RjtkHqL2Kt5DsmpWcZTwtxG
KaF1/7B0F87kBKf5lekOB7hXMhSnhkkI1e1zytnCm8JThSj6ss9NF3BtURTGWbWvTv0VmnPno71q
tkiV+W8R/72xTWmBYNkq6JKK8SqpcIVwVmi8W92yr5lTYpwo5by3JlL6bydNjmwQiLX6VpQJXdVo
Whwo00SeozRANqNd3u28x/OSQYTONvyP8oXpt5rTIG9XgYXnrACnUau8BPkc6n6qxato9FgfhcMo
EyDVhxgpy2SW9Zr7D03lT+LfkIzGj7pyOX1wlKMu6ElmDEcAemPWoQ0OOeM5I89pJtGvyhUyh2bz
30jV9rI7m2GkT3s6bYfdYHwFQTdGeQDJBjvv4bmUY16KGAnV7y55bdarJwif8zmOBdmonodCqdI7
n9p2yDyqBsFupsQs609skZypJNuivzx4/I/irmEdA340B32PwQqbdm59JZxu/SPmdq7S7fxZziqU
0nySZnLdyQKKhSG/96kQBjd+enAx3bZfBbwR4lWLDu9VUFl2cLkfAKhoNppLf7UQunsuQOIfy7vO
vJunnBMA/3hCvfbC8xJ0hpA0GNugyWDoCXugFhGqlePRa/VSIGl3xg4Fupv4C8ehQ89kV77mPbmZ
062lOudB5ZIjowifBF6jAOGKXDhbk6j5iw9sluuxz55VPGWzQ0tvpBRU/FLM1E48dK1Gp1VAuXqZ
F3GB9w4lo6woZhbVaOaU53Si6mfFTi5gNB5UFuSq3RU84HG+e6JbX0LM7vKDKYi3P0pY56imm6zl
2LcUD4lC2BCzBv+jPx6Hxd6VjwfhLTXKwpIN9QhYS2aycyzoefDRBe4dZnw/57w9suETZ3YHJVec
QFiDJ1OImSHDCUVoFN4MHH7ehjWhg3Ilbadg5aq/2A9QTYVolGRu9y7eZHibHteXR0BlvOP3Ead0
abCbDcA8JDBI7YR5pngDVewnIabO5jHg9FPa6TTMX8oTX82AB5+ifJ832JUaQINyM5HIQ8T1f308
pC5htjRKt5PW561nlfWlqlan48t/89rsqTx5c60SeY9Lc6Ml/AOqiIuTYSRG/AHpeDN2vlACTPAs
HLXBVw8M5TMIA+Idrm2C1IIA5flFU56yfe87gQ+snVlSLHP92oUMJTKOiIBvXmSlH+nuIorUDhJE
VFsbQsMlpqTSFqf47PnY+5LmRdfYkjWDbb0Ort+5Wq0QHALYAma/T0UJ2tBQvgNzfij8BZ4gOW1B
5vwweGkpIuVNernjLThAkIVYMPZ/qteOlGH/xSnYWrScs1GC720H60FYDpSfIiWriZql/+yn+/6U
NmXt3lOytP2VZ7DUivaZU2x2lem3Qr7vHmUWj6hH8eoEG19maJK08s2Jq/g6XxWXVLCs1ygc+Ojs
FdAqvwJkwoOA8AVDkeBNy+zKYCw6gNcYkO+LWjofVy6BkpYXJ4JsVLeIqAjd60nEVNBJF06pNfaR
zxgL6a9rW0ZeVStrne7K1PrmRAaBqCY2RQWcSbRmQ4VhfDZEPmK8mbYTCWLidgpP0Hkl83eGqaUO
jSAq7oiKmZ5Mqd59txMCiYi/oD97A1aqro24BWrN7e1v1dCfOCQBOPvherx2dmvcvR2R4roCQA6O
e5OLKfcTSyZaEviJpxVmKu7Vyhd+Q2RnZxlXigqw11VQDQkIePunLK+UZ1ihny+pUMo8LDl1tFe3
/CGo0UCHDsgz/S4v3Yn+3vEZDMN9jSCNUKzKLBBdeF09JU26q2rtpdNS3z1+lOjuI1Jt27UAWD6a
8ASJf82K2+AKvrrppch6HUS5ccJWWuLCpnqjWd5wTax0a790Gqbu3qiJ6x/JwnHGXzBWX3Man/hS
C65Bt0Eks9gUPXMgvEQR9whQUWcdwqM5CD+oLKvMHSQvUA9HOSaJM1CcKt7288UhYKTX9oIS0TlN
M9CPHVrSKLV3h13mHzLdesGQnx4ryXWSwHrdy6+y1A4bcKn6CjE0LOFlzW2Vy2/CD6IHCei5TP/e
/QuheUYYHKmQPLCQ3g/HxMA1kKPQt9J8f+lKtcERrN4qWuJViULWOVWKtF5+DE22prbKrLOoH93/
t9qmE3lh1WGO/Ah6x4v86YM6QNPOGldlgmhViXY3PcTbfQeG27kkbe64oI0rHqh7dGfES/Z2QsPV
BZOEGR/FLPpB0SY5WvCuuvTwRTxqEwnvg+jyP5Vcy6XZGo+d2L7j/aMOmiA4nYhQ6yum94pHvV+I
LdwSePM1WJefVTv9szYGq5UXbn1fi3nVwBJVGWRAc2MHA5V6M5LwjQF6Tsshyqy6/34KtQVmmw7B
IOPtgpw0pAcaIwtN7lYnKn1faFExxNcLoYiQLwdZVl4KJ4OFv3WDbH2CTGvLRGe2ChHrClEsCVST
NYf22arqY+KyNLn2OOKGBD/MWk6dnBWdK29zK87xnI9fufilT4ZIo0uxZRvLUrTXZ4rBGPOymj4Y
UqA44KA6bsMlvnuRCBeqRsxDV++slHdWsSd9L8KoiZ29l5WxuJOpw4mLB/+9BM1GvHgNUARlsZud
Q83uJvTRxgQ5WCuyiHQ8jL9MDoLqCjjnfv8Md+iz7wnnvWMAdYQqrxUYJSHDwrbPm83GMMeUUw/l
zYJ+KUzbnkCdz5d4QpyH7HOpT9Bf4E3sHqQqmNoPtaAqsT5RB1KdCZRIYrdC0OqF5JuveV12itYJ
8AoF4Usa/hu9H4/adPgoJBeak9cIiD5ELdPhF973r8Dti8g7/N8dFyULfD7X4yXKDblEP8DziHtt
D19pLWaCrxlIq0cbahSkpJwPJCVYYGYmt3j1gH1qtbHGVvaz7en0yWU1F9gUH6V8ohsvRZNdG0qR
OV73+roCLMptoC5V00hORdbsnXvWP1t+4FhELd7vgs6dV/zmxNXZH19uhQObOsACsePZyyiZIuDG
/GQ4HGVrNZhDWYvI8q5yl2FZ64uRqGbAK1fc1QKaH94Q6ao0HnDT02lQTXCiEcookl7qZmpUMfQv
s9htTJSyKhzmq9yp4gfIsicBwLX/R4AgBxladcB/L3VPNi3BPqoLNeyIIo6mDmZRm4vVLVZVBkDY
nGTnCIapWW0ylGZF3kcJjGio8FN05CBVPs9/y5netXHov2lB8sA+zuwsruJ6MwZrxsVMIgl4qjBM
Z90PxO97CuGBQz/2ivk8CWNJajyrNWd+1eb8vnscRmFQhnADWYdMXh8JTcv5sBHTfdER6TIKkI70
m58F0aL4dyQXFk5XvE8nODKdBaAvL7D5yWOJ7+wBf8JEJcJ9OsyuSEURIRD2/mtIhAFvym7+b+A0
I2sAgR0yF3L9nx4WLW1yLUjaN2zrpEnpinHz/Vz6/ci8JFOd39mZasA7d+Vaqa27JbBHiXgkemiO
HjUITnLoIAyQEGMx9WTCz6xmyrT+GozMfgvpb3VUbfedIfff7+JFqYpaCMep/Y4BNxtZwT0XsaNd
/9oPerdfe6Unbr0zXefuTHIR7TMSBLc52xn+6kV/NXRFKQC0vTgpP6Zpq3kEA53GDvPlakOpK21y
E95d19Sb9FyGfFLU9JVHoO9IQiA51NSQkJm4/ZjP0A/LNpQSl5Lk3EK/2YCyR2J809DDbhxahwbt
v+663+yMsxLSJfLr5F2xwpLVZw46vSx4QfXnXYUx2Ms/IVcWsf/AeSIUoMe/h6TgRYVtH+r5qPiQ
T0T9BFvNeDdcbURTctYfXvT5CHjoBGkXN1N3I3Y9AjLxjEpqq3Yw3g4uDtdXpgGGNOdpgbceDyPL
6s5NC9d4xzK/Gxf9LufhedUugBYK1P4J2J6VDavfYfImpsV5s2IyjEHT72MLuLxH6s4O8f1wtkhE
jfuv8YzI/G3TyLXZ8y4fe0+eCtB9X4N0pNAn2M/aELVzQVIsay8CYzMiPlfBYu2XLTqet21CxdhB
+/KtPMSU5W1Tyw5/5KJV5dF+dvbd1nxHO7R3x2VnkwipShJEncRabheURVZ87Pzui+C2barJo7fE
X1Z6xibSFWf1kfL8Y6Ww3uQ75sBPwxvgxzk3Q1y61UvcMWoZpsSMDZJw1C9rcCiiGBrqV9DTRz1h
ynMQxTLBgynkjde1z5vsDtr5XZtGoDzfeqb0tXAUyA2i8AB2A87a/v29oY+ipfJjVR7QB0PuYSPt
KA+io3Pu8OnGLbTz6dEYHe9xoP13cq25xlGaG/IpI7HJ3k1G0PCj9tyNme3HyvUHq0d3178sdaFc
JUljip/wmcGUzvc4VcIfGKaVSGO5vQ4IXMtWzvGRD2QOL6vzG1qUnGUjJYOdbcWszAxDUvQC/gqi
TYr05iTwKRJOT3PT6JkLw5TBdzbGFfdqUSVgqbRtXd8af27kew+jDx0ViQCltU1gDyt7Fo5CV9AW
ttc0WORE/YhR2xFBVzSCYWp87M5JjMs0a5hUIMlZ12jIKMLgjH5piGI0+4dLTGhuX582MI+W6Zkm
qT5ceKoktmIbjrjS/G7RGenZPaIeuqV0xyNAchMuKvLTkttKBmZVxnf7V+gWE4D1lo/b0WN/quW+
sc8wvSn5FuvQRtMCbn+z01XrDWChEGnCwTQHGOKWatP9KJf7mwMEwk+5ksRYarxVdg6ZO94qkPYC
jccwWSt9kyIdpafshpSY9yDOx7r+0qPlcEAv2EEhWHm7DPOfz+I5QJOd7k27w2rqOTJHNFm64xlR
0IFpVZEUBjjOOhIWjbLRWM/fAxqVx7w5aK3BiTeMQYJNGdvZJMwSjWo++RDWPERqOt7pvT4A9fAP
MNmjLSTDTrOgRr3neex74nVrR7Zl+yq0uhB+jCEymi598GxklLm1qg6KAljLh7tZ/fSH/elgMVRV
2HVtaFSqqDq0bdXoEGp4ZcfWsK8v53pa+fFvTIR4s4G4ZVKKMAlbSi21pShJ1KI4/n/NNeIvQWIL
qP366LV8zAFZWnYmSygPwGnyqBwbOh72jH8E/TD/KEg+zLM/P9oE//pXVsTLxN2KDNrHBmTLgrH/
XIdjfT0E8XGb0WJljer8YTFjgGRJPLwKsHtzP3wGO7mezojsaiFueBbTjZFYHcAiP1bGhbbCbG99
onr7Wg4ai7ZaJnAt6/FjGlG8AQ4sr/KK5+KFF4j3VzFm/3NF4xuBkECDT9qHwREPIggxG4HiOSan
bJbrNn2KjfQqtrNbb3Km6A+wrovk23NyYgQ8fMg8HfB8DE8uRe8spJXh8lNMIxXOH188bhRB/XWe
nDK8pjmSsBkyqumj1xoeQSI7kf/q7xCKc/UcyfsC1VEH0eDt6viBAsQ7FOr8wpaZHN0qk5qqnlfU
5Q3jYo455bIvMC2WagJNAEqaZ2RwO9Pf30dagU7RaotUr3wT46tFLnIAMxsLw53HLxT+PBXs7dL3
VTD1kyGXVdZ+s8IH2NuLaDmutT0Bh4XU+An63tLXcSzfRzb6aNkW3/v7LQojMUivvj8ue1n9mSXJ
DBjh3lVpWq8Hi3oAmRqx2hX8agT3G0yMSnfr8YqfCFP5oDJZ3zQFfRyVvZ8K4d5MwwtqVVdo8iN7
YKI12TR5ltIgIhF+LRtPmqdUGIGXPx7uqHYEz7kKvMPDzQKTRaYC3cpMkzRS9NICcKQ+ofkGL45H
v/rVOGQUIBid1ssTFY8cXfMy3Lh778dPU3+nSfaX0PxcFuXqPpL6P6U2ih0y2537olx67XbU0fUl
a3jG9mAYfnbQBMq+TGLUnx50+3d+2fKG3Byg5LqJuu62FgjGzhks343oa+m2KfrlEx0MrG3FnoXz
y+eQtiVDA2zW2giFs/aMLjIKop1B/3OJqElWLtI1iJeZYqarRRJmkhsvVbScs/asSiibrZUOLojT
vk9vHHzj3Tboj9fMqAQdtNIvlzhiSHz2uYRccZTDI5iWYKDdbkaDK8qfsRcqyw24I7pJm41KOvR1
H6xzvrcIxTUvyKppG8yeEMJmQtM7cBDQLMUPajQ8mPwe9dvhrSpRRHrliJ3DwsRdmSTiOQD8x3o1
z11z+HG2JDdQSZ2hWQZoRjn5p/qV6/sfHelSTZMyM53xt7GzdxLKmSac7Kva/7tabSlJmXC/MtNa
Giji3YD+8y6VhORm/z5A046w2hA2EkszBg8lgGzgwBrTWNyUt1GlCYXzWcoVNZW/I6P4a61+qFb7
ZtBEfi2lHnq+PtUYDVCL+rsJy7oLbyfPjCF3Vk6TS0BAb0pPqfk4FzvawQFjo/JuvW2OtnH3ebCR
RMztD4wHc8NrKrY4pUmEPEhXdtatU27e/qph6M1qh2IG+6bpSDaFCFFchWIlUEBPvsNiYeGBfqmj
GO12zyxTm7IO6Sxz5RwDnPUMuQE0s2+f2LV8+1pRU9mGT0sF6+I4PHhPNmmGuqUzZjw0zIS3F2MX
axhrsR9IOm+7j9oFIumGLOQj97yviQy/tmATmGBeb5E0F/BeyXm+iVhvR2clRgSFNVGca+voWD0z
zHfI+s0dHzYFYzLIWckwZ69GN8mlgycrNzYTablE9h5eIPzmx7+GA5niZ1UwWJ+koLnv2SyGt9tn
dkqA11HSzGN+6efvlCX9pNBWNUHRBRw1qVDIw1igl4WKuBMk/1nANLa5/4vpOoInxN08TFEp3NXC
KJKKQcbYexGiIHQr/R9owQ8bwe3cJheaoA6pQE0Oq83F27X4ZOJYAKS62jI5F8B9TpaTE1u4PmdU
us1TgufsWOrKxnEZgWEceHvsMJxbVVxuIKeFatLuqRkSay4BoiCyIBw4erAM1iYigjXR+mPZVCL0
k/wMUjmX3yB/Swyqca00Fv5CSiaWsFVLasIwMoTgbklOcLQcJR2jgAiZRYVvSwumarG7Jk1tB+4G
H95a0HEfqzjzUkgBT67LUKAGJJWTrCrkIxvWJJjRc3d+0yzYPOxlHYrJIhrx1/LLsoUZXjlrequf
IE9avywryVwLZQbyaM1R/PItI+7nkZdEQN2LuqMKR7vp0CPmreCjR1wq7/HDWjZRUOJPtKY2fmMB
cMI/3k6wdaWfRkZ3rpyTbiPPLx5ktrZ3uGTY2qpT5mOQ/gz5P4Q7fP15HvYIcUCUxADc9q0rwWJ5
MmVSZAvCJkdoGNbsZqGm8Uls209owSw0SKuomh6e60Ar6DJHJEhdm6Mv+YNGd7ZpD8MEZbjDfSBW
KFs/lM7rEbvos/5oeOcNEEZXbohelsyEuBHfwGYPC5dGzwyspxJW66QMGScGtpXi1Z77rK3BrRnF
qqf7UD+zHTGrp81zHz/svQTYvpQtpHE4xu2WGkACnm8p9Kj55zDaiyTYfRZcbmmqXOy7+ZO2WXZE
AwOe7xlnnCEl4F/81RL/2T/Qtn9En3GOwi7UxJk3nH19jlb8zcU4JhJVnOQNWykY64Qb2fRXrOoN
p4bxm0vKaaEag+B6V9cSq8LBbnNu4NCH4Zsj9t+vkjiwxncZYxMkszVccivAGES/lpWqNgKfNRGw
6GwEfaaPON8QWZj2xwJYhE/t0PePRu9SrKs/bhcGJ19TKzYn9YJWKxJCDxWPzAp7xjq6B1ImUCnR
K110oabwbHV4Safn7gU2WgrzaWsHEihAw/5uQRoA5Z3s27jMlhPLH9DsqVC8jcXOR9ykvdIC91e9
0AWdZutNYuMEu9W9gyshTgw5W9l1L14w+vWWSkMMTvV8K+oNCv5o6JD74ht16+ZUCh1rG/0FDHn3
cgAvv7IGFTtIV9MJ40cihvIFZB4NBPW5j0cJnMVUgMS2QkzOIedPb8XNGigP6gmMeaSxUeaHe83s
jlzmlfqExzZWJ68u2yMBYKu4W2q2ifC6CgWqXctF00BbXiSngnp0ikiXACDciPc2vZ/jldO5ZvcO
rVLDG6EGPfxfzPmfvDfkU/p0XmxxsWrQFqizD+vnbNUMw6qAZC3H1NRxT4j6iozrMyFuAl5lR2Wt
UX7lV/PCttcrSypqO5ZpMvUhX9HmqLRSiubA0NaJri7q1Spo+Z6Esw8aXX72DtFHpMRqSAIQcHcy
IR/RX/hLixxhmPHRC8w/21N59eo/F0KQqLQEy2X4h68IMoQ0TZGAEVgrchGFZba7EpC3+FIZ+lqv
z6UVYbPfmRHqNNVa2+31Fn+NNht11bhEy7C1amDJ7GzmZcVEiRdt3huzrNz/+7yremVn5xDutWgY
0AV3gn+n5KwEdNTvu+9a6zfBj6+0Gy4SL3KxPOTfusT//2nsdaWOohf4Hl6bDjWMrQYAusJb9UCK
2NCSh/e3DG8kKa80r0gSVAUXa9adDZSb+80zJWGW0B/AWabQDDaaJxc5oH+6VcXPobt/FfN79Wgk
saKEq1FGDHfhCGbKKLlny1HNJhICy5m5LU8JBrMKf6nm0bZXnvQR/3adqwkk7MngbZJOmpfpkuvI
ZJ1rZFBPwMJjSnXWDU2OJwKeKqaVvuHv7Ln5zuUyA8ViNWBHNuEiOoHgTVshti8qlqN9W5uBrhDo
4LITSAGa4JOHiSsS8Izm2Lze0Eo7rkm6Qo+LHpXgg6wfPXAPpborfwHA4BoUdX3FXnqWU6y3nLuI
kCIpsAMGqpbc0IgyQU3eq5+LKM82aCtl/PUU0xkHZ5G6V4/3qQ48AutRok3h9q1e8g/5FNxPNwHs
IsUaYT4hx85M2k2yZj0LWWglvqu0ZNtI1wFKLOYdjzt+rzve7vfw//52rGllbUNRgqz1ST4hMxRz
t7JSux/yNgq/gQiZoRchKJDBt5YqLG9Q+4aqpT8I9fd9E8sl17Yjl0ofAmAZz1ijd3C4UlQzIf0A
k2w1bSdhDC51A2+yxdGgUTIbGDwrlTyWkffFijo2BT5R6UDeS+AcROCsRsqOBEydlGZ6ew+hbp5e
rL8vh3GciBgknbhs8zvHKOqWOxBiLizy++PAFlPBeiKGn6v+GF678+UvPgNqLwIPPN5EqxYOQITg
YE3ZzzHBxFp0vMgLI8VripDnRm3Fld6H8z7tBh4XsU7fj5M55+E19uFPIvp1Cvw+Rw/GuANK9jBW
q5mgZ1idfEEm1QfYql76Z//OKDSchCJsZIrKfBCkUj6w5FS9ia33OG/Uiesp2qJNVsTr9Rk9lE3T
O+gTCg2dxUyDNhtW9YBGcETTYZzuj/LodEHrjTfrHRofxbXeg1oMhQpHThBgqgnG+ofkHqswaa+j
F+dLCXVz1GptUHgq1Vvc1qamGXy40QBJhkaradwotjTF2e9XP7+7L4vERRIDQwTDuHYVBNsv9FaD
6YLQoIrhaTvdozLptJPGBg0j5Vv0eaQxEAh1XLt9dakBZSIytdqP4uiNLSXHOWYoa0lYNbNgMz7W
fcOScxjs6ihzJGOR6ZPKkb9WfqLfgp/Krb26+7yje905Qj1Qb7P4RuCaQN/f654vElzdQ0CZ2N/Q
b+ZUCGKvPzAZ1uWbL0baZdLJBZx1/Or7POP4s7BqYwBnbUqn7uNRqsyfbGopwZUmznt9b+jQ268q
cuNQc2w3s1DKzxC5SfBAqPKIqe3Lm1JWb726bZGQQMbIO0Ll1a1eagtdAEj5r1R/abMjB2AEw6sJ
64IseRUeIcvLuk6H7wKBXOTUue3uJrLMhmE8uCGFt8I9nzT/sJMoellbDRJjG6CH3x3ibJuzr1K5
XuOm+rfR/0svXVLqWZ76SLFym/8OgGrCSBiQ7gCOavpVtf/K3DfgRPsALFikO52BX3w7r1hk9q4R
yHYXFNBP4Yytfg3Z8yI/hNkv9nZg5Ydpy2Saylspm2D7d37zNavziXM3FIGTB06QapRfm0J56BIu
NeAafe44CAwuR0pU03OMPo+GZchPE1ixpXXo1e6wpP+gDHcwMpnKnghTj9UQWqSIQzN3LoYVsB2J
plSFTB7sia8mCHiuz2Len0Y4/XG14/Gm3sdWt3Ac9wYuuCKei00RLUxyYYSota3LmxRLHDD5XmiM
jYw2P+RILLhTDvOxHduMo0YO6pwkvO5cLQuisH6Kei2IMoDjWiTApRU2a842yOULsul7UxIkjXDQ
43U3X0aBo+nLPSFtgeBhXO0zRY5Z1hM9gbQEGqDQvuNxQ0bfxlNujnir16BvlGPuQVYFmpdzc7ZH
4FrHLq2TvfaMAqx3qIsGJbVWLPY3XW5aEVEtdPeqZu0o6YL3MC4XbehPYUwZQipg5sfElzXRYgvw
cFYks9VI9sTLx47YVXU+x6LeDFA842vfQWLRuxiOQcU0ye37i6JlYrdP4hXayTKj/dJLPBeBq5FF
SyqYBvO7BkLidqlis4NYK/RTNsJCl6m5UVgTE9sKMS+IGHSkhvvR/ngf4+4BENMAIeiiGJ2DnMWD
boYTmCwloeTy5zSA6kvAGKPGVegnpeYBG0QvbkVSDp0c5yfYoyMpbTIlqFQ1YN3IBptQ6fJTZ9Fx
sGnQxYHrYw4iINUSnPWhB7FYXSyXYYtzfPCyVUcI2EC7xqnAOwm63+uCFG6HSPC0kc7dRJsWycaw
sVQ4bYh5X3vDlnEdWRqQIeczNCu8kjA/pORzY9tt/HYmvMIqnBbIif0CkOr03ecwfsrNX9fGo6og
l3n2MbT7Ts82qTtqe2aHUbOC9NlW6AwnUJCRUQiiZ4qQwJsz+3OZngdlR3W+iMD8eUWNXep8AOFS
sc1yLEMpM7JWrw4W6Fmp2IIA4q/e4W0Pqd5x7peFVbMFofiIHh9vx5upwGqYyhGkBUSNEHqNDtS4
TEF4tvv584ID551yoHzV2x2KJmIRWLlfWFmG0eBPA1skAwgeXc2LXpvSxg616tLCeQLN9e4iSei+
llxXxMJJYwU0FTvk6YIb+VP68e6uSnWlyyoMmta3DQKrjxd5CkrN3ogVi/A8rG0Aiwix5FauqE/8
aPw6iG5/6qCZAUxDRdoPW4N9Q1rzbDrEeBbDJAhL1W0E6Tdsuu3ZS//Wa5R5g6r1cMAPbZtpyAP4
RX8Bay3mKXRVdMAOaIPvQuWNMa3xFGChRwmTm734tkjOkaA6itat8chS5FOiI/Z91xIA+fTjMbP6
sDyAnuJ3DAQKl9gdwym1+Y3CvzK9XBkuMvn/jkyKIt9mKCmtbIo0SEeUuxYfFD8y5pfNT0IHUW41
k/pm2IL35yxrXGArdkp4obZ+APYkXoFe3y9yVXRY9xU0kg+xKosbh+ug9uR1MJgcG+hM+ayubpwu
DaQkySYyroMxfw6AFgS2ahUSaaYXpYWhtQzfJGThZkQyVVxNV89vj1jAAbvOeAJNE/ScRIT4V6Ff
JS+iibgFQlNbbI3k2z5l7fh9BghFJ06Na/J6TXum2ZnJqOd35piinyNa85C8chYdiDwv1t6BSuln
Y38Pn6SVzECqLtL8IlR4EKEvxcIiUZoidMoyKRZUCyH2cKZph7E3y2IzJse1uqfy/Nas7kldEV63
iCHTlFEA+raZoG7ErKX8LkugHvSZd1elj5Af+piPxZ6cOiNqULb9K0Wo4ru/2dyLSJkcSHvNyHfW
jFHZmOOUNM7hyD/qnpBaMUwqe2UycnCWfRfqpcqz996FDmOjef2X+IGNk1jSA33fxyJj2d9tJeTr
RaIb9UM4S0H7up2TyQiwz7l3dLhP6boPZexBj7nyPzx1LMgZiFJ5f6rfYVda92SvR5HKohqLIYq+
YI2uf6tSnbWp7sYYS6ZDgrzw2QF7898/7TvXvOJpH1EyxHL8JBkWktqWwXdv/ds3Psn7J6ELBFgs
AxO+IIzbuFeWP1lCHfOy1B/lRdaZM9tnKOJ0ZoM+saplbE72uSaAVTV6iRiVIPwlgaD/4huA6cql
PEEPkZJBWEwBqQ9dCXOdv+S0Zn/G3+IsBA88NVmd5at+IVR5SmwpN7H/pX38RBZjxzRW5MV7Q+/U
xJ++kr1UjVXkr4ALbR/dvoxl4yfukBplAuyiJvft+TFTvWvVxIiwOZr4I7PN2VmV4VKNWczu6oAe
iNiOjd4cdR87C3SeEPtV5LNiSmxufKKe1OQk9l+F4PrUCDgSbsIg7cri2A8+EayFhCMr6TVlnsJT
utRpoUs/Fsc8ZEUveR0Hwoy6bIiF0Vibb0kBuEM3qBLcyBOW+jcxV/6nsseJGM7AkZ0ncuqkZARy
llwUBcmcmVqld6Hq7sz41kPXbpqnWRlV3Nu7UIqjLxoEDs3uii46aO2nttOvjHjYzixGluijDPld
8QLTzcYyBoH+4AWnXtqu3B2mWCeypeTqmg2Kz0b3jAR9HtyiJs9Or2AKkbANH/qIUu5NUuR3AORF
Xoj0kYtQ9u+f2GIu+iv3NblHZfxZFPqAqA6c1zRsGgTXt7fYrhOZM/t0wUmIAIDMMlWV2yfKth0y
GKQu2mnbIW4miZO6Egb6eVjghKhF+6uSIKHxW4yXb8N6W085+4vWBTqO6GFSmzAC+rj+V22vxpm+
5uXA0CfWqBx0uft1ZQABukOrG8IXdV1YAh6ujQhuGnwWtAmlw+8tnKleewijUDcFiV6A5UBaggNh
c8JpHK9RBtLE0fNQQ+BT9ox6u2zvfus6LqRRzh+jhvH7x58MB3d7Kt3T2XnVRl/hjQf31cf1ndup
f7HQ9BbPY6FVCJ7wGJICxHXcPgdAFEZYHvfkl3IbAr/IdUGrGqojLA4rKoMb5mUY/4Cu1Emhw72K
EqfP7ZvQ9gumsorIngJJkVzA6zv8Iepo5hY74RvubAyCGaVDgyh0HXGWDNp7HugYkaAJm/xOxULA
aH0xxppRvJ9zPiWWzgot69/QLYMU/gzJSUJRH0CR9LN3i7VRErom2h5su8RaMjdG707IZy8Vc2r9
UUdKe67eb41Mn8u/WIiobzjME3MLv731YbgyBbe+vv8ARlCKo+4aAwDU8ca09BW5XPCGgzh3z9Wg
a5RwbWLs5YZrCLKoXJNcyw0k6Mdxrw1ZdBK+KT/Hisie9xdwITr1tKYEW5rJgvRu2s43uAqnVJRf
zXhiBbNdZXYIInYRdGEGmH2V/2NWvv9BZMEcefhyF8idPj47M7Jvvt60/nTtG/YKBhueRJhQAvgj
qxkgMlFWBm7VTX2p9rzHTHIOtC/DPTEqsdh/GADd0HoeDZP6+F1ZC9/Qo+Swc0h+QzdgQIUK8doY
iQOsTakmWiHXRTdigyH+unD0iMcsLtyMDNRGeF9Vcma10c9INGMjwDnJLSoqUhAcIYf6WEKzJjq3
NbS88x+AgqusYu9ZpExOOoY8OBqDWKHfVg2rqAw8J5KhNOOWOA2ouaJRu+Kf7zn0HA6pTk0tcstb
dsfebGLSPiQsHv0pJddchkBd3IWteVxMqh1asXkEJ1qMURm4Hbf82if4Y6qCUx0Cq/bt5HFx9JqE
hsvVWW+BqglH8e2bPgA7fSiuLTPMJCpIVQUL9Zpfq5iOvaVyKviuk0GprfgtBZ+AqRXJBuM9ookw
CH24OjK8Zi466rEcN6DHpGuwrQ9LXH/4fiYOsPHY5wPt4MpgGxlPZCIWYxnb9laDbZaQB6S72rnN
uw0/WNcbIxl9rCLo4k37xz0QnROpKHKtA0DSZhP+bjSBbEqUAtGt36tUibxwj5ZHubV08CQXgQ40
JmQ1YU2ePN339LtYz+VV3HNEP+NiI+a46T8n3WoRM+1MltTmp1kAzP2az0ZDex9O83TdVADStQh8
emndHaTHSPKcPtZLCKusGFLp+J0SB5adOUVtO1IPREI428z2cXeQQrR8W8x5kYLluvulEfSoJH/I
/1BvXzEgl5Hjyy05BCpwLblQxrI9u2u5hgxOa5xen82+o5uPok818xKoYSqdsOTD33HxXdXQrwgb
gf8OEjSmIZbCeWpdDOFfPbj4eCl8Cn3UcqJhyinl0ZWL83dXZNdq3UfxmlMUW8V+Vaj/YF0PkBy6
83rZ25LCIukPO5ILCDJntoN1URGdzm1nPd0PrcbVqQ2N1S+loIDQ5BTRmcywN6Ez0fJVmSXfibN0
w0mi90gncv3wiEivNWReQubmIRHlbdcSRIjfdaPlwGhEn3X0ggbft/VB6X72kZeE4ooWDvoS+gjp
nmoVOa+uVU1H6i2ivK9MZi4tJhsvMqajfnw2fzJaGbe9RZNqSNCwKeRLUGsfGHqjRUZ/g+afpAT+
TFMZNB17ndqYtmtaK8kljjvz8bjeKfuSK+Tsj7R9rZaU6Epg+b5vCg58a+zCdPuryFpK1BikqcMH
X14smjNpogYX2kLFn787SjSqWFMXDzxmuSIjTWaigsanXkfb7YHlEmimiv9BX0GiBV6WSulRpO/F
Kq41BW3BJ7aqu+aGvokRGn7t+e93RlQwUoBPGESanr674xkVG28l+e5RFtkU4LVz4TneInVVVsYo
kjuOX5g7a2Cr+sXfQdmWDR57jZbSDofurAt3BEHZAXq6983peKJhtI3dwZezEWQ9LzZwu5mOEbwF
/Z7zbcFoU2P0iakav3sJTs2UuEg8yT7mRDxzEWItxGAZAXp8/3T0OanuCv2xtXXiTzuu6TtlE8Qy
1OaKle74H/dZj8QtvH9OZXji7t9i3rOMFXoZKMMOquo20t0wInHPcQKcEWDldWdWU5dU3L+sWrDF
JA9mnCaUVMTg17nmvRpIh+3bS1Oe+tLDPgwx5WiEkUTy4XKHGmLL/ByCLBFsua8ySJrJI2hN0qzZ
4i9wiAdeIfitzR+yNYQ4BFfxjB1ctbrMJw4ATSau5aWbixFA8zCTd78pS4Vg2oPlE+3kF8JB4RKW
eEMpchI3csLSTute/RX9f1wnEhGIGj/haUBcf14ZK+4T2OGlRw/qcT/eolTyYsOVDpWFE2NRA9A2
zCNa3qTZDSfZVr1IzdTvOcJOoO7NCqR5INd4P4Et42idNj+dGcE48hDJbNU9U7QF9LTiOtx8z610
t0bnAKNGHEJ9pMuj3yxRhi0H3ef+B4sM9o4mqfpldiQ9sbvm3D7bQMNbCsiKFWCW5Jt4oix7XaPb
y6+W6ljkoqUMs48dWZoYst+1331LkDZTdIvVBjGcPpEEO8+Sil5s6jq7MCXe0+zHwa6jfepSl6rk
VHCfSZn79GtnwsodcJO5xxEgap9fPOxmdvHDY6/obvn2BjA2g3GUxBX2VeBabRCMZhXHkUEJ4Gml
SHNwcwP0AgNfpqQkPZPaYVCyIdzm6BlBB5RPuGjSYg7IFeX4Dvkk5yYXJxYSydtL/QoAuizqNE/d
74d56v25q0QEzZmo0fCqXwC4ZIGcBWM9JiwoGY0SEgwteOHvwRw9Ojgo1OI5U4it2m0Z7ral+dz9
0i7ZDGti+lvE786APRNDt1P4k00PL8hztpR30uGOySwgmM3cFI0KZ9spCSObZnt7961sEoB1Dfg7
CQ2ps7iID9d2Sukfke00ngQ7I70S9FwlSDFn/BZQ0Z3JTZbMl6fBo0kuMlz5aptRMt+cITZA62gH
pr8xqGdFhnQx4RLM28bPb+Kw2qYiuoGXGtgHL3GVVt/NZh/h3FmmC4A07TYqzqaIlcxR/oOy70hb
zajd0sXeg+RQqtWmsfcrZ6GKQJnK95o4QAF5jhqPhPtFZHV4QsSQeLe0B3RjazdARX9tPm+VJUv0
DZg3fY3F60RPEclcSd3uqL5elpsmvcSbMLeQa2m+nUx+6UHfNU4b6kdoKOI21WxgfZiJbibbJSbc
nEnJt+nACrwc63tRWHrF6TPUt1x3HZcIsJ+KoKobe/4j0Si+CbvKZn0iavv+n1SO6oXeFoNfwSDD
jriprpxE4lYYfl2hbscM/6dQFC+HUCKI+OC1nqYjCQJvcESGljbknADduccBm6/BFl5ps/6dIlmL
BHQE87JCX+uZQeEBWINPn8bC28MY1ONV1/rI/plMOMA3lGC0BJ0hUKcj9Zrc8j2pzNTnYFGD3luE
App0YVun5UUp1hxi9pNkzuHraQMwq31yqiKDxGCKUTTKPoXfYAbTNngsKCm68lAP8qUNfeeQjF6a
Sg6dSAKQurprvbZoZ2BInwDtzhIFBf/K/+wiBE15qaUXxMbFnWbOv60IcYSqSdW3cCXbWb4UFlLr
UnlAzP6+gwMvIoceFbjwk7E7IQj6xZEL4OENorkCxWm2B6lWxnuC/RCHqIH1DsdEfdISUJPv4Ddk
fw68GXJb9BZLwHb93wdeXjkjCgHz2YObjLuXX/+qR9hZV4aezAV7vI3L4IAjs4v0nze9KtF2QuzB
dFMNJdWZ+BxvSdHH5MbBP/opNgjtlAT8UxwKFxFahzjv9FjxatRnYNVeNZHsCyZnHg6pfDAbrnV2
TXYTx3ISxRsNCPnn06Y9wxEC84MnC2jYMOul5+h2tebKFO4Tch2CyW8gBwQ0AvIDL5lEXkHmYf5X
QDyBDcrXxAKjOfrR/RFj0+iZX6ToMCV9y9KIwpvpMc5P57m5Ekv9zCKtoFZBZX5O2FXvdeJX59MU
h1/y8xnj4zrJbVy1MYfIhqOAP8pIoCP5udQ4/WaKew3T8cqbBYaGpKFVzr6TYGVMsC3lZJc7Vk/1
z+MidNtoorxGsp6yCnhZmKL/h8OsDxoLs/XU2FggxZqSFiHpJCR3X1jUr8Iqw2f88DqmOlwWqnqb
tzqE10kQyroEz9lvN2uBkl9Kfo7Icm6PSdqwMsouuaH37+cJceAjRn0F2mbpQ0TLBLJjMyUK3hRT
93YeiK6rSwvhpwfwGQMeaP31uAZ9k+e6ES97Mpi/tlsjy/17qcqQ4pVVbMmHTdfNISxL9uc2hSN3
glhHCw6Dmpo3y682+XjQqQh4VPrGiGNYkEWJPge1MhxQwiDfISNocX7iub+tmoZrFdOMemLTWRId
tg9+9QL9oCWlUJ+l1xi0+kmGRAfyY2HZu1S7ryNarJqPMuij1hSR4PtGER2mnX3ahpBXhkabrtPu
MNPRpDu3OC36YAHFPmDE6K13aJzvCHhx4JZzNoHr8VtOQPrZGPtNgAzyXziifQNinQQmVEuD5IJ1
Gb7PEf4SGfAvS6DzfOyPORRUCpZ/HOpdbBIaJduxFrkrN3NHnPZxIIIkgC/n6eJCdNWHEv8STuHK
mrIFAD6mlRginUqcB4uwV1034baWYl8wxc92vrFjOF5bqc+oS4gJJ6pJYkJ+U/bkEI6lO2qTyu0J
zrRoBDECxDcwWcUQqLejEGSjdQUPZRiun/SBIkKOjPdrcL3Z96+E+XEJKl9Q98I75IYAMEue4DGM
QmnNnTWTiBOgnbkRKTFVYfvK4tp22CNa48+N+OUtiJp/Dvvo6PKUqf0ifg88TbllvfNx920qkOHZ
FiSGMKpdmPmLDaPjzOWVqsuasMNCWumnbqS4phx9ZJVs3DvGAegDrmyGu00mCeL3DsLRA9MdRMjI
+PolsmaLObonmOKd+KKISDy2W1I4XhmrOtrlxvf9q5LlJl+MR8dimWZXNN2XNAoDcbEOAh5pxl5h
rVGAnHCXpbD1lXLnv04VYqRnBkjOlODMbxa73v6sis7zHXaf+cb0Ky6olP3ySL6qvT0XBcjo318B
VgqstCu9ZVaNRbHmER0SbqmnUjEptk/uZUTRe3t0V8CKau2Y6Gd7oXsb9r+Kpq+6ihDvcxpqPxHs
75Yr+/tO76csmXzL04pEWKQtURPHHk3U7+aIfd2EnYzu3zabhHgi/yatfT07IuExWP79WM4rlefs
J593h12yBoTr+Cy4+HwKrNLOMK4FIjXsl4X/nxkd8pyr/g12fYtfqIYhaE1ggpy9jDPOG6eAvk9X
R/KOdZcFTjllbNWybMZ9S+hZqaXd6uiZeEPXnKrGj0gNxHLU6ycXAAcLdfdkzV8aOXSntKtu2SYM
UPHteQ/oDm9e390VPzETuP2bUNsvDkBuajyFhEWEsYAFrM8BO7Ii2TZ0Q0ztyjIEFSD4+H05aB6F
Y2HjrJnIbkKS1qYyoGsBBQOn01abGoqKQWnRUeuDUhiGcn5A2w6Nrui6khRzAZVOk8SdxHcjk2AW
NPacNKsMIGvzIrFhVF+/yQtmX/CUp/pPlcZvLH6jn2HYfF4pLDEvwqtFxfF4QbA6BGwXQMa4g4lF
wdZudnvt7oXKMhsJva7sWlMSLOdjd5dLgjMG0P6lqyLccT7SoXqsd1urgFy/NjUYCrSxvI7SUuQ9
r56l8//rDT7ecuShkGEn1XjHK/IQCrRFyJEKgXklheGH+YjXNiakKlWuxxJrTHSUYHN6GnacNet5
zW45INFJmuQgL091/ucbm+B4ns69FjJiralSuzbPdhZTiqKrdSaC9BjVtw8SG27NqjfWpf9d5uK4
VqJ1rNszd7Gsmk7KQUNERGgYcKOfsrZjrkOI0bogCEvkL5O3hZTkQlrT/q4/6j+dBFdfDl1DWvRO
QP1O4oHu614H/xOog+RJKNysmG9zx5Ekudhm+sYhM8/pNpAfXhho5/4qxt9lsJ9/ms3Qx7TsXHSy
AJtuX6L8k5Nq8fIy46M3K8gZVol1AMldrrkU4wAcuK+oNoI4DXB1skT7LSKnVNJNDuII9zT8qQAH
ECLWWy/4ibJxvniFbAt4MKQENh3jkNB18+KLde8dDMnG5EPt9dkWqHGJUerkKQxuirSuOV1NY7Xn
dREfQAMKaNmPRiWNiNITn3Sk3scyO9i85RM//fdzSEyPmBZKvd6Klud6nrsvJieKZcV/9Z2UeJix
lS4TuF2+NhhPimDUNvfUgyjM3q+R9BBMDqSnlExfv/nZvkv5GoWBMqWPuqOWh7+QMveciLjFGIbJ
6PiOY+CcxUBZJwC/8aL8BRWEqStCEv9sb3M5e1+mHPMWiyWS7DxTZiRoXqz4eMkEOcpSBUNzCVqJ
8M/ySKHuMI/623hoeGSxDIMTUXQESQEpbBqMV4jApMc3w6W4w6Pbzy0FugZ9sPcYWQBs0R7E2mMa
Y2ER6+0WgY76mnTzYpxFFdNpyAXouSztUAPaliez8FeafXBLsFGAAeO2ExDmMoY3REQx1LPJWcUs
oUqM0HCWbu9hSiWlRl+Zgp+ipzVJ43lAFZL1WYBp9B29c19jvCihufcDDNolxJ8njVD//tSkXICm
kRzQfxHXPi+SSJteR6lNIrDxy+vsGQrzNTmDJOv0DGXpaCiQPdvzFI/Z+71l0brvZQ0B/B+f6ddK
JHZI9wjZTqqTVw3sYFNh4VFfRZFtM8Uf5PWCzkrqkfLJxosDEmigRG2NMLlK0X3j9xqaOCmF+vui
7nh5lzC8xfWbOTU+uOlnjV+Uio5dUSJlYRLWfkAuLaGGMK1+DPv2VOnMdtXL4npDnUan32PbGzXq
EtHfgKmQLDQEfTiaeObRrf2PZvOM5rz2vcA65Y3rXKwdAk1P6FJfx5Jb9Z9eMMBXMRgAVejyXEUN
shuyvYGsOkzp7nDbzqTy0zqh30//R22O9TLWPuapMZqfUEuJltbeyLOSxPO2GuWK+cS02yO8wya0
u3BovjDIcuNcFbQVhIwf/d24zLLtszznP6AJf3c8Al9zmfMqx+VPht7SJ1Yv+7S34VXsVnbUku1O
AZKOa6R+JbZ4BzB49WJdVFix1fucbAvs8mFLntL7KubpDaAviXylVnsyyezckUi4nqtY3C/kJHd0
ZyExGFhNkOITuBWyx7IkzNTIc9QmBIOl+DaiM+lDfn5qzaLCd8cl979s95EaQIQvigcsmydTfFPt
7fPZxrQ3cB8D3pc/YNTSxSicGSjwAN+vEAjyE5oa+ZNZvxj2EXKn38HsPlewMe2y0a9+/F4u/vFv
PSsIOFEIRRhUXmKBmjgJ1Yr5m2e5RVlQSMof1WZCp6uSYgz/h9jCgMHeggQQ11dk/wV8V1+7FniP
qtz5GpeSxIj3morLC1SyWw8zOxvAE56XtGWnzWT6eNN2niCi9DoeQY8KxjZ/V4NeUSaZJPWuYF/z
1mINMCSWyg7wR5g+9tm82cUyDIuT1l19UHR6pZQfk4Hhix8EryJ1Ygxd2PTJj/YV+w2fCF2qeKqP
SgXyaThZ7riEs7VBJlRM2Z9O/EICTW7XeuxpzQ36+M5YIYSLjvpEwdSfo/S7l4Tr3q10jw3kIHbz
U9YFDoaEzAtDjramb4DVuoAte0Z24aHEKpk3BzVvjbkODhZl3j/TbnLYh/MqfjWAWNU5Ps02RMy4
+2JC09RT8F96r8oF3AZQ7USNoQNGYzRD7XZiQm6g7j/cGYzGjrlpZer2uY/vIH94ki8tVBCKvVPT
5W5WYjLdKnrIkVkpu9Ap9owCUh4z/Jxytu3taggX1FRq/brFdlZdwXQ9byWn9tbKbKhT//O2Y7fp
VSHKe2NcXuGs3Q/CAosshyipE6yJvKYh+ZCe3JsaaVTTH4EymvwzffbH0djDQYwd/aNvgojlXSIz
CK/yjk08YAdFS/LIpsCSPvmo8Q8MAhwSN1v+x/qqAlcF2iIE1RV7vhRBCAEShyf+u3su05WJGiuD
5OOrZHswU8/NrSDsNLR5SOvXvbUOR/FkC7dLl9FaO6RYD0oYzqB1n3LeB0jf7KvWcmJYrzvNkdgk
HV9vbarIhzUOtRN6Tlg2Z6ai8FoURJ7Pe7c+Dbdv18ZFVOXShT2UH0g/1sX78P5SM2kY5In2G2vp
p3pHyZJ/1v9mUtzfo4OlGrShAtoswCZmTYFhjsAcS+ETd2f+HwvRZHDmgifmtDM7159f7R0wfnPO
En6FgIJ1uHlTa7+YoVBSXF8MfxdDk1j5lrpzsIX+15GjzdNQoKyBDsrZzyy6EaqlV3d0rUAvkJaw
GUv1ENEHpGd/p7db6upToEwvGZh+CQRxh67SVpc+RWEtT54MZTRAelKp5wHgFae/lzXF0vnfZf6s
LqsLN85CzyOldJwW69klKEp8eGjVmxyx9WGQd1n7PL3oOF/7Qr8C+5DiRoS8xj3wB9PStzA12Ef9
NTZMZA5fd/H5J/pAi/sEpNgY02bMmViiVlG2rT2iwP2fp393Y+I0sAX8LSJFJ435xrdBbzEmzxNT
bTLT+OL9JRMOXcsibyhCT6tsDKUlsvRZMxrrQkFLPO6j1aWC9mWRf6U0zT8scdnqhEhaznUtIQgt
nsmFFWxmooPtwEU16N+giA9cSizziqj+G0GLBgz/MeG/HgLfEO5QHMnYKEaS1AyXN4X47UTxYxe7
nM9xWM0PPNK7LIi7vQwaY/xZfgnKj7b7ohNTp676jqpTQa8NDnvGn2y5FJ5P+B2HW07HkoAn8kRW
HUBIhs1Lj6i/1vB8lvpmoiVgeWYcBglcwdnfUFzEB94wkCANBEQ5OHRSml67phzIl1aykOo6UVRa
0ctUVGAJqew55DCnGKPz3W8JOWPb2YLzQwqearDj5TPrWsNeeL9NyHn0cmFulQf+ihXrXTTu5Qu3
4l/kRZFoj4/8dNQH6dd+BIqVt22JDz+JUOio0Q5YO8lcn9hS9smbHxfcNftqq3kruvR2dMT2lwWP
ZGsLI0OJV68E06xlLs6CsLMIxmQpzwHWg6X9kEGe4dBNz0rRspbVqeiE9E2Qq/46Lrj7mDGbvTJE
Xm5yK3aW0TaZCXq89AEM1OSEVLcrepHw+uz6ymVDlN/ieegLLVB3rbqj+cDUlAzlYZ6ymhDVRxRK
MSPCQzb2RaAglohTXK7/C2WGGaBJ2V76ZQAO1VztixA7OE093e2RdkKXaL1YwnF/zHg5rYxwxUOF
pkN1M0MqjUP8HE3pIzhuQMHSDhEi07nm7LYOHu4tbaEkquu8Bcih7nUCQP/o/8nZfI+KuAo/Gk6o
StdayvDez0YvWsp0j+ovJWyap7yBGwm+5Ded+HOWtgDcuHkdyB1PO7EKgOET+2EsPkdOtq/EgEVw
qiug+kME2hdjR/ymNXrGilApUkerRPYz/IgNIOwn4SGFt6s9MTYH7FY6/AHQ9gjMIIHm0u7QWNvm
BeFVL6K3p2bYGhLnB5hZUGe/57Xbn509Je19T6UAY1WEi8RqcaZbhWqeBMti6X1GIM7ut5ojw9uQ
2evDqU/HX7nWFovclcoXIsKqFpZcfMPD8ZqoEOXaE1lGte0t6kpsrdnhDsvsZ/6u4VV1bG+BpP1M
GHtZlwVOjDF/S2DE42eZYU2RXxbQ4qEZpsKDaXIAVP3bpnqfSZlXiBcejKuS+5NoVoEhX/uNQ6cY
5XHOJ5kmLSgfAwV/wyCuWEU4NgKNKWvfoa4zm+TpoYZRtHR3LfMU426vzbVxFaWy9RxSi7LCFlfR
HN99JqYNtfd6NJ+jR+pmiuX/bg0KJNJax/N19II78ttu3ypMaFTD4TjrFZMDACXZaK9QwsHx4X3U
DeW34qmscgROZ3JJ+iDIXGi5W4cJDSxnY/YnWvgUKxx0P/CgIOm0eaKxI9jJ5uqTR4s7pBhJS/7d
2TTFc6L5f82ofuvLVkwKTogX+eLUXFzNV53J4e4Df7cE0+6C4PA5RGxFHsp/o3qhj0BjoAAKJrhU
TmCgI44YSKmPN6M0vIVNB9s6/xC3/gSA7SH3YxP/bdKlELAcTIkAERCO5/ffLvmW61UPSHeS/klO
X9M12PnC8CArB1gQViCTwPLbV1eNbNSoKXx+Ha2fz0NDCGuAWk6g4ghMlHOxUv6I0p49ozXc1uVR
wLj8ZmmaSZmTgsYTPo8ndkiCdu+NgEgNK0TSxZMLnw4AwFMj8ODliIQ3Cavl99S/iqy2DTNyoG71
OM6Y1pF4z3R6dbvjlpOwq5V/i0skut75svFKgPX/fnjFxk1yuTjgW9w7odUk5LBE3qSTjAKtEC2c
uWu+Z+ieWLL8nsHgghb2k5/ZHZfL2UbnSPHTq7RuVc6Mg17B+qx+S69644L5V1mcX++ZIRihpIyJ
647Ejr5k1aEc/8lDvp6JiTtmXEe4pRTMnTq8Cxvh39IYTsygTZhwkKSyPxSs8V5vIlMw/2mRH4VQ
UgOenXOqq3L2Czoglv6QDrn6z7R89ibNSJxdcClY+iOZPa8umRWY3IdtrMx+TN9FdLna1Pf38noC
UtzVqXIJjzL+jGvmDlqTbbQ+LbmKv9lLyU8Om2S5gAEyZrwaZPJT80qdC1t9h8Cu2CzyPZXAGJoh
+FzqI0oVk04K6a6tO7JVdQy096foTzK9TNRBm0brEjBhiFoa3kH2S+rchSypDSzOFJGRxqb3qFRX
C9D1N2QQZupCvVEugW33Qr7KMexrUXXdMfXuH299EClkvr5cggmWvyR1qSW/laPr4xJUgYJnfCtq
sg82/L4RwfNXenWpT+Llfj4UIJWKZTJ8O720C1y0ScxXLp9dPvXoHAuVHcovxOjVx609kWwFPzzR
Av5E+GA0zxf10xcBkPEdi0pSgNj8mkRVLf8GgszwHu+5H4lHNcNVim4UjyO9XLoZfOWqjlqRZDFR
pdNO8EVXyhm6lVkB5cITEkFN3qWHlJtYCpcd4unO0Gu3GSxOCm/AIclYqdWJxG9BAMWMp2WlXJs3
ThVVtNd4Y6B+JPns2FwBrFmYQYGaBGsbKKRDxjZxCref/BmLJnVAqu5E9bfx7MxgOj0avzakNM3A
paUy6aZXnsVTIKA3Na2az/eK2XIrBcfTKV6pFjHT7Zm0P+oWRN1ur8kL8kLix5mKwhxt6NyZnh1d
qHh9/O/lenILqRPuGXCW3KHLj6rkeS0s8LrLb0MUihycbGugaxMgf6Xmd9G3rlZxhwVrL9c89sPR
qjs/eAPa/ph6uziFLOvgxryTerHisG9kpBD8+VW5ET795ARnckZV97P76R5bgp6JdtpVdj7kMDhP
AsQdvcQ3ASL9I5R7r3L9rHsD6vkYqii02QWOAL6sCufrXnOoh2RZYDWBbgaw2fz8I4LAbfrAwFus
IBisoqUz9ei5kz7Xy3VrYS/oyM2Bml1Lt/kuUOBtSzcRCLdAFWtHGmSYsW61iW5v0HsOEAvlFUe8
qeCH8JbQvEIeWKe2CaZK4NgMwNha6rSB5VI4onz+Z/p2zSn1dQQYnAedhSDIxbsB98C9T5gbFL9W
bgq+kJisqw3I5vBQT9iL+27F9sGANjLf3m4HmpaylDtcb9XKBti1fwN+ODHYokshAbFYc7BSxELS
LLcBUsAewzI3u1V+RV790wqhKpdYEGD/+D+056ga0kqg4aEk2OF/z8PRKBilDCR6zI4bwo5eN8yp
tCfC1kC5l+T1EbUj9N91w7EOilYIku0OEx+NoHzzlrzrmc9+N+Wt8PpEtR8PmT6xWn2CFQ2XcoIE
EmD2MFdLhtEzis/T+iUDalFNBPPDVMrvMUfSxY2G1YQ7XOFZXqCKhOJoQ2nyO7FxhfGbeeqnbl5U
ypL5Y7FmeM59zqXJSCw1emYyeP+p/kzs9vnd4cuTIfGS8nq5DljkI67iTsGvoSSeODjnQMiF274j
BWGK9IHXKC2clAn9jIvCLwbXR1Monp0s8DOmrv1EnJsYyy3PMt+392qT2D3fWThK+mt8mAI4K5Iv
Ke+bWVpCEDCTtlnOUjSmLOUkTbGG+d+b3S96Iw4FlHzAAKltayzWgFAOv8zAtHDa4iDHD2mYM9E9
pN24F9YEAOaJVw7JHPoaRATFCOIG1mELhdY23J+kFy5Eyufc1KC2kdSxFL2hUzpowJ+VKCr/SMjv
1fnUTALd2BfB/2EFnhX60I8wNLrIbvpOU+gXfF1dAkbku+7ZkoV09Nd0wU4/E/jkLxotT6LBXwvm
L2EJs+mcthoawXLL51UvRQPTKND5o2nSABo/OBj0UdAg6mhFN6my6Tq2qDIZ2Q+GUA27VEyTiufj
bs+gs/rUqHcqLxGR9Yaeh2eCciYcCYAhGETu1eX6i8lh8yGQS3aZQO9Tpz/xXAwZVd6L97wOg+9g
6t4QJnjewoxKLIrVYwXCBsG5KtGcWC6k4FgSU1UIF+OxSDGfCzxSsbJcawSi5UUSA8GAAmhJgEpT
FZh7vtiV+5k7ygOKmAr1/+TwHurLXmzBuk2eCNhY9hGx/zG2wArZPz4dabb6Lo08TBTc/SmxkjIR
jKBklJZs34z3pF7YTrdrzqZvYe2nI1j9Bnm1n3byBVVDKdRLLNswOz/aDvDdnz8+seZ74+Wao/xo
feupAkfyZE5yu8OdsdHeqBpXEqUBecNSE3acPtOeAnYVRo5JkPSUGPd3kPcbroNpkdZOa65Nc096
MOvZQOG2kZOckoM+2xuzznjAYanmROXFRL/5MR+Uuz0KBCIUjUOLnAq3ka0c2g6bkiXogPJPnhXi
z4O0h8YWD0SCc7dbUBCCkamCzPY1jEgKr1oFANFDjPKTIckOQs3wdWP8yIdZTXUFTBajtAQSdfBD
y1VyuLbN7aak6eLjy5D++ZN8KuFKfmZlDYQOwiXhQaqR87HzRcD3QHmvPZBovFWaljeNQwyQIPwu
yTTzQs9NBc8sMg0/auDhlGC0R2WDzAU2ZAckutg8dL6DBuJBTQ+pSi2m4ECvaCYDZKpHJ5VODpjZ
DvSIY4bHU10o3Q9rYS/sRCVIPRHAZCax6OORFEW19ioPyyWKwo6DlUpBA3v2slDhB5jXRz2dh1l5
REx0b3syIoC/MExGW0mgvZ8840YjDgMtRTbiFYnI/8Fyw0HIn7qt/kEBtM2bF7Xz27BiNPSTykWT
WsT9xkDdpFierONVPUiIAM9hh/S1RUwEgCF1OnJDRla3tgGjf2PMZtkRgmL4xpDtC7yDLxxilNf8
r8jYiyeNd9jrjqmT1K+nf8sMWhHLLcUos8KxLlYUtpAiYz9yzzY2mP2d7aa0E59UvldSNCypEMRM
/xwPDJQ7OwIxjU9IP1HwBF+CSNHjdRkYvZoglCTvi7LHHoVv5cZTWz+PyQseLLDgMwipXa4r7kdl
ZnkKI5S3oO+1NG4oSQZZAsU5UV61PXVfpcCJehqSUAwNj/mx9OiknDZZApPi6eJoBgRMkivE+/5D
7eyZGTuuZkvUv6ZEPmY9+nCHiuSB8bePVF5eaKE914MbnNhZp+wIg2O09GXRkFuKXm9kl1rD8Phx
PT/yB/draj79PW937Xat8hhC8rDuUxvzf7tsY8Guw8bIimxionPXBpGAt33vAZt6Nj4lfFbv00Xq
9kWEq1VHjEeWEG0okWry6Cz411F55jePa37G1UfHil0Zr6jB7Ht0LZ16QqjSBWnHHJMYyYz6lF3r
sI+KZAR50QJU4BWLqAY7O+PSe3NSrXYISQg4PTPPB4YNhedrV8crlLz16uYr3tM04vRDw0ARzqG3
YKyXKefDTbx/7RrwqyQdtS1D0MAP3AYz8uwqEmIxbePCEGN33USABjswYPDLiF8a+1AVfzo018mM
TmqgGIdJsS8Gr3ut0uYbq9F/8LHVEI97Nu6ozqHRj+ebHmr3a0JciquF8d7LrDoEl7PGszWGcYjj
9wk0qCHUs/rSoFFoYND891P2feWVCZZTKUgfRl/CD4skXC5eF9CVbo5cjtkkzFPl0kKM2r3gef+I
6XgDxGMsq5JR0md8mH6pxKp3vq6JP45JILB8vXSo5FXchjQmmV/iyMXpNzhThhbulWpyM7mIhixv
MiTJywDFDoWdYxAuhZJFAjxFeiZ/gYCqkvWEvLMpKc2VFW0NaxHAbtj67IKvwH0Z4AmUEQdIUwUB
uCKQ0jedJTjW2oLOlF8J2/7CBtpTsozDDYZD4tAkO9bCoJhkY9N5bg0f53hKnnD+Go7gJq3ZeEG2
6VZ5eK42sQ9aqN5AEjgrd9+N/f1SSBCnrkrLdgNsg+hT4BtGLjG6hFg5S7p0cIXEVgUjzXNZgn55
Kl9e4pQ6Lt7KCaXkPIvQJmsW6pcLJwn3tMmkR3ro6tQV7QlrtFloMppYK8/CmmlL49BnWMY3U6FQ
KiBekFcmZiuoz1eGWAYDG9bGqBy5yiAdWX7X5P1tmhxV9ptEUTzTk0xOzfLWlUSWgVR0RT0AJAMC
/FfKa5NqQ4MEkfanBbai2rI6Rm/Gokc9wPLPCf3UedcWnDhWp7/Z0ZYrsSFny1s/PAz3ScF1aHOb
GfFU27HWl8utY3eRW7fJXknloWY1DWe7Efaff8Cgr9FH6JHiAHkRyHLdCqfsZ+QVJqiZoVOB/klj
dQXH9nrObDR3Vd94NKLawojAJjepA7aibmu7oIMmmDNbX4ohomGPeJHmPQFo7b+7Se8GWVo6+TU3
ogWJAePh2TsJ9zEaTXChJ2Z97zDbRswSMAroHmSK+3AvsOmacjcxnlbxALSlYVDIZrmiVCUHV4xQ
NJ797INeykOGY1SFmdqBlAbhrAyL0L78jUzEqFvUhI5DmFYvpNKndGPlWj5bGzfGgNM5JvDEAe1u
pZ6svI9yi1R200AIfC6N51/irZrdPiyGAF2XxCsruCoPRxkv52O/U+4SHWT1Z8JnlwbFCdmsVUb8
a1tfPePFbagCRt6HeCavhFgU7GBe9wb6LS/uztGh9/Ln88V77izSIOvEd8rHnDllCNaygBWa9GYA
N5Gv9BVtgAua8aiS1gf/9v616xDfrwAMx02mPLcs82UWkxAjUqGC9kXdTJ/PKeBGGeKlqNNyM3+B
GyaanWD1BGUwOrkedfsVGh9QyOjD4ZQpL5FS1+163Cc4+anayInebdlBkgdadzCLXp93Dgsh8OB9
NL+Vhs285bQ5lAjcQ9UPjU4Hra2lc7TPjpwhQIFVGmD8IVHnUBSgJx/hwqBvEPz62gNkpfmoK3aJ
nX/9Ixl9dOt7bAsdCkhAEpln0TZMnFXno24mcN/gDeA7rLP4fmNP3wpbHOkntu2U7O0zu0SkhThA
JvL1Y/MIKAkwMGSy8TaK07EAkf3ua9kARLohOVYuXYd0N9sRy1uzc1mP7bs9Ge4dlZ5pDPzlTkn5
rwDwTKeLBoGwZboUQCgkSMB6QFnnLkGw4BNbjPEi4A2uLS5xdU1DX3tjRP0EVIxgwAv/WNJJfqeO
8UIP+vK43b2XQBfUpWjnEH7ciRUW9uc4r8qcjM2b2Uv/fZIhzn9UKVq6BLQ4QRKzjhoUHZePtA1P
+a+Cx/KJWk8DoKWZqevzF5cyQ73uem9qmKnaZ7z6DXVdFnMxUzHiMuyaqj/J+YWuQ0Dy7xnfvpGK
ytdeWxt1Uvzlaf5i75vtuTd43HOG6hMSKvU04b8WneVrpLpl70tNjaVokHGNhffjpL8oU3CHyafi
qm/8gt66GSRv4mKB2sHq8YnvxRlqbv0kjsyxGIFEiNvP1yrTEDdecv4+YWhnwvkYI3f0D6WkmYdq
o/ycCZUQem0rPGXNe5Bpf1kcKRPw9v9gOfsf8LQw7NnONPuOTYWIX80L0x3sLTubMxek3L1PtypO
kg1bTQrqZZFcMzeH/YXlQ32iqEybhSGWzPR9B3cyo6mV+dz1ZI9eka9i9+5uXwotbtpU7G89SMcl
sNQaY5Rp9cq9peY8SERnBKkvm0JamLrZX54q4AxzFjjxEq28Xeft0rS4N3kEQOR+OLrC6fg5biCA
GXh75UiroAPrtqCFpC7ou5Nr6ZqBuVY68UtFT6qfDPYhIPHuO+OvKpzhNL9Nw+2vmADSdAQPju5l
+/7JiHaLsxPuDk1U4Qe0q4wRczzlFID8W1+GsfzFtx/bZGYOLKlDBnNhBKskjnOpURZ9tXio1AvJ
fdfuu0S6davq1POW7B1HUlhywyu8Fzd8CdKazPEWHdrFUU7eR73WcN4ZK0CrvWxHulDr9036autQ
ZW+lXtMbuRdPP9YPIWJvbkURinhm7NxFUPIovEHiS2R+YwQHe6GAdA3TWT2mV9hoSMZ79GyJ+C/r
LFEBofjr93Insefa+GGNQUyvvYyIszNTMIDI3BvsN2mMNq4Nfb/EqNoIeSmkVcvmAmXPmz3/ZWWy
8sIRAHlcLTOSco3qOnWQHbEOuH/v4GfJctLH2Y7Xitc+l19wMafLD2WQyZPBwI5QM66RqYqwQEB6
Pdgx1ZkqtT+neikBOGPC6e9syjeeZTA5QNYCjpgYk93QArvaVfHnUJAJvNVh6EO6jTmxnkvJeyjg
H9yyTG392ThcF2For0cJnNB9CRo0B+9BJAV3NXu5EFinak0lW1RNEz0FBgaqTKfLluMCjJZXFQWY
RuG40uhyOr7hZ1Q7IN6NLd9aIHGuIKVy9xuBLup/sRUmqZgdqGvoTkBwARsA0zmsuwJJXUWNnhJa
jscAYwZpds9Z1reqMgkChtbngv1qB+RsKFxC4qZIHtUKFHQ3qfWU7t1noN7h0Jg+mKTpySUwS5qh
O+qUuwkGUhq6nwzwcDmEg10pUmXUKt63Yhl8RVeyRTFoDhQAXND7aqE1C+GNk54WTrsev7ng+TFz
fpqZkOR2gpWDbXl+Uw2fwc2gzk18FxUReIyKugfdB+1EXB5sddlYkTMw2kBfZq6KxpxTLP0K4aww
w7fllJJfkEfcltPBwxiYHLjAxGQUs4Ciq0WqketGeEpdRPIO9/gMM26ItMfn+YkpaHxqa2z1sQRa
EhQu8xseysj9iLk5sl2Qgpwj8TUq1izRVE7erL7jVeKuc57yHseedSI6MoqJKQKO0o7YqFVKIqA5
K1HBD5vAzV7/BG/aXLEVqM4piJIovMEdGCHFqqwCfCRloRIR3M4q7/zFDChl++ZBa+gK6/nJxudU
uxhaoFSyYOXkfofmFaZxwGK5ToR1g6GR3U4WMlFhG8pp9jP+kMjFrL8Di5hY87NvTaLN4Jfgipe8
hLMFLf/iYMDHuUFRtekDsItRGrjaNSWLazI1krm/AGZVorKCqFi4aZpe0uszBIpqULo3tWaLdSFD
jgHG0vBQqHhay83lkGBWBWZOFO54kIwTNdbDrbBhDtNZqjAEB+uIvln/Cfjy0/Unzm6de+eQXA2R
xPGJ2S/EzAPKGcNilQZFRtO+uwIS9v2qitEYMgXdLx20hfUrRgZK7hVOzTSGpX7aiyZo0U7BJ0K+
wd/lhs1jYatrMFx07/RmCSc12R/Kb9A26UcHviJzC4SwY42bpjLL3CgYioj9cztZlw88tu9O5RhS
LAWGKVPCyU4ZsAzrMnbOM6bI3lT9NypYWwvjy2RikvHaeunQ1eKJSezE/7OeKjtk+I90j4KDRjDn
xcQ9QwWVN5yn9f6ABmVJU9JV+QC50oBQfweCIyqtqwGJKc9IXY+mQvmcyYIzzm7gGrOtiBPocD1a
a8111z1veEdEpUV8uKj7ROXlLrjgHfN17FhxdofZzZCmZOzawf6PW9WyyII0NqRiMzfhyiQlGIvG
Vp58scG0oQn8TvpNNVrDGT5i5/5vD+J+3ceF+f5ucT9ipqXUYqYQmuqSJy9O72BtEz0kQeSHIGAA
ph4cr+mLXVCGggodXB/xRptcUKO1n7wc5iKTtvHVO7yfdqR4DgUsAKMNK3DQmDOV7x+yh2XTahj5
UYI4xSs648pwzsb+eHVFQOBBCI9S5Qlkznf2EFrMZBJ+l1vWEaBhKMmoVQ+0BEGRDNuGILtgKFOe
GU5yHjdeVr0OBrmuUIvnWH7x8F/NbeMTf5BOgLzhrOSdvkmZA66kmQ2fVWa12rVq0bqMjGMltnns
bt2jnl1NIbZpCI81TfPa8TAUN+EQY91THOQwyne5xAkBpb5wouZSCMuSKT2QjFd24m8lnakO47Ya
HAO1dszYlIJX7tborQlEezOLYhGMMgQD7or8uYdry96ZpcIO4d7FtUcBvvwmR0h4Q5Hr3jtoHfAA
8PBRzDBTQBqMktGmz5tnAgRCXIl9Lb4tQa8jqbRcVtqQ1Vkcl8PviCnrWahgghBjz56IsLn6oxiT
JYrIX5E7aGvawmrhqNttoqZtReD0U72q+CoOrx0ln7lXyp1HKSXQxjPhS6Op9XxQDLBvlqUmK8bl
XxagKN/QjC7IYP5pNp0gBtNH1hY0Bb+t7rVtdCa4Kx4J1axPYaamYlAwCUBsgRg1+9b0uPsPJcAV
Ikr61LAuszKqM2Bn3o40lEmWoSHHuJDFVUntsYOK+OX5G03IKiztEVP/jGm3/b6rRuAFS05L+zL3
n3Ri8ja7xzonM6fiEG9DN6K9fbgjh3WVRSYMKCp/TJKmabQYNYdyLqhj+cpvFrGWDutEPK+0EPRr
6KjJjukSXUalFDXOp4hgrS9eDOIafF1+wDRsQtrkclOe+d8mqiL0e8kWi39XSBG8KgrR8fPDnKRf
Hoai+I3cKOuwhzXTfNwLDXv/MfciL9/E3I1xkd/nRc8OhRb9aLLQ9Zp67DbtK4xnM2x39O9J3sc3
07JbIMNnmGmajRh7bM0oC05jsTeZPEpcevfCxCeDNr7F0rNTGB8lsFh6pvj/LyRFlcREMPzWiCL9
zmJq7RCvDofR7HC2bwfpv3QrUw0hLW33dwq4jHUaqsYEvVtxwOMpjWxYvwHApuWFkobPmT075bC6
7uASwdaMR7KOZCR9dcCBJT5MRIbWdFgg9en+JX8wu9bcjqJ8UdOjt+SfIAH9ugF1xapKHiKHF7W2
t1ehF/oAiM4dOHTAzEoReZXutZYD2zkYGQjGCzhIVjqO5tqc5TKt9Wi0PIsh6m6GeRl0zJs0WrqU
CbmRmWiaOPE8LDkJfRVcu7LF+0a7qaWC1TJPBHrk0WM85g3wcBURAOYKqQQ1DuF/dCgMNAyLBvJt
JcdCje4QuoVR2plpPig/YSL1PppAEkuDXeBPXxHQ7z30VxnN0gI1dIMqtTMoyx7aKSti2ooLt0CG
iQVu0uF1mIQ39dEQe6n0TZ4rlSVJsFHH/0xjtUg161t9AUTJj46Ji2PK6UJwysglJWWVjSDVMJOm
bJVe4+gm9r9Lr+IsWRmym1pFk9wcLvgZNrrLeuLrwPEFi44pFefr4iUef2Hqv/D4shOpmJmzkt6E
tcuWuQ5/FeIHamEyudqrUPsVIfNDD0YmIptgzqFqZTz+/b8UEZdDMdlxko141XBdvkkZgVRsdEGr
mAUsCacWwFNTjwLkRCghIL2TPM/7E+s8fRUbV0dyqpVXTVC4YVpkwqBfcgD/vu/AF4KDmd+BnYeg
cn39ZDmnRjeM8LlYP+TtdOba5femcOwa5oJQtB4t15lWRhoPSHIqe4SErdu4lVuf6lU5mHTsQ5cS
0t30j22E3lkai06VHnrmn32aW4W+azvfQ4NLp2d1zCTUlowMdPlgxwiKTCRSMzo1qt+wimzwAEkL
I9vZu1r7m0Xj9LhNK0dEczfQyDIOy78iBzddOizaFE+gtWHhoGGJzHD3+opa9gnG6djI2P5fqiQi
gQN5C1e/DNqs5veD61Ty1E0gKdap1ZeG+dnDV3TgymzObdd62KnXQb7t4/ZBjdRidSobE55AGXj1
LKuCJmzztSjTR11UpimCSazmMEp5Pt9UzA1BYW2/rT21r6zcjkuk2/rXaDAfC0wsJFiOTl5AriS6
2xmnKvujNiTAO7XvfF/CPZFNG/oq9UQccz9gLr8SSf/BL0Nvw1b5whfQi+b/RV1xsteajzSRIsOh
FPrQRP/mkiUvKxz6VKzxjIVmR0EzbaJ6tLbdHw6PmFU7a6j80HYctTZuBnzGSUqwVVO7hpoPUQXg
LOpNNNaVMPEWWv5iYUSKNmJY//0Pu/SwZ/EV+SGvO10sBiKSe84H7HIirbF2JhrfmNnp1bNeIeTM
2uvTGqFZqLLt08uedummJ+s2Pnj6k8uTDAGeTN7L1VHcP7U77/lLdPYcUJGVgv0qiOR/49S7kbAo
6vCB6V/HfJSzFaNQFPUUvqXdd1dzbZrKE/9C
`pragma protect end_protected
