// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:42 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X/wcVG3KcyhmJb2ZHKZbcHD7GQtiI3XWvehD4wJaoZ2n0MaxWk0SuCEl16Ib9VT6
oGxiMV7Rv91vsKlN9ZZNRdiAwrLoSk6xh1Bqqx3RFn116qsjlFWzAfFZN6ahq1nU
a+avpmyvu4xV54KBKHVQT5HPrqIpbAWabJPRZMTbbyU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7920)
ECntlUhhMCXop/vBGWl9ym4hKb4jyUfPr/Vi//qv8awxJ6yj/PG7Fw2qe/fnTt2F
diyHfbCFq8KA8Fai53YeeyeEbYymlRvGGGdaM8hY/LRQcql/yHLuIVNolClp0veO
mA8B+JD8Z9n4h1Iq57M6TAle5QUEiQLAW0O6bu3LulD4GNjfFR6HJk/IHadfDUwE
iWUU794apEdgYDKVaKv9QoJu+ffWkt4m/R9ZGKA2Zq6EE8fxKLsMC44Q1ktMiF0r
t7sPEGyzUVwqpf9tqoYMsQvBLUG8kpLTxgx03dfbaP76x5LBnZkw51wjcClw81KF
S2t+xw2HpbKI4ousaz+TEkiZ+5cgJNO1fp7KRLfMJ9k01Ut2SwuEibraIHWBzve5
N0w3PNUpaAfUoPGblkf4J8cy6fnu+ms2TdtirhsesdwzcUIsex1WZJHWCDPZosH9
NJ+OugxTfgaR1picGM7ViklEMJRZstwOCi68x7ppwvbdfEFR3vRQIaoy3QXxlsz5
uSPdbSLwDyw0U70IJ9AFVXf9yv/e1Tbz1RK7m98Ksg/gdp5G0a2xARBVOLVCu0b5
lOeoCZyCdyvoXjBzPxJ6dFRlyCjfvkCr2j6lIJyZkysR9yApuIe+YckFDlwSeHTA
Q87TVEvUVUNkVDgwfGlJ7hvN+qAMVyj+0YRr3gRsZk+s4HLM79mDVLUvk7v0+8qR
2Y1HRYNag6dc7bBS6/4OGIf5I8+OpRX6iUi9iSlQFgla6FFhvHRLHF1S3lrKllQY
nmczMBRv/tc2DCV3kWyXm+scyof6Io6Ya3aQiWfSVPdE8HCT5t6V+cxb2Fyu6C8P
YEOuAbzhk0FhQ2K3pf/VbEYwRYo9dez2vZMDGdk0lTvkSLqF6ZOAZ2byUFLGrq7s
+6a9/LKOy91xFD7eaDDGAnoEtZS612Hf7JyutxytSz5CMkt1tV8LiBNacjv/RCrh
6SdlXa9ORY1mHImN28RHYi5FDPDPvQ/G8PAatvgT10sWMj3iXDFCVAxLukYJKy+l
CWJkjQ//QhrT0tvDndHwaulVpHaCNIl+QFuBpElTMmGU89jXzBIU1dWi2Ptd+HWg
e8IL+Fik4rjFLKoRDQJnxQoiIjj6vmuLougGiaXF4/Sq1HXouXOl6EkVhbEilV8O
58QxCUCc70/7rQ+a+PCC4A3aEJyLFIsMnoBa4P6Oqq9Qd9RhIew+cVb6a8wVsqxW
oCyGIievAI7SZLMEe3vCy+9JlR+EL0Xm35JqR+HhqwYgdhE8vXIV6njwf7yM4wC7
853St8mNe2NEOvhAKAKF4f/ikCWTVN6k3t3IVZAnM4uYeINYieqR+wgqjADLdTCV
SAnQVNdyaWLXuJuZ3D06gt5lGisHkpWtIY4Sj0NUChG1TFSpnquCJ9+KAodDCHy6
UZluoocS80m+4dyPXKXCU4h2x97UJf6D8cb40PyvqCOjz84h4l40j3Nen/SNsPeZ
wsuyKJwvmfW5YuGSgMmcrDJbZlyWGIzBW9yd1lr5liOb1F3D6iOQpg8XlKgNtm3s
de9D4BgYEiM4Kz+OS/h5OEby94PBzJZQ1dj06vHnYoBFrd1UrUAEnkouLczQqtVd
eV0PosSo1Le+/gAg+hGDt4RX6FkoFWw479q0R8SEZDYm6l71pssUjkVTSKlKsl9q
jguJEER1wtXJNiRCLdiMZalyPef56h3wMvNvbwGnwiec6lm/+NUsLfeEU2yrdIdO
mEfescws7c1pEaEPAqbhaRYXZbmCU5W+7TB+GEfMbznSIzuv5NBOTeHVbTY0BJ1g
Gm22QjbF25GX74+V5uLdN1Li8nTx1609e/FPw9kyCl9sjyzK9Srz0Wr/Zh+eiuDj
uLIt5cpFM+jtvgcKerNArY1lf/EMjAXDB9FSMOzAeS+Zro/JCOlCGPnijNz2ZH0W
RIO6kETXuNREIElpupZ1vCko6VyEUBfuYkECGeRu8n2dDi2QNVp0HwrDL1lPCsJq
amu7OywCLpccY5A325cw+oecDS43lernaiHcwKLUIrsx8WY30vFUeibvrnCpi9OM
YN5B4Kql+vgf7Um7EN0WRRByBmViJkgnEC+zaf550SNiUI6jX1e80z2e2n6UZdKZ
Medwm1TVp2KFJOeIfhaw1beVTYPOBY2ikQtOrjtjJDYcR+VmHpVRbnJTCiHkDVYo
0THTbiBOPdIUPj/lNLufFXof15M5uotnYqh3vWGt7W93w83s3Xm2s0GuuweL8oVK
sXDk9E6XqSBoWydlcLAT4/thUpDP7iQnUNHVtIiOygu4yRTy8TMJrHV0pdNKaMY8
t2qnzfzyYYTykIcFCjqwJYD1BE486S3Y+DkJ7C2jV7JnpXk/NmYEVSBczgIMUn31
ivNIL2txcy7+9LtA7AhxhcSsfIkSccCH+Je1xqds5HfM/MHF8nZHVLcdkFHTC9mV
bPPkOCpimsUnSQzjngKN4wPPGKOHaZipcXovggv8EQ1czY/lamtMHapbolyQR5Xb
bA2MGgHxEKmP6ofPpA18B9nKEMCihX5tte8+0S2QzNKCApKQEbE4S2NIWtjWXA2t
9tM1KbsT9agtEDB24UnycMxSK/gDSRK4p8Yxs18tbBi8nO/wvLWzfYVVUUllN+so
Es8i20Df64sSE9rgXfteCIcn3aMDei40PcFx7nfjuBzrlM2FIyeO1//uHAlyEL4n
n19XHiRTgkoTliRbCi6ZhWyJsraztemzJNNQn5QWNe5OsqjQIN6sa3wdEaLNWwNO
n32V5f9inVj3Rsa/olBw5uy0cEm4lmHvJAaQu4tyVj4RnTVdr5loYDdku7AL48iV
qfyly15jOEaXpat466CDaBQwa7nk8LyDP8KEmEPNyUAkuWTwsQKoVebQSTGQy7tI
7bxLpm0q7w4zdK42+eKG0azFKL0y9s0jkRoQ5EMuuxiCVxrPd3sFsrNnmqgRYyPL
HhEqYu1gqq6tJjlu0L/vfx2h19FoKZfRI7gTzCHdPVXtZCrg8ZIBpK/7/v/OpNZj
vjRF3ln6OXJ7oGBAxhpqGZRBscFijWT3z+LckSbjoIfueyrFFn3nAXQN9gnCRKg2
yMuIwCVmamslPX3r7YE73i3jCbibIfA5ipyGuWhZQeNnUd8/DcJjXmmpcO8AJqXx
4eXEypXOH+PwdXk3VTwnaxV4C4EV7aS2hFDlmetfLQPLooLy9M5/3NlUYug09ttq
al7c+LwVd0MI8OcjJx66JwFvC6iCobX61f/0GiW9SJlxyrvtU/oEBYCvU/isPi5N
6ZN59HtkB0/QuMBivZkjnf7klj2nAGMBviZi2FA5S5lej7UIdVOZBU9pCvCKvJyU
tJOWCCOIDWzdVTVZ+3l/l07dxdjaNdOROeSgRk+g8aTM6CwRjdW2ofLv1rRaXu5R
/iqcQD6cHSQjGQZLrwGZrukHfGnJvAdHMEyn+hftP7VCH5ndYwRBu3Sbbor3VYWp
73N/XjDZzhflLG9Zk3tIQYYC8SajJhg6Xdt34jyoiSEXFtNBtwo8VHbE/tINnUbe
WotwHsD/iEJEkcxPSHSvmZ9qLJnSs6mmfuMrZnfTcZ/EVIihMmbzw0bg5eecyUTH
ZGuZyFsu2VAmhxBJ22PKLXYaK0tjhRRD2i1JvcTXDt5bPWXaNR5TcMOqIKAqs42E
4f1WaCOxPjMbHX3gSkFTrtJGVC8nArYyTbRhrQ0xCIXtSiJ85+OWEiWdd/DUOaMF
qg1qwmDGDmnHBS3aJ8imTlDBdl6BjM1xxtZzaTW6JWMrFr6JsEOztoYsQTwuMzz5
AzJTW8442udxcBirjfYLqB6cY1m1OVkt9gDgUsdXVD+yr2sbvnykReAWW/XBs0tK
NFV80xk7YfRsPRH08X4O7dYvsC1V602NkfCTbYDo+6P/tWQdcR3lDjyifXpqfF/R
EzLJY3gLd1J+I3ufgrvWTzwfltzzsNPgXhAEXlNnyjtsbC5g5M8Tzmq9CWc8xf71
oKjsoADsI8PrRSg2ULA2yjY0/EBZmtX/TezeQRXbV6PGLjwkxQ5JcZCYXbsizB4f
Quum0FtlyAiHbH6nBPVQMvHzSrmvYtLg9F8r1cvJ2D3y61lVxbjUerudTOtYjWsh
F2m6/d1Jdh/Y4Gdd9yH7Eh1rIejeffuHhyVfFURbjjzmR5mszv7hI5tgD0tY23M2
iXULanDLOPi2u4X1xgDeQ2Txl/MJr0ynisuPkOtpsmqd7k9oB61P0T1P7KLoP0p2
eu/FWlluO4AW0kKMzX9xMYSEegYUDF9NKV1GIKuiykzc9oJoxJaxfGGIsDbIcR+M
Dm8WsCnCt2UZxN9LpBMcjPvLyoD6qWMJONgLNH+B4cGc5ulrLxOfRH+6xKOYJQ+S
Y5R/eswO88Nic2Bm11i9Bgq/LmJgatYC0Tir9X9EYYIoR/kTOGc6c7iZRu/Cg/Xq
4wJdN7GbrgZgafL9l+e/SOcN7FDKnCIzQsplBnOxrAAGYjLPW3bUGt7Pf1gSUgNv
MwoJF44oc0LrzpiHc57Kte7UBRoHJzcLltlUQWaTqamlMWp9NKU88lMmpU/g+QqB
4vClXThCDYSTXthiVD7GySIYYbf+YKDxf3gb3xSCVVP0fT68GMlhhhDP3ea34vtj
rWIP8jYwrjt/o0+9n33N9FDb+iSgzvcQLRYfQavXR/DlCupo6M3lwLdpng9ndALl
h+129PK3SEMeHFvwteKgzKjJzHWDs//neavcNj0AviE6ZvOGrIjIpIQZ1n5akG1O
0G5LKgyqAbuSFSuumrfsELIbquQEeH/jNeUzzVq//1whR/3VQALV09yVJ44d2txH
GHRFuotKDu4KBjjAyRjZGPt8w75jQ5wGvAe4j4UrUssBJpXXagxxVq26SEZF0tt6
2t8pcMHgRrKZDUvqAjjxo2W6uwBiJnaNBI3sOGM28CuBmgzP5hbCZNrJugAohZMU
pxmNC2DE67J8HMoPhA7N4mF2GecyZIXMAzJjyQtHsOD3cs1MFADMqFrgCWsox3su
wuask0+URfd48z/SnYKceR6OPSa0NFaoKeXGxL4fjFCWGJfXXs6qkDbgK3kDGn+v
W9QWLrmluQ+PdvqNt95pu26DISRm5IKVpfH1eaRSOni8lntUlYowL8tIX3qBo4BG
Zox9GbG8QZCb8VxszI7ULR3Hil7p0PremHkuaAWpJ2C/RyGcb2jwHGOe1c7WJpHo
wPi/AEK6a0zmttSZ1EIpm+xFkHTpjbdvasCvkCTJ51UXVdpVLwP8xfuM0I1QuPVU
9n6fx6zwq31XJejR2zNYFZCuSrA4SRZgy4axRs4iYRxRLTtkrjmwYg96NE6wSxsb
eN+Wnl0HDZ+E8+CxoRmx1SaDsRXm3d7hy2Zq5LEPiZV4k3zuxYxg7IaKm6u+fp9L
xZeRKxeXmmRIXIiWaBQbINpxRkfEge5eW9mb6GPGPE+W56hloIurXvz6HPfzBp8G
PKvgqObm0e4DLiEP7tmNOFinZU9n8/TCfARY0lOfH9UDJI4cuC2Gce2Y+jTV+mwh
UI9h3peFJBKCxW5piWlCfk6uBcNQ3ogQ0+JYJv/pEbc/0SDhUNiV+8O0AJwtm6fZ
k769OQTeSVlKtimWDvGO5guaFw+CPTzIq+RlBR14WUBqDD1lBoxDMPUCW3Me6ccN
c5n89NKvl1s+F8ABZYihwNK5uTusbBeMWC4XDKqSp8VgfrF5C4hgluq6ZyFEFo3Q
EcSdT0TAP2PoHvTp95j9ZYN2FplEx4pVNP7UDJOcAaVLrHiVukxGtqwSLn89o2hr
3D/S368HYCFElfiSJQuHQ7AAnFjtCESXPTAbg/KhTZLpu92X/gPUDqCV1lmYykEu
tSzAVdydpvFtcx48Lg3LD++YGjJv6QXY+pgY4c1jGLIjlzd6bDUNU+FkxDgGy/kL
aCgvpfJyTokvmxQK7l+Oz5s/pYjX5g+M70pcuBaeOHL1BwjvA9LOLZLqF17A5VxO
EwFo/yotlfmSrAdmudXPtyG9zOzove5TlFYPM374/0+5kqvC3m27jNh3s4FUVXsU
bazkbpEd/bMweejbyTgCWnEWGid/qKhPL97pMgdqoOKSUBlxBWTLf9uAxRq7Bqao
jhwBKPlROKFfy5hw+t0vuhPpgS2JpAfgTDt+gXvTOIZdkRANmbLgSuN4ZirBgJvx
F/pptl56fIXs6iYjn/d0pWA4XDqbsAIPeDRn7znioibx+jVnsGJObuxHoqAQKXLV
0WQtK4ybdKuVG45549b7fcPlb5PuWiU8KjFyOy+oQ0ksvKo1187HU6k7oNImzJ8B
o3HP2Ijdwnwsw+8BWqYxUU1asRTaTL4fTPtzaSXAQUJOTgcrFCAJvCwLfcwQmmjF
9/9YeUnnlD7jGHUADwPWiVzJ9kDVpDYgRRLiLHl06zgpgU41RkDxWjUepHLCz3Gv
dRY+drFcj366pLnx+8kmjv3lTM0wK15pbpq4wV6GQ08aaCQyKNt/vUke3G6G8SLT
qL737Yrcu8WxHRMzXOXSkBA45IhjV8fd4SC5G4+mYa67ymdDkDJOANUyakFgH8sp
IR6TchK5ENqGZs8jbEOivQzFiAOd0AFKiHO2YOybBeTojxN3Utzf6oadKhWYDBiw
UY88geRNk23BwuGAmL+JyRwt1FPakifaunFsZZGScKlq5Bpu/f1L7Ly6Fw1KXbhj
6bBkl2wfphKfQVArtBegNDOZZXzy/I8Q0wClIMRsNeBgWfzndBLfTTZwKu5r9iuF
B/BasWoZAeiQSiy2syVmZPTro8HhRPP+Zz/jmy90SynxuluBY90MMjqn4t1qKC72
fjUn/BYpVSVQjbxU5PAAMlK+/1mC7x6xfaqeabzAXw4uMDVsY7FY/OQWpfKb68mE
t6oaz+wnQcCZN8tWU3/FGal4Xkjr8OnnTYRxRZAAqN3FF35i9d91d92L8apehUAD
sG5prOIgYOJW9gLYwBE4dFiFMhA5cmcS8YkcKd6r1cXwS+CCSyzm/c79Bt3+a1JM
s985siQPglZ3QlOC+zNLb3ImxhpBZp/qeIGJXiuawUZhnaF1EF3cchWls6xF/sg+
DiIyENa8RBEDLPtWr7ItT1v0+Q6W4fQxsuf5Icu3HVN8D3btLcvTUmntOXer8Rbd
Q/6OjUSktZcZcO4gm1qYccnFDOjX0cXnqvfGmG6yBFNK/d7dA1Rhl5d4hLrF/WPR
AIYWoVLreY/+rbxiyz4MJVLuzWLEfcsGsHzsbR4QZbZYSPC/GuXgcDwIHEJ6TSag
or8hoU0VaLIm1ucR3CG2lKN9PQ/PvPD1tR4Z105nZeeZFKHa54/aTQvviQs6pbko
2OeDerBKFVV78gpcLTfD46iAmH45uzO6mpHNoJXzqzn0J/pLhTc4bAE0Q5j3xc/f
tzs0L2cSh9wlZFjZsMpJGDK6gssYJv83ava+N8cA6nKb/r48fptOCJN+v0qIiUTX
+/Bq0jIWawEAj3HY9rnqgqHSi1qhfOwf4WuiOwpmsVXdl4v8UC39h2sk7HTBSsMv
Zf4lD77jbX8ggHrf+Bidf7VkGjOHg6/H5sT2Tr5P9j+doNx4gyUSucpn+qGP7mw3
IDL7hmGVHCWd9sk164i9V8EUCtDn5+Zghgi8qOKOlFiDtng7VMLbMyPGth6k47Mk
cGgb5R3yAeBHBMv4S0g1+F69qjKnyZU6m7ctwQOCpjEun2fvk4lm3Mh8/rByUX0M
PueDf2WDssItVPv3c8GHoNWzxpVkyHcjSiRC4+j1atZUGdWX1lJBMwpu9Oy9fIqy
ptvFstMrNJnWKxsnrodYGCsnF7JuD2hqQ6Ns/EulwQ9prLEIoazcNioTcpIDfC2q
9RDy5NsTWuqhVEGbvoQxniih51q7+N9CCxAIyxIp+c3mfjv4CMuSzZ8oUobjVSB0
+epi5sD8FmMfRynWlN1pcpK+wMucT9eSLV+viMF1sRdrXpQlLupehyFoH/H7xwh0
uy6sGNBYLg8ChkcAcQxk+JDAFvHZBuBM/J2ZAjrO7SHjIhIM8ZXqpc3RIaq49oYG
fZ8jB9p/8O8oLofVDp+BCZ/AYy5DRznHS4g6EQL30PlIsXOdUIBMD2NdJrQ9iKZO
04GlsY1gan5uAGvg2s2fnwD8gXDsPPTyNu3f19+uRoiLqIEY8Yi7sS8FTSyR+H/I
g47wCfbgvc9zI/irA6OzxJL6kZ8LSDU1kv8zYhTwb/JgOjBGfvaDOGigqw8/pCFh
pgz5kmja0A709m6EltkaoHznfpCFB/2olTEreN9XHHErQy67vMxzVxXqXgwKkiwq
UVCBXHgi+pEJtu4T5pS0wMYNXGH85sC4nED9XWSmmu07dfwJA4EmBSe0O50JQlXL
OFK8C3voshUCNzxEFtRkKvbzeG/iDWJoRsr5YDD2aNqE1mDQhfiHowpIX6mC4s9F
o45TIQGgYRk7HAOh/yPklO8uI+1hznXDvC7BrvHgeEZyHy8Q9A4PgcgYw8D2Ujz3
ZLlaQnsIZ/25on3j1Te74+xc1qrQ29HHrWP/lY/QUIyN4I80BrFpKEXsRv0vHC/4
S50vOqy5pRemZFTXa5n9SAYxkil8tzDsGZvoeSWSF24aThcBxReU2O7Lh61LAA9s
mLocz3mhUmk0PYZPaVb0iXSOZLBmAei1fVYHy0B/MxtnbXYb4tDUo5CJhN60T5b9
0vVPDJ6QEU8p4fVMgNTZhMO6l2R/xEePO/QOFCSa5auQil5pTuSv9WUD8ntn1PX9
pZKyLjbHIOh037gqLHZ/Yxom2G/gemiEJeC2BF9OiA/8nDGgZow/o75Tw3KyPAqF
1c75/igFCd1eAB9QjRytWAYqv0yvXoul+4qY77siuDodd2TS63NF0L82ixGIQO1k
bB89BiDcUMUds+HwUiMtXg7xmR3yd4dknt9QH/ip9QyLUBfflJm7zB1aky/DOqaT
bPmYrZxDWOX5lj0Xh8veMK6/rRTfHptkYqh8KadZyWtHuEy5/rfOxxPLpZHBDZk1
poEIT29TDvgxHs/AxBgGlKZhEqsiwffYAFUNk72+IIrsjDjS2fbac8vMhYQViTGO
mNBuuGD5C/OmRfryzjCavCQECSMy9BWXi69hGnp8aTdZl01gzTT/y+rY5sNlWFP2
FgPhpiRo50minth2yCtjo1L+fH2WkMTyM1iShakpkireJTlB6bBc9wGQh7QRbwoM
ZkUT0+TvHUK8+YisNhr3C9mWjLiP4jl87FXbkgYaI+o3kpPhzDGhFsrAaThng43t
sldi8hp1RudPd/xs5t07+MoBkHQ4DaOLxBstto9zaW7WbLHl5JnRlA/WkBoUxvqA
crlfq3xXWsGxx8tWyseIqsA9zCK0z4VWi3MihM3wfaIFjYfkHCI49Eon8lVAXKOL
p09XbzxnhgC1TId2RkelURc9KnIfynhwx1vzy0ml+HrFp43RPx0wsQGxU6wbyJPV
0onDVPMrtsAPCEVcSreuJLQMgB9alLFzWLE0W8+xOCX3zu8ttf1se+sKSqyN1O+V
FtJNU94WFx2j2sF4KKYYhAWQ52Tr1w3ayJQCvNOk8wQwCotDklMgH+wQBqh/Vkv8
HgEHX+xJctm56gvaG/t6LFn+VUmfl1fCNTw4Oh74Jj2PI2DV2qz+JvVYAb/FFHl/
/P9n4bBdGi9Qrv9ab6aL5xmELHL00NvOfJ42y7Q2s1YxrUyG4rpeHgnkevIrRWJx
gO+p9z47XOp+yhdjtyZPwSMvDySrNmlqgM1HbPoqRyJDhzd8hyozf+TmhcSvUSvB
rAeQTY1qmdnufLpSRAOKRho0/jQ9cRyGRhkXoSznTPmd27d9pfoIA2a7F1cJ3cl7
JhaJO7pv5Oj/NWq2igeHH2s3VZSutsGG5/rCSj7Z9dRN2juLxkCfQdEM3acZ/JKf
Afl703pJi4dQYh4nU+6vUKsDtAA8FPIQve9cqDYbnvZBaZhqp1Mi/n+WYYexZUof
DuFWPWMToOEu4zkHSYYqrra8SjZwd2r6WKjjVfe2YXnNRVrAdDut5NXRHcNcFGOY
MUI/xA3s2Az4RCEyDD1+jOdt2q+K6sJAc8WvL2GAGxuzp0RbZRifJgFs/JAWGUAc
RNGtET21fyybEiRQcVS4VijrN4JR38CVnLszFN63npNBFQNVWZT2Co2rOTFcS7yk
rA51xRl3ibosJjjpQooJO8kimB/xgjnZFZUTVn9jrXcOL08DhuwKfhdWWZJveKnB
1IJwjNqjdzWvrNyseE0PWCyJ6qXx1xkoQemiUqqvluF8Qv/1VVhr1hAWUt984FIr
OND12fxeUBbeiHTJLa9LZjZTUqszNexvRAxzmu5VDG5EB7KR++kQND3XDoYXdozU
k2ydVLl9/s4HLQXmZxQ7UVd7pmB3x3rNbJzgzHK6fw8JsWk7qPB+CeESR0zqWztk
+EN++zifvCmmgEUkg+OzvBQwNZVeA2wnwj7z9umFW91PB65qGFoTcwebONc5huXO
OGRwez+aoGI+I3z9nSbPDbBeb5E9pl9B1CIAgJSOG8pRe5OYxwrv8dlrdWampczf
/KajwlQcrHwQAmLNOOQghA8YaZTO9hnpLrKpwmgSCQsPPH+n9VyD0lCAR/k9nbh/
`pragma protect end_protected
