// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
IG/34P28uo44Vq0K0vB39BrVvdHWgF8c/S3kiQLLKdg+xZnRlFl+wBPAiL4j8hLL+rd+wlTXyIDO
K1lCDDDAogibzZ+oOUYJahog7L3r/YgRBcAYEmHMmHaGd6VNVIcYc3gN8COdgm6oqyvnELF8nIlj
uCEpDgjh7SiJ5dDSZPBI4QLJso6CRMWdYWTpOB+WjyYUieZ0qi370hFs0HrAloe3Hg3F5MJijNZK
mGM1HURHmR8MGxoEMfw6pxDT0W+WHtx+tmX0Gdx9zENItA/XN+wjWFrgh2+W3CR/dTIn2o5f9PXP
5fbdYaEPL9BpGzXl3M8KPmALmH2s9ZC5s2TZJQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4336)
h6GSW3JdzqOtMjHKrqkFyVxJfvXQwmq3c5VpALpalTYqfpteSK3CbBO1d80UWBhTwOnAaxV4366a
M5h+YM1VoMh6YN1zhFPtezjulg2nEUFKXp12VUZApBojt7dLGMiCKXl4pQ4aTquSrjHoMh/yToAC
O3lkqtmWJ0DT2gE96fJKNnDikooZGp5J6OHs2yVRPn4TUI8eGdZYulO2JXacQjcwdvQguJmnhewg
76uutMc5mpsDWHXBNzejvm26xryh4dMUto4P5+sKgNFcM9/RKDIDDaB0WoP2GU8N/p7O6SrAnQtB
6XDwS2WEERO1RG2iUbdi3gdH7rEcBgLF7rxnpnLKktqG9eOy27B6ZYFZly8CTrBqTHP4kwS2801b
O+MiKyoJRp7dHlSdnSEMnmbmcHF+PaR1xosn1vvg77T5jZBtgfbKfCKjx9Z9pc80mwAtA4C6avg1
n2uIfEKgbEIbBjk2wvVkXjwvZXGwMIWvCxMPSSuld465o6vz+i2dctKqWjqygTg7h/TFQPX6KDV2
qj83cWnq9P3qLvXrxOcfthKkvcR603evV8couqawUULnXsTRY1mUAeLbhlYkUKNHUrcEdU2zecUB
bvy3qMwAWfdlktctygAenaI9AN89D4URK7DS5B0tZSQuHrBqyxmyELO7CeC2Chrhu1YGqZ7MiZmV
jxIy3uRNOn6ZPOtTryJ0AooprrODd9Y+g2MqWnLwnyc7vGrEBhRxZ1xWufVdZf8VBacs15rsyVvA
e/ogH1fjqL0s30Pnh3un6tIpICHeAlBT21IfDui9DzZ72AyoJN6lXWLRRc2lJrcuz5Ru0YkAT9yY
sKsvJbq3Ntqq63C+8gGl09mq3XTe/3n6UQS4OPWiFzONrsoSZXOnQTFl83vrlpfiRihyo53NyRUy
fcRLfUrLzqlBEBkIEHbijfmSAanuE56RFxUcOWPcBm6TUEZ1kIT5G4zqsbvCJVDZgnECotltg5KT
Je1HvKCHuNeNdNX+V2rw0K+fgnXDlIYxvjYIKpXH7LrLaRQwREc+Gws8ATgRR50yZo60x5wlYp/J
svfLMNFb1K/uIlL6B4laUS46BxoFur3IT5RVB2ankhb2U58nUhnbYw7Ph1ejnPvQ3tYQ70bpLDJG
9FYRLbbao73OageIq4t/Ftj7Omo3O3yR6jQcyuqUav3qtj5qSH7n7Q5PKZ29guE2khW/31GPcYLJ
GhRKBKDQSiRttlDnC5I7MzKBMNTJS0o1sbaRrX2F98bBmihxt2IE8eKYdvF3HtE0s7t/HJXhyc84
PhlcD0OKUdyflZqLKT42lVcdVYWkuRMctu3k0sa4uv+uPfaSlyEqWPXd7D0wXWKtjlS9fPzJe2k0
yKI4MjIj6k+RZ6H8aXHZ+QTZhKBsmLwSV7CoErjqw9Q7wcr9RTDIcqSJWYK6kUod6GuBGbpYkmIm
jj7ZsvIyTBkl1AKQ3lKVNM1ppm8C9EJcoGzZydIagcyIbrp7/RLSvtj8Qod7L8vr1hykgqok9sYu
vIDACfzYAzRt5Qr4Hk+fTmWlhpA+uUUi2BY2Pdvh6oWAArX1vTj9Yj4Hd0xNf4ZpX1PFPi/T9HSf
qATU/GycCOID7EWzQRu+OVj6zrPSizViG4KYKJb7hvCfCPpgnfeT2/++ME4DMH37t/WOXH4xkkQA
n/RREDoDqtzdmtFMoxZdM8Dz8P8vUcz7TxxgCr6Zed/Z6K+P2dfRZX1pS61w40QvPerthZgVC9mG
L9nrAztA1LsVV+NuRdReEAMfCYJgOOdPQGGxZTYDPu9sjdMZc61S4HTIVe6dskUFuqO5w5NbAGy5
OAdjSz4115bEo0Um0T9dkbmTw6UDyBWDyhkwlu7oTjyKMZ4+Th9NGN6hg6Lb6Bs/mavsCaE3av5M
fCIAk4g6Wkv3q2Xw0zq1i/IM22w7wBgk0sde/kJxPiukWztpgLQDdh2g+ZCE5h+QbVy6VfKAdOPO
tmo0xQLtjTijsL4UWUiwm+e1mSDtgNOWMU+78zoAasKRt5bLBt1jC/KPjNabIN+oZtoPsX0EKam9
71J/sQvGk4MFx2Lp+tB56ncQvXZrs4OpnJLBpCELQ6+EETDI0Y8va8DYluX4R8MwHgHex8qaUMMg
yEnHy03UYPvxDAKPBLSON/SABTV6PRzzUAOmt0PR5JpbTbXTPce+87q5gQmcQ4EzTbunBh7qiZed
yEDZSyMQv3LbAonid2J8xSTjcCxYrH1/BraJOlYXm69q5NRRkRU8r0K/PGdZpZ5IolGUENiTVJOF
uY42I//jwAQU4VuPEgsHkMNKdyfnmrRLl8aMahTrnxQMENI+hGdPp9rjpDEmKffxrGV3YkyAO/Nz
a4WPRhKRil3UkdtsWh4MuRRjWWKaXned/DbmCXhI8fhHKcN5tWW67juX6eSDfmK+nYrdHZVZMSB5
AVusiX7YvYqabuCV//TFilM++NBfl9EmMN2SDhHUpKwgMNwCLDl3lfwHx8J4DoDy80gIqNq2VYlM
UMMCfnkUwkznwWbbJQsgp6HoCxQafkBCga83ZxGIEEBkWBR6SmhEgpyTG4JX45Bot3DbRj1hSGxH
OfDKCqZ9wGWDXslA7KsPm45LLbKRfvRc+rRSSyWUZCZHnmvANiWUmbeGGfKc6FMyBHkatDjf0h79
0YvF9EVzdHoNbF4n+7Ng/3JFIrdtt3a379xLfPemxhiSZ2wwuK78/StzLUNcYvVv3XaCsd+htYrW
D7xe0mWno9FFiKp5Vx55lG0rch2KyI0ExTsJWjm03fmBcwpZ4kCrs3DKRLknEpJ9R9U7aMb2bw0Z
l2ACo+QFbWgycjJ+ipiOcwv1fNAOluQLM9OPGSa+Fh98pCsYCGDjPfGivPLkRiOwz+8aINbBLbJG
E9a3Q+jElwT7UK0kG4vu/eWlRvQpVD2DfsfADrTUTGhlwRfRxLTkOP5Q8QwcDBa3GW7LR2iVH1kX
tdwnfg33eaXp91v7fIGM7J0j19uPYzO1cNqQQfX1yudDbAvvZJUrRGh+Y1xEJWCQqYKJ+enrRZV1
RxSKy7yrvt2U47IdL6GgYlQs4uZUOAEBnJsmwuKfDVe5Cz9vj9uxYTKVxpxyZ2K6fbwa9jTbG1MX
t0UPxPfBOwJRUsa440z8dS/ytul2o6zODUwDIBHpjAg+cXMPVjkktevH7F9iaO2i78tNSl8AR12v
PFcbHjg6fsuVuC7pLaTYACc2oM8FIY/6rO1EFzcLZu1cdQ+wesmTBybHVnOI29s67Nna5FRT+/Mv
XBUIWMMcDr24c+kA7R2N2ZEsPkixOrC4kUELGSUnt52A9NbMYyOe7y5qQBMSBhmgBTOqbkbReZhW
KvVGHgzDBkCIx0+eL7ElUTGBtq73OJlS0/bbe95ddZSJ8Q/WdXb1FlfzGP8KnCEUY5Nbvt9KRw+v
6HpspcOf+2pokOvXS5bYvKB5AHZOPC14HqwUmA3pfMZccofipN6QSXDVukrih8k/dkDKvu5APYZx
zn57Ra2AYA+kyHmlecWNFp8BRd+Q+kquBsYXYrqeD48arn1JgvtVqUoUFj2b/uwA9jrnAsoOHXei
XoVW27TO8e65io5nqkY2/l3mnYq0cmfLtGTUtaEaL0R1zoFKkXNoWbE9Nm4FLmr4lcq7j1WycbA8
tossY9bcRBX+q6P/sdjEO1/InbQ6NoaW/k7kUOPQyE580lV6oDSGxIqLZAmD9WZm3i+/6Raq+OUv
xBVK802WLZzVIaGrVXqztfp2qI7l2B7kY9UdrL66qhfkXgmHKnrADbbhLSNpKs/zULBrvxC5Ea4l
gHdcRfD86v7KexQSe2inlLLaq9swMNQtU99cEbr990x7OL36WulvR2VLj01smdltZiQDhjtt3rh9
DXd9UIl7Uj/8Rh2yLTo8xnojgxLEBy4DuqqM30Rh4+vG8yvNyW1yv7Ru32Nw4dQVAPodgyaa0pu5
8E6UutpsXVDDNH1EyZuaqCWeNs1bB9C+RtsA/PukDc3Oi+HLvSy67HT5A4YCcvkCPD8we3++/9H5
FamviwcSacajXnA95eTmu8Z+3zRxx+PIeAHwWGLNcEacsQXJj7yC92jZ7+pkUtywHh0291U1dG5s
m/yUWbSGVL1+rM5Wn2FMlUCnJBW2R0cOHYtHzMmgKQpIl49Ke46TjK43lqBmyIuJ0q8Zlpbno4ag
r+5NVfZ94t8xBPlGLVhdkEdMiaPgylE8fXwgDd40mczlGIrcTAdlQQD85Ws65CaTkoMoXD0f4E2L
hcY8RxJA3Qb6Ryz6dCjbwTM7WPXP/7EViyYmLoSCEt6oeHuWvcL9PZ345B5EMWeshkdCR3lL2qcM
IKaObTMHvdz3Pz0G1hoah68/ov87w0vSlWaENK7Aa92HrD9UvpSLxyIK6jF9psn+PsY/LpGr8xky
erx3F7wy6nVAADCK65nPa05MLjDUVoYfTZoCCnSAfKt5R2q2hCfJPcZYUaahhJ0jxLxnEpLwrQQl
88WaUrtKCJF4M6/Cq+FL3mcRXqtJ4vUHMgg0Qdw6hGD4UyKjp8ooXWJ7PkJeRekC/I3kg8ukYQaP
8cuA0V0p7eojAl3v8ikIoPtJVRS6kcSQUWK8pXulQ4sXbJzeLoR1hASamX00ES7TSu/h48fjkY/a
TBik41Kuo4qWLra4iqBWtpeGM9J14rfY+aAwHGzNF6zX1sYc+hPN5ym53888qZdRRd2SwXdl4RLA
Ujr5CHzk/8hMF7lPMlSeCltXwk9Bh12nY1FGVe5AsyZtkHnVQeacYTmntbQzqy553cZCXBKPfF1p
DvmCcHKJRrJjXSHX7vf6wH+/oDmKUhbo/rotCBXGgvtFVrbO1kU54vCGdYWuRbPR18OpQtuYSpDl
xtQhRrXkl0j4tB12yLPH+F0HPGkLcok6sajQM8OfImoRJP7MPDQO1hoWGNIdqDwxQaawoHJGkqON
yMvXUCrGTQRUFQMKwA3Sn9N9WlosFZqBs2jwVbzAGGMJjiHJR+IOLCmoT/59VqNNamU4BUm0e+nJ
ILINw4bOSidAVGve3nNF9t+WqvON0LW7R+4aIJLacyL+cyVXyykdEvnWXex3tfD/EB+6eYvhlboT
9N2g8bjPOKoHSOProkV2fwBVhda8alwMBmPSk+dB8FByEUTkbHks2zos9XL1ryDL3olQIi/bG5hw
FhvKIk9EuhQbz5VL+ErqTTh+v42zAAL9AIvIspwymoCCGbZCPQUivaqzMG0tAdWvGS6rNPJOZLKB
3iwTSabZ6gKCS9+7uQrdHu3q/hMTjg+XeF8h+T0c8he2L1z+wB1JBN5On+i/Ova0rMGbloEl8eRT
UsXqzWIYrAZAgwErNEw1Zk6kTn9nMWaEtk1hrFsv4dI4bO5FOFSLsSy2N0GHXT0FGVaOJcZNx57i
XNXLB82w7jeoe24r5iPJdhBIWFCHqJmNvBy917b2lYZfDPFHzGgvZgxMhT4k8pbGfJTwPEFe8Atr
skhEJubATwia3h4VsJ9mxRUUixe7tFkoqXueHx37y1IocHuBbUk0VPhAgyDdvDdUBi1NR9nkMTV2
0oIwYD8e+GqFnt3xiW11USp1HOySY6nUy/0gkDQBbgQ/VmNm9uX05Rak/9i2zHOSOmreno2i2q0d
6nQIdAGXtiRUpNil9Dn+Nxobq+ev2l/2s3va9popfHxNQcZZKoHbaeBO6JdVW5pUIJKNgHNoTkun
Gs27BHStB8ppDkJ66kIY/zG6eHIBHhI2KtcdM8UAlFHX9iaILK/CoyBwQcFOmgSsOYVonh6MjOWu
UW9fMQ==
`pragma protect end_protected
