// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:20 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MhdbUza+yrkXrlpeM7OJC94IpwPTXwH/q25HxQ/54/51Fgj/euvMZpq9RxXdM8/X
lv3sO3c1bG8eeclmNKO0vohV8U/Vbyo9TYMEuQ9Pj4eZtwPxeiCxGoCLZu0EWoV1
5W1JjLPERcGWaZxddGT35r3guvyff/ocz8uqviUekvA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30832)
kCf/9nGEQWKrUXR9CdE+JPdSJ3wgnHdW4qbpb3FqsG9yhf+3li7vJgCgUxptpXj0
CxaIBd8OM/FazGzcwI2VHVMQ1XgQRWKi4QIRpr1oj8Hu75QEKBUdNUymjXso0Iy/
XAxGZwewV5Q+ru5n0Qp2+u6jFjN6BsJ1jLTpauYBBcxBhpK1ZmCFfxbwQsEEZJlo
jIkZ7Efm991E64i/0Ide0oD4hR+BRh1B3+lCLe39DTRouhB1n0gOVhUagjewbOop
E19wzSO75YQ6y383t2U/rSaaejTmlTFNyZjz3MVjWQa/8M/rT3pXz0zCWfxeEf3X
WdhVgINfVlgPGHT4a4SewUEq9UcusGv861F0xciYd0x7C/QiIT85N3McUOfNAIIp
dAxj9agM7W/O7tUlQ+tzzaa1Dl1lA3uyp6ReSAIsNd0F3M3Fhf5KHpcll64nj472
KBzWsEV1vhL2x81ZZ/acKKs350RxhLYDcVzewnpYB880NdGf5/9vSVRane8w5pkv
j4URrdWbl8S/0CTkyUyx6cHNEDEz12AOc00yAaWM8Mpo05UEgWflw3tNk8EPoqNs
xstwGMLbXSGidZ8xcrEbIY/BukLiiKzw0/9kIor4YJ/A0kv+0Hfrr6/lqISd2glo
SeH//chjDzLmGNbogp6MOtBJ1CGE4eLDvZg/rNNHW51n48bUNhoFlVD7BEYByPIb
lClo6zd2TQg5mAdV5JwRT/2DxWJDjFRO/AeKiQRC1QUOBjlgKUG24k1MVT+9ylSg
5KbDVVRqZTw5Bpmxcm46wQ7pXjg3P8FqFlkeK1QRUT+si1CaWVoWresjVeBscoIW
bzDozJV2IZFZZDgaTfcYj28kb+YH5lZHXKIwUKp7WKQrnV2IDwMdsDhKlKzZmu5M
YEXkufRzC7NhRGoko6IEwJ0ZWTVcNp9WSxxqloJ7FITs4Xvtr23a71Ytovct+ywu
9VEYaWVcExkRuKM8GiiwbidOJdDtPzdzyGQqSrV0T6J26p0zG0CY1jGFQ9u33rTO
/PQXwY8lT0d+vhW4aD+LNfYFr8VKAkOW8l1ne3fnmYSXTwhib5fJmdKzZS8LL4h6
IdkjiwYVagLRSnGBMm+D21PNu8H78w89LPkeXcjKH5BXdbp+YrWFdA/Q3js4+cdS
cWv+/kSmqDdYsJg2Pu+nFbb/lqBL38DBM00OgW9x+2XMgGbA+4jqA5MDB18O21za
2EIBgB378JAA9mLuZHPqBHiHN7bTeuQhgW/vDt4PxKZqJuMWnf+yAk1WoArzwDzP
TZMLlkAcAB8apoGKPk25MJ0x6h8Z9NmWVNSKioGBijWjPutZR2d1UzINMOAAGZBi
5xjCclGfSCfC4PGpCd/vSBQ1s4haw/PKl0a3DEMR+zUjR5RC6NO/GIeoUHrRIKzh
/Dc2oKURCuExsWHLWqNUDtp78I7i9iVc56F+xQt5CeOfGJ77RTXeHPlyJcYFE/XS
PnqXbGL1lEsoH0T7O2E3VEKUxIYAmrl69FlXqcpBrZKwWYBaqDJOT82BnEHb157b
ncm4+qLCuQJmiXKFTId9VUrprcLvbfdZwSoJtzjs/R9PaX7m0hKo3JbnlOxEZu4X
NwJK7Sx7IQrJLfATzkVO+YYh7LX71kpITQqPk8pWrEnrnHERr7qlGi7EJ05agL5y
0x4C7HNYccB6AQEj6FkjHsfeUkYvJm3XzNj/gGwuI1FKbK4j8beCEWqlM9uErAdD
hFX4LtNb5ZlrAwb6zHeaDWKeJ8ZLhjMT1QjzHcNxt1d64gnob091FNi7DlS1FlNH
J6bIhN+sSHb7YeZWnMd2/Ww98coDR8BY52x+psiBnIqnLSOBHphdWoUdNMGQhK0D
JeD7l19zalBUjBMPihP+sqXaxvm4jv+Cj3CoWGX+PAJ7hD2KVlmZAVAG8zQeckgs
zq2Z9gdiJZ96cO0o/fT6j8VGboEztQnO37Y6dsJB/1xjM2EGx+AUojUztOQZc9PT
r4T/CnloxFg6fPtrExoNOaLKJCmT9arDQASe1vbYPvnbN00WMmrKlmpkx0zOMjns
d3nkyAHJ+l6+gmZrpnNB59+29Y+qu3brjwvTPUI7haA9bwMY9+etmwbi1J9Q6NCi
3GPpJMw0IEUZpoMDFQpR3/Tssmsxj83VyPoFpkdjIAnal689pTJLoGfveCbk2inS
UyAI7k5rD8uTfHrGPbr6YH7aZPYsBH49lzKTDfkDSMYSb1wC94uvny/lSqRRlTcJ
Wnv7rGj/Xv/3XMr8hJ34ToGHvNqwH2m1exJT9rLXC8q66E8Orxw+zw4foB7K9mpT
q1iTqs8QbFHPua5DwVRLOZTZcKch9RJzrqTBInOJU2N9K6ucbC1IVlJzdCTVkBBy
+qUgmvIznhcRUKBOOUiBczc5AbmKkoX4S0Pe+CzwumIdyyh8i/FBmAWn9+AOU+Yy
Rwvi/bIk1H4CKvZyeXh86noZTueAB1Po7Jxh9yVdBJzQzk330gzq4OSTwT2Yo54l
ky54sPPkx7OWNw83AT3TVS7P+ZNKBUi60xvsViqVM5PEzpwg0EN5sWcS13VMxb6f
0TxrYYdd81LPf2Kk5cNghIh7eXeMifQywMi18qJ63h4/mc9opB3fKad4BEzi4osX
T2PJOLYBPq5TNYrGVjBRoZTaP1Q0iJ96v4OVdSr28un5Sj060cNyjPmqs8P7syyu
2aGVtCnWc0JXJ9wGwJZXVbchJ5UbzR7h7g4gyRTRDNwzMILUXowrsfvjVcHFIgVF
q9gSsVnyp8mwykYW+jn7FgkAzmVKW+Rfth8YgH8X2TW94Kh5KcBImhtBdworw6wA
Ei8JnK8RgQYzQw30pLT9uZC2s6mFDp+lc2qPQHQG+CgMvT5afR8Ouqi3fcY5VPjM
SCX3CnRKdySJHyN/xSrKH6n7R04BRvfJFEsSVuUt58DQbCjpIK+u+Vy4S7YUwFI7
kR3YhTPss4v5wGStpeznEpSRz5Cv2Ipd2FaxCCFxm9h/7Pwc8WOrrSukD7thKjSC
1uAveQBFpZPkXnBD9aGsKuQ+shdx80ZSkH9R2k+h4eImSWqsAhLp7a/UwNIG9rpW
WV/wZHM9uJEwMwL2jyLDlp4Iz7ALeGVe4mOlD/1+2OnwQsBnrqeO8kdggHIPzSE9
5BWFzI3uG9K5Zs8Yi9iD3osrwqTx6wlO/9gIaDe3h8OMI4Is55n/3v9Hdc+hgWpE
fxDnjAQNzG5ugFdRDCwkuBnuPsh9NDXgeSi7tcpn/hpyIWteO2UPSosKzQ6SpRWD
jPISLs5s9hwqxsMJHYmm1x4S5HkxaYJGdiqpWjvWiIAax3fcXfhxlg9SQgKpC9G2
g7IQD4TSuly/Doxcmj+9HZO4KvoordExLArHY8yHPlAAT0j1zgAlGjZ06mJhwagq
4kbQFidWRorLenC1ssEOB6xYLsjhQsYAqYlco9yYGYfcNn24zrWTFKVrNNMhXsAP
LOWXVYM6W478AQpfUchCN/GWSU4qHDNhQZglvn5MaYrjhBpK1Zl8NAt+e3MV5qbU
2Qu8Jsdmo6VPi2+8Sgnm9suBsNPi8g8MboGEhNpnNjA/94HoznNCI8ATq//Qdmc0
c21So/T2aEU0O8Aa7Z3+QLh4zC8k2FjN72a/El0DMR8avOYYTFfUItxXZ9skEHUU
jY2B9tx8CoizZxiH0Gb7/YoqEhHz6tSvfYl3KS+5Tzh0wcMU+J8JUeC2oq3OFLO0
XzqvldGx2UIwo0Knbpgsy29uOzVBz252UUIvbjlQrB+Q5L6A9BQqyBLRkzwboiLI
J/38kYpJcWzv8JKczKWzOEC5Bjkh3xa9lXlneGnjNoYVNVLqwCMsQQ068+mrWxRr
BGwW7dD1677L/AEzsVnMyjn+RGNmjxszEub91TBGcOGgXlv7Fhl1j+5zmmWcXkHh
NovbQtstU5AqLf8UsdCyrPsLMARrKYWbq3+ZDIzHW88DXgwEBZE4R3s7ehJb0a+d
EOgCnuSXX5npO+Y4a2M559lNAndOlfWmtqMijSsNqMu7LDip7yJk9xLNMd1WwA6l
HHIMsIon4MztPPZcM4f1UFwHDvKOu/Po2hn0k7wUWdn57EIhgcvjHMsaWvwC81ya
kw0aIhCm2qyd0UZT/OawcAFZVSx4PbKjEdFh9jiL/ltM2S57g1ONmCdEc4GwOTwD
WsDBo6WP5oasTGW5Yy7JiC+dME+D01TnTAOakIFsRrM3aJDPfpEwqQMOevKTG05b
jWPREXTI6OjnlhN5jUmvSNmVCc6BBAujGWbPFgNgRjCBIUlvU8psmbOFT8Cd72iM
RN4pyW5Tk/xIo3EVbg7UeL6jqt++gonMh73CUhofEQGuVpzLhhSxgDbl4UrOvogz
T4RPCxhL8l6UfFVLLuehdhzpkDfxm1cIdh0obApu5esQwIOgNLitZB4MQKCTa7QH
IuTlLKiw2vsyQP5oDiO6hDikYH31XxlWPRPDDPcVDkOu+ra3i/TbFqhbpuNrfCK1
zEbL7xN6pEqJpG4Uq8F/LaMQcME4l7YR6Q5aOruJWtRNM5boXdWGhY8W9utxQuBY
Gz26p2NRXBikVMPgdyZK8gFjlZuZ5P5D2xGPqS8lDnsaVFkgfcRhWTZ9dT+xwNsr
oc6hdtDUPV1DjPBfaC069I3ozmOjrWfgOUvQk0oATT6/WeD8oZ0rxKM1dq2326jB
GX53ENVxSp5zAZt7npIRYVxyRPcXCU99vCHmCTZ55cI1WkuLREy4yrdpejZcKfy/
RUjsqZtXi8x3TGciOfU0UgPjRLOHcL1GdsFb/MFsKjBLGnde6cA6RKyzMZeoCWMs
B0z9schjqV2AqLdWC4NJyutwCKZ0Z/DYScy0zqPEVNSBlTqo3ONYuAYFxkuNzWV5
3mgIOAjpiT+kSPWq1xjqa8Jk0JDfVszompBtjHjoYiASRHGJotXjQobLKF+u7L6l
hC1+rQ8wmMlUveSU5F69qURTMcXHhUnsG6rT8Khszc0+ZPOJ1kmb9pVIpw5iy15C
3aiT7NEE4uXboUKbc5UjDDKIHtuft+XdHVFOLu0u+s5D9YAXNNjhIKvxN0nLvmyo
8LgxFJheiSR9ecWaXnA3XXPOy65JZUgd3urSb+TFCdo5V9NAo8IMip9Bz8UGuF4W
WKs81DIcvd40aJBI3rilivfs60IVkaRcXH4NrCNZrllJ37SB4/5blkpjjTBvr2aO
58/11mE36ylWV5CsnpdZQteswABQXmHVA/TpC8A/sEV5nN7b0Om3OY9XvCN0tM+Q
JnhoujlZ3voK40oSLRQr2tZIMuhKODcAs1rf9jmBPC+6DzTbTa1VmdnN3wpFRDUo
t6g6xtsKgnG65/VFIMjfiGCJDaKgqO7UxWKKDFTP9sv5sHMiftOyifMFIIBRAcqh
nIpPVXtaP5dpKjD9K1iCU18TjHOFbTT4khed5dHuljhjJwaLGkerugcN+rElYHGK
bcDsoJK+gPTTnMhT50Uw1/Lg4a5YlmMBwRzNIybZLUVnpZWJ94igEYOUTL+6Tp0K
u941jk9TOwWXNR7bZKp0zJkjpEFU1fmdx6oro1yU9+9hKpnCqZ1dM4oOocjj6zKB
xDafyQgkBnr7NlZE+MhRoVQtNYvQsomdj923t4HePtDs4wQAfqcLOVO1DivzASKt
iGdzNTIM7d9LbpwEp1yMZxASajv+8y5XftX/MBr+UxxpkPN8wEuuMGLEYTL3z4R0
fVQWdmv2CgXJZA5wMibMfnOdrUt0gT3W8DnFqk1Ppo/FXmiu3YWj4a8rMdEii/2K
dCdkzyvJWF/5q3vMu2PoRbMrTjBAiNg/Ux9aJw6aaNPISSliBcwaGrMePHsAYPhp
9SzBeiKex6yOgaDaQ+M2ABSgKHgjZpNSJwpYWfFQdazW3oS+805SKD3Tc1Pl3i1P
LizfvA8NqwFjFCMh5pGbq75VU92fO1Jnth7jBia4wKYy8/hbRt2DAln6uVC033tV
49cAW2vgaAJse83ETTyvlY/aml/Z1K0/MsbfniqzMGQKNQq+uKVu8NqgKYSuXKm+
flLQrBWcOJ9XGXr6JyInLNvG1np+y88HCkrQuyi1vKiIate6KzzWZxg8ImOFJGnB
gYSYwsLcEeB0D+sYzDHypQyRK7EtZdo/pVRaE2tJ6WeQnqGd4jIB5leHKfIqUV9C
ay1Eq0DrCN5+AaduKh4vO/PRuz2y2pvope4NLqB4sWMAEvGEqkHjbu3+cFxKgave
fffG+j2SivVqDvmFEgCgLDYcHfsVa1H6QXdEa+AKbIrbRy8J5peOV1K8/8LqqXs8
LECiEdeEK1eEpJ+XGsa64BcvWVMaV8uQtcekuCtkVcZ7CQf1pmJNlB9sR95Cl+rI
Pf83z4t0cWuA2Qrna6xRRpirR9JTyzU88AtZ8xLsAx2Kov9CHxW/KDpn9wuf8rcw
A6UED5mVAaH1maW/aUMOYIyFudjnPqPvWboVE7SoyQySajaE80z/5YJigL1aQtka
5Kzj9/RM9at5NegCa64lh6XaSfo7XWi0T5E/nOuDd9ko50/Zuoykcks47UIs9V+E
Q1+nO/8HKIq0U7tbajbzVp0QzxYYKU0KJ6Tzc7dtjQy8YxdRGBsb6YoUN04t8jZJ
FSpLnCYcwCza6Cuz++sIRCblR+nGYFQYoFF4GhJjofjLYXaaq93F3pXgPdfQjhMO
rTqySbR3RA5AtYZIfb5dUWsMSTyQ+HeAGC2ZQA5wSKsPU9IjBvgj3vBphsAGXTon
Pu4GREJbCpzcihiW/g8qQ4u0RgL7NxHgZ/WHLeY1WEsSKGX+BfoPj8HaM2jA+HqP
I5PTVOnSz0W+mkUosvjDRsGZmxpyVF8hKPriUPKYHGgbGDsNg4ZEvWF701Q4yUMW
DadcPH0+gg7BZlrO9aNcb3WhN25SwDYGctLHVGGU4jbiqp4ilt4OICY228wxQ6Kl
L6zzW8geePsm5OfokqqhdLn5F8fenu7hikgMKuTpIRaGUxAgieB22qs/miqBaeGJ
YDPzmNqW8sayhFWfy3PguCLLiMS7IhAYDOsphvHeJHPKkMCZmT6ZFLBsIFEclVVe
lcGNBuKAZSkMNygff+aAMGPTTOzY2nMBWiUAQH/eC8Noh79canU5Np+GvsCL6g/L
UWv/zaK+FMI956K9W4pdIR48us2HsPGF6TMljSbGZR2iSbocRcLeZviKQmzNHycR
78LnMlK9aiMITg1oFalUSujKgkmG+HZrttxiUrA9FumhXBgks1fnUip2zxzaNWGy
HMsX/9SfH11FMb6Bk9p7red4pZLr8Pxxj550J9Rww6DueUl+zE0FsV5ghVZ+hGV+
sdL5919J+2kW/8nQuqgf0A/0H4poQR3Y200c0+7WBBuGP/AI9aWXsbEk72wKyBmT
2hAc7nTVnIJVfkwcIoztZKtoyr3AIJiAZsqdqotOtxuMxTa2HRnMTV/2yO3hCMaV
aC/yUncVASr3zydpIZ6lNqCDrri7lSZKZiYA8MO7zpDfb1P89oxcpdcMH8VEJEPa
s3crpCt+lcYYt7NTTYaZ5gHdrCNCobZikXVRidg6O/yL9hZXwE0IGFxHM6NYCf1K
jCu1d1PYhnpMPhk8wrTNp/jeBC47sf3Spv7qLu2JG+NpslqrB3cjQm6AkyOArK0i
Q8+c2rGW3SZKbKWndScbYn1YI0TC9zk3+6JgVpXPWzE8ewIMwr9VXQW8eoWWT+tC
433XwvoZrq7Dfzn+4lTrBnYujCuVKHyjX9goKjQ/H+NlP1w33/wpzWp2sPKaIVpe
4R62g/MjHhzeIWFD7+I2yQvqSBU0PeiC3ZeUhCQvt6+1s5Pl98YGkM1QIw8jWnPr
lOJQpSPhJKvXNWsSgd8cM4GHlE+KN/1ed76NarzN6ORxQjAb6VjxMQB4OqD7UAe8
HA+bPZt6QH0tyzSNk1Z2vHLqRcZEJrDHOD3IPwYpVlRp6OD/ryAdavhDx23S7hul
BEy/qQIoAir3VgrCJCOMuEQk4HOv3LRPiS3j3tUcGMrPzLEqIANbF808LOxE5/gI
6wWDrOnFIem76bDzUjzgddVNIOuZ7gqr9odwUWlWke0WJgaX1N71C0g1QK+YiJc4
+GR9Zxiu67NGQZGVe77IfCvHMXFgTUQeLSoKOBR8rmgQTYRuKD8e7mqFKEtpYJbt
X0hiTRg6aRB+gseVyKUGXdwzT65JxgBKIIWrqRDCQA3cMfQLjdPBw3OBmzqjUk2q
qao9d6z42MHl8/DEOMrPf9Gcy87YWqxNgRW8P6ZFNaXHMM3iZQE6nD/Gtz1i2EZF
dPo1G/CEHSoJ9Iwbr7GecpQ/nRje59zG//AGCv2Z8Pr3mIYIudYSU3Os3Akawp5G
+5bgdtX3cW7uVuHdlzk99bauBMB9HBGOwYV3S6eqX2Sz9RiWmBdy/pFzeVb3SP1c
f1F6Hyu1bd0VDkWhF6RJBbyjtxamAYpsEHV2L9qaewMvX9tS6ni8NddWJwEEn/02
KHERvvhlQQueWBFqMktP2caNVflVEuZmT83SbUZ+hGz5Wt+HGtP9/IeFgrDIjR8Q
iBinU6xQIhwf9izz2eYJguR264kROZLI09DwWfC39I/LgwN8ayj2j7y87AxpxVDW
0ecsnuAm9/t2fpoScULZ0+j+smxBSKX4OOU+o9KGzwLW0E/pTZ6togGNwiuV+Q85
8LI2eyDMOnIXCGy4R8A3gJlEspbTNuf27xYBXIszfDXK0zWpCLd6DKjQBk4qAHis
uksQ8dFwMHvsFWeh/jyjwCB3RHA3zgwdTTqKZrbFGUDLyHE4kmNJbR1iS1tclSno
jRAqgQqTKI1xCZ+WmFG2I0ejssDT5gUbtBDF9A9S4bJ39qADfBQ8pdzARnxbYFI+
Ebw5vwUUbfAJDvzH46k8Sp3W7EfOsZZRrXchZuvAIiH6laNqkvzimTU/oPlK2O/M
QTiMJe8gjimmzid+mMsu6vzLcMBI6OKxhca3zR6RpDCcvR6z7LCwCH8IDb3hKNG0
g1+78jnLXTe5Ue+4wGi7a+bR22pRDQxXi7U3fcRVICLubPjmyiyXWZffgeHerJgk
2npyt3X+GXoNMsOfPTqH0ZztKfzKNIFue0ScH1XbIu0nGycgM4TnLmefDSEGlPrt
aVILKBRNv5pd997sAjlpKZXcOn8arOkc6a62vJZQldfEnjpSAKBmnv/K/5I1CjVu
D3bO1JkR8VgxfKTxDV7XrOg9dV1rv9ig7MuuJNBucOKiHRRNi5lt/CiBNvLtRLr6
381ZmYUxqiAaTg8jza3RM8z0j8AaWQV0OJWGfJAiJtYf4+sxhPhRmxAFGWYIBebI
KyxUyyd5fJq5sxR1HQoXrsv7l4rtWgLCbNrEs03XAhOwfLqfXrd2xxfKVcATqVHH
JoacYsnjWM94+jI+FstJAzZFv5juapYOOjubrSTK0gLUw53b/GaM01V/nkx0Vhcf
wrrE1AGvpoJXlte+j3ptDBzzOIY6Jdp0GkSMDqsEXF151Mj1BbDsKBK9sgrmWEuv
D/G5J9OBvVWh1j6y08peuE8iQKvBW0/V7kqN/YK7MZkH6KdxKnLvnH5yMgGzSBnE
3UOzYRnxiEMPDrX5HlIUA6zcQQMn6YgYoQyI0u2tGlg9IB17A/bh8LHdnUHaaI4z
ViDdLXfnlh9p8OlQInvfvBkF4M9F0I/pIROgXKfNvss/0xwtVqDV3veUVgfVSij5
ANI53RWPyUyrb7c/KZGSgsJz193HTYFFi844KFtDr97jAIaEcXCa2pnZeNw00f7H
C3xLgCBawRSme92s2G7wDk9DlsGpAWOvgMG2nUnVOfprcyWsrITSavSPx5WRXY0K
iI3wN0DaWbLzC3e5KrUwhG3kHmFZyqwhRcxlugEZhzfTiUs/tZlGONIwycoEToKC
a2uYfOGvjoBAI06kMn92CjGKIc86zJtm+s6t0e+EJJhk9E5atAVX3oB7SYGaj8n4
M9KmB+gCNr9ehgq6R22TkA61EVyKeRzgdmxnw6XBlYO0SYs/kiBHgLwug32F4lDa
YK+8xzHUj5c3KpT8DytMi06291sbZtwTlwrOw3PBJVdvvCP4BO/l7EtR1VERTAsS
pTvqwTg8UYIukyOxVbcEM3nl/zxjclAiF37jZTdBMZcNiZcbHiGU+b7hOcfTwyYb
aqgInFPCh/hfVipm4TqVnzhDijtPl2VZT8xAv2JO/m2gFG+7vhWNhdacIZVB+XvZ
kcv5toJsNUFBuJ+8I1gIUyjglPOlQR11zvPv1JHUKUNDuF9TDVXxsdCfWu40eiJ4
1T/MZwnTDcOyMMUXOK2HocyM9Z7CIPZ8cKv/F5yeCkhYGo7EI6i2Bj+uz9Z0LeCO
oOJmJC0HCIZOvVa7vrm+2V8AIz3+5Fa73Eo2HoyAEpcAz2wgeBtY0XfqBPMngz1q
YKm1pgR4mBsO0M4ZkGzpZWXfzT8lrxZbQJSvy/YswiCdCjpMxL5f8vY7ZivOyfNC
UXHKGuPTghPN5nL52v6IMgEYmeIlY97V3Qg8kVIy46hn3jhiyfetHgKuuFX+lJkc
f5dOL1UpSJOlR69VkF6fD9h3nrVccWaQwiboNtks8D4frj+tdB3CR/rYpt+qEZhQ
NkIoPEHS7t2kMaXY2HIiEJeM4gbGos9yMkmWoaeDXSWL4QScA1UhkaqkSe20rORA
6CLWhgGKn2NtIjo4G+jzLEsC5evEDN4+ecfVfoUH8xfv84qHk8rT5Cg/8gXhdYzR
fnIUTRES+OVoppm2/8WJ3aymr1UVctY8AsZM+cnFUAyYN9bAuBQ8eTg5B6LF+h22
DbABLlapHzmQ2ex5cPxN7lBV2HujFFDhdv4eVzSnGDQWYTrAZy08aaiXMmEvyx4h
gLylzY7Jk67I+UQFUoBcfYe1SfqtqIZIZXPf59zdY57f9wUBfze3baO21huJNay5
Q5yAENOyKSOYqwPYNohFQm43iL6fSnRrRPCgCck83n68sSP5e5piI4ABxNMJ17X9
+ytnVC9em0Q10VDSrSSEnEt/kk2gRpXuU+LyDCaO9iDwI5PEiIX0PKQErAA9G1uZ
4sZ+5Yf5CMQuTL+hDyVVc9EwsvNXBlnQMGBlvYBFAArwos12NkttLtOzE1ZMknuE
BBIU5/CWWoVdbww19w8fj4rUWsw6oyN7pgcTWy17SRmpVIsfCUAdC+LbEHtezm1i
qQD7eUgwidThty00MfbZA0G5C9zIhWVo00D3fjBvd4qmobEw1hyE7/tzOmwwYJXZ
H+UtPkYZdb+bs9fFBzk3BR4jN9RPkI0YDJ2o79i+EI6bWd/hH3hyGHc/BvkKgxKt
tAhYoD3/Uho4DlGLs+VNjowc6vCLDXtHZBbOo/p2MwZfj5+w/ClnCLqRzKieRpwQ
XeQUxAr9TGxtiGsuhQNldj17GCm2WYkVMjeSSC3k5yUr2r14xGX7sGGL6z2FOR22
I8+p1HSzBoCWRawlO5Z4dA9iJRkQHbacrSvwdCbCDWbC5Kh2CCKHyt7iXgBxT5G0
JDXAXHtlAY/R/GY7B6EGiu0GvmE46ryvColViDNpOji7Qv+IugiofQulVJXH8I4i
iIJr8kMHm1gtojZFO0j+GfcNL8LBM1qxDcwYb5jjY9EsxHWtROFjKYCAtIUXahaM
dwZhvUxRL+VY4VtDdLk9M8tF4ZI6ETIZI/BlkQ4l89D+8vi6pMcR/IXbclqO2S6A
ZEmRlC6ELeIskhK/Vikf3pfnJ6WtnUZi5GWnhJa8+0MIFLlDODoiY5AJ+bF/lnpd
cgAATfW99/UWPKK3Y2oEoNlvAKKM74JrRPKIlM7KQuKQi90xKKEehgjQs5sK+39l
+Z38OCu5TxEZ3Eneq9KQD9wKTZM+wPe+B2rSaBUvVexXOY8AH6nWpEYSpmPdcy8R
EFhxVjwhUht5cjSYxcfeRJziH6yb+1Njwk9ati8Wlr+0g68lFXQfqSZG/nuDtEpo
HJParCPEsqgimvVlpeSjz02ttYVNmN/7pk2HVozK4hafMQKQtvVvX+MaboQ2Lhk9
bVcNCb2u8xCxR9cK5XwYYs7zOzRyR7YQP6KpW6/Oa5oKGIIhIMK1WrWJvTJFvttw
3PuTmLu0sJ5EkwhUlHbg30vaII1FWN7aYl0c1QSmNbVySAMQD1ImjkFWNgmjPRFb
hsigl0iZYOiuj5CsZ9KKOti2QfgzWJLjkCuwMGIZoI+M49mAeMRq0YVe5HB7+Fsl
noAKM3zTj6eNtfF16juofUVpPq3G8hNHjqKgvuemtDre6pze4h3UzwXKVuVP9og6
9hhdtEik9TSyOkJsT3PKJAXMV7ceZWp+fC8btwZsk8eK7I68LHc1MB0HiRkFXR3M
EJkaq9RMqoSdZEzzG1r+jYs3LxUi+PZgbax7Kn1UhkG9veV8Xz1rGOUowlgYep+5
Qk5gtK8jNsNBAUZJdfW/hfsM8wVSaRzo6zkYZyOmiBLYYNDLPDAO4x9ciiWmacSy
dXZ45PaSHl2Z/cm7BzVW4pY9jBC38ZZOmkRxWZm1Wg8b1lXN8sOTNN0nOmqepU9p
yV6jLcaS1HUHqN4kvXHC79qFGf2TIYI5T1O3raiNYswH83vGAPU8a3/qD7uCcv70
vZkLjeJ1kgUk9nv9JSMKg6waUwX1SKydvjANbEnV8v6W/kYRqTEmV6K/AEmwFu8/
8UUY/or/a2ICACYMmH7iE9FgZFhNjVa/4qzGNpFYbg03BGg6jQ10L3oU5YDxGLoa
A5VAw0JVYKOJTMDYM9h5rTAQK1sYUOqgDgOaxjhY0Wg+2GiIq3xQW02n0LLtGpWd
QEmT3SvW3KQXv9lFSUwQok1EKbv1ux7veqm5F+uAUJBNETPIK+Zd3vbvErH/rUTh
WtuusLayZ4OqbiKhuK5kqC2Oh49RCL+zs9NR8wXOCnJEP3TqEOEt81n7dyGX3FEJ
nRU19Cw00yuv8k0JGWpNwGvnDYaqSEdppJPsljyvy2eI4GWHkZl5+YyLjwutQQsv
8CUwoV3ejYM/j7ulOh1jcIzrCrst3GIGzcNjqt2LG69XdiBiqI3e8Nmc4bfnQZCp
QuSrANJF7PSpe5n4dsGqrNCsqiDagUbxKPF/hQFZSor8Si90o+CVFohU1J/X7A2L
jRmYuOK2mIo2IuJiZVJLvIZIj81tn5qUu2lCq3py00tXXi7ViN93CWYOMRlTuygx
RK/8sX38ErrJKckYJN0tmX2NWOOZdEH1WbJuuDxDlM5RsrFw32ekRg8JenDwTL1w
KsGcB5iXmJy8XHUGNE8f9DAY1u3W7dNA9as0P4EJkEqTPpp52Z5eSk+wUhOhu0aN
dNszYySr+CD2HgXFAdVI6/gGhE6JskZRbzZsyPGu69pvpHCZuvwaVIaU87/1XXPX
ASDaUB7yd1b9huSkEcw1yp0aTXQOOwFkYJDSzu0oOA9FSg/39JPW1KXLHwa8lLsY
ww/u7Rycqq/rNg0YiLKw1hKkPceZ9AK9ME8utGmP4GDOgUz6y3ifU9mdtkD+BSGl
+s0VU8uGQGKZCdsEHzwvk/9wuzfuMpJu+3ZXu3h14QEnDOQ6TFbXRM1PuJmRsE7e
gt9O1Yn4COzVwvHWToKjdxVYtSE0sTf0wVwj7nAys2MNZ7yhhhJU2rW3z3S2nYHT
jf8XeLdN7pYUs5Tpk9WjDp4ENH3m3tlzCUlIXvY0fzwfQU/RpYdVvk2/pFPjp80c
RW+TsHVYuwNjr2EeoAZ9bYb5Cy9uTWryj5EfEIWQT+tzJOlzNGTYBls88w/xivjz
jpQ8TsVGp0H/zqbf9XaotrXWiXuK23yHvJ72YMR/KI35uxHtR6zWGtlvDt7RPR51
CzNLBPWSEXdDo4Z3mORV63wgezP3GmIL4NXem09bjZ+n7DCGG7zQM0jeN1Rvi7VD
Vn7nlxjhgsu7O87uZ+0nsfTzCO/f+6uybphwdv6yddOEkdgEFAneuRVpg4VXTE54
u4Tk1GZeC1lYY3sMMu+fzQkqMsqEP59D6O6h7tuFqh0Rta6IVCBpdsrXWkO06adi
iWiC08LsanSsPDAgHtIPZJi1g7EnUio0tEjThX67Y0GWZFM6omCiM+hkOpNAJSoP
go0RJGtD1sb0usbWbSEDH2XuXJQCFDretJWh3ha6ny83DGMl1MqHOCdyJ2qc+goE
fMFNxvtt4MfLVK3MXCJyqruJ9EKSorFJKobcypYqcv2xPTwngtWSx3SWIDtZvyib
wmnBQA4XKzIHzpsNjtAsqNnf4sNDa1H+wCYhFglOXGKGNda7deRgUqwgMSciIePa
a1i0J3mC2CER0OsXhfSElUD75M0yTz9DwPDCrMp+RCSiC95MfjU/9DA2iiSVEXEs
Oyxq5odhqB1Sgxfy6/IVkReEOwTTFenZE8Z7DGNUDM7yF6goNAh3RGwd+ufWU4Hi
CwJW0dL3gxOgmMVUrga9/N36tvzxUGXY9zB3nZpZ4TkHU4N8tLsDEKIeV6uPBbUb
ny6Xwc7oH1ZEIA7xj7nQJD0z9bJhabHVNVDA5QlrGOpTF3yffKU1xdUwQIbg6uhs
MplJPXen7Odmj2jxK2qdE6jKBqm3ZvFBIfcNxcX+Rg8xwoy+Znk2TxrOFTAMlCDO
ZRI2dEvRydiKLugqqwD/SeazSKLu/ZLgnHfEnk5oxGKcDEOT/3/XsctXIw06Hn6Y
WdqnAsnFrFrkDLyZ7m6eXl99o1vN0KI7zQLwFLmpmSmNyryS8w0Iuun02yuh0OPk
T4dHlekmk5k8vW+9//kGrhiGlqZTSLcEMFEx3xWF8v67duDO+4JO+rEDI9h7ZOY5
eEr6ly8xduD/U0f3gUpf8QIa6I2qNWBpVMEakQZ2t7LsV2HfvUxDiF4+pKPF0+OH
5UcgS9TGoZwqcsywgzVukNpnRRHh5kOGch4hUsH2Tinr1fn7IGQNotk8JZPIEXPZ
JKZpFUd5nyozFj9bfQM6vUmusxIL9If66vzgo7cnB8K0LZG8w7wVpwzCHTIleyxM
TTnDhb3FcW/Qi2T93i7OVyv1jkjMsT+3bWct/2VN9K1GY84fPjoXXjqrRRl5bzFh
Ph0Ilf+R9NdwLMH99CVATKDNW1BqWrYWhCZTiP0/hbtbCy8RCZ8gbDwLBlrVkR5z
MomxYtW5Qgej9dcHi+/T7oBW/99KawcZa6CRNUWo6fBQkYBlZnilh+NfqNjJ9zgK
gyxMK/UtvkRIajz9cb2OU2+vbvyx7dvS76B0Vlu2usuJdpD0YGY2KbfhJftvKztT
AHE2+/YBakG7fih353bRrpSq7bSHaWHLTDypbU/etjLsNHdjh25R0npVjhiltyPO
JZ18XAH4mIAl+o+iOdWQqzjUIeQv9BLAnYKnCS/hWhvusuLudLSg5HWL9t1fvt8y
lksnhW/FFD3kdx2kE30sMfAq5FUxDXHUx8CHQK4o5foyfnA9CWz2yJn7AcQ5k4O6
mAgGQ7G/INpK9XZdAd4rhx6JNPvZBI+MtughYP5KnbvAPgmt0veZai8N7iIoErvp
bC+lrHKhfWobbek+nwt6n3xtC0617ODFCkIOREUSgoNmiwybe4/O2P/y55Tb2oaN
sw9YA996vYyBO7ZGxhRqX2xxxMGPnlD5dlFm/iSG9Dv6K3EK/tASBzzm353CGCw7
VpbS4oMGAc8SJEnXrGrbjh5yx8Yf8AB9pBaR7dd22vh90pWVg/LKp0tadI7u2m9J
YpOiffxqpE0yLZ9l3BPgU19taGne8WfLzywthhRQsKqwW99gIA+oTPuiIcro0GFw
dY9yMMZsR36eqhgBIcqktHyjwS1GiGJ9k3YsJgpidngu/6MIE4D0geQQpDjIkRvr
Vt24im/2pX7QDzOSVoG+j+KYrg+cnMbiV3ryyIblJf6mKWgN/VFhG1mz5quYtWrK
uSYDvmQnir2K/PU9rsCmL2MwqYTetHn61Z6KOichBiDGURHbwznX5NrBXe0I4RFg
1HogBz9IHNj+qlrivBBXrc/avYXZ7qmkhbxNtaOxF7IccN1VEyCEWvJ0SREp/4Eh
pP2JrLaDr+7vAg7f7UNtVqR/iXuxRZl6xVbLtvJbbD2r6TEJI6D4DjViSA4fvdks
HSWQVxowXiD7FK2ifHWU7R9AT6MRggXB3pNfUt0qBPiXTLsrhGGFFtNX67xNbg7r
9QfmW6xhnF32VCe7RdwfxJPPG0RJzgLyl7Rhj7sR0+CuOBwbSOXMvLerxiD3utA5
hSRxLk/64mm/KV2/LdLkcOEEISbVrHUmF+DQTNo0V9+DA1JRLB2SOFPKsh1/h99l
7MgUV1dBGKtxNBbrjq9PJEAjDBP0Ehr2ABFIdmhS19D7sjYrtHAlUGV0CkAV/z4V
8kXDOEROf90HHxBl6HB87fvBaxMffBRLfM2UpBv0JUIZF5Cuc/26EBIZ5gW6Su6t
++FTLkFfqraEzcitIHREBhIUDjVsFjH/xPDyhlQdRQSV1AThMMHK0n594kQOSuL0
sT+hMty+f7pujpyjYbNejP/8gYHDpnem01cDWzA/Glwuj7o9ccCZOqls0f2K6Hu4
ypL1sUhVC7QdMy0WrlXMt3YFG03E5SiOlusWVvsCpAJsvabECdVxS/VpIRVrAimj
Gtu8XXRSqMkEZGBxqtyVoqNGnD1aHT+yotlD8slqlIYtJPc/Gx+TKdFLxSHCGteD
pz4wo2d9l6CGeGtwGVPHhwQX5p/Jy6Dm3/IAG7gBS5yKwJlWzBkLOf+vDLQeclb0
bsmHJKuAzG4IZVywtW+darrTVUk3fEWk9iQFUhs+ZAeCpAegDcWYWn77a/S6zJze
cGcOh5ZkXPTmjT6m7X22b4MmY5s9fGORIa2iGJjYUJwSxBEz2ydJL389DNDuIkLW
4RUQlS/846MBuOeqCH1sGISLaHcvidJLbidop1PgSHd5nTWPlkIlwvbdo8XZjrWh
z177US+DNJHeJMYWKP3Bv3JGXDqm1JBpBXbI7HHP7N5XZ0pALS/+MYZIkmTqibiy
r52EycGXIsUdysO2Nik41EEgExTJwfXrPJGi7DWHsHZxKzVtPO6ncazXS80n0n75
HMvU5Rxa1E7lBYpQlVOXSfBjjgqAG8KBwAeq27+stK5BrPGWQYoQjU7tW2krcBiC
0t795rGfMI4vORdC/i47y+Vr5m/a3Idzi8h5Y6SxLGmhjax9SKGQfAJCJGpPsL1j
fE4pOHJY97OVhE5JdUq7XyQTdFOvsESXVdMyBzRIQgrVTJXTmowhb1E14x2/UTu3
p82Y4gUVHP8xcG7Fii+ttE25+ZRkGUWJ2R3PFL+F/gf883NuL2VxLZYWODnZ22ku
0shyrFidUcVCAEQtbvthY81VjUw7Upoi4gvJWpCRbeUpphR27Ik2nZmrcfrbgqGR
6r+y2vryjZN8rLwaIMHOV3BekdQGHhJ2WAOZg/eLOJKFzkkePiyDYTOk9rSnCE6v
S31jYdo8w3N7PGmhPbqtdufWdwsPFHPe9B8gQsPb/O2w/IU8KD4goBA48Uy4KIT5
gGy2SCNzDDIrg0bzTI8l+B9gb+NkkvwolWTDTDztMgt/v4QV3LHWtU+wkBtwmJGj
LRj61k2lwK/r9YCTmWNE0lisX3c56/ELadSrlcQRir/8SV2MW2e1onVH+6WVGKk1
m4Djwji1TQd2z+8VcIgQ4DASMAzJ2OMnBDDSdSMqAPnhXPH2U/k1P7+CwP52HFkv
BaWMqWbP9Gwjzv4axxcYcnwrgX4Kdt+8pkaJ4J9+wtIs+Po4M5uCqtlhHtWkx8E1
Tk3WvuRXB6tH2j+veYnLr31q7S7AmHWdSSMu76r6S167yUAvuF/TURGeYGFBf/G+
XmY8xA6VKz8pzgjNMtuBVzSoqPPUz228ybDqNQN0j1u7ce/GUWQRRXj+lXSE3cWJ
wqwm3HF/SdER0vguuY24+QWixlYzsP8xiTukebdx2KIaQUYOnYeTXCfMHadb+tC8
/GoSyz5Bt7/7J9+XlQfsir4SY/JQ1Uhfxl5f8abIQzFC1cQBYJSOa1djDhBMgHsV
WXK/KLYzCeLN6nYX9qmosyffkpq0FdwZqc0+FDIzGIjeMOnWSxNYXB4d13OwFBTu
1OXnH/UZ0jnk0qwGbNuU2uEWG+P7QJ8um2mSCOPI0sHgXJ6/FTz/iUpqWZuv2VNO
Cnt6aEJl/c9/53WRo52fMQnW8dSGH+xpefpfIT06vaKsEHFFfJVqSThK8MXAWwEJ
0/QWP3GRzdCjJuKT7aCRCxzwvcna4as5eRVsm/5uWhmzC2ONHVy2Spvef2XOUM80
8x9vTEWbD0ccq8sZdKN1gf0OFVZ2ySSqMcGwV5p3qeFp0Vr9E7QkC+rcZ/Qaf4me
3QipHPeP6IChLdecillfbCdI/uK/JTkXBGvIfyLjZ/Rq5c/tQ6U1sEooJsdC6G7n
aUlQ8UKNnAvw0vqwzd3uGdchzoWZhGF6DpBPeU/gebuCo5BApkW1od2eaXLUVs2h
IjQymcdI13nz6MZFWT624I0yYwLBUaQHDSfammNXyxoG+v0NhG9kLsHN9JS94D/C
l3BmfbUFdZ7U5gxDhlW8h2GxplkJ16S/okvyH1PWb7RJx63HeKyuv85BQBZpJNbA
t91yER4pGBk6iMVWpEtUQQPyC2wDjfVtOG6qX6WNUboFklJbz8Xx0NpPXfIG4Ju4
AtfjeoiHY8cfEsUl5yKr9PCTwqQiibWthoDjpZk5tlZa53dBZxki83cBtprTljdr
WruEAmM/WOtES97CmEi0b9M2TKjkAF/rhvNDTiHZZAQLG2pD0ovregFq7Vb2xTtt
j9m4iig+/ESQJsDvuMXIW8mFyMHsknWY8cEu+SE9VnUAGSthrZuyIt0HTSWCRrJ3
tZrMLJkoxI80GJLW8IABcjxCUsRMPfpSJbQmlKc72v/3Gj5MJvZjFugsBqIYiHWZ
u9etZ39L50MXVoAEVCuMJG8N+zdpxomq0b0FAXZnvbu1tw4Z3jU0Ym1SG5qti63S
KgSn0LOLWPYlVHvYVPLYKi8CK/fxNzCI/yAsptPQyifwl/rl0Nm/J3b+otT9+nR5
iRmqoO0gp6nU0/owVcOuyAjQ9fdqO8aQKY5Nf7mN+f1qUjhvZD/t13aXmWmwmIb9
n7GFV0KgbYOtpV4yO/nOyaSZq1vxBK60L8F3J9E6GlPtVwrhTJ6rd3pZIlJ/lyID
mpPgGgDZna8aH+84bOTivxW4lpSQaN4AX2YvBZ/3BOJnH/7cc3cBsYGnI9OW/0df
PomBRHpTZ7JqMml1tg/wmABZdlni23ZXLWrFrAam9py7fTmOIP6yPR14sQjwBgwO
ju4qHJzYJPoXzuKcm9GCOwe5lZvHkCYSgNcUpXWnMJmul93dstqDpo8TKyXhe+6U
6R8A36rG5kAMfpiy06NPfDt40mrWLLQbay1YVFSy2ar6Q6LV4fwOXVOg7vpCkugz
ypMvJzsb/Q2+CBPNYdLJHlx1KCeVf1DUVQGedETcy3bSP8SmWXrrlyhRgafrKqIO
Fzq8Ey0L0C76MCZSsWkDy7fyhvR0L+LoA4rpZtuQ4rFp7MkxB4w5o+0y4qzLu6mU
6scZuOrZV9wdqx52yVgqkkj4lmpDGy4pqa885IEebJVvZbzmDksvRQyThWC9ZRtM
m2/iFWt1b75FsOVGsx6cVatxIF4y95qAoryqZ2FQ9Oh2hjOj6u2VKJD36gNqHuDS
dA7OwuuP1yxScVGzJQRXh7ieDbxIs+e5KN8iQl2CbRG3VxnXHuvnduT6mCBdeM/A
u2Y0FfgOQQTIfT29xw7bu8V5aKw8D/7JebLzVbJ3p3duZ1NfwbVzEQ0ZKe/x0dBX
z500pkTaxbkJy6wYw6HMl1mcicLlHNHtin/bYGgB8J+AnLIFfESyKXU0pDKXnKae
zHFnRJoEc8nOOLb0sYDxrKyZnid3RkEzyO8NDDJnPUM8uGEfQqfypcmeLzQfzAhI
ayXJXR0MSXQyyQ+cuOlld3ZHggJKj1S9zDcmTlXL9nD+PnZW50JK4qLHlxUWo+FG
PxDg9VM+H5Yica86lGLrgURscf03QKdyywffOhK5Njpij+Umvpsb+fMkMT02dnkt
TE+m06D0tPugAJatJjajUT0uE32+y5yop+t9g8Qjk80dRr9d2Mv47xylw1CpSEX0
LG7iOF/Y8Jpm/sNRDf6jFhPTAHzTb2XRudIyDLisoZ1/UczKNkEWvX4ywEvwp0RZ
QIum8IQw4CDDq6cM5m0dzFFXqdZYhMMEJEW04YijlQkaM+4i6m8akDvWedObOJL2
83P489MBHZT0Drh5GlfRjy5fDJ9q9qSBIv+ggC6DOrOGo5B9rZibkhQQVrs8nG/7
egiqEDocRpmdH9b5+ax5JpJaLyU2Ie6rRlR5c4IL2TBPrpl473BC1xf2bZ00q05g
s5KvxzOgRlRSx69APRF1fA2/FNgxkMT9xKN3UQjlq6p1ic2JDlMzkjX2lC+nDW9g
PSnll6fxwDvtxG25k6tC3zRWLRAgzFipcEDxXcnajCn7tOIH47U3bp85uPJXb+wP
EbOZCR9sS6iO+qqn6ChINBMCxxcIHYbZUFKsC9si42rPyrSUWLIuxKOT7nA1rqbC
dn+vx3surjA6soaSQRn3A7e6COY97FGmaPSjhTPSL20/C5lNTcG4/fsRpToVNdMl
ygF8JaX4TefC6wn4GGyNQOflguYLSL9GwP+vjlPFt2AZ+qD5XTJNBRNekcdqLIe8
vFSrVbQsa7NydtwKUywCv0E1ZASHDz5U20mW6NpPM/zETLAHN2X+ZxkABdSsTkEf
DvmWvmDC5JrZ8+fRvPmSfSeI75YWW1dhI7QPcbFu3ZDVX2lfelAG7Ajq9H9pf8p1
oYlIPFqgXQTkKzZKkL1SsYVMSsbrRjjZOSNVFpK/ZpkTuIEQB2AasO5vsSQV80Tp
MSaDNyTp+Tl5QOMVGwRq3vW/CUI9zjWz00R9N9T1csfu4sfK2dsdx6Dvdt5/Q7Wt
pIQycplL3kN7HaW9fzqSekYsIZytdyh06FzeBIA7HLpP8bPV3XILYNhbgInDAwbA
lNiZEImsVqT4rXLnV2Fu6PD1bC6InLwzo6RSNyPqrru/mLqLI++a2NY8Ej5EChdb
gM64evky06LlHyVJsxPmACgCnUU6AzhCF9xiLmlF6R0FC1GI7q6lsfjeH5jX8zQR
iyci7SKBZgCIz7kF6TCBvznd8xmAiWnVfUrZa8cs6uW1+DJdCrXfhzMuAITd7OgX
FNGVlkuA8TmA8ogOq5PC0Fn2Bn4JLeunwIWDoMlATxyMb0UtBGLnL31/pKT5FKl+
vPHWAiKRHvXOwFcN6JIFkIgH23Ud5/eK6ygWDcOcby7VWoCtuiBGdhhBdvJywpo4
X4d+H1O61F2dcjiCtYYc1XRRkvPPFoX6hRA943lS7FUNmAhceL+vvqMYbkAcjBbm
pqid/5kj2R8TtZ6tZj1HoWoM8LQqr53MnYNLDhoxB4VEYNnrTKahihW3RzxnFhBt
ZNUFFj6xWkA9iioa+s1CSwZ7jJOaU0HmzohlGMrL7yDcJ9w0BrqsmLQuXlZ9ivgL
Gw/g42MPGU4+z2/2yxdWab6LdLJTLjpifZqAcmp8mKvgT+f6nSgJf2Fb9nrFL7+G
7irAe2G17yWBndwYbYELzDD1mba+piiyiBnefDWGgz27mQ7s/TIq8/S+sz4Uu54j
A4ZJ7VEJknAKIFXqVnXeOHIfZBx/G8MSwfcXg2SY/MDaNPZVbMulu86qP8NTeY9r
7rigwRfVkgRBXTu7bku/Gldxlzm/QlA+1NV0J89f7w4eGoshoVkJGJ0b20Vhzj33
JTCPTIoPttobFPGs3BJbuv9MvWKify678bYqkZVDkBathtHzAi6zt+kBIhE+1FOL
Ga17CsoiFNDxG4/I1abNnG/P2XtbLf/fH/npqMpQzJRdV2PQ5p9/wY0DsSd4V0nC
0+LIiQHyRb9sC+btEIIVr4Vb4Xaez2RKt73eckCT4J/JCVT2NXIT5hWb/yZmyo9d
XmpnYmQyd4VwH1bOVlR0IS3ugEiCW4cBRWygArzHdsQDLLMKqvq7NIVBy2DQUjHz
xlPWnCEoGWIT5nFiJ8GYWiPcAbbuJ+P+U51D8KBCobvPIH0cVykY2ZM5g1zBVsZn
9EYt7VaX9GvtPKnLxdFnuv6Uk3iqLCamDQCfU7qHVlYJiZ5mKhHSBE/xXL3fzB2t
UxThHmevLxoKwEtTkrkPRYiCrQI95YKcNT3/Htw9C77ry99ryLDJh8olovkmYKRD
mwdp1zD/U6qBn9W8CSm2g2hzDLATByMnSyS4T+9olMPNO3e2x3TSOGjiy2omSFng
5Z/8T2PEsiJEGIXtVkH8QWRjE0oLqfgjsBN4KJKNtZzkPbv8na5TLWtwe9KV59p7
hhA4CqEjeES0UDxnTEkZacrzTDzFjooHGFG+F5etVDew5meBF3FsJ71KXg+tL9Sq
ZQtW7crbk2BlGJh4LuBOJ7YvVMNVNxoee/x/K4B4U42i0m7kR5GE8PXYv2UFvGCA
eO8JqjUg9Q9ig5bGyRixU12flt3FWxdxn+lJy63eQbCCTOtvIocKqJgbE3Z8h4Hl
0I6q7UHL/2iShvPNtmDPje9qsSELNRP4bOVzF1IKudclat1nx6sUZ8CCou+Xqc86
AKHOMGqPsaTTWHoNFezCCCw2/SHrfc3bUB7tfTfh9roMdKM9uWvf1MLVi47Mv0na
zkPpSXxqTMj8SHJ0GE7+qrCkfta7CA7XDisT4UAFP+esln3KrqduE9qa1uTHhQ3h
QuLzkAaoYFK2dbDMK/uNYPQ/lTrYmQbeQ5z4iQxhnkzqofPUFszgVBmxb4h46nsN
S9lse95kP7uL943fBIEw0z6+njPh3xgUJdhmqYzUvxJy8XD6m6OsEHacLfT4jDy/
+PtINoQBQa7K5gk9MvdnHJscXNxKE8TUcRja0NPMmk+2VyUgYojhcyn8eDg5wf6Y
60nAvV5qLun/pH4QO/AG4ti76lQzQQo3YJTbN66sDdg5alzlwJvC/FUrvRoC9lnb
52OU6cepqnHL6h00Xwwm89Rl2YZS032ckndRd/wTUTeyT+Epj1aNwkGl4JbFl0oi
zcwlvd1SfzylHa7Bwa2XlbEuM23LYt1UoYbzlI1FeRp/6HfPjgkWPm8Ea5OdwylY
xVZkPfbK+NoAuAzQ8euBaRfNHoSt6ywOjGKXzlI5rFZd6x4rfyTbwtQDWPpq29XR
svaA84CARNRTrMqx+obeWcEQ3RpdomJDxw8VWvRV/oeidAs1/Xsr0WC7SszaBKy2
t2WTfAEuaFc/UsuKMWjtPp36SDBgp3FNMhkTlokCziTlpHjsos6KcEmtL0FfwTE9
Ayi2+lrd1vBCJaEVW/8nKTMLDruYOjTuTwaeqCQi6OH+EBLmtwHiC0XnvXL1vMli
2/T5N9A+ez6cNuKLFQHB3FkkirN2UW2ckDWvHtzAJr5fu8dkIFkFpFps/ieFma4/
SjNMr/UCpV5zHIqMShYsTEYCsJKGABrKdVuprcTGY8mtuZ0izrIfi1tcRhEXqIbY
jYo3C7W6l8H8Kq1QlKseHOrbj+3XaoBZfengCQYrA6l62ZGZE7Pm9RTZ83IDt3Ht
sFSs+ddFnA8pJA1S3lvPSIFrHeh5tuGeQ0gk5KiyQ/izmBw3NLlZ4SdxnV7fM5yp
led/YqbEN/6QGcE8IqhelFpxNRHGet04ZKvbcvexDSrFnpUDamSC7yv8YR0Gm9/g
MJcgFmlZLUO+xgy2psD4lMplsipUMlxrH/i8eY5mdrnuMheIZw/NEDVFa6NQnVtO
ksiRS4Oi/f9oo3tvJvEG7QvMWOl15vvZ0cBypsH+HCKJIH9+2iJmy9jT2YvDzynI
5Br2ByPmGUzChkn6dtExKpgrwMRIL7Jbu/bZqU+X7Scy+me8PoY8SEyuwr36gV4T
az7PTLhu1eWK173Z+YbxpYJGPlID7W6zq+OWt72p1wmUAuUO93Ih0XUZuCbNUx3X
6Adk2PayLjPLOKFD8EVQ4NnBj0lPBMok7qxogb8enFmFiA96UGvLn2QvfEfNkqgK
txhWMw7VvNlvCPLIjs73IBWcncaabCTgj/UWn1pmA6TQMoY5szBTvSDawe1aBqiM
9N42i0l/JO1l4g5os6jCQ+nUmEk9JwtL6JB5Zi9cYdI5U/jRqy923f2j53wgyaWv
nVQMBULfHiSWMhSRkETeg9wTKKXVJ9UNO+MvbZSRBTkHu9VY3dI1IErAj6LKMOb+
0wc4WMj4iTFliIiXNRTWlmap5YwKf8dQ//haso7aTQ8uWyzgQIQxpwWy6St+Wzou
xqjpLdV36D1K64eI+fmwmJCKiniKYwCHtwjNUIeLKuF+HrORjtAoWW6V40v3x3j2
KF1/VYex5lnJRVwqlGdnLBZqlTpJLcXZR6x6gZvFg9rifd2gWzUaKTtr9wql3PUX
MJKsL5SfV/QP+Wx3jxtjm4TyRIuCYWI08gU6lR6KC6O7lguw/X93znwdApGg1BY4
h+EXwROH2IuxZf+hC+O2fLocVvd+Gx1fa6jshquYGKuuK8C24UlrXfy55Lp7eeb/
JPd/0jaZtOkzTQ+vS9B3T3JB+rKzTe0RYyiktcs3EMVy0GiVDGi3w7DGjYgAufqN
c3vLZC1sKUv8uLaakqvYtDZ06/jV+ul62hzWCc6M42i9FFicigpm8bw288wD46SL
u7GlDc9qtMZdXtRZDXCY90L7QssLKI+KVB2I/S49aGryLCQ3BQj9oBSZaXOWGmn0
kTmRz5Hp3auaXxgtL/ctQw/kfDEKOE4+Z2AdypXze2aXKZSjUVAh8Eu02O+ZXVbc
dr5I0uJ+gvwXoD4kR4VvgD9o7mb4p1gRB8WTeMFpBLDIUcJQ/svq6ve0AH3Y44o4
/ibXezctIxIxn3h07rrTuLbwgVeeUg1gHB3m6/7cEXwkwCjrEhNEArIHi3ovsoVY
2nIB10pFYfAFbLzYWAs6Cq/JsUNTNUv2zr84fciCs2teyeoKAoGIMFwAnfXkR29j
SC0HdH8n1RMg0pqA30TEmrzm7HKRX39lmLxt/bv0ZJsBG2whO+75easImPRuKGtO
qX/oSWTLeHBFFvabEawDZskhq67w4MnpMVAnfKZsPNQvzfrBV3CnEYNIkClj3I5k
zaC/2vvIHkwJKoNZulW72rmPWS25bRB44sKgDo1w4G6XwblUIIi4t5F4NDi2zMhi
wq68IbyfmWmFk9iJntAqP3AhYkssL8vsRWG5GEmRhqtxLYjG7d5O2FS2R4qkaUG0
9actly4JWyL6vodtFZMfP61WIWSku1hBVJUO6UZ+WyN72IUTze6qRHwizxc1wiGk
CAsMzBTgbPAaLyc8YETy2YK5jypnD7TUKXGVpyI4zd0zg779i7K6khZtT0GqqZ1I
G1e2roXhMAv/5qG9KDQ4rY/z2xGUVJcF4RUgUVUYVR1MZ9TdLbi9AlxG5K3BxTQt
elxwjFFVWiyhitPEmvQ/kE+b9AaTAS32DhQXUjKfAVT/i6HYFq8Z9x48Rl0X1Lct
09kB7mDQ7PW6DxfCZJZ0gzIuABeti7Z7XeE53jElZLt5zqG9FxILbtctnKL/++g4
YECfFoBI82m8K3WgBQBzTVKTs4ayDtgn8tErss05qZm4HhsdDuWjRieBh6Sww6w7
MhHJTlNs3KAsZksnlce13m7u3SFPJYCYHG3LkBPtdYIl/SR6XcXid/kaHfng5mBA
vUtb9qNbG12ZSwJjSP/o1DgjQuNkj2CF+xmAnobjkRPDDYI2S/EbuhnB3alwiqEB
0VZ0+0rX5ESw6zYCCOYB1X/4Qr2GpN2tcLVyhHToK+COpfCAZEBYhCjhYrR19Qyg
JbuxbAXDYL+iorkctSIOycGLasI1juCmdzlKOMoyaHkahAAYaRxPYcMzdZSMKPtV
0pu7iPN5cbOKm5N7VpVdyNDBIF3eeTQ5iE3NBU6GnUpn3LYLdZiXWwlu53bP6pYW
P4eVsQmmbdgL0m0j1aYC9+fdyCRMJ6d+vYva+GR1WK56rlZbtpPpr+QZLkr9nlBc
yOwJ899Hv5+dmxqOoNtM4EUHGBZPi0XDpTojbI2lIpEurxMFCt448YiHztrtpCH1
EA/aGlWBVK0SsNcVtKqXIJ9u9E6piZBVeBk4rH75wEWBRH5gSiMoq5+GgS0x3QS0
uamLCImnZbVVZ5t5Xx6lxCmkDJrUdyxOtRKOhB+SOlS8rOZMar/isZXbemBCgNXj
lxsVvM+9PJmAmBJAurs1isI9Mrd7cNtN8NMUDM6QrU7ExH/3DsoyjqtkY3KkfKXy
3ZqMkoVqkDggPUXPlwPAO9IqGmGdzvVXQaIlRXch6DK13imBO27WOHutj/ZAHcCG
SDldZXokOv5GDbWdfhIfRMYeMUUR+ASR7pFkLFKQCteZiqsESg8Z44nDxJ6ihRFa
IkXcey+Q0djIvacxfDYYXMfMPlvhPKSkTA/dtT7TCJXJVdMwIHxnJkg8S5RKGXLM
1Mz5sGMTQkK8TOz/1Y/jxZ+aW9bWGwP6R/fWhYxlhhwm0qrC2Mv/4ia6eJVuycEO
LoWpVV1sE8+q4u9OdzpexLQ3FUz29+gLcktfPfdA4kGKw+oxzsvZGF/U5xHSRjiA
pLZvgkWmcClD+Q8kfvIhj3qjDPTaS3C2FVdBQGtGNQaFNpNRl9BBX/WIg/NArHJp
J9fQ25V059h+yhFVW8LdA6TbR8EvAL18IwtqZz+vZm5N5MCwz8ZDxhmTaxUpMxYE
Ho1V8QWNH2KUe6dapRDC8HOpH/n1YLZNzW0H1lzN/SRGNWSimpOUi5FRdHZQ+cq2
GAishJ/oXTKXWV66fz3R3Io9pp+CpIjcsP9hdnDMTiszHFNqZ8mUEGbF/v2uNU7Z
4HXGENedWnLow3l5jN06+Vse0+dd1ZyUbP3XT1bZaE3vzVF+19de3cIm3rx29lbI
Bw7IJkgdh3wUCBnPYK+JGIgwxFARYWl05NBlOkzdqZ1ASlMvebv3U7ca7PPYu0oA
CZHrVLFUPPocqn/gifzlbhptnE0NItUsm61x18ms+bQuJ68nEwJfnF7ZSLjgD+18
/ss3rYULsEPmUAFzDyOREHsHGUmfGdtzQayJskzThICQAFcW8NVWq+O8WtL+MDcx
29U28WuKjiCjGwZnzyTlbZkVSAhM3+uveBRAB28XZyWfRR7YPmCaTV1aw5zlxEPU
QPO27+0VKjR2L/POp7ZgGIBzfk5vW497ZK3/YiLqtOttmKLO8TMCMB3kf3owQDiI
VNneKRprkQVLPaScU1oXzuIsjtdtD1GFzByeyATRo/wVPLd+Dl3Q2zHo8LDsMpWS
hb0wAfaeqsNrhrQGepm1JqECIfqoJpvLGrLkxTR7qoKrcs/Ki5LLemSts9xRy91K
jonX1bDiYjnN3GWw+DBBggYhY+/WYvbKw44q2q6NftZzNHmsWRmDzjqCyLWkTRJF
2zw3jqTwas1ZjICPDQ7igKrznuXfefhTWKFO/BEVjUhyN8kbMuo/2VXZ2uXfZPVR
vsNTWETngEYCdt9OFDIhbB/xktYh49S8IzNYuJHnGF+gVLmdPGG3T70olutOkgsW
JZB6AIxmzsOyh9vSRtL33sKZwCQaPp5XzBjdyCYYsNGv3doV3hTaXXJoY34iX68D
rBjKiQ9hPiyu4r8ev+ea10UqSDHUFwuRDPR8uB93hDMu4KaMJz9Uq/8+dpP1PR5r
4k6sTuZsqpzeBEWC0w4Uzk38ZiQInwt+TEfNSJcpMV9oe0uvilE1wHMblVtIh+gM
jBChChxfCf/bWf1+hovlRBEQAMAd+UHQ+t8nr/TJfMZ9ipOgIZE4uZ8sRoFzoPVa
Xx3htvAPslRj7I4d0GazcsFQW4Q4gR2KYEUig9jnnkxsqKh4fF93dULwulrbYcRv
gHe6ALVC+tXo7ahfQvEGudNc6vhk1hO0WkqH6h1jXYxyFYLR42t4nlfVlUdBwwS/
uJ7sO3tWnhTBHVZJAfIimszVuM79M34G9qcE1fApVHJn6CWv2LVFsSVzXZDGyjka
yTeaCCmZ/ZCecRo1TT6WmGvxFa3mVDWTX5n9pZd7OLCOXifnmaRkfQPf2kgERo5P
JWf0kY0vt6UPo4+Q/BvKK/xZ/rMh6G+PwRefrB/qgN406/YxGiYnAMPNDZPYbxX/
tUptjB8en2k5sniKBbzmvTo4rFFnL7g1G9NBkwFUmA0h6BjYIwWiq8Duc8aPagAe
4/KqBWZbh6GYltjDCghxK0tky/NhnPDg31SmSncTnIhSW4uM+wX47SHSf8HCXqFJ
7SQ+3CeM9llnWm90gwGfSSHLUI8yyqfSAixSO/SmmvMioFPnGAfVFEMQbfwZY47i
OvCZvArXPep/sXudZb7rMTinqb1DF6UsVxVlqgTdslYQIlZew2SNnb6MyBpyg1W9
6U/BUsmi7Rl9Nizxih3nn7NpgKaCckjCfU7gkw0eWae+1wdRoB+r/JXxzaaxDfkl
WlyrEg7vGzIW2FKl5ETGcveggYsbchQLPPhBKwuxFcgbKFq+icuI9JPXr64vYDJE
jvB42wzhr37PbkXo2dx5SGt8VZx4iz+83XpkLZyUP22Nq/UIQv0l8ULUPEMy3fh2
hf5RzIAoSabv/XkfqxEq7fyVX6eo+G5FBH9F09cp+PI8pAcxkbFTzo10f28KYc0d
LX2FGEL707TKE2c9HrpCOw44l/MepQIRYFxbvhRxxfiobTmH37Dxphcu8VShWVEa
vvl8hNQuG1e5VudRx2olDZ4UqFsv3mA1aisc0f3SFunakP9MtEI4qpuiohpH11Rn
6hRpCgL5PX/8vb4nnLweU7w31KkDuJTyyWJ6p1MJdKZfzCOznAd4QNPiL2PPmLLD
EubNQ/tUGSPWz+52LsyPLRO4UGwBdp1s7kiU76vUWABaam/Z/tjJJNvw72GzI2EX
NnGo7PnmFsTsl18I+rf+47dNJ3z8coN6PT/Ur1WFgteFOxfnGXhui4px+0Ry59/x
OMZRi7L+j2P5MVPmTQU/yG7LZDH4qXjWaTGO7f6xsptxtKCI37myS8Kt7/ZBxHjS
0GqWpwU24yARVkrlmY/33fUlD43F/Yg/6OTlimes67N7vnLCwR7oqNZfdHk+cZAX
WgKVQmi7DOKuSEjWzf/qgyoeDKuyoMxzWauCQYDx/TwU6C3vW7YyZVjawzmTwHhQ
NMeKxp0KyQO0F0y9BgOwgnqFoiugMVkNRc34KeBkRjEiSVdcN52ZOg+/UmtbDiGI
/czh8EgQaZD7yk0NHxApv0YTomJgUwxa6nIEiab8ZCvVSNEMXhV0xi9iCpHz5phD
XkruMITNYDk1LhGuiTJbSbWKfqOnUILU864wn+OJ1tFh5DoluyeYGMtMzmKQCfgQ
n+KvoLyWsHBhPPShbTi1sIPA24c6UgtIDYapbt7YDUfDpDRtyi3CiWX/QqHQkks/
D67hxzgGFEpoksURjBKchaXjOBKoyhi8wzjvBYY8q6t7Rr3jmHXn+hKftej2xAUV
eLWOA/4tMtMJYZY8mTmB0oqF+l7IRXzaHN0rhvGkgPL4yIF9gDNKR9Q8FkjyU819
/9H4KpcNvfvKNnuK9QfViBOqtnV/nPOtXM/oFEidlusONQ4J3zRUjaa9ns2DzETF
V5UkeTs4wrz5oT8k6/dWKOUsFcGQ+N8CzK6/gdt3YUmRNHlkOBRG1x0XvTfptnI1
4mfX3MV7oz///dBeoqKCtc/gh0YfWTMkH9+92TEKOuGNVKuPYPdcbBBc3hOT4W0b
CL+GhvqS4JDoaM+ak5e9wXzp6wfW/xvvjxkb27MJBMT0DyHhKBN8DyGOTi+DjMxM
YiEMYtJ5nmeeTnYiOwi4qo7OaJqOhL0oFyMr4Qsiy5frtm0Z6tRyWyxj4QmbI885
b95yk3iW4rLsG9ydZRNP2B80UmbfHl4s0L3BFZnC51wN4nElZg+qGwtLGhkrecGz
iL7QHX782m5D5/PL6jzo1iu6c8N+7ZYS3oXx1fW1ThnhU6lFr/gI/xcy7lB1aQpy
gXjVguknO/O0tIkpjwCTIAm6nkJm+wKhHxbzSV1a6fpX14s3jx6B84+cyRfDAAb4
xZPVqf9mOJFyxgwlOVtIqJtwFMY/wOFmaS1dU3XjJLTjn4j5g/ijoOzsS8YfRXUR
EliAgbhnGQuxvhHGUs3wohbUS9AEy3I/Gr1BRlCG/RuMqMMmLVzxa9o94ZupWtTS
e7vcF3Pz0SIpMPw9eD/8M/ofXqnLXWqPKuYgNMBxu2p2nLmtwkoouQGd9chYW0yo
u5fkEgDnJTFAU74YsNA4n8znHbYWuPOc2Kn06PmSaqNSrcV7PbziVdDbJcvNo2p/
GxfcADnObCCp0wDI9OXou8P20b1xl71f1mu77OJ8rj49FKkzbqCgSUY49zOsPYCX
ao9v9e0BVj0ZLGWMpYrnZS7rcbOcA1mlNMSBZSj/XUUNkB3zd25uDkHH0D0bWhdw
SLEMPOEQUQfue7XCw2zCOAQhyS8oxaaC6j2quDfuCcMB7eqN7iyWdU9ZbPk/dFsP
SWOgoBJ44yRwGpELMwa1L6V6wYe/e3NPjI79p6Xwz88+bRC7bGQRyhw//zoxryyj
oRvRpvxw1N19kfj+zv2qgEE/LFWcFNLe9J+1tixF0qLQIq+odMk6nT7PaNiet/0N
lu7MhGLav35o1WuZHnc89vgwfOKnlFDRKlmzAumvElc0ks9QL7MaWmGw8ZHgbk4f
e1/iUu4C6YwKEApVkSj3ZvmeH27I55J7K5rKeOu0RKTjOGdHwYhIMQpfj/OCqOnG
bclwbeBCjouQZ0CG0IjIJFtTucKqdwqoJf454aRnHIL8Df+cOHjg5aXFTjuJOgGa
RH8cf1d02cnMOc8kGpmYVcwhd2hI6u0H0uDxR9dNSPTTiZ8cHGsIP1tfdRunprLq
6o8jDDt3pekTboVgY1cpPTzpMQIC7Gzjlbyw5UpD8ikMLngxSuZ6hD9x0MiAWR4a
8ET2EeZMscTvyLPEBwnvjFevttMLf0ubJA6wilM0EoLshnDcsjGoEJJUj+SWMcXw
/a6czOt0ka7/aAcVyDrh+pXPohc7DMEc6r9zfDg1VG1dkLvHECcTSirUXHDLKWlB
9FtR2e22P3DL58dKSHlALwmVgTFV6IN4Y5Sex+lRgfam1PBFYm4Pc1xEIkjwucV4
7BPe0S5d5UGb1doXSFfFU202EM2KF+vP/z5EliVXpuAoVwkyNHo/Wp0mdXtlpRXP
YNlVbhN7juJz5HMadCyJOxtAroZ+AXTbP0eiLsPqgDZQ7fr9dO42+6gJqN/Grbeg
miNPxu5nmqQrBNSyQBMcCax/3tIXMSUHn1m7Qa0ep52rvfH1Hp1kuyAOczeENMzM
Od0ZVfi735FPhgHWXkHqZZAyoCbSWD0WWAmqarJqbyFiBhb3HisbxJHQEWh4K2Go
ebvnHOWdo+qqKB3MV5FdORrDLtd48MAlcl0Rjzpw9Em+fRWWYtBvWTH58Ay4jyWG
xQOd6GfDyvWThJ5Y/ZhabX6JGqDj5nYCISvag7aWurO43HouwoheO8Pcp3JPDWnc
D1THOXcPRZqGgX2n+3bP10q5LSnFjVvdP6EhWBKa32QCn7b/McsksFsyAzUNr7MI
y1a5QXb4Rb5dBOAWDH0AGMMULcOFLx/om57LmC1BCUBOKi8X6TzxcaWeQMqy2DK/
dOHcAt4vPvsfQZ0KbD0rcIXWuMHo0sawTMvqisuUKEksUmbyJ7cSz44a0a6MdH1+
mkrDndgiXMzIl40zODnptjJoEi8jno8WxLI+f1Y5apjNARb6h88JwPb2l2WHF1OB
rwMZRF1z488dxRUKWqfwiMsTKD8Gbwm4kWShHa4TuREXXxSOQCvl8EJ1uweNM2zN
DAQX9PGfpeBih3xxif3wuwZxaaOg9jfJZSZ5yx0wBKtHWrDieGiy10yHx207nO4s
vEBrW1AX16BBjywAqDU4dyfJ2ciramB20m121nDwXKiujhbdJQWnZXG54QN2vWgo
BsmZXU217kVk+VKf4UPOZ/+rXCociLsODYIuGPVieSsoWNdfhpED/5N7a0ZKz6OF
8BJVELFVpF2yVpouh5gmGwNeZq2/4B6qQfM9czIBHKIAmG2JyjIkk1WEd8I9w9rq
BoZ+fsmIHzgHsBFUgB8Dtja9NtkfblD9HYKb1qyvwzGDaOTGKSVWyLhxhDleKcKf
lHWe+Ct1alR+wY8Yx+fo6JguwiFKmjULw7GsvDwKWGpZUZT2ppMJ5VofDpkINWmo
awKwzAt9YrW3XjobqeiIVHhhTbEyM8MOiCFLsSYLGM7xJbyccdVGGpw4wOgOMLqv
yzVKqb3oc+qJuVGOHMSpvxCy0U7IAo9wYibgGDIHWgYfzwYRlNBjVJMVWP3zDP3a
F/cMiCLtENsaIxX+2fL/klzL/VBMd6zjNvGFZ6dCySxrTvHVXTfy2iCvYWjmW/ZM
DR0ehEaAsLE5At39pESqAiyL2DYsFBZFNXPpMCl01LBBYu0i3d0aCYa7n7j3r3zT
oolJ+awaQsrgUYB057Z1PhFPSPYYN1yp31dNylqUrgKPRzHZPMq57KLueB4Nis55
/d51HQAi1dNSe2EFw2X5Is77p2JQhrLxAIHtQ6EXAT+e6efQH9uZ1TFQO7uHxCL0
p5bQMs3q6kDsaXqLEUyIjvA8egmRaME9tQio+TIsi6jO4QNgvi4fKE63JSww9eno
cyDn077SA7pFO/9xNfBZmzMgpjMBAyhyYjSTkfjRV/9uYtX9S8wG5xZz7VTe74vb
bD0IHpr0rmX0c419plNHM/dGUtjKupeWbZCa1wgcYe+OH1rtGHunO5voUbBuIymy
oSWTuzAqK7X2IUWB8ngLy5JahvjnJyKT2oe5vObXPTFkIYxcYHpHOlrvuyttHlB3
/jl7yp/1JP2qmiSB/6x6mERCQ8dkz0kCu9h9FTm+cKJTPzZJVLU3QuIt2qqXnI/m
ro5oBvUniAuqU6S3/u7BH/Kveh6Wpgt1WZ6YL8Be4V3AGwx4exlEr/Fx7vzb+a+j
N59uN5FtVN/xeBUSq/KcJ0/Ow+iI5+IVZPh9sSwd925MXOjjjzz6d75KprZCYFT7
Gq5/Zmg8jEeCQJVViHNIBSqbQS8F/BExH0YYhKjcgrFjZmNBQx1zFoIzGkElGoYu
igV/UcUtwQbjtrk/NX4HG0EBtx5KfMIHlf3PmVfd9n+gat70VpQCvsT7aPwaFSaL
HpnOguJqj8yO3ZjPD+9Q+PLPqkxZ0PaoHOeW/HjF66BaGjzkYjjX2+gsBEXNAGxK
M8J4/zBXur95xIn4HuAneM/RsRa96jY9vGW23r875QYXNsF5kW6glktsF7mQ2UEC
w2RKv8Z7fh4RnKyFFlGvW82xA9iBBWaRHnw/BEpWOGrRJGqujQKdi1Msvq7AdhmS
L3nYsUrKU6S/0IlLYzBjK3ICbAxBRAVQKdFpq621M2JycvTVtiZeNdzblPGlKJZV
kfo22rvb4PuFeP8niAAy0g5Nzi/G5Pmbvwopm7tFjB1kADq0ir+Ze9bEkbrs7p63
76qI91ym2QF5ae5trxuBAQdZaWSuP1MNXtKT2aBS92sO7rLV/2zkNgo/eDVGlQB4
9tmDEK3kTZkTHQJ9IBBgItYYQJkSigUHlNDWFmS1OyKZUZVD5shqINMEoFSFR/tN
3z+tVMuexG+AVuv0v95bBfQSKV3DZgsMCHDgtF1b1pstnEkHPk/NohQEij8SaYxC
NDCiQt+0ys0T9I9TSIPA/7j5EKS9vZE3kgv/edBdFbuvswqEYRYUyIxySrZxBYeW
ygmU7I/ebbiQS7SMn4yk3sb9TU8Nk/d0r21zhVMZ97s2IzcAgrPWMpnMh1XRu1XS
G8vm89GcWrf6ar79b7huv1/XYt0zfA2ZNAiFbbFpk8ho9X+CTleQHFlNH4/8MZRZ
kGAgM6TH1eZcNvtIUnfdX7XwVFlB8i4fb1/76nZBVOCIf9HBkShPI/BsCsTXY1tE
H+VDUGIlVcJulErUxMohyepeMO0D72lyxW/q7+rXZWmZzJzEc/+E1OH3yWLqOSGB
kZXTTlL0YeWwFgAi5bV0MP+8uP8Zzq5qDeR0nFBAqeC6s87X+ELO/phTV7KpB+nM
eisya8hg6Rl7y+0ywL+PqCR2kSFbPYdLiaWZxylSGL3C2+TuBcgzJycIArxCugJ1
bxjm5nBc6RcQvoadc5m4E5KmbKp4hfUvSciTbDZ+oRzKqVFf7JYiknJfgCEdhlql
T0oduI7RJYrCBtOK05cpj+5nO10vZDFTH2I4+qdAtVUZQTORwrZ33acGK9Me3w31
nYhDpiuyoDrGw+iAN/xGtkkL+dYCv7Z4Y3Unx0tp5coloWabQDl4x5Cllf7PrYuc
OpdZxbKiDVDJ/FiDyNBSNJyM/2yYgz8Hd5eJ8SKuJJ4iCX4pZ3TtWo/6KTiNV1cN
ILP+tMMRd5WJioCNSt9kRA2ZrEpFXxnJVHQgNPY8XcRQqgG2NaV726+mp00j9zdO
/0+Qmv50hm4fpsPQIPXWY7waTGjHNDOdnILWtSanp8CEbLYG5RFKgWXOLxEZeyHp
cZm7mv2fETATXJJwZ7yW4Qg+lhNV6Vwv7rcFsMO+xNe1Jbb651+Phg5h82cIZhKg
N+w7qkUquVDxD8+BH5IyOZP5zXi38YRNPly0aDZJyROzegWUnOte5jK5c7JmjP5x
p4uuaUcT42u18U9S0uDq7t8Hb2WfH9J0H5G+MBRHxbaNneBmlvdZ9m+qk4dDE1Rk
eVOOPXLvh+Il3Hn/p6cliwGgAqgKPDCeUghHiEs0Gach6cBzbzt4GXCarvgQhoNc
6+0CUB2zQFnkA24FcldcPSeVsCI0+TDIBNTAQA+fCforPRaBFbUnJKNvDlJhR8OU
dsRWImgjAWYLjGhyde0CbmhZ5T5MCZoctSV4WQNvnH1SkueIvMqw6I+w2V1xwvrc
Y4Crj1fCwzeh5VTPvxwXIYYz49GFfHc0fF5dzUtJ6BzmOz5sXMtI2w5CiS/0A01p
rEZzAVXSIQbgjLrgKd50G0j8VpPvH8I2d+aN8YwzDYG58ssFewVWaB6ZImjIMVbs
I4yehwGJLI5Am4tH7fHCBFZhkV7l6rGsaCm9Fr8DGGczf0xQj1LxlyJsZ6rpZHVp
M6hDNo32KPyZIWOsdDeH1ngHh8WL7pV/DEXsRsGfRcbr7tAHRF3cMLb1nWgQvJLQ
h/hBp92wz9K+lELyD+MZ4XUQNzNZs3LJ0Rfz/IXpFk92xkmVHtCfwzSpyCvmuLMt
PXyNGqjJgoa4FjtVSw8UciCIQhpisMRYJepe3dBkYkXnlOPJXHDdWf6QDoXx5C6D
J2PUs64yMoCcAxzsITTK+//V5Kd+HOx3xLTMWBDysnSDyETiLLd0hO09Bqv1WGa4
mDF8luPoMlx+zWix2fGFR1AXEZC9fRf0Tw1lVK+klLT6331OYoPuvIEk6f+GCL5I
v4qAj6KZTtuRLLREQrmiGo2/ayUvNtSOO6GPDIEugsLPU+H2EOw85JiXfk0AzxfV
TmUhwmcInE1okyDxnK8NlZEYM4Yy98b2k3B0ZF5RYTeFLqawoE850LkPUvEPXG+f
V52GxcwFgfh8B+8RVzBNpaInh+lOWvrc1MSGt9otqCsMB3LgsoXiPSAP5Gz5ywVj
GkP+z4bRXAt86eFyUG7/G13138HQ6YlaArwtpdood8RWYiWfNfk0XbfNIOrKVQHE
/E2TzcXPmpniixD6ZOICAuuyEHQDb1hiCgbzA+kvZ/I6iqZ+/kp5+4URu7BW7Ni+
0OPGSc/UwWH97nkWKG4F58MYkg6y6kji7iAR3kVlS80U0uFdBbOFGNffbsz0VAPQ
JNKLdWSrPG0sBpRzbmHNS9Z2IiJ82iikI5WG3D1Gwz+cCtYKdy9TDX64uhusvY9W
bXfev/EIcBW+oY70gnyM3wXHs0PXPIqOh43tQlpH1Rhj9OiNCZs2AomY2MpOPdAY
o/tuFlquP+81erJbiz7VWGPvrTL9sMQWLe0oAYZRoesT9vG3CtnD2drz9ir8LqlT
FeFVY/Am0Iz7Hjac9nxWOY8DFRMZwHuBWm8duBb1qL9LOqDKe/FD6eIM1x1vUO53
xT7e/ySZNCHFJbLItZT8BjWVGKykAyNxVCYI9514/ALajsl3shNCIxoL8CjYJ2x1
dZ9qWHMmlay9kWfjg1R2rrapIJDNMLyBRMpvxYPypREG+PAAd1UpHjsDcexF90Bh
IrQ57Wn2Pje+YeJACRD1DX/CB6Z3HaIze+/Q4bfCH0gPuSmtqVrfTLm8/kte8D9u
DoBcQTMwCeHbd59SoUMXQRdgVBbp86RifYmolWdI9pfasjLC2t/WT6Fwc6W2yZuV
MXMLZ4lZESNkqF/05jIra+3+ScMtiBEpuRJnmfn1nO5CnxZkbmHm4eEv6o3mYb2C
9Fh7PaE5DqUalx+ISwcBdZS1ONHtznyoDzOQi4IupD9i03kUACW7Y4JDgv9ZlHo1
BqcEHsk9XKG7mLm+jff/39/kCBPgf6lnQIQJj99R/2GNHY7GoGD4jwpJ6fsRm8Il
YMdxdI3JfJvH7G1EIgZkbAGJAO5dsowLlK1sFB5O9YBlzrhfIoeLlQ6SQvH8Lu7d
nCHR3fGp072dCsI84F+doxt6MtDqWSOLCQB2Z/hcnMXj1t9w/jr785dHpc6EnOPs
+ADg4VYuAoVxdrFDarIGMiJh2/6TDH6IEC2AFkUvS02LvH/MOJ5+zUslgTAs8cU/
H1jc4NnsEaISu6klgct4hxiIk4+fuwj2YIjsZAKPDmaK5Fo3xAL0Ob5AoZl/A7js
oNI4JREAfo1a7QaTZFz5KPVVorf9YjPSj9NhjOn05ETmjmwIn0yF/dlYY9QdrtjO
RqMTGSxJ9UUW9YacaoTQG9T5swwD/0tG/FelM+d5it2cDBsOv1oHiA4gqltIGM6s
QTz6Hbk7QEx1CnoTgcyzi4Rg+mZSDFluorV/1ETGvmMtJNev9PdGGUYROax4U1Lb
93oEcbojV1UU3HoWjv5C0L3MYiiIdY7AAX3/tlYyj9xuU7SoRl0+87ncBJSvwpKa
+hCxtXE8cGRC6Bh6KX+fijY8o7xt833mXvCJjoadZbe7vP+1ZidperIDl7oxBk2j
7Bdq3NDGIgP17V3XsuBYYMHCb///s4PXDmsX7ECAIUxyQ8Fz2eOiNowKHEqayAiO
d2t6fiY72/i256NOqAwnmJUVq/CnnQkGI+kiqNWU+5pE5PIoPgIqm9O+yguXv35e
0ghcXJuvcnJMRPQNK67EqtT/JVb21FvUhN/YWxFRjjYx2SYN+hjdOgndA9RgEnSL
RAq0rz3nMTVRvnjUTcNxFsdFs4KpVz8SeEoSRGOwQLo1XlwpoSIOFJYF5icrJqgP
5OMBDLwJJ/uwno/h90WQKvk/mAkBRkeO9WbSSHn7M2UpI6CepXduzJPyBZdjJ0K7
NRPDr5d6FQQ8WtyJrSx7LulrW9ANKuycfRmHVJfHINr1SD4gMZW+4G3sZaLm2vF9
wKtZqa/4trO4qO7OoZhrbIesPwW0lfuBcIlfDJDqxX6m0OupJX5NJO1yHP2H8P/e
MZWgAYrN3TD4iEUPfpnVVVn2fGGFlWzH+xMj9OY6n9K6LGN/8AU6XcQo/W3AJef6
2TvBSudKHKNqoI/0JkZZQK3qIqwtwJSuYLb+wX73R728SLOB2Hr0icfj+hArrUqD
NFYxc5H3wSKcyCYxGwNryZO0fgLiUWWIG03UaUIfd77/Zeys8mDUtzv9LpVR5WmU
chb/va1AEOWGah1USu8q2ICGA4g0DsankO41FHIupG88tlD9xAA6lVNF4Lp93u6z
XcskSlTjOJEEo0lXp0IERUluC65632mnkYIySlLUmjXuIjc030W2fvUJnuxAtNXQ
KVfukh+8C5yll20N4xOLFbq19/WYbj3+dQDBtEEJAxSsmGIuHzE5YRh1rr4IwNHM
nLecV9ZMGO3Qc5h80G+Txp0Lhxf9kYNuJxp6IhZ13fZo472Uva+Mym8VY+/rfUYk
D98zcJ8/jf09aKbuRr0zd27p1yx50X4JtdD35Qzg6xcZbQ2FOi3pk3cu7RBlmbAA
9EsA9QQHRnE9KiNnkg61UpP6ldSbFbeSllZQAC8o0c91zJoK9vr6QJ8odnpFu01D
yktpaAZt5PxP3X6LxynW451HeesXzG0J/It/i1325Mku4pV7UbSD9838c2dfIn9Z
FTXddE7dzbXZIjxccEfiwspR3OBJifOb52zSNRl/6HlUNwgVsQinWnO2DbOHyIUj
N8sClzdK1b9CCR0FgnqXB6ZM39XVy+EkHs/XmgR/8V6YuCKuBPVYUOZ6wUgcon3i
zJJ2Q+oVa+2tCpIEZY051yMz1/v4mxFTITFpK5Kk/OmrB1I/s1CcVGndTfyARUcS
Ne7W75Zmh0Gwxq3pLNUya8Whug9M03tjm3rChWUIhJQSD03BnTQoTADEDgqZnqhH
Iwep8fyflFqRn6zJRuk6GAe+kXtD3hy09GsdtW+Q8jyqtW93mIfuj6iNVN4WEr9V
gjvbOikjcQxOtmygHww+YEgCTuWaXUkVd5bLkWsW6xVM2W/VjZkYWtXwdQIHU/mu
rQa+rAeIiSwNgyVchyRanIY63hPeoxkGFMno1p3swLJxUdGVenUT9loNVffgCRDJ
6bD8BtHRaqiJRd1kbWGZOn4JFvyscNVy/11q7/e4bIDDh/aTL0Wlg53UPyWwg96m
bHuaC/dQky3eMKkOtzktoyQlG0rkU16M5DurANlFAWTr7ldHBWDgchcQDrYRCb/T
pEpFkYRZvU0nyvE4CrjpNQnAr355vrc5c9Ik0cSZJ6w4kvlcjVaYm+akI3P52PS3
yAh4i0al7hekGw+/CK6gTwP36jSrpXI1QITKmSYFispi7lg5HjbFpwsSNh1nPx6R
cJNsMoQlnoTEE/lF+TbRHc2E8eEROwTz/qJWl7zH6RvFcVTyPtRLHkMO8V93bdOz
wPEb4MKneatSzSfYCCMaOewL7kUmfPVhsDSIU2sXaFHN4Al4h0LlW8bZZgHo+cJT
RZrApVDnl5Kh/VC+DXoy8KlrXt5llXe6rTV2R6gCItSDkGUpB5INxdOXruWS5ni7
COVSNzZ39sIJ8uc4CX1Y6N7xl4lf84qc+SSN+AudEwMgFSAK6Pym6fsyOsBu6w04
K8IboRKzApvFMbGJfaJQjamygGmGjmKBaFwvFGtVJcILhMM2XBajhWWGtfW6Ouox
PZRWYSRUTONKUii/hbY+GVrPfG4GwaW0FwNI3OPvttyCKWgP7vAgI3JKd6TgitF+
piKkzYUgSPRyJN8clNPG4O6/tFzp0VDk+y/AgjD0M/3JTVEL8JuPBLmSi4SiHiFf
Eb7h9zi6ln4LPcBHnTCbIldu3yHSIXBPsoV7zjIQ3bjANxF+N9sImRsN7s4fdMnV
h+9bbXJi/wpds4ls3HCQOvWe2ftm5QKThosqJT773G5MAslbP9HcSkUbRS7Zp0bL
jxtweXdfd9SdglR+UtFCWX9CBe3vG0yZBk001HX8sY/fl2WqJ8eZpHNMqiYoIYj1
FMdUunUnOIkrFMnTuCaVsnnrD1tsir2koXE+TOxQST58/dudI5n/3HQkMAFZ4oBV
9iOTQIcFDUc4b1mZrNXbiowcsJOd/J5PR5uv5+Bjlf+ET82Kpee1dQQ/HaKTFTLL
Jo6DY3JY5KAy5WB4wCN2wR5uFuDhq7S15ZAoN8MCjL1Yuw0+M6w2R3bvqq04RI/B
iE9pjG9BgPFhxMvGlArezL0TScB4g7vpV26Chm0IqRCrg0IA+h8YXipwae8FJEmr
aQYsJ86LZ2XwvtnAaH+DsgAM/wGIJEYFx4fCRvBlcHzhnKr6DQ+HqcMgtOFjOYb1
DXhLwsrz8z8ZUWbZSUXinnuFGD6MgcpgneyS5cNwchi6kkQEiegUh+mnakcYZL1m
IwWYa+HozcbXENVJlWblbF5jxhmqDtrxDEk8Y+4I+OaB7+CZLCXM44XDGz2WRSW+
93DEInjFi7FNxjDN89SBLWorQW4Hq3cUDEiTcTw1tdjEmEHYQRdbRTCIuZ2r92P8
uvtkZ26Ludh0c2IHsue9iAcgHPNPiJ5F3aEk2gjsasPI+e/TCIfvMwbhguSe4TlE
x2zTOoiXXTyNrwXCsMQFXeYfAWzV3KwTumFMMGDzJmCfrgFCxv/2lmwCiOMH9rYJ
//HcMcAvkuVW+SvL6euvDJ4zI1Hx9WEiK5oAblg9ecuhMLGCNl14VTtavxAJnzox
x6DO6MKYjtxDnuSeFaQteQZAhbleCM4rVNj4vW58xEOlsgHBqtv7/ZF4/J9jBoC3
4hDLYYayex/rMwMVgkSe0FoXKTKorxcUAEZppqYxL3Sd+/jsKC9UsOPAaTjSI5x/
nTIkXysM/tLPx9tFytQEW0nr9dxLUNHsmJFBRFUTOEoH9lQ5Y2YDQx3ArNb+03m+
5cnInmiNj2iUm2nyZMQMbqbAHMGNMVG++VBcdmy5O3rmTOEAhr6Ht1CrBsNbcDgC
+AzVrVA0379YsCEkjAxTfv9KiiqHS+wfZucDPohnbL2sYbWY1M+UJU5org+UUWt0
Eo5pgP8C5Bp0z2AYpj0J8SBaB2h/Tl8JvFEoo1WUcVKKuspn4puilznOD7oANOWe
ppbJEf+yho3wXiJXIcu+hISqmOHpa4dn293FzMjrStK5u5OBOV0fnPTR1SjSfdtz
UJRqV+PXsQDuR8L8rJKr1Etoq1pCXh8xWMaD6R6gpb0IaoFs4oHh4KiLupbEqcH3
wk4n1wjJcVRWLpl2UDWV1N3TpPCzpuzPiv8L3L758m3mBNDKx0Y2Vx1INhmkqE8a
nWOv3XpUewqEiBiKrW2wBKMbSx+p01+XSmSuKgsNiKNiFoH7M4TE2TJiqCk3fMJJ
jhvkQ/YJTQGfLGUWimyo6lmIaRU9BqY7PcN/FSK2eMjjlv/WkfrzrHVC02ziAZFC
0MAklOphzfRAP9mIuCB5/jbxtIlrjxXrBm/wOdGxLodAwzbTpD/nHVFR/WkcejP2
3YcJ6fYccTs+0lNH+uNQRTvJ6l1JlOMKL+vDMmSUwUyTEwg4DNmJ5MeP8zV9Uz5S
DoFpQaLBhvKO8ItE8PQLvnAR6V4itfH+qcy/TJk3U+w753UG11yVT+bknBheXuMz
wEdFWNXLMsJ0ESA1bWxdBszwW/g9vf43zWwYFivBm9aj42uTD9Zq6/Ww4GTrFp6w
vHY7fVCWqoMQoupbVrDWzQ==
`pragma protect end_protected
