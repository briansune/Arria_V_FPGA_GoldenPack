// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:23 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jMzKHuwoBbytExpNC1W3iz81dMvstdAScdIi6oXsI6sSzOGjGqtbyvt5RDm6PRE6
yYVf8VDmqsc/9jFj9JGHoyY4AoNFvjuGaIxCbYQymnii8qmh68IpJRie5Va9BDly
sHB6LiNc5Sz9UvJix/dGQiB4UQBEj84MHTszxoecmK8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3312)
tSU9cp0mchTlcTNrAvi3U0Gkv9OoFdYOdZ4kpf87aBO/e/lMp7JNzTGofviapydw
uPodKy6LNJQaaxSr6HcPj6VwVKEMZ7S2xoRIBh8qkqxKB9IWshvMDNkLTLX3vFQQ
NxxgoimLpezq+010abG+JB4VoiARTxueLEQnJLO3F5mi64sziD3+aR3AaiWZOYhX
+tw7bLQqyl7qfj/n/k7F4zFrxVPJAzuu/aHXumttkDnKGn/eoXDwVjrGz4fDoaSO
ZCIvdnurbdpdMWtzgBcD0TsYG94/20nwytRq9DnMNCTTokbBfBksBtFH68pwG4SH
0YrgeZb0scon/AWUItQ4H5y4ROde12hHvKcm7yq8iGRGLnP/wz3J5mT5ltb7ubl0
zd3P7BltfpjBMpP8Th5ZOYzZySBONZHERMcH7cMyWkJ5d9BwiIBPIAu/fg10AsEk
vwF8XUf198vDmFz2hVZR7qGpxOnR4RHEknd3TgbIswDsOslDG7C1bi4v+EIMLjPh
Vq8wtwrXrHSL2gs31Bv/jp00v7FNN7ipQcWKwo8ijjV3+ARjpJvzuNtkE3BPFrk/
yM6Qwo/tK+0z/nTuz91T3mdAeNOOjwVhsIVJL9k9n7BtBAyPER87Z7vuM1/cPZnu
5V3lNXHTKpHH8+4YT1/l6Nck8D/Jxh+krSD7cYL1XF9vdAC2MK4RrG13xNEvQ7sH
vTbiVcCDL1cXo/Rzr80QOhf6v7iHlv9dXqymAXfY7eE/J/MBJtEz6LDbue0CaKBF
gF09ClC6honuPyjPd6MlEvIL9dQcMc6g3gEa7d0Z6y/6iltxYuOGMyh7fNGZTci3
kJxR0nN9o1RpBbbh9/Qmeil9iNV5cdjmlKlxF4u4sqqJRsREIdagDJG89tUmHbG2
BpoAyrYIwGLVNMBoGjYn5HME/xtgI7HnrFm8KIctjtcgY/vrWhox1Zq/HEPQRxv9
7PUvA7RjQ+Y97JapyodIL/qSPRSX133VgTnPNBxtQrCdeXS8OeBf0aLg0ur3Xut2
NJhZmBuwtLLH9XcCtss71pkXGlnX48pFLvneN/xLMBiPaGBYXJr5EeEKmxxXWWD8
FjwGifWAeovQyYuG+DsX1F0hMEDkEfVsd/2pqV6NlsvRCzImzNCBXlysVsv3QpZH
B3fPpX/QQbrd/ZjFSwZj+zR7ygU9+1FJ0vCoDalAo4POpvCV6A71JqjwU43q9+gg
Na3C+6gvje7N4xxsBYpyO1By4jnw1Ynk3UTnhxOSsUEV+QJyLIlhANMQXGDJ6oLK
p+d2PcmPxy0PI/L65yCH6QwOHiZg71hz2+Ul+v28jpY3h3tYizi/qKYZcf5o0K6p
b19TZyIuxQm1rTLWNpzdfNmDyh91rKvq/z+hEUEC/4RLYSFbOvKNcQlPlBvEFbH9
c30yeB7fkrPrRqWJFdPMBGcxWg4ISQNMNKqDf1xmi97GndZ1sff3XVzwrnQ5ZACS
XyJj6eVHxFj+/f/gOLmM11pcYzx5/d2e0X4PnXrJQGjX+qEX0wI2sC8d5EdPVPZG
5YkLRjVHqJwfxnmWJn10k6O8j3WzsHhfkWsn5c9NSC1QgS8Leoq8OFzhKmxelysO
JxrhaGT95heR76+YALT41gQsHLqDTp2PSVcgIi79ycZttehnIVdYDmti0ZCA/RTX
ZE2UX0xfR65rTuONH75QIiTWwGPR3KtayHFfeKl+M+BlahWTng2BMWnHtBAmnugP
UCwVWFcu0m4LYZ35+vxMXgHJ/CN+uYqK9wEUntXOQadVC7krrC6crgsAIj7MPYBQ
HKHR3/fRVaOrBwtD+vd3cJ8SxeC9NYCoXB+sofNYzdMDy0O0AUvtF3TblD6bClYt
uasOZtCbLr0xwzNiSjpOA4jJ5pnyx2n4Izx1oa+K3OGgro0J+xA9Hkgn330qNL1P
CMZs1hmtJQxxQSSZBRncNsZd1WHBkiqWumiZnXDUTfUgXT77+Rliq4xX5XpdFfJ2
5hlhU2tUr8DiZIhb63pYXGC4ysEdP2fKz3LqYXNU7sPz6PX6EAqeEtU3y8FIJrXl
WdmRINhV/GLX1/VBuKzXUOEmr9zJXQa6lvYMWx9S4nNJcMqbGb8HH1+O3yXsDHT7
YeH69R5ftd41RmTcFwqZbeVdiozXOC/u+FGcqDCxKI2c6bkoEuaWVn3AZMfIQT9N
nX6HjGBZnZD1KvewrG6JUP+GfrmhOZcCgPUPHr5PxTxS1HkLcrj/LsXnaTHJGChm
8HfONr7orvAc6jZnO5XDO8uj4anxxeXLI4J42cQ/9lDO0snQLEb85oChgjGZXaiw
DR80S8nob4YHp8aQICh9X/DJjeyrWbCuYUSr3NdguAeSNVUfSvJH6SI7k7SkjUxE
uPFKKlWIqLgTWve9wmqx66FO89HtF1RII5fJct/QpslLTWIsVkvcndebsDEgumET
63jvDcdViGMhKGuQJ2Asy8bMJNNAwnkbv6qS1+zrx1vEAIyzzRlJckmwERbbBzKE
L+PAGGJ4aCXfiVYe+FldMcuFDvSvzKljCmBO2XyEzkCwFvRpK69S+ZT+nyWinz0K
jNgu1Bd/fKERR7zuOKs6BMVlkwEs+9v7J0ijaOAL4FldgxvrsweyODumQZCrmtvB
UM4q71C6k+RUBlNLRkAQ3Z+y2gyweD+aVV2VBiRyi+BVhbZvJ7jnLgV+Hj1Xb1hD
oJbm01tfbkmcZTqeZVZ8FfKHqG5NkcGdqebBcXG2ovT5K1LoZ1LPpLYaStbduxRB
MsZXvzYfmAF++6NaSN4E8KMOvgHd28P7HXtwm+O9Mq6UWHudDffgK+GOP9mqElhx
yUIlPqusLJj6eJpHvrjAECNWM4hYTXu19UHQX9NKoFlhVjpLIYv7KHuXjTsDYkrv
ZGy8jh3O2+Xf2DwfrSn7wQ/Wyf8+zRH1d6WFBIkipD5lfRnmy6Xv3Fyek2cr67gm
k5JwZimw5sSSCHYeIhZ9So2Nf1SpiXHBTzLtVrRHbQ2lya4LdGmqfKBizkXAF2wh
jT8ff7RgJC2i1WVTrWk/XL47+Ba7H+e8QumDi/V8mQAxJlxg/BPTRGjRQ7YcnP3u
gmojSOegMRnkRnDehpB/oQ85oO13/3wpQXIQ6yr8x82OJV7uANq3ky2w/QnP4/zH
y12WtpJfZ8RtRN3xC7qt8ByYdd8Ucm5mj3bXviLTYzIBTpQuGJ7ChJB2myqfSKoJ
H3NPxrnDWVjzxnUzsE2i6KkxURTT4DzqFJgHu2DWyKG0erdSO34FpY6cStyZF/jq
iMyAgXJDzQmh3cqfSR/2fbvN6UXNKAr1EC4SYMDfpSswIMrZBAfvmPR+UIFNCxxs
hAQfm4CqnMTceKIzZy6MykHlp0DauSl45RP1UwFwpXy+0HfcB8lcyku1KedtL53J
PZRYpF+BIaowBXwT0/0bBJd2ihb321hG7S7Im5IRyOyCrzT85WiBu7/wpOX927uB
F7JGX3869Ibtb2s+9C4W35qJEkvVcW3tE/cYugWHpE9YghMBoxn0pwJRyyydXPpr
HzA+gJQxtW7pSEb+5q8D430aLwnSYJMgJlDgU3O4z8Cwy5Ic/H2b1AzhdLXX7M61
cRLAl9BD9WNI4fmOH6qXaGN6t0TYHSEod8IYHr+YUWiTKZQYyiD0g0XwQM6vh7j/
sQQIL/yTPkvyu/P2y+SWV+0AoDrLmK0htfqTDcYmTwwvWzNwAgixi6yruSuAfxTu
Qn1khIyQ4q6YFZVg2YfS1Jp9mqlWdsY39Z+85UwdStzXE0gkI4VC13CgG0XXhnHA
mGeRzqdM+mozy1mLM1gyUwdSDykNHqfeFOfrf/28elkSQNOebCzx98A7IzvvlQ1W
Ukwv+e32muCZRSiw8D+OcXrLLO352waoO/If8LdSstLgsLvAw/1OMVlv/KBZc/Zl
nkgp4S7GVl5wZkibmgOrN6cFaz6g51w3B2GEGP+XkwowHAFZ0RCy6+ftBYqA/AB+
qH67fSoVivPIR09Zn/MFuy/TY1b5himt4+yAToM/SK0Fq0oRFS4PkYjTdBSgtVeU
liXRy4+MeCxkw0F6DDU8dDEQvGaC+Sst3K336+IpBM7L5NdyduT2z3Y7X451rThL
8Sd282uXXh411ygLByGIp33Y10nuUwA5nD7NBGmRcwv1qROBgOU9pve3ygPetfLh
UAZEwYTmoXREoN+iq1JNYeulRTA8n72/Mka5RHYftPOL7fDCR7NrXchqQHoCuhyz
RVhZ0AYV+kbNfX1h/bDmtamv7wP4f0rfv1CL5YJ/MFP1Hl0wabeO2Gt1bRybLAU+
ABhoTLZ4U9gGCtXQbcXjpJOdfCz/z7XtIesVzNp7xBKHPR5qxY6bRPAX7dhySUqS
oOK5Ge4lEZmHJ1cCUFHFu2ZjDpuXqGxTSTlO2PAWGaf3xq9BqrHBb1EpsC8AEzZ2
`pragma protect end_protected
