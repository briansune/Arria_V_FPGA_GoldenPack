// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
VrBT0FYSNbeTpiHWLMX1qVBGisf3iZQRyYQh1rc5EMFKHVXG87bpIuXiYo8o/qjebswRDaKM/idh
krfsUG3bxz7Tp7BD/KCUddCUUXHl5wPEA6bzbYjjKM1lN9DsICWgocFuY+I2/AOlb7rK5tAe+KUR
tW4Ta8P/4IFfiqHqn+3tlganvgH5CSU5rUQRG/HH2RKNqVZT+ojBiRrPZn6NvpqN34Z4EIL4edUF
cTHVugy6mgIfeq9s0fc0h+OJOc5DU/TXb228lhd918cuPMyQkiuDXChLlKlwgHjhHxqSlm7b1jne
zsUd2feIib9MkoGYAPFib/VPh7wgv8kpMDHbow==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24208)
ughwY/q6TtfA0Y33xQB07wDiyzaiOGaB5C90iYUiDYHtZWFZ/SCjyWJX8y1mDUuRFOnAyMcacoh3
jq7J6+bHdUrLH6WM5HHGlHw/lns6tcB8OE52zi41VM6WHMl/LXQG/BaO/yrjMqU474qFPJbwPITM
4IEisQavrwnmRXC4EqiS+LtJYulpbVs/aBxji/7CqQUXY0cK/W3WN2hGKQ/kdG3a/6ZQEyi+M1DY
2ia/p2G9Kd7k6fEa0lO3fHds/ADIkq5fQBx5059Ry/J9Bp5pK9gDYWmUOJMChMB8jz2dIR/P3MsA
at2mrZlqFwI/hgICWMZ1og5ObV9M28FdJ1y2ye0noqNb/NCwvCZe0Z83pw7tNjD+VNnhJQ4YYNNp
tlYi+vH7j1yCDA4CAaq5Lo45pN+XL0Rr0KZtHfKMyog5DooOKTjNCD7yd2JwZ6+H97ggrplNUMxT
1LQ7jZiMDLxLPVZdDjyJ9prAkELNGmfSe38NpSyTTANaiOfoU1y7N3PC0LPiuBxsh/233dC30te0
b1G7trEC9sO0vGT7XfDKfdHo7ZgH9aD8rQMhLacdn9NPJTlckrgK3kV3YNguMHQGkhpTmUKgevcl
lAugrosxqY+lyXWpJZW2HKDTvJHu+pKN/QNKUktovoyLTL/Hr+vYzFoekY0UqqR0doWlRTPisEGx
vdTtI5BH30dXceKDh3/Tr7BTH4CSb8ExcoTDqrYFSbg6RWlQUP+a3uxReP+SGA3kuBXsuZAHnvJs
auUFtX7TPNnal/EGzX1j90htmTug27FDuwyx3uTYG4d0reziQ6TElS1mrIN/xm6FqwFWZheyRuw6
bJTgGESaKy5BtMmWPj7X5lk7b+AuNYFfxgfBjSIB31uRK0JF+sO7WwtLLB1EQTKzKWXvePjZA/Re
Ang2040z2/RXH/hgmHm6fSkuDifnd7xbyghE0BWRWePnZbn/azIVLyMafX+h8WbDkirtRVJLHQNR
Opof/GxQ2CBu2DuFNTGTN287Bl1qRu1NfpJpY5Z/Cj0F5FFlOiVCe2eKldoToXodfDwKgWInrbQ1
e9SftHsxAwZn7dPgtud3FgyaJIOapC5A2+fZx6sRUjNww0z2LkbLr/l2DPlUfiEpa5yIvqhZNX5z
Eqw8PHO5ON+6PBnRphzl9PiKki7nSpRuwKPVRPY7arEGzRn9el9JRExsfbDLvOoWWNduO+KRepBH
daDvt8J0S8TKlIcbl0StXqs3n/Ta2g1sUjIKcYLNA5G1zB4n6Rg5lUnY070vRo7Wts6t/bqQub8B
iumM3lp6h+eazJrBlf1u71Dyi3hXQ9LJI/HYx6aAsGCk1vExUC5HvLcUa/bHNZGCrEIkDdT5UXTC
+Q145BQmL7LnSQR7HmMKyYzPfDm+dtgp6y669VdKQs2uZYBPSivD2EdmvZd4aYEh5c6GLaFg40GS
EG+ZjhgHSlcTstvKk/56g8jGeDDSUzrXZBN1pcSOsBZnNI8PqZV46e1BnN73YPRKkmj+Whx2anK+
RfE366jG4SAWC9Ew5fTAllP3UABBMbqp/1/Rl6ai9I5MkauJ5lmNwXDV1/f4Agc57+tmxeEScuSM
/svikxbkbdTF0j4agApVhIsx83SUlz7PDm7AZAN0G1FNge6EmDGarvnPIrFEw2l795x2fMs7Hdf4
z1b83LY3wmMnQ32a1hcB1rLJ171Cmq+jg41fnuqhk7bAw9ttlmGITYO+BVy/aqBQ8mCHzIp0AOeR
n1brztZ59ICObp4pEthMTYXu6c6tY0gfqrhZQtrTmuVNOw/f3b6b1AhSF2HUJj5fTKMA7uwFhQKP
QF8yAUfTS/HjiXlobCy20rVF27eGCW25339CKgxxuOfTxWan4QonJ90JhZmbmTuXsj0/VcnzBxsT
BgrA2MYcUydr5bH4EOF1afZ/ho3Isuh0SUj43jx5bB1fk2S8GrxIjUqPSy8uFIqpiP+0mk90bPCq
ra3yNjhsDqMphkVIuT3eQHSI4gnXdwn9SqCLgWgiCiE1DSphENIngSUHIiNPVo/HlSa0QHn6MUG8
TFSFoPrEl+Jr2hGhzhnocWcTJk0fAULRBquRMT6GnJ70kVxkxV7ydqxRs2VbY3zxEg8ozU5N05ua
TFX0zVn4Rw/ursqY2TKNG83hfJbSo7gp7t8ZdxZetRHR/6+Qi8yL/zspFk/EaX6bSRBArD26srKG
oMWq3vBK/R6+Ck7G2kO1yE6qYUlpcpQc+sxiXeARCxDjq7NA3eR0i4C/kNvE/2vTcrkb/1b1X6Lm
WZ/h2/tuSr0MvVFnsNbNfjKREnczP0qgwta7tYY2u8ozYSOgDo3pxulGsv6HUUzpEHQcNMsSusqk
841mr6z0NAsE1/D3RPhc8qdWpiLBYJ+1u5kZ4bxCZIRW1TJt+IMQUk/+IXltprYR4VK+m9PogjOq
XEJ22a1WvcF7YiJv9I25JCgfMRkjt8MHJOzwXwtja7cnOwf8sbJ4W98C2+4wkMHYrAIt+sZ6BzlH
8GundRc8tx7R9SalygrUItmHhViuIWPrM4M7FaL10j3sK70Qx5G/jVYzq7sG+NaiPKgRGJFMT9wN
y+JTAGp2UhK8iW7EOKcmDTyXhZyClIbrduocsNO4MZxWzYngkpWPxJ+dOtYdOiTs81nGO72ACvCI
g0PKbRqEfkxOKkEL1rGdd6+QwkCyRPUQybKJ8dyg+CJSmvqN4ZVsNiYF4nEyW44DZXqfWTMNwUad
izD8BZ5ffCp6Tdcjo3o4rMXwZFbb6XJq6ZzT+nyvvk6dghSkTj8Pch23yIu6CoExJSg1MPyYVGXm
7VLAFLM5DPhuzOK/cYPt9gpoV1YwwVKErDA1TaF7KuXFU0Sx4lz1XpmrlzmVL0ME7ZwTSMyljg9e
19xFaa1IGHwwRD0aoniAUO8MUhSvwlslpBadkbWG7a1/Jx4w8dxVBOHhGBRkaaN75OnQFEHr6fiY
rSOnCLqiH6CoO10d+YtRREWKD26NfYSBa/3ir7rtpts6qKf9AihWDt5DuO71d7vFUef4IGrRMooV
E1sF8u0qb+2gbpLyKT4RTl8BFkVNfK3UU7r8MNGN6xSLnE7TYqvEo79BnyS81OcUIKptWL5J5Qkc
uYWZNtZTDP1JfUbHTo7ef2ecA0CDpS2Xp85dRF+owej/mCKsLCRAS8Jz1yy6VgpgINtM0xnS4jlK
i1mX2WARKFPTbEhzybQNhthyqqtfKQ7VUWvBYenp8wLLXCv3V1xSh0vRmFyratEcLIZj8vw+9siT
8Ra/a/ABd4qwot33uWO5hqYGG5d2y0odRbf1vTU4g6MEn/mABe0QsbvxCMyi5aEK8o3ZfoIioZWz
LdfoI4qqghA6CiwQ6kAr5A/sVN8dY6H5Lz/xrfzgp1MvwYfZLEZF8OQ8M0slOCfNRt7kvLWvG+qM
tt9FEzNdMTYCZcw8RvG4Ul5OLEx//B1jBKj9AkIDzPxAU74D3ZJ9Xk15EY1xKSk4WuDPnVPKW7nW
r2rEyrhG4wmvAWoYIkcgxMRmdfFU6XeVnQ3n8cmNu1RnRf2GNSBmVyXNHnYPQVPSAEJCXz/EgKOw
JLhuM2cmG26IgbHEqEHqWYBlcYdX4pRNo87DZfKgp4iYzmh4PO9gHHU/Gfkbw3+NsicOvAxl/Omo
e5ER3PC60u1hw5lMr8MP1r37pI8BbGG0c9KPBCIJ9oXROY6RNi11h4+aTRt48I28AP3YlrlfoA+w
9l4OBkD5NBJ4/DNnoaB9CzS8cm8ra1u/7f7mH0VafPrwSNZMpUUVVEN6p/GdMAiPslGjB+80jQie
rxWnsMXXbwSGv4E1UGnlTLwRqdnLTVBMI/nXzuRVpjDmNZ6tBnlBB1Wf2Ni5nVt3Uu7Y8kEgrdeU
0e32oulVe4dft3hRSnK5GDRJ9Gdg0Y6S7SMqdA+WRUUm6aHoPFp7ul20plkGLp3f1LHQeJ0lCjOd
iXOFICl9Hc5QB8cB43hSVvnpIt8qMrW1JY62GQ4eSKhunUgbl01uRlsvCnZ7KUn9vp1vM5ru6wGU
G4mhhY+jM5kI0+70SKFSNtZZ5K8ooUFWG9nthnlHnT/n6flLHjzTxMnPioo8lexinhNqC9quvFDf
JBosD9R+PCuqlH9SzuCMu1OLvhWAJitnIQdpxu2o4t9YC8K5OmuVRfIXgBPAi3ATgRRTW4pOyxd+
NZ41Q146ya0iDIuLhQQ079uGizGt/KmXW4RCb2KOjxfDGYahu5hHw9Wf5QgtbYtSd5iMizCnBlrr
yDj2EKkIxWc33ljsF7QhXoAiofLNcOFG1kNMitU0vEtEEhRrisTnxzzyEi5LbvSskiJvMDwVg9Mb
fFPnonuvkrWnLjjnpRaREqBCfHXHDBHC7Zsfg1PlqLvFQeMgWTJMOCPmek2Cxlh5LXXOSHKNHGkw
IpgqJUjFrAAS+2og0yuY1vaBTYlit/h3+M5lsWF+NDFJb3dvgC40D/6pJwZ6TCTGi7IZiInTL/wX
YSqpdpzZljcsRJQ56kUvoh8dy3rZ0LheRM0bSwB4QITenabkM+X/6rT9h38+Rv2u1OY4Z6qOQDyO
ImKl6YK1VbcdSN9J+lk1FYCKH3Wbw55jNTfwTW193qoIzBcT6wmkBf5OcvXZ2Nk8mA+eT9W1AWvo
EOsDr/sRMyfQE8ezwEJiDIKWS6lU+t0SY6l7GszUmzSxLnsXJNtgeBucQ/yO4WIx+GpSS0Q4xfSL
ICrF5t8CA/I+dHqACbj5jK+GdR82OCcf2LGC2fX1Wgu9/9LPZLgnHlJo8vXXo627VLoGenT3pzAp
lhBDx36oKOT31Z535rKGJoxQJN76zHGIfqhvJt2yaMhiCSO6CFeXLuoiVsL0XgpYcX+2C0NJQ0fi
XV6QwpyuTAWTQWfe4eNBg8hMD88N0nFi1hkrxKDUmgNlbKeJmYzeBs5dWUCEovi8viQwAVCBSE87
m1QddkWN5mnWDjGOmSWpUQ7cAEBNXqrzPqxah/Cbctq9ucPPuUedv7VEkq6WCyhvTrADPGmaEOhN
SllyqcO5uYt5/H+nisEIAYmaa+HilY5TGahn8+kah67DzaiWMXdJ2p7nCH7XvDZhMHCl604u5eq7
rKiqRdPbrtRMPbuPLaQXMByiK/OFIEKoEa6wSew7slGTOEhK3D7x7XrtpHm/XrbHpweZkvFXkkbM
cJ9wtfMA16ief2MXZqh8w9MGUvkgCwOGkayyBGg6g2HAC/7L+2RXW0BxfUNjYNdgZJuu1tF44yI1
Gv50rbG67uRA91Wapxj2KJ0ZNOxYj0SvtI7YGSF9LC594rzkPeFuBD7KfF1IOvecJsbYEVqANGg8
nquGY4zG8P3nC+bcnbSgZPdNZPz5jI+8kWM1DEThFlGEZGqkC5jo5YG09fgR43IxvAcCKasa8fiy
GFJjfnZILSREcYlBDu2aNfKZvR0FOnvdRzOe7rd4RKWK1DARouinbJDPkD5HQu1f3z/GACX2iVdH
HknZJebd68csJHmbNyUG8nOFqMlMpF4cPmJVWhpQjz0igVSiDTNBJWjP9uVD15DOeRLQV7goxzwx
t0OYs3Y7qofbiQLhLYMnV+xxEslB182YEB01KnmLM/zS86G0uixdZRRJ/c0pWWobvquYYi3wP2OX
BJtthVS4NE0+WbKKFp6yR9tyUlLrmsA41095+pTl8aXHNnvFlruhxCvnYN55p1GugqoPN3KvDgO+
kDbeHlcvNNSUpV8T1d9ewLmx9xUBYX6KZ9riO6PRDOajVw+pd6i8XqZauR2dEYDsqCBbOUWVHRoL
I01G5U4jiX2yW4OK94tNz3mmVKNd5nX/KWt1JDCQKUKyHKMpoz055zt+nnFCnMpOxqG16Fy01T8F
mq2Y4delG8A75FYnoulgA/j2UuxhlCEzwtE+GWEdDSZfe00BYX4ieGiHig4hSSqg4Qc2fcGILq6+
hqb7Hsfb1PZzkG+xj/ZK8ov/30WziawG/G6dtOwROr9OlW8GHRiscimnXVqY4IIt6cwl9nMh/jE3
OZQe06vfMv59HAyPtHBs59Pp+cM5ModKa1X9PtK8JvyxsbcGerj924PUQvV0XBqndBL1kguynwIW
IsAZq0hsDkzx21zzCltcwrZg9AhbY584w9aj2aAbHUEGexgFSja8qPRpXryEEr6C3ByGrV2UCiWQ
m4uJEhcaR1lQFKOLHhbF64Uxm+Sy7Mu3x6/sGictMkDWiCu97kFvsYvWIOilOPaCLWkbFGL5AAYN
VD6oxJvRbBlTG/7590noQTOyPxZXOSRDDp3BKdoG0PufW1VjGS3c/vsPjMaHIpwWTiZWVSfdnpA5
rPTA/zCcuX+s7L59D/DOZ8zep8iZ39sNGnQc3Zc48ZMbemHRK4A0AeFIEE+0V8iXZYHhFWyWl0cq
QSwQdmk8BiOy899ui/0xzqSJT4W81XzmPEU6TQj2Thmk3a4WtNLHhzDRzk/bkBecRBrLnO9fBupg
HaBYh0edLO/z71DpotP5AOuFTVbqUZUyopF7uLgGnkNfZQy564H6aH55JjpQg1CCME42RhjAD7oC
KBM7HoAUHqBOSSl3ShdBivMisGNuHUwIu5eHmgr7O1i5hRdvzgHEkTb92KOObXaQsP8iMTCT0QnG
E4wrwrH4uKvLKuSEvev5P0S6b4QCuGJXCkJBqvUqjK6GLbCUiz/Jl7GHrFPNEjcRymjW+3zCBgyk
oGiwG4kI+hS04KdY1piZ14xDFYJSgOPNc4KDWDRV9P/DqzXzJryPI5rjAxas/lqW8EdRVMxF6nZi
3PkXMHr1+Esm10SDZloGZpygwrwvUpUKRZCfLJ24Us9MfBMzRZNidiTe21jWgjx6nrC3WT2auIeZ
WRwp4vnDTrVWfTQa3qNzeiaQnd1TJDoQuyD3/+DnVU8Imw7ijy8ogMw6nQHTXViCQSykD9P4ur3U
4PmJiW5UKOx2yrZj0qVrbz0BxV/iYSgCgqQBsq/4DmpJAjakTGb6uTChPfKIMVZV/UaWoRtiT7ux
y4LdEtADnhkX8bclxsfhAQDwvni+VF76ejpgu8j3+wkCdyTvB2+DcF7uVPh3MNIBFr+/kmoKib/1
7KhLRkz2SH5lft5jmG3KGSgaYsYWNzqBSajGMKroJNfXP0HSO3laa/RsE8x1Dwn4U4cW5ryetRyb
j7wWu1e2LUCO7yREdrmg4xYRjwDW5/mX62CMDFJHxK37XJZ45D1LeRffMIk7Y/BI9JXKlX4Cl7hw
JShWnYMDB/WDZedSCGmZET0cENZYXBapwVplZWjRmc78lFytWYcbbnCL845oidxd4FnDTEKIlHBT
RAfajSWsPLl3XcyGZuv2NcaKdXnm2B12EWBzDtnG22lIq6WL23XNTDZ9FIe0HX4zS9AcybrokBKB
hv+tG7Q5wpn1y4Hn7isvrCCViEx2M31iwNck4hmAJfJXe5pn4G6Jo7KOzTyW4Ig8oUwZNrR63fqN
16Die3jrpDjTLPSh0EDeZ5d/TDD3/WOO6jLVA+8pfxO6bo534epPC9U7aoGi+Rud/jmFliiC6yXm
grtuL2P+JI/GWWHUMfbPezhDGjK1Ye5hu+FPGrQzPZxH/O1pqrAXAJdx0wyRF3pmhHNu6nIPY9rY
BSj7BUF8nO3o2Zf4Tki5G88CSFymikgnbS3BSUjcAnaE5sijKVY8A/iT2eO5uUCwDn8JLoLIC8ak
6UJLzlouEpOLexz6D8/t6oZwn02HZ35AUUuTSq6SPHcfUqNJUZ6HsnfYzVNoTPhkLmF/Pgr3lg+E
gQLGWQ0OU2Z9RVFfSzzrjkGdji37uZkTv9EjmRWP3BIISuJIFwoGzveMgb0WpD02u+kneuX3FZz2
E1ZoMa2c6GpUFiam3lYJwP1qglG2yFLAn/+kiREWMyparjCvIVRCisJ5Eb5C9txkUK8ZWvh0kRj3
2/n3tbUQvEkLIfqnnuUqx7FjKigL9u/ZloFI0jgmWu6dbTTJmTfgg4LkaPrrRJfK39cNBW4vOtlP
zsdBZAOsDNdzUTcZh8XNsaOlXpKGXokztfG6I0p8xrlkxI9pxMp3wDs5iG6e/IIxv6HbhxD3hc9A
8WzW5ltDKMVupFSV4dhmJEJeUH0LeGkMMNCeeZ9oLEiyBwbDVp5zuNnpLDfsURfQwCoaQdPPLQJL
15rKyqMaKMDLDrguxWqWZV3g0hZfsw+uFOLTN1JCeaV5/Sf6EUvy+5jot3yvrATKEaKAkeZzuMNN
DR3TZViKL4iwPsqSD5X/jkO+1+Syk6jEH1lYv9AVvYpFEuQCZ7893BJznLGd6elrtCnklscnaXCv
Fu2cUZCtVKsC5a4ttHtYOwPz3CE/J4pO7jrmoj+iHsvL31+ykAG7s8ONREBTvMpnFwe2BM3YbBZT
slNPLJnSvJAmd8vS6zMyA3KpBKDqW7Z9bxrKRch/MowCs0zFfxA39Y59UkSXdjZHYf99G5+gUEEa
kF6dnqARqVIwcTTmiC+4LZgpE69vq/FQmp5G12QHkaxY95nQ7hBen8igP+eqxK979Y0gxtD6VcdK
u4FlpYSgEfPJhwbk0j/yDupQ2wXfEWLOzFrKAqtbmiegylkJ+oxMMzK2CLv+cTlX3BOEPUZowu/+
iKL/v5cGV1TF7lkfwYJvmoihRAYVFItIm1aTkl0XZOsHcOxhdD3AkfO/ytaDPuGasRuhHngMvtdF
jHDuhI9QakpBmUOWTKQS00Ny2KURYWRbKcoorMdIp7Rpwunutz4AlfboOFYaCzpVfz9mj8tqffWM
IFYbDE+OxCqv7yViJXgkyrg+wtYkPCw4UraabN8aOZ8je2Yq86EYhWCGak7HPh3x3007m9H3mm6/
feaOe0uYcGmLR/0u0+Exkuf1SFOAhQvUhvEyCHAADQzHRT14EsQ3wfaJTPiN8lPq82IYx3PROAFE
4jHDnSV4KtPrGNLOOWHWfsX2afhsYvpeyNLtiUc9Qb78YEtzbsyDVsm6NndrSccOMXA0Cc3iuZAL
oD0R5TW4hnFipNoicZxwgtU2jRwnYthEzdvcp176GPtG+vANhs7nPQgdK5GASx3OIzqGIgbZlxq+
3z5LWa7z7y6q2lghS/JGJ6GneFqdN+Up6J+SoreC+FOkNoile2XPuIxPRIQywll76eLIXBC+6QyC
hDvfVPw/ZgjfM8JB4I0DNojUncHKryDXlPjdfNzSTIx+YS4vyk/ufYpGkfsV19sGq8764qZU/Vyh
4YE2ZLGkFlEi3XYlnxs9PTWqS7qg/Fe33zYGWMaMQt3IlNKB83vhup2lPDe4B1iqy74VPs2xMDIK
Ed9hao6//+pTYgvRQAIVo0uJEryYaLKOMoGPQ4be52PPbNfgMKhCbtSOlD+MhcAL3qxOXdMzI582
LttCCC0xXktYEoDLh5naCeyDyzkCo7OPvyTegt9KsaXCJQY3wWcG7SymuCCSmuyuk7e4Rq4LbsP3
lguHb+3D58LSAqdIctd0b0bE8KjLnqHwCC5rhhDwIzPS7ScwmPspHCApVYDNqpKrLr4FHM5QcfVb
BToGeP7UWLHFbv2D9NQF8U2KuzA2849K53zaizxtoENfnG1oZU/tkTNxi1aeGm9r92UQB0XMUPVN
iQ/DBS3utDzbhj4orDG8DfcXtWk+kNEe69wDBtq8r+9sgx1S6U1CMbV2bMtukLsUqyO4fjaG3ZlD
VylfaqZ+DXADKwXVjzOujwDb/aoGkZN7eEX4nvIe4O3GP3HV5UMb+wvGyvPluLcuLiKpYjbP8Lpl
9E1olGRayoT1dOMmyvoIgxXLaEFEcnOHHJdAnJ3Rnu2VjzdmT4JDTMKt51qKvjyOGf5yXJ9aNBan
yGaX+HyqrQTEIJGggWp3qVgC69NS5Pvcdynztfau2tWZ9JYaVtlL+L3yWX0IsOXoWMMiRFe7rFw+
dA+hvfF4f3rxIv+mMs1CoF3ryZuAPftCGF3mR+mr6Z1FAzDYkSkRx6gApW2n97IS4SuqVOrLcM+j
mRcEQzzabczudvORdh2EuapQz8I5jrttCxC9qAzkI24h9dZ1amEuygMeRg2BHuWWuTUgPH9/aPwx
6Hzf4Ou1OmGNmM5DqeJTOzbtB5owAaePlFgwAmAd/d+HuRrgaPhBbAFuugohiTJWq16dKgmPwtaG
r5d/OEgWfb9BBaq49mYWBDVnj3cOLxhD9aoZRZO1uJAlzyKm3fktZwTP6/Qry+xX9CoO1K41gdCT
NBKZWSnfUHprQK2TTgDjEGM8OSU0yT+kLeZhXU/d4Jm/BIDKQjzryKczBqOHEpneQn4txZN+lAiz
B33JeYhxSSBTOezJBsQx2U+vlYxBvTDvh8Wq2GpVnLBUVKVAZQhH1gD1Y8cKuNw/KrQzbhT4drry
BgYg6/8TNqDe8lmL8vMeKcQ+AEHaCUWfSx3nAe/vyv324HXwAGyaoCjDEWrcYrXNe/rbcNKRoJiY
FpVU3f6WzduZn4S1EMxXjpFfGO4qsYiRgxoxRMr2V9Ws4PrAIuqpJn/6pWC9EsZ1ZYztFvV9YpzA
Q3TRpelR887YcD1E+KiMKGvTHR+awcoGOSRpmhhrUCT9z9T/p7DbHcRMuIcgHzceqi4tozR4ctsn
b4D9qBUfGMP2RNfZsmeVDF3ZfRgbjyeiL7CpWdj63ze6B4+rVWlm4gE2g1vc521JciIdifhgE+Pu
z53Gj9VRAH5W/wftM/aaUcPOEwb8nGrvbqgpkDvMANH86uhGqArzd0GZHho37pO1j6tDBFi5/+sZ
O3+WyQGuCV5551V9OjTPsnM3SqOWF2blYXIRS2wI587E3K2D7c6wZsGEkuViHhjNbekgeweVPD47
lpuyisrwTho6NOOkoMqym3qZp5BYJeEHkdnlYVpIlE3UvfnOaxfbtFxf/3Q/+FxnKwWcvc5a7uC6
H4qmFk2PjQAjHDTK2bDkBGZpgPslsgtX4/vOqLA/FTOj7cylsAb0pRi9LzyfgiYqbUrNbtsRqisI
Kwt8YI7pQNmqSm/HaSrTzPZc0dCkh2l4ZU/ZmoNZPVUGsrXK9LTpW96xxN3fxoiSD2LuU8FfCjfu
n7XhSmGuJ6sRqAQis47f5/vQnp7AmwWF4ARTjVh6l1aEVOe6qVxq9HFo2bY+Bc48dfdIBh9DBPX6
vwYjEkb2jilKQyGFH9oXNvedbe6Pl5ebuMQoID7jCuxlxpD9BCpvxrS8+6kHAdoMqmHXxusvViZF
YPoyriU/HVbf1MFlZus+Xo5DOuBL+rMVpkwcAftFXn7bVAx1jY9dkVY50C1dBH1T7Q/eBfWqmzEV
0ltfOjXjOE65KOqKKjqZ/0mJKfFLrw4pxvIX1/3toUcUH3umboaRTwPa8GUxUHZGeeUN+GcBC/IN
UPd7UV5/6KeOpbgBwU+PZw5pxZVLqwL55JtB2bA/vK2WoM/NKKJ6zpvq4ngPmEnZmCKaib+V9xfi
INNaG5AVZSDRcLSDkMHnb9LOzbICBXkaesoQ1MYvHKfrRhzIH2x+AI7jPCeiFTfw9y8+2ducGiTy
d+TVm58UXKwb4yf/nd6q5m1AQtd62fY4EK/pPSU1iRDpipTRkDRQwkGo7kZk/4KSiRonIbEmN2F0
7s3msZClnkgcYjuxBL8u1e0/EbMqQlKsMHJ2TSJ3KyzYqILuoxS773AtiQbRXa+eyaOCsxNbfPRy
9mtfDi1ER+olXpHRalBrMRHu9Q+jrN3cpY/huk5ucFbp+/JPh1nCeST1/pKOXMYLMYEUWnGVrF0z
jpfaqslNKX7MPd8f2AAlvPCTyvx/M+5HhCudKGMmBxtP9/mMFCBPIXT4agjZe56m6Y3R07UoMpKL
z9Ha5AEOlyzhiJgoKcnuPXJQyTA8eqsEaAxBff6Re8mIp29Xzl8IB0LnKMIWUgDDw7pcj03DMo1e
dgF+6F7kqpOEYeJcz0m5dWZC7jbNVA6tO+Mpf1G0tBmKhg2UDpaWMc0VOr7NvSHXGRWOnDIHxBYz
R3dXpsoUGuc3EpwuyXGBYv68XQsN4XO+nfg3hK2Y92M8OyQQOQXDIecnP0f83DCl0Shc1X7ACaHR
jHi+gDpBo4GLCoQbUvqgZh7azYtUDbi3DZeUVbgs3RySRGcIXJekYX01gyyICA2t2yaz49pP7u6E
NPckrcFpKFMAbX3XG2V0hr3gO2PpF/dcIL6jzI8PHOdhJGuCJhXimg3WO/Q678IbLYtabBDOt2QR
fwbLfqZwVw1fQ/qN5sKFR2YIB3UsY7CNyn8NKVK/JpPHD8KgfFrBN0EXrAT2AcvFYPwqRNXAtFdb
VzXBzuEz6cLAziKfQO6Sxe4Fk7m4cQb7MOqJO3453aF4+uXST6OOSo+JAjcTfLLEJq1K/oc7hMCB
rxunxyjmR9FfndWjS/sAvvwjoozwxMvjeNn9jag3rq8ML3MQI/7IX8yMxrKPdYzr2ejTQJUtjoMY
jaUCtqDl4yzTiSSmWkHz5K1mEQ0EpkMdPlIKatrCLUz1FuvQGeq21aIuIo838i3R6O7HqVtRUTSr
6Q8+PIeNiW4d3TOO1m7xPLjbLTTLfjXV7rKvZoiIJDbCFCk0sonYGiiVLnP7tYUcYwIH6MNFA1UO
NcaWf+n4tMFSDzJ2MksQoCWZjdmdWU4+xkQSaD9Rz3f/nJnHTSietAVwByImegt8gBcj+lTt2LmU
MHybqJ69UKy6zx3AHFK0dnWqRZ0SnC6zq25uWl/4YKJAYThMKk9Di+7awitxLoXAzVfsXfVySdj9
pIcW6Ea86/oHykW8H6+uh6hTIOO0MJi6BCb9baApSbcWyalWKAPfh2HXN6nSKKr1uQTHx63eur2l
p7HuxBkwT9CfBdJC2GWz0c6CPvx5xLbemp2u3U0mg32DCXTgU+wjP0mR7ulH0jzFawhFgyYgZS/x
rLJmOSsCIUFcOGQyagt/TcQhw9jNnTSnDWoT1y/91rtW8G2GFd2Ifhb3FfjaNHbteGqQljaFBMV+
HcbH0ggUnKtl+x8SKvvTHtQ90BAd/wUxpKne4p5QTPrFZLYsgMAlKS53udAl7Yxx0vn9Rj++EC4A
ha1XbyjJhwp8k7X2S3PZt0yP1Qsp5n1yv9/Zus2FHQ/TTiwpRSjOWxh5GuIcLTbILUYtwDCafRBk
EOzFXWx0rPQTTWTWMsopM1P24xT/ua1M/dr9vdAJgXNqIeJQaIWTZjCdMVPhTdtqAtdwYGxkkh1p
QQcCqzNMz3vK8v/HiafyET+TD9A5Cqx31dn1yIQoOZMvccTev33Wx2Ljawhc3NDNm3qREyHNeqYH
8cyYbjWzHfVk7DpvgWw82hJk5X11GshEP4Ty7uV/loLqN2eGXBZOXUrqc9TZxEqJWa9q7Up9VaLi
CouJ9NGsFuQTSu+VI57zFPS7TGvDJyQwgqk3HafBYLGquwvR4Xvg6Lyh8lk394rcEP39BAgK7DwS
j7KTi5oJQInUnJgntChBy4Wa14Y4z+B0OZP4PWp4dZJQQ7JSbaTYpNg+Q82cCUxWPCorjgVJSnP+
UXHg70+qtcZzHJPy2/WskSRgU8NWKY8XQkqabe2aQGI9tkDsG8D9juhi7SfXxKZpKM3DEs9ZceUE
4JncJowQQBlSf6Thz9CeIMylVYjd1BUn2VBwpy6Kg0mySRc2Va1wHsSmKVPq6PsEGxqXIU/E/RXU
PCi8XYxaz2Wg/XGLu4V4x25q6+d1VPTgoVt0IoGDHdHX2CxTp4oxnb4/p0EReQ889B7LMonpPBnv
DlB7wL0iKyDgBzFCtiSvmG/ItovP6qGBCKrpRTppX73W80rUi2NTHgj48dedHrZgaoKyX4R5HF64
74oZQ7cSLXVFn9iC/hBI5l6TUqjABl7IWC7oiv6lNp42xAgDTfv60VnNXDvzN41pNg2CXA7FeicM
E3OODkFlH1M/2wKkhusc+U4+9gQmkjqfo+/65cyAhSJuZTpFr6FX+hwIFMmEGA5Qdx1WortIXYU9
PYNeX7nV7UeGFRrROQP0javEF8cnaF7hzUjpRYv1IZxwy7yuGcMnEx/zyx4lWtn75Oczz7tdQhP7
hWH3ST377hxGdsTWGmILx7FYe0WYztm+05uwDRapo2fXY3MBfVtJbXvL0SjBCX8E0x3gNgZP2dqB
v35usyCGkK+ygaE3SHyQh+8pf8Mxr7e4v39Yxr6BijkW8MhT5RYorzsR/F27nYvGcZpTvnWyMeQf
307r49EQXlVPModoVEeQ5+CtsevIKvsu0GKqj5xIKofSPvu5jMI4bk6Mf/IcfIuyyt9xc3zLnxOL
AG/qfKAjTAAXtL71hGUC3p9r+B/P+YmgEGycfbtdEoyrc2U6++sYKxmjzDtqd+nVQyyJ77jbUbfl
J7kXqoChBTxbe6lvpK0f8GExVxgAr0Z+K+ZzRyvyzCPwETWnc68qIfLa8rMTzwyx2Hqp6CfPVh7m
xQ2maZp+1jJ/V1m7+1pwM64WoLF27n2/eGWQVhh5yaVSsN5H2t8JaD8xAnm+pTVfjpNDZs1uhoTV
x+wMFpTAuYArAIshSpbYxzUmDXyeOiM0y7LNe8HLICujJvTjDuuAIoZtdVswm2Z45VWcFS7sNVyQ
V/Nwam/qJhFcZO2ifIwOZYcLRLnnvpXiel9dIdWbNgMYHiw4UCuVlPRj/bpkkvX7n77hIeC4e1/5
dnE8wJErG6/dplE28ubPpv4QzPi+XIT9HqAp3c1Fp2LNyQDf4SKVIQRX80DhtqBcNCUpBBYiQaqJ
Y+n1OKVlHTramYXuQNCsEQg8AHdZcpdP9WIJEJiXIVgU7CKB4wLm8GSBlADW6tqNT3uJyfBHV17E
XuB2cW7IsFi8y7v2+hOkLFuPGXzjGLLFOhfj4x8Pm8VvxA9sFKav9QukU5v+IhQkBOqKZnO/xhJh
EoY010x8rboE2TG3QeANscLTBG3gxNqAfIr2pICBDopXS4Y9BeYNV5YppyD0VzzUDk3pNCIKNISQ
ndCoAkQIP6lsMkniEFRGzLGdvIaGr+xELD6bfFYXfvRYoUXn/j0Dt3LkcSp/ZjhWPYjWZp7DHxcm
qMxQ90L0h0kiLk00KV/FOI4RnUuYZWs7HHYlgpGah6dqsBWPpO8b2ogyA+JWqSDcmILQg7bkmeB2
//KLhWPMgjjXSLH60FdByVj7iYX7E6wwavnXDVisjcN8KuY65qFbMS3YruKNParbnxeZ4xeC11lG
wDGCsAMzzEcaP9svxH5rzsfQkJYD1vV4iLTole4mMaaS51dauRqbEYiOvHFiRWH2Iu+3TNCS2phY
KHoKrrcnkPHo0IWI+NwbEwull+uVC6eqApGhU4vltkWkr5kFmA8Adt8JDCt8zGNGNyB6j2fJQL5c
RWQDXCL/pyDuAVJVlFvbIj4nhE/HNZAxLkz9lBcts5jn5vgORd+xOQ/hcTaU+O64FXoKgckKGyQt
HI21TmJehxYxu/mCJrpHewk1T1hVahQ8cBsZkjDgB61E//eAVNjOkZrA8ALZPxLUEcuPfHbqxCgs
6fr9IRNva76RIWTSgEmyTj2w5Jm+PqSvZHwWXRFwjzxbRhrkDA2uCTcIZuazuEzEOtvyyGgaErMM
Dj0IO0nHtrbNBH2GWu4ltwm+1hAy2jX+KhtT66t214jnFOHowITLw74ectsx8fJq34CqBxD85vvB
6Yuv+S0+0dmGGt7SdUoxnt+nLEDkACqp9RJpdAZEegET0KpxJPftc9nBUg5xjDIjxGkQOcKBQh3b
vHMIWQ3aeCFSW9Q+zAuSAkdKa5TUfoMEysAl6U78F3j7MOA9f+7hryWh4ksWnncPDUUctNsvx2rC
ubF58Qu08RFJlEmOAngmIs/ix9f1IdVgrHCuxutjkgbHKORtWZmZ5shY81GY8Acw6WIUpLAzVxwM
WIzc4iNZrvUm5di2GWZHDZ5DyqCq6bAVvy1ta4a9ZVJ6NuEDIRk6Lg9cvB805cBaaVBL6nG5mLeA
BjyEEoYOJ5bwv/D0M02e07r1tBIimS2jQbni3N0sM6xVbl/dKmyQJTvdLNdNkIj9EZgHOjJsZJOv
rQcsN4Si5GvKxZcxS4/4DpW167g0KgZlZXwbdKb0bwjHEYqJw7JCQoodK4bMFu1A2nvgX+JCOgkV
OEYEC5q3wXHbNkLArEEecR+hB9tgqr2eXdW0/7E4EklHJq+POXWUjGGO9P/416vHOUWjOhsNipqY
XzOeHYo9IrpkFIWBuagoDoe9axDy5ccCIflfJlWY3NLwH3tz7WfxpVX0gEX0msWDwPNu+lI2CWa/
oNo4lH5aEf+lORUDdcx1PsjsGRCKbr94EVkMHaGCb1mWo5lAtBlaV3KlTXkhtL8C/usJ0pCWeFOM
PIyaYScq36Wabiu9lmaRzMWv6qaCcl0XyRfY5CVxRwAuF3HCVXyXPkhGxIhWN3bg33AzTWR7fm0d
Llorets98ShB/1Zv1spwguMgNYhesfxNk0pn0ISQtz8hF6ugRw8ysIDrSXsNBMTNA2biOdG0yPUW
4aWH8WVMTyKnCtMkBaUVfPuE1zN3Nkn52Lhqvuzhe8GQSIpvZCHv1xg1srA9UzZBEcJKQ4MbWK4k
VbCFUK8tus8oCnoLI2fZU3Ts54MH5WMkmpNfb6+A7yUWQRVRTygUqH/8QkMbovFrx3suK3waX0FD
WX56/wNsMJ3UUPDwXQKbe5a/fuKpuSlDCXNAqe1N91DE/d8eFJwvIIEv5A9TzAHZFuwQF0ssE33V
NVq90Z1QWznYfQhnkGVDCYKzFYshCcpE037nd32v9y6oLI4IR+HNAkpEWfYKvk/HrpCIFvw+ygLO
U/Xg/eY3LBkwoTaCrpxHzmDIaWMdLYvlyc2646SlrVROzzQJ77WP8OMkNUSEcPSybnFJe/4KKAqw
INiieGPaH5k87gJpJi0fr1MmL1SzAeZlsCEYvUfpIkEUfU7Y55xfu040jC+weaVinyY5PUWVUIOS
kxUG2D0BivDKz76rQQzrh2D9AcqNFlurMVGnF4qZ1aPocTCGfiZMffDGSU0ciWHD9NFbqeB0RwhL
JO3KXuhtnR/kRcCpXGGRMgTMN/i4f3hjAPn9qXJF234eZTpC5xdrYC2Nz9sQhXIZB+0pRwWe/KdI
yh6KbtD4pSZecasNoBMwpX1xiXEJDxDnqm1KP+P2bYJplo8R0F48yUh6XPzLBQVkZPve2F324XHn
cUUaE+qMT1baRAsK2lRVyvsWGkNvC+FdjxWLaacYIE3Z8ipu/GRt3RMJth86p3ejJZvgPwfvMfWF
U3Vrr5sil0eUnxygqcXk4GWXv7Jp1eR7nqoUJakzArDtYWm51ejjYx09rauTJhny8v+S32SioQ2a
eI820nVfHg8ajt+XFcJNk+yyt6yU5ymVq4DF2Cc76W6WKE4QqcCfSvTHRcU3H3sJ2aERIywmb1UF
mSdoDJHi4jjqFFI/585LcxwN/7NpA6kw991mGgE4barIaZ7AQKO1zDidrCQM7r+6EHamUOhFpZlJ
JieYtoDNxscguBu7xLSGd+5cGLzKRDhR5OOLlqm++JBwDM4cfUuWo9R0P4mtHpbFEpjX12Pm0yJs
/dioRu6fVfXz7wzPhvq4eJB/lNr/qe5cJIZ86QnLGuOs9zfNjdiMZmtpFyjYSnp7z/ODKWsTmFwI
40MyrEQ5BTEgfVVMf1Mx9qKWGDerAxSd8rSHNTiQ4E7aarEa+jIWwnGNe7aJevPre/p7H5aJt9bc
5tLUczFLdML3FPfhIez8dlqYWIIhwOuR87NYS9fJLTUroNsQTObnLy8goB73V1naNOYLI6sFqhXC
ROq71XqcKM8WJaaWM3Voj1zRiL6ahA8lScbZvTCaQ01FWNrzBAzCz9bQOnfFn1R39q/XxJ7HGe3u
tXUwvQMU24K/VAjXUDN/EWYVUkmfYJfZIjHBIPcgd42GT0U5ub1FkFoPTt5UHccxES6W5+wOTBZ1
MjP7k1BRGTcKea2ZAo4PhMxb8p/s93j2BNdx03OuEDy97WPh2a75H1TaJCTLwGhGdSYIxoX8+NTD
2LR+9jLNtYS2NfESg+MJJ6mHI98FuTugRwFxY3oy5QiXcs0MnbOkgd0Ni8oxFLxKpD72yCn/lu7h
xcYGHACGvClEIYIIN4f6sVCnmHmdzS3KD0GSAkTymOGI6oCoTEKVTsV5sAHlYoCNYtbaQrv4Qdh8
bYmKBF5srByB38dLsdaIeVUFoXZ3cEnO6KUa+d/MHMYeRLLmySlZ8kxLpgtz0W/75egWXEM2pXo3
LJg2efDciLab+0kYxA20/XFUiSPcjUJU5uPhzDpwvrmYCbKtNg8cvNTGTDvkGWQy2U8UZcikN5aI
GM5y/es0uundxEKborn+miuKKLJzf8LkTB4YHN0McdfN0t/8hLJGr6uO3V2ZdH1JmTojHT6XkcsQ
4wrxXrzD5VmNeJB5tY7LH/1uRIyPxUCgBejzXmFMwSFB7YdxqaQaFZGpmNmQfN90vQliaQt9Fz4T
RNgmwpGCIyjRbpO1vt6TBppO9feo4Vzia2rsYLpAqF5ZLNBeVuao1xB7U/m7feMPoieGq8LxhSoi
0jfpI3C9dXFnaXgxwQStT5MDr2pS30tkjdqFSOlP02xPQQ7Prl1xULFb7EI4wDfX1ZY8L2V5pLGy
nStgWg6WWofDpcJFxWBv0g4anY8I+Dsee0izjfqGFIkCcfAf+li0Eh8hNTmoHQhXl2nZSx83Hp8G
VfTD7ElEvEGqgQ24gaovcaJTvD3jZ3JJzWvEWI0S5BvrqmstU0E07KHzd16nCjK0JDA4o/LkRTOX
Ax4YCD3eZVTaCbTCpRlujhGloCtm+yV6WC+MZleDrSbQK0BbnxXe0IgSwxICiK3mLo2FOFnbFF5T
SGkHOrJ9PNkRz4hVlg8patOCraQ0Sj0lEAkJN387gxWvfqFk4yFT6cimX8vi/Y0n+ztwU4Zn0fCh
VxKJHAbxsysvEBTO181IlGA1JH7awa8fZDfDkPheHBwRNhkdHn0zIMIkScv1upYPaE+N+a/ZWXsm
a0daSOfdxbbZO/kop+SEOeRUDNmgo8OPTLgBxZ6ZxpYXHoCze0ZtLcenlXQVTtILa40GE+WTmR8r
qi1bzOsfjeTQTZ3iOZqSaelZFSR3Q/BVS6YkKgx7Tv1gMQOXCau+IxigdIzjO16QQYFgiYRSL6Jd
6FxrvO0LnqKZ7Lp75Y07Tq1TRmMEag1tw4CZwO5Bwc+PZES6Ne0ZvdJUW29XC9CwtcFOY9lNKNU3
8slfY5e4oGsGi9Gb5Kaqq8QbNK19dT8gaS4eixZ1fe/lEhoSgHIxEQbH9eRcz7Q8l7iCDLqOmgRb
O0rO+emjKMbTH1TSfQhrb6PRj/rKO/WNzDNtBP/6CueR4Ua5lvhKVGSHiHJvRVx1mGBO3KzwcASl
JHf7v5d3545qEHx1HVeDKlxREv3zB5QEThPLx3AQnHKOd5wqBu1ZtlizXqRUMthAsLBbxNG9Co7A
I46KS1/BYq3StS1mEji20nNjQsro61fPzUzwHKVCF7bs2mSYK0Ql1W5s3TguwPnztKqS/HOo5jPT
Iz8t0NDvDfGFO7gQOClE5Qz9N7lphjFuizUQbCXVrJIp+A5LKpQqoYseRi2++qdFeos6HcChchGq
muYQ0PJ2P0BLyHiO081dJhUoD0ClT0WIPy4ZdJGDQrqJfEI1aVxzSlDkD1EiIHaMgorVMCYZhG/b
QLWz+/F4l4EVDNGDy9xIQ3/+vXk+ymC6t2yH6roQ4pVi5zC9xZu1Lh4JdzIsA7CfGSwzDjjSmZ19
ffYpCHlJZ/+HEosJRZ8SXp6XzymYW3niHT69R7eGkwSqH+cLzYnIYmff8rSAbkV6Xhf3ViU2wOGO
ugcwWSiH9C662KkM8rljFEWTDQqIA2cbB+GjAIc2FNVDKaxsLOeVThZxuhzNwiRVpNmqn6TKQxWR
NhQq7Dgw3WS3JxdeQFyOg51agUzbsKP4JPz0yN47mhtsbhrn2otmWrhHs6jXMc9putCipBXuSJiz
ZpRob7onXc3oJ3tcLgx7HIonxIUIJBuylf3hns+9Iyge0+vzksWk2Qvz5GFGRvBKDq6LtDLi+A7C
ULXWxngiE+uwpP0cdjhTj0fkR5y0ya9ErRp7zmwPoUk6jmgdbjPaJJorN7naFcFE89VALa6/nX3y
JTHhE2v5Lfp1YqARVhUNbQv+Qwm6wj1sqJedsJisQGA0PTTJkgtsONNJGwlxznMSrE3Ku+GMexFM
PY9MT9w6P5r/Mr4AFl4vyUzysF0LPVzgsbY1AhxcVB7zvltTDJk9pz1UrJgJDe8I4qkgLpC+IOJM
bF+wzjF3cLq5S4UR+BXfcGtQfBc3iNFUMXy0DSCVD8b7hWsOvQnSufJTmsSjFKSv5N6I043GLCgb
BzEnqCTKMi7/VFs+nIjMxNyAfPPx4hAMvJBBic+GfI9LJXo2bVH0EYi10+eIyBcV6mHPAGUaSapN
DHbcPSLOdUsEKSbQ1/mde0PtfQ2SH/F0UQiHlN06NUoPy8+7Dod22wM3P9uJCkJqQX2S1WFxr76M
JjFIsTNHFgqQ7Ymqkk0OBFLfPOl9FfWKdSR9+weVNVOQiVZP0A9HP9WgXskRQuOPjVy9QOfXICrp
H+tsC7RR6cZK81C7Kpm6DtI3SzBkFoCXHA8CnuuyUWsRqGkra42LxSfzwDLSCFAi1vOxsdHecr7W
ulfW8CyoPs6fwrxd+tTy+0uDYMA1T7tMN3dGV5cQgsAmTqTQ0MoYhsHH42SqCOvZRd8e+bZd/FRH
Vjdq97jOy7tKp7diLNdFDxnD2b80LkeuV2H1CliDBGHMulmDIHjR0Qff6buixgA1X+YzBuo5MX82
mrpaxLbqD7Ual3EjSbcqB7571p5kMxAdXrli91WG+c/hHNIKMEzX4XwxKc46twKpRXiR9hK8qHEQ
2Lp6P7i/R4SOousLc+W3aE4jl+/c2t0jJnRNhfJ9fRyDPUBXh04QM/uU45S1sTe5RU9JT2V5UPQV
SSKW2qaoEkURGp3llpCpCvmeni9yrE0+OY6tg362XldNcN9gxUurtgKEwmyh1U2BNiMZZdQRhNWB
nThJ0sB5i4VffaZqopLxv0LHXOrGeMF3nN/tz6MOpbN93WB0xevUkqQWX/UStnBi2dfciPXisbyI
AbqfaeAC+u3IAH3ctM2Fq00U5mmuN1t+McGBVzR6S2jeW9ZOF8I7wsKx4DOdK9cPMC/UCnLKd1gg
6nwW6o0MTvTmCOdaMC86jsc2yWg1wz1lnmL9UnAnAjIMjj3LjAEsVfm/tvCgTHjh75wL3Bw3JtKP
LWk+yC9C6G9Jn+xEUC1AWKz10aFUL/sc6HuuNvigXMYHCx0TyBXhjWxPvCjRzYJhVoVIgEFPueAg
nt8+qnM2qJpGFfDyoYklezfVef43/Jz6lT2OFNSdP0Y5LhEU9/9LEE7pl6gdD78T12E26vvz+w0R
E/z0bUUR2k6p545R+8+R2qUL6ieXAhg3objYioQwkXzy1pjSmZg6sksuji322pG/1ajbax+fFyo3
UF5E5bn613VWnmR+E98TMK7wzkSbQiAUP/NT/rU62htW49UhnKK3fSeTW9kYxyMaulvfr4OrcFWT
fzxU0qKDwf4pByB4R4WJIZSfg2I21t1SEntpA4aXo/Nu4ItYeb4peOQM6dPeQ+RBYV6xi67zHOt2
3PrbP0Q/iu8zYzIJlm05F4lbK27sqI9a1bBSrev7DMb+LSnRtr2viNOYJTXhsGeExS34h1oRKWHR
tGmE/8TofMpBhFC1T839leKjq8P5X46A5NFKrYNzqaMAM80z02lnD+qq/dC7mfLEdl3odlls03LE
DjZKiiL5vZRpb2/phVdgbHh1jlkogJquDkbXq5moRzwQi/isXuF8tIMU0ibbCbluXF2RxDAJ2UGA
gnOXd8D+LFdCLb4BdgdMlQSS090TPZX2F7p+ga3B0M6C7Y9Hh2c0xGemTDE2pXEzEZwlcEjv/qVR
nJgMWdJUA4CY9jHha18ex5Jg2LUYjLdvFi9AIBDdYU0EjxBvu+vQG3/SjP+0JNwjda1U65slk6Yl
yvXTyG5P843QAK9G6B1a9fkAA5M2rTmR5i3cfnhJIJlLZdrbiIwjCzFrSW4mnwrRk+JU2q/6HNUB
AXaJBhihqPd8F443G5HJ4UPSqizWAtNlfiHunx8lVZyiuMDfX1OC4pMGkfhBwOnWI8GRskNfVFz1
qO04xALQK4EXk+mY0jeOJCb5q39kArbI0EklVXWa5bosgcKd+aMLwjsqbcYSyRxNtIxyHv5t2BQi
Fpd9RsXOStmBPGkEdKcIxFErwfeO986xYDZ6AkP682wxH4U6HoPfiCLIJcF3h4h5iMVHh+EwJwAj
TNKPUIxL6cgxT34/PY3qnHVZPR5CKTgkjWMJmT7cQQvMQ1+x3y6T9ngBqSBgWsaOwopZQ97eEQxy
qlnzuWg77ADcQuHRHFNGvMrFXuy2xWpOd+NsRo4kq5I4+fS1kDnh1BODnC1D6YCwAT2nfSaMev5H
AyQjBcXMveg5Ys4VT6KoCZlsNAIxsI+pR0rUkEdYWaqKJLGnJ/ucvjkLSbnAVBB94N8vV3zSQFpd
LO8WcSktDao20y8BfolYtCJkOhdLpVEAW8q8fmiai21nm95I5vAbAuRNDlmFX/7Pw+8QAVDrmU2C
WyryoDFzg/Ie2zXFOWAZI2fQ0HSTEalO6D44Su4Zut/nrMRjuj/6OmJ7s7LYrDTBR9mnwHPoZrEP
5hb+VOpUFG3kjtvTmw0dtq7rHCgMaH/f4S5TDhNn3+WAsXic8n7BYWxyvjCSDZ+YNgDzWKgwyRCa
Z8tcaOfk67/nbeJT50GhkhEldiBYoB6tBBeMN6R0MCXJFfOjPAvi+xkPrzWB+AQXqibATpgcPT+S
05NcpR0iK40lb/+fxuNhvPBVgLxHav87tkriCMoGm95Bz9mRF3CvUjAf2EwmF1mKep6aKT3/beXk
SKiRoWCvv/K3h/UlTF1tmN+g5Ci4PC2GmYLwmqJhqwJ6U0RDgLm4mJrEWBj4vSg8lAFgBTPsuB6h
/0DeNHhaFKLlCvMtmlKhICzfNMhybwrMhQC6A9s0iIEUXZZmgIKFeh/wKRN8dPgxTAaKujCmnJsI
qICiRLvVvrI5ppHfM+bYjfUyYHTakQ1YRzF+glnNaqDnt5Z/wC4YDD/WgUa9B/raTSUdQzNvcuPT
xnJcq3LowIcrK2XcoJ4SVgTCVwpuizh4BYB7Ue/A8u28ywRwB9Rghy2cdVJJg9D8YKtJ9zchE0+r
Xi+s4cICh9jLHQejukzpLTeqQQeruQavUhUJmbVW3B3uX6QGckGB/ibOcCMMqri04mcwWe21ta7N
megGotCnsTXDd4uBg+LJ1ko04o5tXZEN//pdnlGkuSjJRyK67jahDFBpJ5bUZUgavnVHzXzTxuwc
EGYZyXi6M/XssSpkORHRR5cpBRn855yqi9pFIUAQtDlCUAUubXG3Kd9SFit6eLwuAQTSIXsR5ZbN
de1jnB7NlHp5khAMJZCR+CwQAw8ZPCAk5hEJyMM1jMMTcya6O4rOTJ05hJr8O4fi6t3bD6qMT1je
gd2FGySTRrj+mP9goJQBG+IPWlfVoQ0bsNf1Vo2I7KamLOhGgrJYimi75+WiD0YH9ZBtxjTVIwXe
mYWcGrc3/CXTCmVwRylDYXW8msLPY9Wi4T+e8IQEBgjZTq4S08znUJZb0+TtHMJdq/eUBhw3WfnN
XS459iydPqEfl2lh0067wG3eJZIO+88kIR8pW+4J2EMQc2sWBZC2zxQH+l43M+5Mv6zHG4xe4Eij
lCxC66Z4i/LkmGyJCmfGkwixtH1YQ7k0optzweC0E0Ts37O83gJnkuW2Le2/soupjy8zRhhFF/AB
69RrSfgNsCUQBgrNnCbJumTSAComAvxcLrdzVcvzu9nBl5EySmnMoeVeli72J19GQaKynHZrTs/d
zEgR53NFWCx/eZVtHYeSyPBHVPBIGeaKRQ2bktNB7hc+43GdZN9nUlJnl/uY16RZVPLiLTzjlPNZ
LnMwhYY+0nRqGjzH4pQtINRyTf81inKFFodFRUVXPLmW6pglrQaPNmCnn6j4EBtkPHAe39kQo6Tn
Ld2pczUwmIvw2sBScJgDiCgVo2hXcqV8D4Kr1WFDhaq8ixajLZ2sKzI6q+Ue/pivBFmehOPv4BtB
4DwC02SoinWV0s4QKhbU1sW9DwjF18B/4XliCUczo4S5duCPVM6/afVDu2Cjl4MTOrN9BYspJUx7
RTcFJqOTRrtdU+TwNMkOyqo0v5ydJ8GnjF/QMY85ibtKUzZHbH+eh/OguyEazFQvw+JsfO1275wv
OlvWRlDiUx4aKoBJ0xVxiXMEEnjmCgsEHHvd9M5yqKjRYznIrvVCv0+oxqU6uulHkkn5T9l5s6At
7c/rl2AU891IH56Kd4TE44/UOZG6I/YYDDz5b8cGkR/bmIYTxd5GIc82cwmmdMpzU6XsJFs18DKC
OxSo3yy/YBQiowhaLdnGGG58AOuq9Ap3cTIEoUHXRJKzC1POWJFjJH3y1McriXVx/f0CfHZEB3Fg
60l6ynVjKJHl6tOBjHLV3zrleQ36Yp5n/M/3k7u+1xW89Kp/VFyA4B075hj+MxE6zl8ulkcfhum1
FNdzHgBCfiITZl4+aFlaEJvgGR6t5I02tf83xTj+4Sfswkyzhc7g0R/mCtohXSAcVPtvol/xbFhu
rAzmTFWu/RkR1rbeLp94xincQ2rs/eIEvN0vb8S78Ley9+3EaAsLLPK9V+2AcdPZZvYMjSmt73ER
1T42FEFwKKPZgfIwmr4z1fPBnToFC7M4zhySx+yWrDjWcTiSeVyfr4l3DnH9dXrLYK4t98I2oQRg
5tzi/c7xD/8z38gbnqDoxdiPZMNi/tLaiEdZdmJ5YdLNQZK+KYaJQEp5JpwgE0vhDZLREDXFJJeS
Wdmy5whEA3HedspSY35zTlikuQWBh8CTW6faj/l9Yk88+UyByWNQQu/ZqF76yRCgrWKqt/mglH5y
rC4YXIasYx3r8wx2ZKRW2Goesngo/V+0hObHui8yZ6KFaRLsavb9qsd++3hNq9vrYLvuu5/tKVx0
U2HrNdBiCDkaNMSL9tscg6oD1T7YaCpwl9aKJElI98FsJSMSEuBpWjSFhEVAXb+LQuNWXYip3r6u
VFVChtZwnKVilZek2t8dwtMSvHOlt9hgeMdXFpo1D+VT8z75dJBc3ycy3B1FflawFasRI4wyzS//
aKhSpYoiaGxEHZijeJgrf1+IfAL0iyMXHXCB+tOyKCAv8qu5ytOpfLCTwza5ZWOZkrnnDgXY3aIT
snt8jzjWCU4wQamvSauhftGAQ9codJFoXVXO5w2T5WGqf9XeQTexbmy3rbef5A5gazMUFQvz4GOV
dW/Ce1TByaJb9iH+YhTuKATKqutghkPPqJYalJETBodfyJd3VIkJn8Qc6a/FAFVl1upYHQ0iY9Gt
n4jHuTD7jwH9HP2quyrSvSYzTbJGS9wx8cbbvCzxSIiAwlygAe4IVui84ERF/0Y8BYOKxWMD7bZb
J9KVmUehbilmdr7SqFp1atOggObbz5q7N6W4/w/5E2PDsJ6fCrOMF2dhKua5xwIUJ3WM+mBihx7n
jMdvaJYrT56KK+l/JOGmG9XQbbfd0Zr4H1ycQ9pB9KHvM03NutNsmFui0wWTzzuMWBM0zrVWPIKm
8MASWOsUmmYaNuzz4wOVGgtbEq9fnLytxj0KdLGIp57D2NnoivvbCsNCkat/Uft6+XY2wTbXdvn/
4yKw2olDqJI3/Sc5HBsgVLLh/J/Lu161KhjpTKlVooOJsJNZPtBZybUDSI14fBkhC4+LrQPn/uK9
ZHXmfrO4NQbRlaZYqFBn9W8gU7yIXvX37dDpIBdfvtx3kp84mQzS4Y34N0Rh5GZk87Pbsvp6lxh+
UAaLxTatmUiUR75t3h5oplSmiIPRU4PqXGiJxI9eANbC9zuLLg3cQQ7+ZE6s+rP90dUVihGTS6HF
xZmPOwOnWPyrZfOMSqgIU/wV5GxkpV0nIU4wdUlN9+gSxn9z0WKzWpfi6eFVBUF38KvDKbN/d32d
8AbtiRQeyKcOltlFotk2F6St63/ADNYzchInBGBkWXdkmj6qRQx4aGUlgt2pN9QMwKfpITdRFuJ0
YBsiaY7T24p4+tqPDYQ0F2HY/boDMuQAAlIuf7z5HW3AXBufdVbnTqjMosXVxrwIFbnKX+g/9cXw
cQR5wvAMIkLmMWCS80GkHKURN8YqiRlesUoQJqO8tv5hrUec5esQimLFd4fLxMINPLM0X4BtCc4j
YM+qngFUc9dp/dVhnh40fbhGF10o6/lG4wNGW5efb7gRnBpy4/0riFNnHckSVxjnK/dBdRyaPGTj
RTkn7uMbOX26Tkykb8gqVDAwNvr6Sro/Wau61FnEwudeoaC8DmT7sLYZn5hC85gYKzVKOQPLKhjB
feAEpi2f1YkPQ87CEhoMt0/Y3vSqf7HJDGFjaBMaQbsFtld+mFN/qAxeNrFNxOcfm4QRf08jEdU6
OUth4CiywhdX7dAPhNHsoMXBfitid+HaXLnxKnWntRzGOWxkV8LD4ZVlycFl4On3g9BiBDrfaFsP
l/EYrc4ex2gY2Rg7xRMqeLvj7bj8Ihpysdgx54lDabQHeF1eccwhnTO5bwR+EN1IodSFrWkBpgqX
htr1S2dRT63h0LOADwIe9j8aeqKJr24ksAJj9sBbdDyMDPCDVFNVzQAPfR6ZAwM2BLfp7GC6J8vC
CespuUZEaajLzbI8LcEGnD5/zE5RKFC1fKHgtf0pU3gkLojsrJrtzULqMoPl4xw78b9eMnjwi6nr
puCmjByV6jFt3dkUGYKklABsclyo1YAl77IX9k9CbtEe2HjxMVkNFbMs343hjVZbSUxBM7RU/B+8
UQLs7Q/4opMawzKSWKNJQCjaEWL6x27Fw72KC+GVh7og/8u8eEyjYxIU9l+XgtblUgEUDaZ9oG7r
2mOXB7eQJYQNJSKlNO2EI5yZ9WWEHTQPjGTCf5msGWkYsVyGSDkg3EK9fAQ1oqyuy6iJBcPjJQ26
3ONv65+0u1OS1cxh7Cn8ZihkmUGCRX8RPeIeZyyC2Nsp1W0Cscw7nAfjwqMzAeQUDsQjZVyoEBPK
W4VWCcxjYsp2mKXWfaJxbrF7PSfWBafZfq+8Sfdt5hSY39uH3gkc3Q1xPwx4413vI8JVaPOotgbN
KE3EZLjWS2aWEYRePxm2u2Mcd7h9CsauBG674aMN8Y6ydZoKoFGG6nWAVMGr0NRFeSxhck8PezxI
LUapeHfbloyAHpPfaqK9JIt8J6bhzKlv5rRhZS2zjb48gC8a1TsyIrHGz4OW8wGEWBUEWxcQJgoB
Epeq+bxQU2Chq4Pyb4tOwjMuIDccUQlWmtBFugbeyypS9IFlfdKlCL+8cCjq+/vSYmxDYwS08RkD
kH0eBjOpbizDigqNZY9jmwFnbJQIt8kUWgYuYjmjDbg9r6FEzBLK2BGDMDInwPLrXCloBz3wh8xg
M06rFZ8SB8HxAM3rVb8TH879o/C7WnSu2g6HISZJJfLwZvw6rTPipof0SoHECNMwTM5QxGwfxoY+
AOlcHi2bbXG1jIQ6UPfIdAns1H9l7+PL6ZoRdcl+oHRei4UvEicJnYVzOCxDH1e6AEtibh/1TC5f
HR0trWsTiOR8yBiDbXJfMyckTyGKSba7sBamEV6nR3KTdKESimwBQr/gAeoeXQRF+CQPsByvbH87
AE9VL44ZS4znb6cF/yg32rQ0qLFnWq8xzgnS/tFpT1cGW/LPX55mq8oTC8VwaFErcm884cv9IIpG
/6yk4zWp/dv9wZvVmJnylrDJ3eYs5fA9FQdE/LU4Rb8cq8NPcWpc/0BxKcCPDhjeoxwi6teyiErY
dMHpnWzW00Bm1eVzZWOwxGBOVcp2kHD+DKZ5yo2p11iCIuv4vNb2o05GoqNwWUD2TU0UOLoSYEK9
x140a/FMY9EfNQE6U26RNoKa/gOLfAPQYlUJd2ir47xTCbinstlPLvVnhX/IcDMyi/jyJvB4x3Ec
mGIa4N94SqUQqSIFhMeNtCbBvdNYEEn1YNQzxHHeah3luWO2ziKH/ysqQ5FOIBT9o2vQ1I4KBiUA
9klAan1ooUHjPE4s7fPPmuyJrYidNp9LZm8DKFSNXXg5yN9eJFKL/r8uk/6gy+eNpiDQRg7SoKXu
HC/CC68f7+/PtSCROTImBSGaXEh3rnC4atyWTu0V1ah8m9RdNzHLmFi+1zlrxDKDYlarYd6VbEnA
2tz2Oyjyq9ossQSQHtzogAJ9+VRUkNA/0ZmM/xJrjJwpjTq2tbHxLr6aElC8rJkxYAs6yVSxaEuq
8RnyRJ8GswmW8GzJuZUYgtsgnIETXKObkFYxHqhlMijyOAD5FSAY2tvMe5UAZCfoTW2WrDq7xgo2
y3QBsNY7W0JoQC4s/lE/W5+SEqzpzxc7Az2evoMmBYakZXd27PIUZyuEqHDy0e2WA9w9vXM0cPvC
9tBBr4Q2ZSgMjMUbyh8XXUGb7wjLadlWYgwmpAqGRcKtCdbpaF48m3PzAGWRJHMK0nMtwLRzoMrk
XgRwvlcKzKrtmvCLOo8DkgaCi52k4GYRnm2O70x5dxOwF7GcvOerbXmnQXk4y9qqquri1ofsznI4
4gbUgL8P5tgh70nJ8vSM2spAliVAJrTz8tK6FR+N0pdA3kXfqXxvLRAe1vcE6Esyn/B3Lq89F0iD
vl9ifn4DF1VIVgB1qKmWMSdsYw6SUoB78c5zTc7MF55hFIi164u7C9P8JeZkhXfqa1yYWs1fX+Zs
YNUYAyYyCYFjBZLNPYqL7JcNoLokvVLgwzUnktHHZJleHvBdkfqhqD4VAKZ3iU/lP0Bl0vWPxbRV
xt/vcDlnC4R597H8ro7/mZLsfN/AM4HNSRDW14x5SnRRznkVOXmW7C/Oxg/ILUQgZ9yRLihdv9Mf
P7ReNIzQK55LfIEp6+Ff8UiKmmGzlQzO9612W4i+e9ZjY9F20B7hWARXmuPCXiUcVegZVlZb3alZ
d+5iSFRffkaHnH2WucA9W5juKF8Xk2ET/c9Y227MDd8RRMZFC9fdsfyzW65b3Vv2sRbaxUkqItC+
Yd8/rqpJKkTWRdRKzXGQdleFoJvCK+mnDSR0bdcPWde50vYj12dLN0toKTBQw24tc4kWZvOcTGiw
Rt1814BrtIblenmV7wnC/V3FJBcXrS2GRLFrJvu4sfu/ZhsI+fzZ8eAwGgTUjJoGw1gBapOX1TKy
57NalCmFXBetyTwEhwWHPlgdcWVPTQNSHMtI5KpgqnyZkjHDy6z/N24uPqCgJpCB+z4TTE4vXvIl
6Gg9MdQ99uaBuz5FHhT7feM+DJHnztCtXfa0N5buxE5H0rGoJ15L6EcKrr8zglKp0vRCkFbCkAmD
1T9ii9sokrvVCgNRq7mriOkQqxIoki813FjTMMm31BGe7A8Qog8oDh9zHenCiEQmtQ1Z86420DPj
kKAMa9HEml2BqtFPqXVIL63JodaqDfpm2zjhSJDXwTbRGP1L1Lris2IY+pXIkWkU0f09txF2rG/Y
ypojvF+9fnJFYlFvTDG2W+sONY/WcG2L5PFc1KH22ovVyU8uEG7u4nKMPKAn4m+pkaFt+vFiv7EL
rSk5UovPYCwwpIZpukeJRT2NjMViCnGjhqDvpIyugGJ0DdoLD5Pd1SYP2odms+lzAv3szduqMCEE
srf0DFpFeDqnPQkJUGccxt/15xQ9/J7BOedCF/L2gKh42H+S/4P6sDH42V5Gb+dzI8Ym5hz+ONZ+
rsbmQSHVB2PlUmpJcWkx2X7hTOWi0ohxfBVA8xR5XKezQQRmUlrrbpPhPkQj405OyYR0l3voxs/G
kssn6qfS+JY7KW+hZdaxYO4byjt3M/m3oLVc20Hx+NebLDhVVOgPdY7p8PBwlqwaPIgXCSvzkCEv
lU1u8x573ugWqBqvewj1j3ryh5L+AgCbzsD1p0lxj/8x1uo7SfD983ZWNK8Bwy8rfYebEDC5M6XB
+iW/l5RCiaQlduvMZqybc7o8scXXaUIvsmNSKsXCv0SI8JyfVHPUDf/KCXgM4jzH8rWvAiOdk8UB
OF4VZ/ExNkjLmj/DGSDwx8fiSdLWcmAFNGU0hReKx3rRWEiDCEJrnTpslQ4AwACrH0MXfh1X7zal
QILtTWwizmKAmE8F7L6vKTk6GdkGIBwh+8qAfbvDoWyd/Cd2EpO39cGVuFmGtwTOvsVh1TKl0yW6
MdqLAzfVJZmeerus0nXpEls1TYanc6DaYx0mI2QGN+F1j9i8Y/1dQENUVkRRUHCR6e5x7oNPjd1r
juoX3d4IZqqtVhKOurBeMj18fGoDLjFLDxKMFp5+CEJMQEyNUm4GiSlyNgxx5j5NkBXBBdJMMtIs
QHTrP6pYS1meGCkutB95cPST5Ia/Lo1DRw6LotTL0iEzLpo+FPHNmcwdzGOgIbkPRc/t9DLha88W
lTj3ZnFcV/S/DYiyl2A5s+zml2aLnJbA8kvPLyjdNErbVc9PQk0a2cfbLExoGuhlcjM52fRB5bp9
M0ZjF/18H34loMhUMN133d4Xx0mxi73tvBY7u8YXH+3fvjg0AZVSIhvZ/NEk+Hu7G9DnHSRNk5it
4c9LGAUV6KcgRcVsHAyWtre5Pu1h9g3rc9fJPcPIBslvkDyJ+/Q6xn/6+9VlHYKeVTk+XRIiWfp9
zDvZY7Qle0CHMLOVBaPDoTL5qPHkrHiDcureTL1RSAaD6KVUTpbKUNi+m6EtwmjcEj0ezsKxuKEv
0OADtrj9akVpGswEkUydYDmADXDSJG6g4OcTZplIl/yahFSGOzpN7Gn0ZMnowPdqzqiT/t4WbWOv
HsOfNLV4/dUsJ0UgkanGWBPWVwh6Ugnu4cdIB0c8PJRD1OchAoGfRXIfZAj2z7dwcEAHvpq1Wwfz
iVcKkpYG553n8h1rmDfCXa5MF88/TJwPEExPHLQQrNh/GEyG2Tqq2UCMhP2riKhibAu9taSsKTH+
bU4vB6iwsNFGqMlIP/mTgqtiarMQEl67RMibO9OMVwo/bbfZOoINSU5gHMjWRyeFvtJhWApsanOU
gwvLI+llb4zzypb2niOCT1oYkOkAGNcOgvH4OTTlGWikAxmkibC2Rs56VtgewhHUDLtv2wFwZ7kb
tkWKgW4mR8qKAC+JRK32x9QtPr3HKvvAr7omQ3KQctoWWqAfq4z5t0XLjSZ0a9ewD7wkGtz0YO9n
L2l74zOtycdTEBBI+1PBh4JmUByfVbKqLDCNnOxzOe0lyJTWsaDiN7A2yObpIdE9+WX4aVX1VUeQ
vpn28FSdI1IY0eZkK7KqKfYKVP6KsJSXVpC7T+h4webQbAj/3Vh+MH6hp1eDWWA4U0lb3VLUobuy
CHJ6fhkeg5N0dEwaQRmQDCtBDIWjg5Of30VTj+HpAUH+pSivKlfUuvVQiqC3l7JAdlkXhEt2Lmuy
F1ojjYfBmXwzoFvXtWwOBQrbJwWKLeumBnJ1BEpTK1RQIG637zGHn6FHOp13Hrj3NDt5agHYiHn4
vONgtlJ2jm5KLINy3SlGUhbghJaRl1M2fXhClwgdj2cotVQVewTT6jtEtmVTK1mI4uK+cfNEDLvk
wpYKhZ+MqavwxxrHnoqHVzUefPEHETZ8oUctKNZxexQkDmkeTKPJGR/KssQvj3ZoCvE+0FfS5it8
1a7sM28MWfoz0NZlNsj4TAMCLZSSPvxYzwHgd1V7FPadhlycbCug1iBXc2vyitMoQkIMKlt8kDGB
D1sEU8VRKWw5V9LzlGec/pas8Xadaw+zvzopV231edJKyWDs33/rI/dc4fY1firqxYnH74wMfUZw
5ZHVmvyDAHkFMNB+AvN6I3y54eiZBMLwSOD7WODWk7kPqN79Pok4QKgd3EOrtTMxh/5qupciurKj
xhfekdcMrq9vrL4p42iviOUDTuDWDSbKlHX7K3itXYLCmRDAV45OcZdhgD6zQ3vnPP/lsMeQdxLH
XAGWk93mbsT3LmcAyBynQ1aSwXE4UIRylDSO+8Wmm7Bl+ybaf5GDJXqkVB3fHaQHZ0j2w3+RFRVv
czsGr4Rk2sXA1RyMVuO3oPhfc7iYdzZQR+aJCRG46ggCCJGQGQz6mxjg21HGfiwDcBwbrvZiGcuU
vFUZm6ItzQEbgYAlIR0dvW4rqqaqEkwGo05q35AkKF/AU0IuPmjf8+bDLCF6mU3qJll+btjRbfxn
/SacYEjHXNWbHh3jBvq42UTmxfLm+eIUMRFtaPn65xhfya6IvH4i+hnuUKE0+L0ToAJfGz1kF4pi
cH2Lwe8YM9hUiq6sZaAy3XXD33rs8XzXPHp1dtAfC9VDyoCLF40oAA==
`pragma protect end_protected
