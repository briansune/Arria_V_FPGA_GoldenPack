��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)���vG4��NB*v�^%��_�rG�v�2�H!�W��m�e��
W�0I2̵�_�}���
����q8�Ι�t ".���c^|�F���uY�����UA�Ύ��C�F!�'��3����bj����ggcI��I�ؽ���S�c��x�K����O>{�N#�M�lq4��OV��b�}�� �d���C�����f��T�٪���7���Zi��.�Lua.I��7��B��ѧ:ɇ^��P4X˟[OF?�&�u(�7�
�$:��A����S5�dȽ��N��B�(��lZ�ȹBd�Ը��6<��ȗ�B���Lh���������1�mw��T�Z��i��r<�E��e\Q�0��VAPF!�����JM+~�����@�6z�t^��ڲ�_1p`�=3�ZY�X�{>[����� S&qb�����m�L��E׳�2���|-��BH��\�=/���5�Bpt8Ce,��]�ҋ��-���~��&nNj+A-������C|�4x����_�������a� ��j�)ء�H���V���X"��؀�
ebȂ��m෪C�67�ш�m�	UC�N��@d[G��1�J�H�-��m+��m�t�� A���9�ĵ�bk�9rip;���T*�wܼ\ �On拖�Pl�2�����3q V,�Y}�*Yq��L+�ܜZD�3©���Q�~]0�����TcS���9��=�a.���z��<���#���S�]qY�X��K��M�^��?�/+�Q� ���`�cm���^�ӏ���O4��6�����+����[�!P�E���S���t�ڰ��o�i�b\�l���s��b|�����DY.���t���l��S��O`:�O`��hm�*/��+����w	=Y�6�r4�v��כ�v��@���HW���+��:φ� 9��1\���	a�Ɉ߬��=Y���r���e��\�0��Dg*LŅs3�����.kT5[�
l4�(K@�B��Rʨ1f�RW���;�����w�=p�Lޣd�镭vp��2��!������M��*v��
���3��@�~���U��|P2v��{�����"��\����"$��FlP��[ɪ���ɚi0���5�$�ș�)ˋ���%x)F��r��q��ő������)kS��5����	m�[s��� ��8_P��10	j��C�R�GG4Y8ߋy����&�}ќig$LG>JE}\P���m���C��"�(K�=�"�-S�*�4?J��=��n��l��B�����,c��O�[)��G�:�O��:�g�l);�|�̕�E��1�z���ϲ?���J����~�6�=��\�Lՠ�]�$z��܄<����!oM��G�z�M̜M�&P};i�J�`3YF{xy��`���)
nY��n?��7���?n+�o��a�52��҂�++��"£?��"*���c[>Ɲ��<�)�!��Jڤ��տg��_E�世ttQWG�"�Y��i�m� j�ių˚�q�6]ŒOdh�%B]�1���*Tf��w|S�߲J��T�B蠘c5��C���yc;6��.i��%D�������A�m��6�H~���׏�Ra��뢏9�5��Z�� $�K�Rո ��־5o��vh�&�J1�w�v��93����>j�ng���5�V���Z��f�������gBv���fyM������ƽ��=`�����v��G��������@�E��M�Ծ�r�����4��I�w�˜C2����1�� �n�k�m\���8�T���i��Ϥф"t�R,l�KwsG��3#���D�C<��ƃu��bh
֗/��gR�&�Q�wo|t�ѣ�".`��;��ϯ��i[��Ka`~�O⻩� Ċ\X�g�$�}&sC�ž�+�^���q8�%j�+������lU�h���[nխo�\�W� W��C(�����tz�v�4���W��M�@����ɬ�ަ5���](���˴c.�"U�A �f&�T���0/+Få�5��6`�H���f"z�w#����c5>4aЅ(�'�4���$����d_s�W���u<�l���p�w��F�z��q����+�ɻ�/��ރ?�z<s]\]fo�*�-Vy��&k��q��X��YN����CF0D!%N4/� 	�d�ۚ#4����)n�NnF�U��s<6�r�3��%�N��&sQ�����jĄ��T�RF�.���.-�E4���7��Uc"� �\� �O00ʭܬ�+��1(��F��5w�v�I��i�A`t6�h�캓��c���K�^�j�oE%?}CB�����1R[Y:��Z�e�w&R�����$Wyi���g�\��a	)ͳ��4FL�)d#�U�L�Cu�|��s��x�$n�E'  �n�ؠ�v��S�V	=Zo
�r^��CP��bq�c����o��SA!�8�;����[*8ܟp��s5�E��Z� };@�hO<[V��#��A{��Z'$f������c�3�2rkk�Y@��g!�y��
��j�4G��ΔG3mhŜ�z���L�ژ�:)e���s����_1��erP�] 5�Ĝ����4=zC�w�X�܆%�2����	@ �����nğ�#eC��i��������<Gv}��줐H�����(��B^���S��`�c����m��Ș
7c�C�����r��S��w�'�u����-��8�'bX�ư��g�ϒ��.k�n�,�Vywa�{5�U���a #z��@ػ������m&��nz�)���]�r�W�h�ʱ�T3Q$:	���Q6�e��!�V^������(e}@?�:���m�?��U��I;EX��M�e��n}ǔ+	}+�)n_ؗvk�lF�M}6�4�Z4j���s����T~>��/LvMȃ��.�WjS���f���F���
�vb���b�&~�g_�q���|8ŶVK51��K�PrS�Cw}����gg�w�	h�c,�3�8!�{t��P��*7N�P@;Kd�u/uw�)�R]V|�	UQ�������F(n�k��Z|k;��)0��ǯ$L� ?����~�s�!�����\a���P]F��>��n���4#���أ�c��y�i�[Ȉ`
VA�4XGU�����a���#.5avw�����$�$����,�W���.?!�������c'��2ph�4aSD�+��ڝ��U���M�Yx*+A*���%�>�bT�����B�h���>��J�J��L�|��C�K��Џ�n�*I,p`W�EM���u�ܠ'��Hy����+��'u��s��7ߨ���yn�k����y#�����~]�ݛ2"G�2�L�F/�J裌���X�⋂�5W�.�x'>qF��a��{^��S��9� �n~�}�g|�Y�����v��[������i���,g ��7y[�,CW*H� �����2�Ӌ`E��^�X�j�h��Ss�"YCX(8O!���+�~�vYyF���rm���������u~�Z��:�d5?���^������-g�FQ���!'� �V�5��]~K��t���.�9�;�,�O�{p��!�*���[}�ff"ʽ�bVzfG���P���jyqbh������Q��?#�s��k�aAq��{�PΉ)N����.�$ǫ2�FAI�+�Y��ZI�s����<���P ��AӒ�Qc�6��,������}j���=��^���XQ_a��:+�O��^�u#R-��Biښ?UayWlD�C'U�\��i@Μ�l�|�\����r9L:�(A��ӄ"�Gݪz:;�,�.#� Yi��C�?����� �wDۓ�ě�0�_�lwj��d��[�Z>X�B�|#(c|�eg���^G~�	G�s
���t��B��L��f�;Ik�7�.�]$c[�7��޲ɂ�V��1��W&�!6w�@6o��-�kŢ�a��t��Ԧ�8�� o�,e�,-\ʇ7+8�/�5�|^L�g���5H�l�[�23UH�0����$�0�ӆc�Tg=6w�z�g��QiM2\nr;>%:�T�<$'�g��jιIT�9H�X��-����
-�7~�yzm��6����!��5����<E�8�-c�ڿ$��O�7����?��wA�������w� ����h���R	�* �����F���M0x"�;ڙ#=`�ZŐ��4��	:��|cDp�_�.�����+���uT�G�v; y�-�ɓ��n���O�v�V脾T�?���_|��oǒ��2��a����ζ^	I��Ju_����ɸ���l�yC�n�0$ΠDbk��+�
���۽���v�\n`�&6���=��G�_S�>�9����rJ�qe'>e�b�8#�{��_��+|�S<�s�2��;�>~E/4��$����A%줆�:�Oh�߆�/z��f�g�*Sh���b���r�27�t��Yę�ֳ��E%��x�߯�!*��W>Y1.��x��/���`.�L�Y;@���K2NAY���eZ|sAD��!ӤԒ�K����m� ����eq�'�:�6]>8:c��%e���.T� �q�a��ئ9�
�Y_2��ѵ�ð��*�ۻ�����N�ٕ����~o��^�����<�A&&U4��`��mdZF���H/�K�>&��BU/��TJS:nS��0؋�����nX���$n���{+�X�<��}搅 ����jf� \���&R�nT4���p>���fu� �)n4�J�iR��*��t����� "�->�E-=R���'7��F"�!��B�x�dv�@�]1k�G8,�7��P L�>������C˚�vx�x�_
e���An�39NgO�����,����P.�Q�q����i_�Xa;oM�b��� hg]�(���d����y��g��v�?�-�Œ+�nlT9+��������~���$:�<.�`��H�wJW���2Kv*��V�~�5]�27Z��,4�arǧ)b�4�����yP���ȔQ���4���9����_X͕�?%z�/����e}�t����5
>������s�ή|c����)�+���DߏX-�z����(H���Jw��HmY#69
��|+-ܕ9��-�`���:hKʆ������z�̀�P���Lުc�Vj�E��n��j{���P�j��g��+7Bs:�O���6p"�a�?�AИu��Z[�jQ�/{�h������1�r���q�I��! �e���>c�쾏�h��h.3 3`�a��da�vdI�Py��b�_��Gus�a��P�L�������	�X}��u�D�7H+ғ�H��ۙ�Io�p�� �c�;5{f!����.HTk�tj��5�/�L�|��m��_D�8�n���`��U�(�)�*�G�34<�Hҩ}��� ɝ�S����c���l �L���VG��kG�=�6�����	��*@���%��tG����(���nX2�>�S���`o�:�G�3��&e$��O�C@xs�۳(4��Cˤ�Vڷ���P�K�(d��c8����/�M��E��Ao-�c���x�𸻗�}�2M�_�zJm�zPfY�>u�jb)4����V�A���8Y��vq眪�fp�5ך�8(���BY0Kz<B�S3������Z��Kw�v�Z���%�;c�V{�����t�ܤ�D�eyȴv��U�Z��G�po���9:,���Rk��>ܘ��Acf7&��I���AۉCsh�۔�y�r/�p�=�PM��u_�F�]��!w�g�b	I?]������9K{a`�zNM*o�;;� ������o8x���6��	5X\Q�Bǡf����[�l��K#�Lh�K!^F��~� O�q�p��)��g0PK#Q*H��(XU8	�M�O�8D��Ö �{���`�� s�(�X�>���Iw��@ct~�%�of��Є;�L_�"�He&	F9zM���&������-��4�v[I���]�9�f!�G���[i=p���c�ɞ+ۏ�D�E^��Q6���|/0�/��b�:��B(��v��@0�,?�H�R��7 '��*1���bͻ}=�8�~��h��x�&#�4ҭ�Td�m��pS��]׊�-���qMvm�Fϓ�w #eNt��P���/"�m1�<R�!�u���΂�_�(�Pr]>Q��,�$�-��_+�	˓�>J!�c������՝����A4J�J$
1��/_�1Q��~s<�Ƣ�X���]J� �!���"6uƯ���J���Z�������ߡw�܅鞟O�Ϙ�b� t�y�$u����	4'���|��ЙgV�Ml�XY���>=������R�����*���&W�)�:�e����Q�׃�>U+����6���㯳��pd�]�
5�1>�}��sj1�8X|�
	Tbc��/e<�o�[�Z�ݼ �h���	�~X&�߈�*�\�n���f���@��V;^�n��?���U4�g�ž��@�	f�O���8��_�%qT��	�	Oe�=\uU��Hmkt�̃l2:��P:���5�pg�#)ĉ?­� B<i���O[�q$.w����������N1�U��a�~uN�'���5�S��+2{i����U��t��S噴�!t��~�1��+��Y���k^^g2�B����bV௺�4��urt��R7���5\�1�U�R��������ўd��&��)t~��㤹rGB9.�vq��
6JQ��q *�u�݅�E��̀���m�n�l3�Y�����流�٨B�n��)�f؍)����*��['��4'�sC�Vj$�wBj���+�{�k�I�����U^0
�nFnj]QG;��>N8l��T9o��]����[Y�O��T��Ӌ��-r_'g�..s �L�azuV�GA�ՄX�!Lf���r�����X�d�.E�Zs��.�]�D
�y��ٌ�RP��#
9�b$��I�����v����*��K-:�$����w�rIh��{��XE��1�jD���ƘY ��h.�O�d ΆmBJ�+O(A򅴇G�A�Cn�R�]������p��^����w���P!NnA��de�Ϸ|��M��y��3֭�p����z�Z�_m����'�f=�A=:7�^�)����r�o���_<Mj�]�wH
�?:�����JY�s@ղ�m�
=l{��~ VvE���e�K?"�K8J4�j�b�׹�ب�_�H�p������N�Nu�ִ�{�)Vu{�^�5?W������ ����f�lsm�1j7֓����T&�/Ѽ�TX�C�W�u[Q}r��^MB���e��aԜ ��	��1����6�"����F�XL/�V�`hNvhϮ��j���G�����vI�����_��u}hh���QV�(�I}+An��5G'��̾&��9�P?�s�<�(�7}YA�W�D��j+�G�m
�1�NƼ*�
3����5�A}=�Yr�N<�[2�~��T�O�9W��"/���O�;]��F*���]e�4�_o�I���y�\p�������j3�.�i�������5(��z��c�͐<��I��ˆ��r��m	�~O���0*�1��tS�D^�h|Q�P��
PE(�	� �r6F<����O!؉��9c:-)�O����6��_m�2c�9|[���D��pu1雸{ U�[�[�KJ��J�5��ϲ��8{�|"_�N��Qp�_"y�Zm�D�B#�C�EXJ�>�� 6͠�����<W��_)�^��E0��k�������_c��^@��U^�
�jg_�f9��A���@����sV*ܮ ��v�T�z�n���d�����St�I^Y�Wr���#�Oa`�i�Y�p������"����	[|��a��l�=�l�Kh��6�kLQ# O���v���S]�&y[Y8���z��#4]'_4�-/3�ո��^�H�ɠ�o��4���݀~���4���>��{	N�d`n��մ[+AnpE�J˘`����Q��LP}E.�\z�/Nפ�˒��$�.:��<�������<�К�����)�9���Z�񿌯0Bi�2S�.e5�,h���Y�T��v/�O~��8ꖁC)qP�.���W�kX����4�w���Xih�&k�~K�ۗB�T��U����x}�?�Ą��_�����t���S���#ϑ��}����u�^`_[���Ӄ���ƩNvV��#�4����*�G�YO<������u�p�i���Z�0HV�U��$ @I�໙ht�.�Ԝ��w~.���E��%�m���n?v!�^A4;,�r��J���H�����o����n�SB�]ɍJ,�9er�w��ie.�A�����8-�R&� �2i��Q~��,������I���e�2sL�L�79��y>��&1=AP�t?��Ai�pԔ���xq�Y�;�\"�2���mūkrt���A��PS�B}�(n����u�1wi�L��A�]��Mq	ݽH^=�WK��c��E���՗�td�%�Ԏ�Lb��CJt�ҿ��UN�O9U5��"9ܗ���o�|d��������S�p����P� ��~6s��,½�<��s8��x8��훍�M�w^MwUړ�1�_�(�<q���+�rݖ��B��3f�,G�X}x����v��7��x�7�q�b=���?m��M�l�Q[�-�k�"�m��ik-}0�{pm�|Lq΢A}��!�73W��O�m(�/A�o6�V ^"�1�sW������|��#-~��~_ZQ{�
�]�7A�_e��H���2e�K�Z�y��.�:�������#--�(pWe�s�|	��IR�K�Nʽ��ao�'�[�B=����H�И�uu�c�iس����4J�ܻ��m�e���)G�g:����\aaτ�A�����@#sl��@C0#5��WµR�-�h�`X���"󿣨�oHm�c3y^غ�*W�񢬧OO�~[Sj?�b@Bg�U���	��SEڿ"c�I��7'֝��ܷ�;�<�5��(XGӡ⋥�! �7(���&��yC|R�ʿ��/@�g8��&��!��� S7ݭ�ye1�!E?�̎
xS�KM�Щ��:i:F#Nlb�7�1 �O�[��Ce�Ʌ�B=�*_�8��h��b�΢���D��Q���=&�;!��ւ�H]�?�a��������
�%�0�ͳ:��Z��Ujn�m���z��������w�}��̃M9G����A�=ܮ�8tak�%+��&�W~Uv��]�q>���$�.�kK,���=K
�w%eS~�Tk��W9G$`'�4K�?P���nK����
�7kg^O.W��A�Sv"z�
6X���ؑ�?j��{qHS������Od�_����2��~D��p�`L!r�!c�~0\q��'Hr��O?�Yj[����տ�>�}Zc�[ĜX���ߵѕz�l�%�OGT����o��rp&�;|"^@8j�q'q,�;�@��(���W"����XX֋���ka��>��Ҕ�SYSBέ�Me�u&g
���FG����/خ�h�]�4"���S��]�l#��F��b8�x�g�ͨ41�[�H��kVMH{�w[(��O0A|D�F���<mG�����k{[��D���jFB_:ZQ$Q��m�1޴���?U�c��t4�IXcLٟ�ԗ*�9d�� e8�p^SJ�8���V��ާpV�Uͼ�;d��Ss��}~�b`yυFP���{է-��k�ZY�m������#�CY�c �w`8���p:s�-ȏ�j�D'$6)�4����WΗW��wEu� hEekA	DmBИ���V��V�'�ޮ$�W���b��k���`.��!]%��t{�	�__��PO���t��d��q����kӁc�T�����&�k�
�I��*��j����g�W�l?'�&�䁃b4��8#��_n<k�mS�g6��$5�l��b>�{����~2��!J�����"���%l��8CL��MWc�Y���ml���I[����d*�[*��3����u^�`�tK���r�v�!�\����S_��8�T?�f�=��up�yd�g�k`H
#�Zn��-�������ڋV7+���=��s�$-o:���y;��LDm%"i��lfT�pb�1���x2E�s�@����
��uN����׋�G�}Ik��!Z�|O�s:^��sR�ˎ�)P�	���l$���X��T]l[����D���ߘԾ+�$�J]9��@�)$/��Zp����SG�[�l&�G��^C�(�%>�σ���Ԁ[��Ԅ�h��I>�� �Lf�ɚ��4}�*����-\�24X -�aN�������6ͺ��8�-��� Ժ��6RwT�%������CE���LZ;�d�'7"�š6�@:Y�g���[.Pwr���X�UK�a��c ����L\�b�&<ȕ|y��o̙�/�Q��H8S�qy�Y�:-�]��eb.*��j!����툏I?j��/�2�}��[lIPe��q�|�/��/�� L���Y@Gs�}���	��,�L���!f<+Nw
 $�ЕT�|6,x���6�|fC�#G�����.����g�yRU��q�.�vm�����2�)�*W�'O39⢊���}〢�o$F8����+�]5{N���ǵ���B9���T����x��&L:�&��
�l�_"b���y���t(��3��]�q)YW��Q|=lJ+�x��:-7��8u�F@�+��v��q�ߛ�>{S><�a�u�,��4��gT����u��s8���]�T��RPںA�Ƹ>>��#�@��նb�7cζ��ь��C4[���6��R������ŉ266)��h�3�:S�̞��a_��꡵��MB�t����Q[�ac����2[�o6�m7�L��DH�ܪt�Nx���}�����~��l29��Şx�g9��깢vhz�ϥ9:_�/H����h��s&�٥6�_Ae	��l�M�jS+L�f4���Î�
�3�����U�~	T�V3����7XBcp���Y�4�	�
�G���5`���k�G�E���H�Q����cEay�.e(��̇�E7�uQ�|�jV�M>.נ<��~����ęa��o"K�Z2Y���r!��l�������јx���_�� �Ƶ#�8$�U�m�~�|=��E����|�C��v+]����B��H:�W uu@�|�4���m�	?�/�$,[Q�{}��{^Sf�Ӌn~�'�\���F���q(r;(A@(N�6n6`� H��T
�/��X*o�qT� ���G�K��X36�{ׯ�%V\�����-8>	����_��-#�\G�('\P&96�~	d���%ܺBꅬ>>���T��e�f9#K���v|i��~⾚=w����� ��{��4� C�?���Ț"=�D�z����{bRb�cĄ�[�{�>��|�>z~[�������4`�iU/���F��k����h��a�떧#�w�y=��x�mlٴ�*�~͚�x���wP��K���S����2Hig�Nnb��o74�ю�]~0�{�X=[2�D�G���^���u�.��`�1��T�ش�8�E_
@����!z�qt�����r��&�W����I*+k�Ľ(^�?�Y�/!KzA��]�:�0hi���rO_��e�2񻩬�3Xh�;������`���z��W�G�ԥ��%�[���),q�ֶt^h�v����h,a��ģpU��#S���,(�M��Űoo��/�'/������R�Bʵj��&m��~1� �_T���^D����QНR" q��g>��y�|(2�b��z�l�P-x���nS�����3(,��S�	T1�����z�2@��<�e�B&�mjt���:��t�g� �]^+n8�d�W�	Q��b�"�7��e���F`l�Ր�g^�RL�l��Bk����CI��-X�=��a��C�/�ȯ�����Q�P3\y��n�_6��S�������v�@L��9�0�:���w��5p�y�sGpc��i�Ӡ�P����.�>���W����������vF���*2	vT��Ge6�����	|ױ+Y{"��)��W����)� ˟��v��4�X�|��	<�f�&Z�v��aO��b�oM#�2\�ۣT}��n�N(K>[o�T��d�?�v�	�&�i�i�h�R!u�KZ6z����z-�3C'��jƐ��u��8�S�w���$Ь�0�n�II}�`��3Iy�Q�Ցi�+��
B�"����u��I.ay�#r�4O0'�6��~#��Tw�@�0%I��b������ ^��2Ԁ��,�_0���f�؟ov
��s���]��<~��Z{tj+'�5�bL�uw�i�
X��F9��վC8�yϯl(����DJ��b��>P���Dh�($dwR��uBd_]�P��W��� �6~Oe$��#�F��k{nn蘖 /)J<i�(hq�e�	���P\���{�f�bN���b��'g�s�p����	�Z�0��᫧���W]�ب�7�Nq䋣�i�nX��8��R������W2:a��i���k&�p�$_o�%��W�5��l��³Z-�(��/�xi k����;\� �j[U2g��o{��
�
���|��lE>���ûF��,����md�~��Od�Հe�L/�6���6�Oݟnؙݕ:����5.�^�F��G`���2<��ឰ����Cυyc_�m�C͏�,H�t#�c��M��";�D������R���>�}/�I�����a�e���7@X!�҆����$@a��a '�ž�5�U�����搙�F��c+����s��>����SZ-�TO��b�_��m���E��[,P'�� 5螥0� ���.��I׭5G|��W���#2��ɎI�N��x I,ή���Z8o�6F�
W'�E�?�)��5K��=��F�X�ά�p�5d�͝�~d��V������dH�3�eH�-�s{��m�ymX�@dgU%��s�QJ�������K�B(��;a()�JG��{����P ��ZRQ�ZG=kE�&��ANYʗ�{$a�<�a��;>
�,���H�*�~Z���>c���/��G~ӟw�������#�jw���aW�阂��T�YA)#X8��
fR⏏O�>͈�e�y�pz�� ��|1�F7�K;�C^�����9b g9��2J)��Sa3�UT�<ڜ'���L��M�rVÛ��#�ğý=�`����Nr��o[Ⱥ+���jRb�,�B��$����sy��J&�/�����R+,� �0���4=��8�_u�&���ޱ��vOc���c��x�Qa�����y?�U�x���2�<�u�C �dj�$���A��M�F�gy���٣	L���L��d�j�Q�Ў$�RC�)LN��FP��kLlj�{ָ�Ve_UŁ�5����&EV��cd�y���,��ާk�&h��gl�M}���.Ҟ�����{4���j�wuЁ&���R	�S��K��ح�H����p�xT�Hі�#���貫TcD�u����0�� ���%�M�^uРQ��D��azv�|�����#K�8�0-G��ړ�ҁ���� �Ұ[*����I3B,z�+M�<iU�_#�B��[���_K�����n�=�� ���{+�ꎣ��){�	#=٧��ȳ̤jݵl�& 
.\:�(��5���[��5/�����.�������ga����L��4�OԤ,a�8��n�`��ς������8{�s��_�{���֋u55凊n�1l���	&?�����z� ӥP�����6_�7�{\�(!�n���}�O���3��K��+C4�'�
�БɊe��0��ȱ�{�}���xc!Y��5�H�uĭ|��]�Ν_;�=,=�?��R������`w�V�>6���S*[���[��kВ�p��Z�".�I�f~ ͽ���Ѓ�[���r�y�]�P����:y0&D�+�=Z���Ϙ2�������F�����o���s��6"$fЙsr��]��Gg�X�ݾ A4<��ʲK��ڥ����E�k�=QuT؁��w�*c��ǫ��H<��W�ϐ���p%�/A]̎t�4n�y%��-���t�����o�Mѽ�j����$L+t��-�L��6�h�;���8��V��3E��)0��l��h��U*jhu�ӻ���ʡ�Y�j�\��l!}j������{8w���-1��Ik#.��'�[ ���m�pLv<7���v�4��'.���5�L��R�}Z�ggaȶX���=
�����]��N�ͱ�d�孬n���_��ϿO]�; }\��x��H�� �Nt�U��UJر���v�����0@{ω^��j����)Df�U�$Z�q���OO_��/�l/��ʩ�?�Y}�_�qK	Q�d��^��͓m�?Ep"�KE�w�&%K���ؾ ��Oվ�K`�� %Se��.,���@����:WMH�@��Q�&�eMj`�>-7x�	g!�!�d�u�����Bŝ��~����@$�X?����9šz˟�"΃dj��_���@n�d�o���J� �"V&t�K�A���8���[�u��`s��I[_����M>IP��_��w�l`WS�(+�t�;�sc	0 �#�`�{�Ü�������rDB���Ϝz���[7��s�?⾤��`��x�i�����e���՛����V���.jL~�E�,�,�)iލw���Η�k���\�z�W������"�Ņ`"�e<c@2.�[��S[��1?����nB��������9a�dd�E�	���&�ѩ�Q��,�Q͓2�G�L�x���Q��ٰ��&�Y��M "��Ꮿ
��nũCN�w�0�-�!�Al;�jN�~�����s���=�(�y�blY��:�F��O/o�`}�4�(���8X���
�휜t6�gB���|^�P���6$%3፰�2l	��
+�H����h�!^IM��1�����ŉ���L�^fK��:'���7�V���]gl����
�s�γ����e�%��,隫�/��K��2G�׵s�5�^��슐7�e�=9�T�1�ݚ���O�u�4�9�Wr2F�t��!�#��4	����"���j�u�D\+O<�C]��A��n��x� �;7�j
��i�t&�: ��Hc�P]��5F�� �8�!݃@컍�#ϙ�ч��k�^{z���|Xq8w��M�{
�B=�Gb��)���񾐂�� 
5[j�9��R1����q��޷Nڌ���H��ʺ<��W�*[>�U���J>�Bd4�R� �V�ʂ\)K�rlϧ��7�8r`��6��F,� �u`Ĥ�p(y�Ĝ�y5 kv� <����=(�s���1Ǳ�{�I F���?�����;���`'��-����')��L]�ȴ6m�%��N08����`ӷ�x[dW?���&x�>�oW�ij��y�}g�ș:��K�Ǟ}��-�7�X�Ă!FBf�'V�"�.x˧ĩ�<��R?;p�?�Ŭ��t�l~����_\߯�)��K,f8����Z�����F'��j� �$�H����0Ր�iKʊZ�|�t/�6G�3�M+a����?a�+���,u�򽅱R��v�W��9��ݡ4�Wk �,�[ܲy�ύ�v�	8M��T����,��L��ͅ,P��z�/�
�Fț8ϓn�����溂����X�Sd7�S��ݢnًtcQ���gd,���!�\���^K[��)�M4�}�S���L�*!�.䌈���R�q����)Ԭ3�w��(�ּ�@���V&�z��۱=pE�KUQ����Ɂ*�҂s:ܖ�5^s�7lkN3����x�;�R��c �psg�����:�QA{3�a!�h��MN��)��!�25T�<���C�h�o�"�\���mU��J���{��O�]X�=����T8,7�M�ؓ�Z.���j(�0��vy���tK�7eKe��?����L�MÜ�U6���T7�g��ϡȻN&GyG���;�֎�T�:m&����DS�r�t�u�5A�칲4�X��4ɓ:_�� ��=�J�#�K�f�ډ�tRlv7j��rۥ^c���I$��u���Z�b�p9(�*��I�Z�}�A�宩%6��9O���uO�`�ic!�����`����a�e�F�}�*1���u��A��~x�ؤ�Wِ�+��1/�4��H����z9��;"5٠g6�T��A�.�W2%:�|��yw8�W2�l��+��BǦ&?��6lˮ��0F�
��#�6�ś���^��6�`�aF\B���Г��)�ށ��`�� >���:� TSL�!^_�v�|9�Z��K�*����}1w��`8M������"�S>[g�>J�_3@���蓇O0��9��Me����Լ��ȟ#, 2�s��k�|o����;	��+$�%�����ʁ��7y�xn3e�A�dFJ,6��Z��oZy��_��ӛz�8Vv�v��dF%�Cp����#�v�|�ejĔ�M���۲�F�����J�¥{�P�;z=pq��JH��oٲ�ϳL������F�w�AJ����S�G�Րٕ���K��`�GHB�̉��G҅lh9�"��̚��wX�fX{��"t�k�̋{�Bn��YNC=���~����̓�/SRV�E�MÝ��x�I$�G�}��a��E�S���-ۂ���^M
&�ѨI܈�.�@=G'��&s�?D�Uk�B��#�d��T��k���7�_�f�,�z}Js&���\Jԅ֔yL02���
#|�K����O�rC�~p5k#� ���/�V���]oZ%tb��ސ���L�~��]��ݫ��]?���|k�.���~�hm������xt����tK3jFq�'AO��.m�q��?cճ�#ykg.
��F������4��o��[���Hh�1]T�q7sέrmC_�E̇��(	��[����8Ap�d2�E Ԣ��?1�.��+�As�6�@�ZTî:��ٰc(#��ї���U�Ҝ�w����D��	井�����-��r������8d���U~g=�3�q�<VG�,
q�:Q�a1�Ӎ6��
p�ZWԻ�#��X�r_�ԇ�zH�^b(±�$%66|�Q֤���)���Uġ�}�F?��kt��%'+�gR�dnϺl��8�)�C�h0�����V��&@Iq*����NԄo;Lm_w��;��WU�F*������ߎ�& �k �YB�b�����M^.�n��/Ȑo(:��KE"�Q�"�d:M7��tN����v��
g+����,z9S���x䠔�-8�La}(�+�CT5Rf ��b��2GL{�4�� �3�mF�ߦ�G'	�(f�7}i�{��ma�p�5j8H�W[�[��%J
 �"P��P��̎��V�eS3�54��5'F���2?�h���l�Baӭ�A��(���ȧ�ȿ\F���#�~Ȼ�l;~};��q���>��[n��ͷr#S��A�V*��V���ʜ9x�uu��Ч��2��Ɛ���������1x�YmôW9sl��KvFe-��
8�x�%��qo�Q'y���CϘ��}��ddQ��L�"q��R�-j�G��տ����؃o�Ҧ��Z�^g��ɛJ ��f�
cf�Wg���x/f�~^^�0�H��h"����Q�}�u=�b�Us�����4YB&>���i1V�@,HO���O�ΗR���Nz� 
+345��V��x]k�{��tE}5�ȵ�6%]�3ȴ�k���{�K�O8��O���B�4���a�y����t���f6��7�;P�������H�!%H�n-����խ�����tt6E��άs��|�i6������؀~L>� v�2��_�4�[���L���cxG���x�r+���%WQ��(���aq^�%�����t>\=�:�lєm�{l�r@�����$dJ�;}K̅���ҡ�3�ʴg��٫��7�D˴�%!�!\Z� ��2\�6�B�Q=�G�M�B߉@8tlL�s��0 ��34-�q���A�:�H�C�ko)��c �~�!���ؐ�a�P'���Ok�]ֳ��a-��
���U�-V��f �E�mݰ㉯k���k��D���+%���^���nVS�,��Q���҄a�'W���0��C_��H����7X�����Gk��ơ�'u�Q��xS
A���)���7�ee��׍:��ult=����ҹO���_���}	�=���g3��g*_�'����*�duV�ݨ�ιԩ~M*K�F*�G$h���Y�@I�9Z�>��y�Eu��\�.�Q'��X��66�/�A�n	�PI���%ej���
�w�Jp���"�y����j�
?Q���[T���<�3�zl��h3��|Ҡ����8ސ��c�Ewc�BC��ϵ*�E�/����E�<����!�i&��l��[ɗ���d��v1OЙ;����%�!xe��0@D��1�cѧi�-��v��6*}�5"�*�C�'vPciD�r��f���l1��9%���S��$�P�w"�-��_���g��Y��{�n���'Ov��f������$�O��ᜭ��5�{�!(J�z������%��~�G��C��Sex P���,A�0�����Ў��ts�X=+��d�����XU��.�������=,�d��K߻$w�F��;!�|P�<)A�V�p,����S5ρhj���(���PVb.9"2�=���8>�������vm�}�#��:dr��c��rIl��r���eF��}'+�Z5�X�C�{7�4@D*���������A�]]6���W��jҫl�c�y�\{g��H����1��(��<>{�E���2�Q)Km��R�>��y'�0����&�q���!ب�&�-�f�$ӑ!�M17"�6�|��O�ݓ#�xquW1u1"�ߚDV^����t�S����E��gi�u>��;�8n�T���5h�5��9V��TW-��a)��6�7ZD7���CVD��&�W/�[�y�1��R���i���f�.��9$�����d*-$��B���9l���,�OF5��	�
8�"K��.t;$��a�L��2�*h�bRs�%F�����!?4g���2<�����F'Z�突Z�� @��ڙIZ'yh��q}���wir<���j�#x���qW؛$�F�!�_+�ݔ�D����0����)qcld��Ȥ^=m���e�P���3itxiR��i����v~��M�(Iځc	2\���%��Jz��>���o�����-Dޯg�k~���v6��?��A���»��
���ˠ�G��zK����?�٣l�~�^qv���x��oH�A��9���(�]`��ؠ8F	Z}8:������-��!؞6��x�v?[�r��a�J<2��A���W��Ԩ�B��\�B%����L�_I�V�+��5�곦�����KR�/N���Kj�ڴ4#��n�ߙ��DKQ��&��r��ɄI�V���H[�U�x)@�y�J��JE�ν$ݘ\��K��PW+�q��tا� �s@����iFVOJEq���!��K}�~?��.����Z�����r�ձ�0�t	��� �� _�f�Yq���}iA�l8�I�u�����2|����\Z~�V�������CeܹمHw����1�y4l͗\&-|�*�̼S��<җ_!息��.���[X�8T��eX�̞&ت5�i�'��������2�y�����h�����"�<�1�S� ��:�ű2�Ż৵�岑c;sv�`��m�M/H���eF\�s� �X�p�m���%�j���S˲�!4�E��/Jߪ��V���ӌ���䠹 ��>�H�+��x�\�6��]t��w/����X�VL+��#8����0���FV���DnK\�<�2�� �~��%�0�1�*�1������z�����a�q�s���޳�����J�P%�Y���R9����I����' �SP�?�a�`���;_�;]ځP\Ѝ�O�1��$1�������č\1[oz�F�̱m�s<��Hd�BYH���5c��,��j6Zm���k�\v�p���3�P�����|�07��b�
f@K�ȉ�4�E��P��#k��r;�ct�����^`�T�*�l��8A��� Oj^ֹ�Rw�J,FPS�^���W�$<z�S�棯���>�eC��ԔU���̑o/�$�pH�ʑ`Q@0d#�!t�sc�=�X��4 ��s��9[kinh�@���<$W'��F֣g|�������r�|�}�m�f`�@�C�ݺT�.p������_9�6���M�c��*�wǟ�/`
�
�N"dU����Y���_�^ԓ$,hœ��ԃ�s��5�%����M���B�=��F@B�z ��xq�6[~] oIYL;ơt��ǯ;�邰ޗ�#�	�8��	����&��%+(x��i4��hH�"A�g$$�0� 2p�{Bn,]���:I%\5rX<�WZ����7�G�U�Clt#�la�)�e:����f�ì��yϏ��VY�S��5�E�t���'	S��/�_Sg��]��s��*��[:M$���o��¼u�)A�3�w� ���Ij��V���1n�D(���O8XH���O	�Z }��3���)js|b�I�A+��}Wt���xSJl_��H�7������۪��^��Y?���yPݲ�adR���ݖ;E��hH3�m�_Q��}����	z4S�����D��L+6��f�c�&��("�C�CV[���hσ+�ڈ4�J8�K9)[Xn{�%�gKg�ƪbpQ�p�D��s����n���D�%�7�v-)�,��A��d:�(�vz��J+:$������HƄ&����RQ<Pq;�s����PN㼅1��Z����}D��f6.���~�7��H�r��+y`={x�����u=����2��$�5��Z��Y�M杮dZ��_�>Y�U��y�u����/z��L<6���R9�_ۑ_��1ñ�M�6�*p���E�nk�v���������K��s-����,ٸ��	tFJ�P���D� �����N\i|e+�X��� _�%���ˏ�.F/$2���zM�">����2�=����Ic�$�KFƓ�����]K����8A+���:*�����N���٘�H��+k^�gS��FM[*�6�!�E��׮�IX%ԅ���%q��J��J<$���n��*���~�̉��'���8w�B>�ƍ�n|�i���ss��1� PM��؋��"� u�Y:�ȖQ�T�Vy�E4s}��4c���*���nL�O���
�j�������Ub(?�`8�o���U�-��P5�r�s�y� e*;*4�'���W���������ђy�f��xC����-�M���he��������ʖ���ߞVt�b�"L�29�8	���ڂ�ӕ��K\���:m��H�p��8�,#8\���ƪ��6b�1�gÕ��ĺ#�7���lgHC�� yd�]�����FZz=zH���A ��YCW�on�\f��WR\�K,Ի�O;��0��@ؖv�j��	&�V�x��2["F�A2H���Z��dpC]�|0gL�$�żD�m~'ʞu�[�5.	��%�a��Z��F�\��.��	��&�61#:u;h�8�!C�g k^�%�L4���J����)�5��oY]:��/S�vq.��<

����q�!����YY��]��TCg�/��Np������'�UjtI�L`�����gdp��3;�����WK�rE!Bȥ��������Y�gS���z���;��15��uz">�����M�G���RZ�\���}�!c ���j �W�38j��S��K�Df�>F J�Ke�
�HDr1>sE"o
��]� �-z�3(�z�7'ۯ4v��,b�Ô8�z(~��s�;�t�"�n"&RH���p���տ�Z��&VB�Z2�}6�V��:ߎ/:��.ig���|$�IB�;�ӓ���˹��K����%н��^��ǣ\(�x��2P�g�tX��6P��:��#�J*���x�X�o������N_J,�B���į8j��  `k����PF����5�a�*�~*W����k&'u�p��,N2��g�-�
�����z�4*Z^̉R�7�8G�� ��'�hN�3��(/�<L8,.L]�U�;��[�