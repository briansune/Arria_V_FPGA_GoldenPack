// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:17 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t0rArzRSlgKb3WxSOrje1/d9WMnfzUGk247ONCo1AxIC+RnbgOeAVkKylRgiYklk
zNi6ug87mFzOppMN0tL01cRLoZITEsWjMSkZQJvjb+PbHc/LgIPhz+iub1DK5bFY
2CLZd3OHqUzxLKz9LmlgDGcbvB6xUMi05cJkorPzo7M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21904)
cSJcCPI/DP1QH7sgbcPmFwOd5La0pO3ftkcEln9hKQTxVTJiST+/ERNhMbSBSYCB
FnU7VMCBCgEukICSDM8JydJ6+AeaGG0Hmi+VRhXVPztUjbTpG3ubjImfHgml4ixj
GKeeJelaJgeGOF80SZPELG+SiZPwBwCPpV2h9giDNW81vdaE0MFtKXExawOJKR1T
1i5ADzV365iaUogrFMlna9EBwjfy2gOf/mC2lWD69FvPfb3Fr2MfLvklFL1vJsPA
H55JgXdByZtYZB+l1r8fPdKrFRDznnd77qLcAT6nKP1WdHczvYBgr5x2RcGVuiFn
YAUlR8gon6LmEoYOlgsIcnb6G5D1dfEeNbn2tDMT4/vDudlJH7Dc3xj1Ue6ZkWIq
UQwh5E9NPwKOndnJAz9blEIvUvLOuVTYOmTNlGBsuMQPPCEGXZpMvFoLh0FrVa3b
RwHcI0sPy11wPMlcO7hgZLkr0tbuFfbQLc8RFiV24dCC5xdWMUKiL75ZWKxI4fXG
Nxxukecoha71BmFgaMMgNtS6Y02DxddCQBZzujKQOv77ESPnhetIlfuUaSwMQDZR
ptVZ644YZVH67THb7xjdyYlUVerHsc2B0CkcTydr8QI1b6XV5y9mh+B2M3lv6QNC
uf0XeTElMrd1gQR+/x4BQ5+TJnL+FgkWar5+1hl3g45deLaXWC+u26dnBsYOxCOx
aZytdixmLx+r1HKAfcEcY5CLJkslpvHk0HFjTyVAziQ1uqkRh5z2wW5ecHqA5cWf
YsQb/I7qCEmd3VABKHuRVk7Fg8VHpO5kFYIJYfrBdW8saWr0LIok3ilLoyP7LLbd
OysQh7ALs4q5urADfudTsxQLDKqqAZx4T/9dotWSVU5l0YgGDuDGR93TcKqdE/7Z
arN8a1l9n0kCZ64yAdYr34WpC4LKLNvGkexu9s1SCKSpFXACwelRLeZzu78eZ5V0
hMIxuWHNVTV4egh0J7bV2OqWzmAuddDdGnYvhHpL+2+iRiiBdaN6qw3WEoiZcQLk
3Z6NMtm7Oh+zjP0ZabEpygMJDOxeqFdONH7OLya/5SGsMf/mtHj/lWKQWKZZK2wR
AwAjUNDBt744SdOBZOFLxNrawbNjIHFbwMBST0WO2sjl6AJI8J0HnxzZBj4JNgfS
6dTbahPpnC3IgQ88oRhjDJGiyiUBSvRH0OqD/pUvIYNH9/VrZ/50X/4H/bq04w5L
e+NkjHb+dhpmISVv6FL4stamng0P0dsQyDdPt9jsdhXAIgEVY1rbqSpm9jyRzlGM
PVYWIiu584u68uyI2IDWM5o+y4c+7ucRrWHuK2q49oSk9sNIXzZCUEEaXBor9eUJ
0DehqgCmg+7u40QuyJkWM/MGShIjErtYk8YBdGyj3To8MumvWaHEM7+3mS4VDh9y
aLPWaBortPWW4+DXwdJlUpeQUFSo7/oUmgNFJDCx7/7l27cL6nAZisF0cZGUuYop
7K1blNiZTL0H/tfSxSwNWuwcseHFJSr2OE3YA5NWajFCz/Vb1h1CxXMbWOFLNySy
7eNFLOnBiHlAicPYZVKOIfRboghA/7R1O+AkugVJH//26lP5Af1pvfCSp2vKucB/
DOVJyd58H51zfFT5Ku2JuF3daTh7zY5C4HnDwRe4curyPDttwZEy691r6/1aL6vX
2f/8tykAmcWInx5xiqRWKZ/QmfDDB4xg+7mbyq59Okp2iXSr+abOn92buimMME4o
VfvcqM50XmrXOLrgn/GCWHNGmB8pN6RXb3y5Axl6F3J3zIWu+W/RKj2MsJ48gexi
UWWZ2VuXiJaGKte3Kq8AoPW5ejuke+5eNAw9h3aXvbUuN69YrKkdySabsgoE+e+p
E872ePYRAtYCk3okrFNy9mlbeQYmJNTRUCwFAVKqlvYzZOfuHyAx48zypgj7Dy70
Ryx1YNpufoKhoM1MM4ik+ubJ2lqdowrH5CfyTtxToJEUM6OyjS3Fz/BMOMsVcABM
JBifeWHbnPzJoFTuo6bmNuKMudBW2pBOW0cFDDnNxF6+UdUUESJB//NLaOGFv6ib
+ru+y4wm/IYPF7bGuSwIJmvl5emSTh9XujNEToQoTmLNiV9K/5TFRiwWzuoFWT2O
VNPupI7hmrum0z6ZEpC5vie5btmp1sCAtd8PrcqzCtcJPUK5i73tVNKgQzEvPCvL
C2PeVEgB05zdDN0ntyql7yYdqkRGRoTnZIUKp6vxkFtipWmPmizEsz87r9qe07Eb
7zIfZOa6vPkTMbqRqqB763joxYGph5aSpEIBe7hBCp+VzirLoIgKuQyjmwI231Sp
oVAy9578MGldCNvlRNNrpCoP1dIo5gdtZSJ44Wdc0ASKSa+Gp0ZnHzJxuV/QzI/L
zqb+9jD8tAUOn3BrNfmTFTbVan1xwp/Xbf4eGXWXktbQlLtYCeV/c6C9WO4BHg3d
UmbFxSmf5EbUiEO/PltnaY2wRsnW+GyNzmpFJkly9Cof3lzm71/gOVdzzWL0fvQ0
1ICj3a6JSo7cuEOvw5Jtjpk2AM1lrS1R3JMN+ofVULeKLQfgHFtwujREiphOtuke
tWJ3Tzv+2/Tt+74y0DDdtyzBfLvvsdRALcJQoav7q8yCQHxtsjdmRoJslTyyS1hf
Pve580GBvOBj/ljFyNMThTapGggUYBYbtd/dUsh0pF7PIN5eyy4PTu1sngeGvBOY
WHrxGfgxN5Xf+eZR//rVIFZl514QCASLUBqdCUMlTEoGEaWvhwmQY9iFRZfdd9iE
qis7qtIIvV6E11xpOxLbMARuzvuLd+ogvJf+ZUbHUWUxUOycjrzTDJKZz2RodgTa
S10b1pIDMWeI3JwQXrLs7J/vg5YFyB8M+PkegJv5jY0aW0qQHJQDfHHd8L4q+Ai3
Hs8JJjnI6VYm6NcXlHXOOjcCjXBHyLd1P4PgHU2Q2qF3tOW2Ux0bqIEXwZrYcxKH
CA++PM+xH7x1Eq0I2EqipTMln10uXYM5jWBT1Bq4lKk5HnGLn3Q3TOhXV+cXqL9J
MmewW3sVZu/9vFRpXWfjSB9o4IzoryuXu0FOMjFe1epx/KClFC45AxBkQnCtTjZQ
WoqvqZkRYMPN+GHo9YSwi7xd/ylN3hEn2l9Qn7NyCgorSyLWZlmjzBXHPEx58qY6
7iL+VdBlgw2HzE8pOCm213cfP0PaGrGG51E8uf5yISQHgkH7Mzo62PsZpLGT9bAI
IPJSy+FB4GRZc7a6PaBubE5jHKKbelUbVPvOzoF6m1rj5Wehnn2EhqHx77PxpDel
wBNILPEX/vVHPT44UqDefGR3Ta3OsR0hUkgsGpO8DLqvJMG04DpcX2yZ+EdYnI0M
GCsr3Ivtic7ZBKI784Ur5L/N/W09WCqp6DC9VHUQlRT5HOUnEjw34WRMT2JaQwdq
xizNbzYvnmnXChwsPifH7rW3fGyycdAdQbSyt+Dql9rZrhoceW+gOPiCxJQhiiFL
jljAGMQc46lxuy6wt4H2PscsDCRXlscPGjEdkTM0oDNPRJmIYkgaE9uXkHU3KMem
DODc+f1h0D/bx2wKuv/Loa/WJVl4LrBsxjPjbA/ix0FjCzJKwtlrQlEbxry4r1jv
qoSyuxGGymk2jYWwiYqwfSzPuFW9L3y4Ip1AHJzZs3PBY2b6mPetoud7a/g7eVNY
higjcI1CdzS8z0NOza3328mZ809Uyn5d2aR0ue9nFnFM2WWwQEXpu0IHKQ9iJhoL
2SsaskhwAC1zoCAlM2drKaGDjYjnypkv/PQXx5oFw9yOakAhhpULwlbaKVLaFEjq
XUXNzT8zqEkZ5OGK/8ESSx+2O+40sqhbBolXdg7ZxSuh98peKpgWQLPJZW7b8jl/
HuJu4jzYxHyvecxRmGzyEBQ3Xf5ZMPOBSuZOOGAt3s19redlmx2gc+h11gL01FN3
veCVreSoitMXIrgmHAjbA4EKs9wZ/4sY0lU+KrI+A+RntpZTlh34vmjksUGvCNmC
KB65ayRu+3b1wR1fL9rmBVChPEMPN3xBTungiDsii17z9QEtAX2BITgSAVvzGn25
B3zPQzhkktlok8nxMwyUL5bOrOvlAqe3FJCbMFjsC04ORBoFe3vlCTYbQjQJVgOp
slCilsjvv2gzubXym3MxJ6qQ1bVG7/ZOrZiAKC0VS9GcwYMshOgqUBTHEYjZWDLF
17iD3YIxGNmjwdx2WDGmVSQuzpFMZ/F7s7hFjpQuR1xzp6Y5M/sxPXZDl0MIcCOL
MotA4sq33a8R5EoK5/DgCTBmgIlthZAKsSEL+6TCPgxLqgK82HhRdJywU1Ba1gE/
xp1ymIVVaOeqWQtRQbKHhnZR7W95hLgtjV8ty2aASQkWYgUYV6ag1d3m9LzShHG4
AesgUxYN84u357NSyPegRix7SQkdGW3fFRAiSDrbBEujoKxC3/7196WhIh0MWHpK
7FLbbTmRAEHrWHo5ntEHb8AR/Y0vfgwx0V8f0Zq/AgRnqW6sI+9rf3FnkPZbLyc1
ufU5vBI9DFmD7UP9uBcqTUBWGgIaQrEScqzQIldMik7yOzfSwJyTIGG60AmHXZLk
5yZwU71xQodMC412Wl2Kwn8BR8GlGGOofNJSS9hOfNN5WypUJJ93W52M2YqC8h8X
DYt8W/aLADzdY6XPmeeVzQPkig3eontr5fpF4pXdgYAJdLb4EFVj+a7TXJ3PpRBQ
nJNKoHcbQ5Ifdbe0wbdQTXlgw3MfF89ETqGE9Sh558tqqE2q0wGfKOCwofMk758u
yS15mfNDTAEDa//1dvxmyD4SkPYv1e6z/FhbTfkUiqVur0Joy2GbBH4PS55tAvkz
5k+IuVYFRl5Z0rEZuJW75u135sqhkK21wIz3Mycc+1V9ggSBeTogLR+QhVWvqm7X
7fWhdFDLTYfNZSlKHWpRnv2zDp8RFGycwuWpZrYZxr0TfY/mEIAaVNc/wNOlanmw
JsXSxcpIyuMMo4+4gf0AXvM5ckVwCDp6cDgvxzkcMbjPyRNZFISYVV6M7PiXzBc3
+OmrIiqlN8aRk6jKT54Mdr7S+WSlNI+zufT8/ebRrRfdwLMsmuvFbRUsCqesesQM
QjQBRERkvLd6VWryWAznKpTbHyQK0qO22/xCM2vB0gbSVAGkXmbOw6l3qEtum+Cv
5ssbmI+D159yZtwOJDdMonbbFo1pFdzvJBHKQzSdP3p+vTvYYFb/eHNxZKD25wFC
HBq011lMcyOtRqq5HYGFhCV6r2QeaJap/hNpG1OTFkRgKupXxyAwihdTDhnkvERh
a9+cyESdUxHrulvz8BF+zkDrMMUzhVVmHs+psaaAnsAgtw2mzL8HZpUlXicPlj+d
myttzmRiYSH5DIdw0vZNJRXlw5tUavQdR5UCzaOlOUlbfV2kjfFn1BZq1Pkatx5d
HDtWKVVJDdgMKpJaKMjOeyXwhW3n3U2rnakwSLAF8yy5qJYLdIAi1yhzaCFYHDzx
qBZUT/6kKsaBGqNsvsVa02AcCiU3s0SWNMiYWSNvd8jFk9f3fPN/tK7FshgBOxzu
k/2LEPhmKZ+aAJZbeJgczizp9TuBWD/d5UUB8myb57WAaLtsdtCEL3hZOKp2pgIY
XV1SvRm/OaP6eJ9Fj0cPZQ3OdeqgJMyjyd+Bae5fPTEGv2BpJodv3uIZCRZiF2yA
T46JQX4UToMEpvnzdlJ5eMAtqNos1RBACe7Qay0LwQS7qWqftbYtj2Meuy+B9Oe7
mB+isWSv8ZU4goUAVlVeUsxzwbLWRhUjlrL6ra2WrPSttOD5AKtPh7rSfH6Y/oes
D8d53bEkTKnygaximS2ymz/qajqroC9rlzu4QED04mbzRGKTOawb53mPFP7ktqye
K3SOBu7oD6JhJDzxl7SdefIAS+OnA0e+8dQsjIBDBesVbS0ZPuV5OjaaO80jStdv
RZvp7rXirPNhveRiV7RXa2GdJWkBUEP6PB+JeLhG9HYkcrQ/g+X+c3/ZnMp9K7/m
FOS0+mPnMghZLogLPf7zcUXyV6u3cDMw1u7iydeNmwUXQE0KnLLFMZDcuN4s5WKw
tzB8slMoCQSm4gSxhFgu2kfrChyRfe0+OCpxnpF8LD3qGBBivtiho8s7EXKSQUIC
ZigPZlE/4WcbFRltXF+N+axYZVu+kisgtclfQKS21F2gWkuH2ooiguMBHX7/KnpH
J0KXzuveLgWh8Q3Bj/Bsc7s0h9HE8j613aGSRLVC/ycneglfcSz4qEQspWDsDjT5
t4DzdIEXYjrGld7ktLRiCojtHqu7G2H0Vhz0rdZk4YUM/lT3RL07Vnn6q/wmObEe
EZsUaQ8gxZagMPm2WKMvWH1HTNTzMcx0NYYP2l9Hi3bo9KGYo70c7z5/dyh+ppby
EvL6BvPj6ndqFp1m9P3MwJklrklot+a5lCNQgY+2EunbDnrwNeEj4lLKlpFG2eHg
k9XW0zWPmZg46G/VUWK2CPL3KSBgYl8XMoecs7btQc2OFcTKy72k88xjyeY/3PaJ
PcqfesAkhEjEiOwWjhgNhQr3oiWgfmRcuj1H2NfG4Zkul3/PLrGha4oC/sw5fyS6
0IRJFJ+E6d4FzfqSuJ4fR2gFPARSgkwDKOMmmtw7yoMYZiP/vNlPHqh893VQAFFH
iT5dyBwGukDIa+52ZkiUUYCGJ7KHiTYGYIDaVCw0XfGLcipI8XrkPpKBTkIvqb2n
QgmOyL/rNoTosmVQ0uIsf1DLPG0ZDSKBJvtHfdXwKnHUJR2egkebySK9yAZKQZcz
1Smqdc0AJ01rpws5E8FP1EExf1cl0E5IhfhybSQkEaX6lHaYgZv95xtEgJI7h5RO
0KnqMR3oZ9OmGQ7Ast8XTak8Y6mHH1Bq47cBxSAkK14jCcUfBVwt0pqwms3dFX+s
Odh1D00Tl6B27dibTRunK066jKYunGi57IahrFBUDgldqDYR2Qe5le2xR/ZeW4kH
r0OvZjtquBZVoIHxiunLuUTEN3fHdvTYHgWTClEtn2LkLMNHuxb3nLoYw4qSR+pT
Zq7puMdwh0t/3j/tViMImjgSr/iuSGrmu3NOuIqRIz4dO7Sl00WDToMjn6HTM+Ck
uMajCqe+0PMyx78i5Mym34eDuCAxGDJc9Btkma+ZK4ufrl5gTi4h4rmWLIU7940X
3KIACcBZxl2Lz+qEzqzf1zdhHukwpDiNnHevX5Q4ZU6DLXkP5RI/lLYi49s69Ch+
M9AYLWMSecNpJow6UfnfUq/3DKvUY/ifWveHDjNcPiaE7bQ4uYKT7OMUS2HHIcnt
NemSJMDcAuggBBWTjBPf7FwX8TdiHvLE3BcKTOPbFvzEo9cJoIXL2aVXC/lsnx4q
3nv71oISkTV7APMNoYgYIvyl76SZo4qvjERUTJj24FhbtYDL+yj2KdaxiUY1LPW0
vGWICMhRhrwTg+Z1q3mhlQF4VcQZJdD2MAaYDLhApAlaSOW+nROQkVKQbaE/5inH
pk+Eww8+i3aD9vnNs1dg7/PNoOx5t7HFuwHc/FJCQJUjvoFPtkJ0/iqDyAyfQyTf
YsqWDxaa8eq8G6eyJ92mPD9Rcq4gmc6YhJDnKwBypyHnRGwIfopIGLvtBVcbRxDU
qs6V3ijRKO1nvpoBcSbQC3ZmqXzo7C70wIhmsCnvM00dTjxVcCrQQhxwntswPvfC
v8Wj/LP89chpFoQuKLLcXLXsqmOW9OMhxxxQKX9Zy1XWJX+Lr83cKUZoKjD1uJcN
16W967LxJQu0Qvl5+EaeIPCk8k8zF5oT9dMfytfaBsA8LdU1dQYaQhXKKYwW1Xuv
y5InTA2/bjxAre0aVYLmnvxURGJPSCPjXxO6NldmYLS/nkVRPewxHSpKk+huM/Zg
9WicaK/w0SIDDdJUiAwkvmU2SrGzvbIN+7LPRfnWelWFCelFX54RduknFUOSBPiy
b1FODYoE1fUXmFYtQCZaOyA2cuzVRYsXDaOjMi/5LXcbJyuJyL4UygE1f04JPi7M
jAW6Vf1HfehuCmf/APIp1tIkjPMhqxQjIuEWZLUWpOwO727HHYwpONbHXP7XLh5I
+/3ATSkF1OPzPyjizFTyxyWK+TL3M3Tnb6+Mr0z/JrD/sWBbOoLRytn2KpanOoys
+N0RYegVYDb4Y1bo3aT2wtdEKbrES+56pY6N2qBj4x2lWzBJNGkYTnjvbNlhusKp
clXnJ77Pm6cJneQ8/ORcdc0Ouy+PqtSj9fJ2nacpP6EyKKcWYvwKU/TaIvHrX7Cz
YBLwUX6X7RfpGtG7EP5kAflXKNx3dJjf4J64HFirrnZV6QQNl+ohwSDN8dLIrXS1
EUTHLs9THdeZZZbw7uxFhwHdJ6s63IwlXZGGZbfeepP9T3VI4YPzbDEvMB8Z/81f
tf1dVvQNL3hcn8blzy1dwoMui8Pij92I3K1Uh1wQPBpIYTUqgqGsuqfTnzOExN3k
crJl7kRmIe6GBsFkjGE25XrmUrye9FYxjhAeRgOFjjGoKPrxiUIrg8Gx1Y3C0Rcx
1hNV8Zy42h6rZL7sOri1zL++rJ/2A+N/FWDKEg+HB6ymlNd9B7zzlT1HtRMTOVhg
WrpGWjpErh2ZdqK3FivOZDWBt28RcP9Gnz61beCXL4ixp/z5CkWxl38bAz3dPMZN
ijxhSN1Q1+5q7W3+cVPAoCaweVrrgbvKoFjDNOHRUdZwNDZeTVfZJs/FvQtSbzus
uaLf2iuiVFcw39CfzudGZ9CpxnY6B4S6iXkN8KiL6ktgVunNjeMtOWkbNe2TEgw0
+8OCEI94zmAyBIvm7Tqdzh+LKWQzYsVWy0wBgBHZkxi5SppY0YCV4PxZZUuiVkwZ
fkUqzdCxx6dcRgYJN41mI5JnD/8oEgC2G00NGEzB4k4oAVWeSdXMhNxX6QHhIuRe
d8G/DvM9ZWqQ5Xfjfk9q9yHHqy2JFHFgVvxepApkUB4mAwaf6bSedOh1HN7yqJGj
Yie1Qf78/KsUPhf0EGzU49n1Z1wCdxmOfUhCj6sWxhh9ry1VZcaI2NIw3KhSQvtn
vHzbbmaN3NoAZqwo2XrtuHEWg2RBXeo08rvYK3eDNDFjmw0O2NAl+7uO2ndAXBXy
vRIbiSwWxO150LEo8yHjctRe8Wwk8cC2yDvbx8P1VbQpaJTMgWfiBat/q17eG9gf
BFVzCTp7RYdx4PpwCWjQ3u/p9riOysRo+QH786xXTA3TuKb63UbERQvXHxy8WRMk
A5QC2ahmrC1xoOiZ/pLAfkAYWSpB1ksciQ4dQwDW8/p2WCOjmkrbiucz1T1OWKeK
RYhxDb32mRbRjYVvBtnf5ycCtExGHlKlf/Jkj8NzoK0cLTyKBf2BM8MPSJQ/ATxS
rJRGdPo2M+KCC4Pqji8twPZ/uejJWl4qlN+GE16D7KjcdxMpG84j90kYiAPaOzYx
In+jU4meT3rSA/YHHByOXzYTWFJEOrTu7u9YUMddViSt3bdYL/HXnZaPPVFU8d7a
0AI1F7k8KSylQC+z1075lHZhCR7IpwYLcfPtLopQOBVFnZGqPRPXU8H1ffpBcbkA
BUKTlK+pC/BIF9THJC08jKeIu41cmsQmlDpeysCKQv3owi5POcFuBILy3k4TR7Eq
51nyCWVTP1kaUkemrPNQbfJZAGPLMIWMrgde7Rd2FRTPO4SvxG2aKuNFkRskemRO
p+Nlo5LGmN0mZVPlD6GwDu7wfzcuT+bvg/yp11VK9ZU49Ghw5P/phiKHAch7qnN4
SOddknSQF8NTtzy6Hy8ghPTEluPg4qf2LhccQiieaARpeMYCL/xbKegs5885OgKI
ZJzVNsjxSUYrcUOOAlYTbgiZ+dKnZiFP9dxUrsSJio6Mas4H5E33fbM1Ie5+Ajmj
eo99essnp6HR68iVCSqLvEliQCONk/EY6m9NU/cS51Tibaw9/s0meDGW9X0oUm+m
KYjhGCjzEM5c9J5YlmZeTpszCZWB8cE0zmwOO05SayKvpuce7Jq/Ukt3W8IgvqOo
vBc8kq4seSWSNXKCbfJe15LDg5hiPtUKJRXNeIfeA+dVQv3SqcCrmzkt5jhTb8Gz
wlQoSmBpsfrpZFrCSVyfOeQGci891Ao9yetXjnCkNyVkm7Zj1hWUFO+bDcJuT1N5
/X5Ij0V/ftUNIwr7/D44xhtoH72YMnfosDeeTwu/FLRwa3DxLJcPcIBAkcY7ChcR
xO5XYzktA8/P9U/wDI2uovrVlKt/VvyOETQ+zuTqVjQZ1KgJ7xZ11uAUSUie5xkj
yViQY75XsQ7aelEpVg4SEHykEYANmSEFg3MCsAPOwgSD/xz2wvUP0expky9gieJU
hsJno+a8hdrKwJLoDRF0ug+CZArE3oeLdcoJcdkIT2M0auqceHdorC1CRGgjxggZ
5bE9rSLi7dtOw9iKeik5pn4bMJYHoqh+DidSmV2alXZWjJymRbK+w8hF/13U0rJf
l2067YZRXmpNCRryeOwBJvhTaM6yDAZnLGurorPK2/TOgl6oncN0A3PKraHOR1Sp
TZkDms57m4ftuWeRUL449gPRgCUleKaEzjZbPiRANOqxTchnEUxPDtRzPbmrpSmc
7s63prZuj2EPZf3jodybfEX72D2aDUTZ+Gl6w/2+INwqzK2ad+7D4nImALvD6t8b
Q74Vm5apZirBjjAL2nF6e3J5qJ7/R2FVKLmckpqSaQHwS8q0UGQhUDEHJ741RAn+
Nfo7Cn1ch4dpTdfaW18zLU6mh0d4/5cIlclEDE/GZEfBaA9cDCV692R+gBbRUTj2
ndlrrB8YA71nLsw7MPVVTVwztG+IoqP6amHhWCZAvMjskh5BPx2FH2Oh8RcCJet/
sFpbbqSGB9IBG80ysT47SygM7DtqxYp8VNglEvhAUkfcPRgrMkpHVXjbZruBWjzW
0Jovj901r5OtU6OHV63/ge8WnEWJEcLFmpZi57wLujENDQAygtIBhr48qHNk7hrB
xuw0Q1b0a4k0S+9Z7RraNRv5/pGO8gtgjoD8lvYTiZF3/rCSV0Pa5VYnNrPfAcrN
j4Cc9cv0xyLdwR3y7ePGjk/sMsTtT4i4umJ8n5GybPL8+Cvm7TQtHPVB0Eli/DIH
1umI1YsZ39DqfsNBPW9SIE2F7Q8TygfdBU6JRkKymSoTIsVUjk5ItgPwlgA+JL5Z
mrA7K79TMTd9x9C0H+dwx/G0D91pkrGceRwaD3TytsE5rV1odn9lVSZwRYMPtYqc
K94h5IUCqN7t0Ga4/1eVzzvVTVhWlFb7JBje9KhSrxyf+6/WFiHcRXN86jXDtcph
sBxzH2+GRKBqwuDVE1UMR1m2V2d1hVbq1m3V9qstxrfPrYXpO6yCdunzfBE3VRd6
eK/mcjXLKtLtx23z+UsIemD8mR+vH+VAZjdOZE9F32+JuIIlKdUAvk2UNk8faTBu
qa60ur5nhpPYBPD0eSH0W3wlfTQae+avofWYwqvzlRB6QUxwemjn7JpdXU194V0B
HqCinOSmmduHO00x9SW3wlIrlizIP3kJ3ok2bdquaUWcREvs9KdHQMgTNS7tq6PI
SjJ0+pCd6srRDpX78rmFtdZvNPJRrwveMiC+lGP95kTFxjuuJcuDz9YXjYoYCYi0
MPfsu4RXx9kUdJGLFzrUB1xcCzIF7UdGx0hmEzZgYoxARjqpPuefBqgC2NVihMMV
8JVfQOvJa3XasK9AodGF19GpKI+ZGKNsfn9FnyE+EbZhmtt0dE9MkbGsFQVETiyx
5PMOghreKoSR8ofoA9PlfWWYCnW8wBY0pFYpEOVxlprNE/7ASDvD0JSLCbJ2qHES
53AWvSXo1wkZsBsirFdJokO70ILevJzcb/pq+Uc2jQmuA4Iej8ywGOUWblzP/USB
tWoDI4RuTMg5DCeOJrDjWbZUFjPw/N++hW29VfKNwSw1GgnJLENU9/YGZfrtmRCr
0P2JNxnHd2wyQH8IU+f59UZ6w3C+HDA0ORsK1YPW+0NPIGiQuxCM6UzfDVnPtGQJ
APrPSiKVpygDsRnOVkmSbnoRUt1wMegNobfHy8QA4/OMy36cfI9K2Yb3zB92+jNL
DBKWPGIfyjpB7sP+QIyb4OX4VIaFwy9v6+PA9u+RQG1EIKdR9i3Y+QoLuOgUgEhO
wNht5Ii9NKztMhnSQbCt6u4R7fCkC7WPtyO1syt6xYJUxN3/GAJuMG+GUHSYvMI9
JZlYaE6l/B6OKU80AWRkfgPz7EzSqvbSgI7khNrjKQLe9fDwfwEZl9/TW58YqGhb
vxN01/44MyGh/vAFbqXw88o7cmewPiVU95/9A5qJUMbZ0LkUJteB5Z1dyP9Dcv9o
IMa0eLOI8l6gbdtsY1F4LmSYfOb7M7YbSthWxFzlwQ8L4OSbv0RU4zkS3atRSPCz
BbHdG2EMwS4MpRsJfgJZjVeyMbtpJcgBJ19OZ5VLGWaF7Bh9Wa33T7LAchQI9R1y
uTm8icpqUyCwSQO82123N5+tyGg3JtTu0KWdgQQfrPOgfmTFTpAyzR8AajJGqS7P
1KD3JLwCBWjoxCNDG7O7Gqw9huvbPLhFO/3oN9dXT5f40c26vKUFjRf27Vt1ZQuS
498nQ8Rf3gUd5QzR+NauTD7fhMK7xk2WnuUuoejUgKH6zenqvMICx70/IDQVwhVp
Ngyz3r1GcyXGvIk74oxoNr4bZSDP8XqTVPXFt22YhgxEEah6ZtsCL+sOd9DyOU3W
H3sZ4o6JeZle/Lp4JqswoPvKc9kHSawaoSf9RwJX+5U1pYZ8lQOHKZjDkFccYds+
nKYMxQzMK6YXA0dWynp5sGejNzXREaI7dRrTTkfWzBXiBHCyZ/cDrrJevp1ubYDR
XkPGE1196i9jSVekb950wV4F4Tj5VCwISZMuWRJw3ecYsRz58BioyzJtjr/jsTDI
dNVRGwdlWKNC/Era4lTrOD5yemBciXtaFmXZortoc4zd+3yLNO+ttjoMB9Bz77gz
/9Q84+BNMKZvlJz67q7oEDKJYqMeiqPKyQ1leeSBeQKCqWQKTVs+fiurIZ23FnpL
qOGpEynNme291ghpN0sFbxJJTgNbpl9BjOb38fjlP3uye+eW21g39YBLxZ2JRxme
oyvoawhsJl4j+eKlN4x/fp0+VqqbS1h4AY0j4F1kU7icZDk46UreTAODX1blP8yy
zvRhFqzG8f6a70DJW9hjyxc/oTNt6BtAjNeXv9BzW4tdBvytO0v/eG6kOYRHevcf
Ox+QOLMgCa93TSapknFwixoJ3GZib7dtfIUUjwMQruGtWoYUM4upEcbyEvjmWU7Q
t/DyiKLh8G6NBQA+s9rQwRuvgyymflqlzWy5BkI/3XNLBiV4uxKG0HOFpv2dWqgV
NfdqZmqFNbWGNrscJCQwa6OAwoKJ1eSg5wW4eMgh0mSJhuSXa5RCQ7nwjYQ4Bi4P
h8IJUQlZ+78hQSeCh05w7uhz5CuAPfqVGtafC/7fHMbjRupnTMeBD8XezHlyRGgQ
12YVG0ANpsjTVbbF9yPD2YaeYDpyEHfl+tvHagg4F8KQtg2dgp84t/s/zV4j9q9d
XJlkMjt8OTpi4+YXduz3aqFsT6emw3GkCknRrFao3qDn0pBtJmRo8+bfMRYMDJHp
Tgp3HXHLWqNA6hOLVX8+x4A6MeG8zWrljOgaN5ZfrP/tewRTfgqccerdONzZwLpM
EUriHnvfqz4SIN9U+h89j6tVVuTbGdPz8BD5O+9tvRBehBA6D5MV4OUWH/gq1Ppa
qUQK3ONzTd6a+Zy84kXJ4yQrrpNu7sI0U5IQXWcZ3HE+BBeq2l5+PNXLK1/ZUBfA
y6Xyc4GTkczbhXtWSTpHxKhbRQNMRiYsbywD7vetensK9ibLUdzLWuTivkNYoXc/
vsHTl6CleOwZa0XXkpk1wPx+DgrKjdXYdUcmJ91aaoEPfHWSQv7FFjcanPiMD5rR
yPCxCdM22X5HHibP1fajA/LZaO61Re1SVg+bQu9TeSNe8Ab/7adIPzt4lBtnNCzA
GCU3bp+tf/aj+gQQBowkiVU/TVn0kTAmfY2eqRGQhfjd+R5aZofkO7Wwp/23hn58
6OGjXpFJq6+H0Br1Gai8KfszEWSDWAzFAtH+az/58vdWDmRYs8X6pJT8LYHrL5mM
/EGhdtX19Eu9dBNqzoTNKIu2j2TdEtJx1LFSjLYEAcbgbI0lC9l4sm5C3nRo3Xiz
3LkeZdqhPmlRHKi5Zmxvy63ZfpPOs3zsbp904kB+bufGVWT39hDq1ax+EWL4Rnt6
kTg9jABBEC1WjTDLbvLGmaDiYDIwCk5EGuFHB7GnyE3q1slZ7ef+rbzRmXDBpSQN
u62dhBOai/dtVNaq1KLN8fOQY2UH5xzxcSrpf7+kp9q8qgrjHHIhC/jnDDjqajQ4
oqtboWh87+h6SHlMSG9tdsoTS7ARHfVjb7pD4uwEmc3DsbRu/zh30NwpJDIvsz/C
O1NYWZ8iIYGQdBVi9cMloTY0abuNNIY0HxTl1HkwVwwxJsKnHxu0G6D/uNNXHHPk
CzDYNgVKoQ50N/cH9aa32wDJzSigdilugTnZ5gnq+tcQFnPYiCGah/fa1WF0uvaq
nCHUAKU4yXrfuqwPXnfylHdxQpXyRJ5cnhLA9SzmiYMbiPAsKta3kNFuMmg17pSF
LuYuCCz381hd3lBwF0ytuVRhQDwkSdNTY3vZWOcFPvaif7aOU4CD4bqa9f3PxKeU
YF/H2UpnCiQy6lAsflcaFinvL6UifgPO/IY+xSs67kE5qkdpieoKdYUoMzOb/qEG
POw115jTnu97BUSqkBr6jFDw44U3iUb9rO0fDhe85nixb7iGplR0RyNtScpWR9at
dw8qHnsFyBmlnO+iNta5Hj+uV6M7LRV3TFnZDq9MJFVA37LPjTEKfnup853NmPUf
1LjNxXOrhLl74rTNGlLD3+ypguJO+Vwt5mVSsxKZYQ9E3m+M0VGWEx0gjyerw5vg
7A6TnOcExAA5u8f4MmBt5n67UXWjT83PTzAZxKo8kCH5VKN0/iypgD5fZNxeSKOQ
pw1PM5EFVkjvBHGUY86k05mzX8RGBlyJDiCgkPMnaOeuPMxS5ESOr92xd1oay1Ly
/322UFM5K8X0XrV21mTvinbPX0opY1t+se+2gsAqLa9j1EGA38wxthfiq+FttNlZ
SSSXeNHH5V6xgddHj8agxsxDgsj/DnIdEkpDEDS2IO+VNuqvTuuSfTA4JW3n9rUt
YnZcMmIqs65gisxO/yFxp/71ob4hNDdiIKehKZh1kED3/xvAVLbpsKnUyMTpboS8
lvJvSQNzWxzbmqVYdEtTEgq8PDjWPm992I3f9c32lEO0sKHTgCsRpDG5is/djm+Z
tQAukO5JrJ09UH1EkiuYnBrdhcO8h2wqRQlmEuqLKFeZEEfY5aCV0cfDteZYS4/O
janU9QRHPvCyiQiOirf//wYnrlXSfgeL1Tg7dMUOmORw5QuWHk/a4tbQ5EgI8o6k
Hj66Sj0mr72i4VNUFnokqqDQ73W7IyChfe4KwT/N7/Z3QDqa2JxpVlZ75ZmBiqnH
eXdB5mcXGl1mo7/Ic9S4YVwPJKGk3c+ME9n05aZOpPGhMWvBlxwE36tN63TaAKVn
wE/6niY1rj9U5msHh3DpMRDXbad+ONeBSrsW00G/9F8lOpJyRIYk94XoigWo8ErK
rvOHvPE3VA3d7pH0/YeqRtyCzN601pSc9aNDeavDQATMyFG+go3sCaiS+bHrfyh9
BsoUMmI6xE6syA73yQgIABsOZ7W2TSKCxEvB+fOY6J0Xt/ggWfRsA2ejcmtQx3t0
Gafv+e4SsB9J761gNpsFYUxNpOFErBxnQ/5iRHxJbgUGYM/8Ih1ftbrSpu6FKjjt
GKgEe+k76nmA9HsQJJtkyNpxNMSdkEZS4NCaErDbem6A/dnhIS5GZSrW/J72HaQ2
vvSPGPmb+NsEpXEloudBhW7R/8mRqEdyUN2//BG0lwYwAf3VfanjeLrJoUQOCacH
YO4ZIVz7OSEhSRPWK5TO3yax5h8zEnRt2Q6iBMcMz7IeIjozF0QD2AVqhmGMKqW2
Z3ImKxfKMkSSo2JlAhMzE9pd8PkxaJ6qNYcLZRkB90VCgiKNSt8L4zueqieGF6/b
VItk9TTYD2QtQ/ubiEZ5+EmSn7xl3i/rIvcqOWliY5/gw92gwdPsw5t0JdlkVmom
IhhCnpBEM8Y6rJTTqNwRToTXjhC+EJ17LkAaID8uq+2Xfw2Gcmb6mod4VdCIkd6s
nG+iW/+q2Ymqyk1ILgzBX4a28FoTpKjF9JfJ/9BQr+Lsc74ZfUVW5jpcvKLfALUk
BQ2DHwWFcVZ+iPpbSao4wkOk1LiSeL5FIbu2zqs1CwFVBvMqy8uo8/hvzlvAofzD
jhpHdazujdmuEq7K9Pq94xuel6wMk+mi4vrEayIaXn9EIq3UqOkBZ7NCY0rb0pwU
35eht7vnFN8Kzhxe7kEzOne/HC3xcdag23MpK3WsBxXGaUvpSvMMGLjcRu1qrhqm
ekXos06ZrVrSszrcp/mE3N9LF1SxV8TvJapoP2OzYpbJxrt/2gSS3YQZCbsf37yh
ox4BvldU1qXuTjQIeGjDpWK1X3eJYtZpW77OWFW6UZWjHqby5NiPrF/N4B0AOKsz
hXq2UaOsZSx5u4m98a2zD0ejQrrvquEApm7NdfguXAmHikVvC+U+q6uULcc5jans
o1bl4POIeYUkHXCcOETdQGUQ6B5dt1f0TihNw5LJ3AnoU4MY/gpULEmwOtKZQCGI
lQ8Ncht1FW16JZbQBvasSJu6u40diDRHm6AQo0rN3BK5NU6q99k2DSE9c8cO9Oov
k0SF+Ap9hAjirSoqfVmIfWTa0nN1sWNftYqdjOYnlor2mpE+Ko1dNSkQuUvHcVGr
JybPNc2WY0GuFBGaQF2oi5CTNMhvBd5TU8vBS9Uhq4GqLoge4rELrO0S1xrZTwTK
0I9BMDFq1lzOGTt9dFe69AestWRKITi+EdyB+eLaWl3KL7VPi6ZL3DnLLO4fe3GP
LeeVE4RKdcHCVMYX/SJyobJWuTvI0P9xX+JHXc0agoJXEsHivDM33MiIltVppjh5
2zDkQVFPbzkmkXkwyh1Xx9D9adwNSg2PDRbCeP3+ZkNzkfLFNq7lfbXB++wJs/+G
5sFdSXSOQGcvlX0xc6WRZq/puCaWpDIFkDbsVpuEbTsVHb2edwjKUlLrEAR9rKt6
9lARM0nuJKhzaTvdEJvkyiCNRTfHlhhBuu0BmxoygrAYe+I+vRMNgs8EaXqbT8Aj
doKuCiq1pvuN/Qr0F2Q53OEv3a7f2w+PXayUhaNpOGRhFhIR5l+LdkoM3IVrsCD0
hNMjHNHw261+Kvocrye5oVOBvq0c/vP9vxkpdyOuS/nztis+1tczNkv93AGoN8Ny
SlCetUg/2tMjco86PNkPKx8Q0ny5aICRdYoMbJYURvZOy4ItEB2egmO5i/lG82g7
eQ+1MoH5LiuoJA8LHNIIwoz4p4l/wWPbEAO5Jk3tjDIpFg+s91Xeh3QK4bCeLOUa
Dxx1rDBp8wIvLEawq06wV6EcrztWlm1fiPKQ9uM2WSC4GNT4E+Un5UTzyLbloxIe
T49kWq80hT79sR4CXKbcZfeE131amqfWAdObrLeGSsb/cccnWwJpw0Ua6awFkqqb
HzSQiFQr39T31W2TwdhqP5psbGLVSq+M3IooMe2Xlu/n0NiHNO2WluvTviHC6+T1
8V+iwAL/vQDvzmRIXWGlUgTOxQDcEUdHdnyAi4ZCfVTWabA5XoXf/B3fWXaAyFYg
DNS4mrlsSIfSLt32FDM8z3OJkz20N+2AGoBg6rse3KKR6k62UCP2VTNfGiI36cbt
Yr4wVYLOHjLLQtrmS1tPq/HZ4gKzyJmUGdwDBlsOtSI05hMvtIZHahxEMn7fU0vX
fX0Y46IS4c4g5KalOxnUSdzYSEd7l1NhUCD6grLiZT7T5VQ2rgPU5Y4HKj/wbbRF
0O4yJhR0Cz5ncBrqdOhmIkN2lRWeltL0hw/9Q6jmFilHV3LPc/Y/0Z93GIsKploz
ZtLJvjEFE0gmZILCgCigulNR1TgOE9Pz1J5I9Jd6uc2Q/XFmEuHs1rDHWLoymD+C
5kRoWuFC7lSMj/4sIgZgvE4uK7EmnShSMbh8xIgNu+5UPmcBrP6AzEBVks9R1Xud
kNmdaWhF7AQKJKL/M09WJWalCVZ429QEeAeOyrfGOAX5euv3f3dQLQMvdXJS5uwv
kqMSchmfx9W9Zq7dCnMN6xb9/DkAAWdCTBmkGRj82F/wRLmwAQg0Ov/9VWLnTb19
7H/H4lbDHP0f3PVc/Sih3dpW8exsBZBCGDzWP5qUCwmVhDuVKTgWP80e67baL3Yr
gdipRsAkb/2pVRVCOMPpWtApJDPh/bgfmp09qkAv75SdG96c+k4QME+zA/efVpni
pjRfXBmGRh+i20DzgmVcsJ7eqfXLFGm8BtCzo24aNTjmv3yQkc1/v6vY0Iqhuw9h
iXQ39b7mxpd82lItYMCmkc243tv4r0y2uPAJBJ0U1HwNMnmGfNhlVjZoCnQVyQHv
WgbPWdk+omOHDa93HVHVf893mX3u8FZRPK3nYYEszXM0t80m3ro+uxkTUPlf1gHg
r1SxdOoMrSgZQeczfEyzNsvSxKaHTz5AxIAXvg4U+0jXasO207n9mA6WAnrQzppd
SnOlYP4VLrhZBBCMU6awzVd8Q2y6NRUvytsw8O9J8BIfbUVb/ibY+QaQcKgkvSIa
7cLe6H423PULAUc2uz1v27WYXZ9Qf9xOgCL/ccnhxpgMfeHRaTAO8bf8TtrzYxdk
wuS5c03r84YaRmXJ8fJh8xTAbqUKmRXs3Kc0F9njDxWGGnNI8SJa/05mg9qlq8fk
kZU/u3+SybbYUTARrL2k4eK3Q5Ab84cUr53F20eBTDZReMSagXr5/vVHQi5/M8Iw
Lk0bvXZGsEprGzlInzzwhnuZyjDWBnd8/hAHQ29KWgMTAQF16FeZVoBoJ2J4Msw9
lAsK7vZvy0jwTeAigXkkooTm0QgxkXbIvVtxZLGRSyiVNlIU8YbO20CNFl7i6JWY
u7SlpZuCiB/RCcxbBDUK3mesZlXX9tf6kJVD4g7qHyT0RD3S1fHHDIygGimtt5Sb
BqlLTNw1jf1y3AO/mUsn6FhP9rNow6mqrxs3cD2RENVQSVxcKYJS+yhRdDhaLC7W
Dn8ut3KmZH5m82g30hZROKyc2K1Gro8LlBDBc5qQRAiV8zZ6GbbaYh6abE6y2Ms9
Jq/kyQUeSeI1V2X27gmm48F2FyygO/J6U8jzCuZBrywSju0fmGLtyDQbFFnlmvge
FkA6sEF0yGZBpm1/0/BYNChcr1OA3q59LxYdbn3p1W1kh5/lal4YYbF7out2DZcB
VEpan0vxn7VDo7efn2y9sRVXv7Kwbm+H70AKaGoQTiwM7/k+2X0GTqoCHN+PyBsU
JUCcNV6gZwywODQmVVMbGQuLf8PQXgS4yzJtzZtmyKQT4X1YoZVruQSIMw1OHlzt
U3yqWqJP5TGAljNeOdFT6xppasqZLU6Blm8cbDZ2p9Rl3H3Qtcfl+bfd/HvCVWEm
BdjJ8Rnlzd8uKFCrsZ8+vbf2OFJxOqaOowVqf3shFeJCB9B/K+46sEfBvl7/LYMH
fNQXYoV4JWKf6QXMsKYT4PAkywYWtXhV9vqBvdXOpVO8md42y9AA1GHlTchWdxK/
CLZzDd7FrLPzZKx4RgIA1QvsMUvDSbcTlp69baNmI1hd1NfmqOdZBvaexxVmmFoA
sOhhMJaNHLmpLuP/NPlBALt1bakdeBxXERZwxwlsYISSuTq9JeewbSSqiXRCcYJS
HMa11HsRsWuf4+XDlU+Wj0A8t2LPKPOwmw1DKJ3nKsasPagI/gYPU7fBP7+htVro
ypJLQgKafeMftngjQInRETLFAPpjnatOEPZPkNhqdoBpJlADTNyAzJu1W/Xkt8r1
UUmCdThBspyIrmYHBQLAgD6B/HMTgwPrsDUPTZZRyjOoyPtNQzHQzlOzw+ZV3lwd
RTKNa/M6u+aLqnTLaH3gyVmbO9BbRvLv+KHHmBBl4pJY8ceYT6SpylB/jSYt9NNk
Bv+tDaDFsJ6LUNIyp8Lo0OJf/BQKGLywxHLSL6P4yg9EskQaDhmAQYdXq1KjAaVf
inI5U7+15VP4u66SyhrcGFNcLQlWN9Y5jkGKKmqxzuNRMXKcpatBhzbgTPZWn25x
4ijVaV6c0bWIXmTH6DQS6PKVeHTsNe5hyTP87YW9Fa/IxyLqht8UIKAkc7iNGrl6
F3SvrakqweHv1x21XDuC3wwRJgLtU/jhRCRFZRuHiTsu++vsrU5zh+rANPxgcqjh
MZwmwwP2MBzTaJhU0l/eVhg2Yyg3BIV6tOsCuKz5RGMQGON4Dg9oFd+DUeyXY/8G
WSfGbPTPA3JC0MuGPscCKlz5anwkaqGjLUQFUcaGxSwwMINah5ROOP46ccwkjqmG
AikoYvLa5AEOFgbKqfk8PXfaRIV/OcWy79MF/1zOsqYjepAfogNlYHHBf2ogNd8B
muE/jUC1MYpVk0I43f1lIKR56PHnnRoLbl84CLjyLAAFXi5BrzpDlN+2x/hcfGU7
xQ9Zh8XUaTXQ5zH1M9tglqYP+OdoqKFa8LZCKTrmZZqJF1HmiiWR4rPSu7HRhyv7
wggb7Y1dlv1eOlbka7dJuoRW3FyREbJJVL8TjOXm2/NYRbM6OvUjD4nQ4Vh9VD2h
S3PxVTOWy6MRQZcQDOVUKbAiNivhqKRJRftYGMe6pHLVOXgErVBEmSSxl9Fxksj7
/TnsByP8LeT3rsePruLKsIfTq6ln3f3oJvA7e2hqgymXSBdOsXODHWGL1RMRJQVm
HMzptC5x4uZU3vbOgEU8QWSOHrmDk/ypHwy5OLOWjpIsCkFeQLXpmeq2w1lyAxid
MPpXTfukkOvjj7CZoIwSLs0gy9T7894pPgxpDGLiifI1Ac1/cnpx76ORBonsVH+b
isSe70f2tqyqQ0UHYEgVC+5ctlvGqIc4jn7CTAixTVgkPp24Z76lnb5iy1VYQSGh
wzpVD0ZOeuKPYkWaJNoHW7KY5kkjgLKG+C4Rz5iEJVD2qCnD0n48Tjx+GQxuPAot
U2dV9289LvEhGtkthDLICQlKYngMxQWMeuSJp/QICTDZ0k5gFaxPAEWerWHkrzYV
MLx0BJfZ2cujStrFGL6FhpP/pc36cWLfS+Cb4aEWHLY2EBCashOn3lFxySCNTBWK
M7rI1uRHKsfyb3otxFyyBavY7MZZQl+tVe0YlPlekfhrX9aeFwRVFNF+wcqsjg/U
iPlq3Px7TGnnGrsoBXb9Htn+VUXnikymnFbvM5644iDOxG5jn/KjGxFdqw/QAwQ1
59HwYATdV4WfVbtO91ROFk4RpQQAfyNYYOGvGwv9gX4GReuIIKAlLZIrhgoFGrwU
hNTo5hvcrFHQiofsWRjJ3n+0PcpUK3pdjwy/1a7c0uwRjRl5CaTG+9E3xrbGrFXS
+XojpxKCBqyxrJM2HSX7eSJPz1ByQm5XhkrzWtTY23HInlyc306GaK+DbZwmK6O5
I9gKE6rpvWdptX9lUri8LjwbB5nhRVWUK6G/jpIe3wfr/ptIBqC2EjzbRhUukYUS
zKIgaEVJb4g6ODNMmIgx3IJ1cKm8e5bvmoZ5bw4IpTK/WgbDzpUeAFaMR+O1v27T
FvIw+t8xo8mu/8OIL93dwAq0+mR33L8x2B4yU7GyEwOXuv9D7XvaeNaulox7Y+UT
kpWLQ3iPHLRniZc7QzYwx+uzA6umHI+oHb55mVjzC4jrf9SKJLqDhWR1M8DaDlDM
PK7lRYQYDSRUgwCuAWJAYzQazJAlLHXmMyIax2lTGkZ5w31v11Er8Bx6gs7hPvf5
3tTIpXXyjYKDgTRZsFBsVpIS0BTO4i+iEJmxY6f+Yl5K1iDgGs0OXghreCnrnAO/
rIUpV9b1Xv2mEwfPXGvBlWjMoV1hAGnbDaIQEVbEtXN6eITGh/uPBUT6Wluof/+V
M3KRPRMB9QigA+PFJxn6diMcxQXWa+apOOm+aLi0vIBEA0GxzCbmKfJKowUdMppN
rcSYMso6/FgE+eVPISx/1w6VAuKH47ccRA87K01kuJiIPODlR9lahsAQ3e/wal+7
HSGO7pAPUmAv2lM2dbIDFlilUPdYJPNB4yhOn8gYGYOeo7Nw6LX5OhJd6JNxzz8p
W2G72MTaooxGhT6sD904SaPAOp53MDpsjAgEiQdceFAnmgTtuc3n/+SBupfIEmKt
EOJgrs7y8Np8NB/YloXmO0bDq+UTRVE62N5Nnku94WxAgwQt7o7wtYbcpIi0Xfae
NQqvMpX0Xzpff/ZevVjwlWDF9W5bceAPRTsD5zpR8vsvGfpM87qFDnNAHe9vrOmY
Xpn0nTfuIuTrvaljVS3tCUBbCEPVfKM8LzJuQ1mYAByN6pSDfxjrBNWS3DpiLLJY
q3Ig4GZ9GCPVCU+s7dNX/w2PqATUUNri9yiVe/OMpslZf8oRHR2c6pWCDWMJpFcd
hJOV7fyAHlMz8iPnfGda49RkCWHMebIcxqSfR98oM93gsF0msbXzcFKth5fRyvbk
rzR9DHRNfkaVJs04rWnkgfFIQC8ANP1OtZFvja6BR89niuwNsocpEPESzkxZtNr8
3ufq626QJ3fayczwIIRN9rYrxS1gSguf5VBIeTuix3nysgC9bBuTk8dSf8JxU0I5
mctvjVbUVIJmPAWpE5uFQBtHnd/OpUrZQB7ouX93prW0ACKjWLLLEROX05gWVEpb
rAf7Df0fymr2QuPMcjxGKP+EC+0WGpWjeGEAxw0EZEqEWlvGN4V7Bsz5B+hYvw9T
I9/+bLWQHQJEUQ3B7+q63lfk7GO6hryqJp0BRt+jSjvaFzel4XaABDQXOktFDp9j
IHF08+vlZ6YLYuN2MIsxVHYSfNH3pxgV2LjNa5klRTwrNcFD7ttHmb5owSwHD9gK
SlJIjWxpiSTw/oSgzxwMH9sXpNiqXxzZnG7ixEvNvKdj1kpN19SIa1Y2hKSCD7Uh
ZDWSDIGSNawrSNxVFdCLWCcG39NKu0/T22XChUh4fPgivoWCX2Z+GJCERYcfbGgn
uITcnHFprD6p1RzQ2ECMGiZ0sut7vWJAQHZZBSnWolmgTZOEPIJOhwAmT1z8I8g1
1Snk7F6DHs2soesE6gKn6vMkR05r+HsahTC+ItwknAIkYexg7uSPIJGAT7wZLNZw
jeoeuee3aON/FkLQxXXSavBA7p+AQJMKkLw0Kd04xROT+nu4gLEbFmsgqB9ioL3a
YFr7/7+rY00N2Ytluo5lKGLdx1fYMsyYcsmk5pjOH2yRmeXxTQYQqXihkI9Gld/r
l18BOqLK+ELqloOfonN8KCl2vni0exXMwaLH/Anic8It9ZumzR/8kybgs+2MDiNH
W4xCHQNyZ0sziYMD7krumS2HyvKW1RuL7dbt2/l+RpBeZEWLgofXl9EjZ7WKfawt
0hSRnuIzzSsjuV0I7qEsnr1krDAHhSf718+KVvHBbmCBSQSu3os8SgBRz9NG1wf4
1JBJOW96G7uiJcuZz0Zsbf56hjK92Qly83BDIUSzCQ3rr7DWGLe8lcUjuLWNOqBA
pL3Foze/3JI2rPopT1wk0SY2F1UgiccKGpOCsFrxlbwGVSCQuHSjUR6P7PkSSaMX
DYDco1D1WN2gXbX73pFqsY03D/XBQt57+rPXY9nWANy8pav4T4W1SyMtaTH3oZTh
AK8/WueRiDp/NBzAat1YT/CYjntAlgGzVg1Fs93d9GT2RcDontR737xJl+tkZC7E
D0RIgfoythBAExQ7eIYq6DRR7xCEwSwus3RYzv+b+1Oo9ov2zprG1LwAroRs+Wkv
Yz2a1Eeb7g4Y+54iUkWnDt9s4Tz7Vlqt5+e6zHw7e1pCevLXTe9k6dvkhhnWYp4N
LRJnYhK9ozSixu3Rz/vg2zpZeURIwbDzKinNXqaFAVsZhhYwvwMVlZNYTOqQ0U6u
CEOTxPYMIlndocKT6YjIX753xt2An1fYGx3osZZ6ZgpZNEiGFJOA3v3YN2opyaXs
9WHhGtsA4n1U4yanCQPxSIrc+oURujx/HI4hOQ1GVkAsPdW7Rsgx98e62Qtbc7Mo
9UzYRuDiNMLxK4fmi60CTTMlCDRcjbHeH6oescXvXP6nDwHXlht7bY0teh6fR1SQ
3NwmGhFgn/PvQVLFD0U/+FGh4UhetQmZcSYU8ITei0nS+X/Z/77G7feRJgddwQrx
cgIMzsO0ZZDIy3qJrt4k7TGUtPZn7pT9MAnrR+1+/TSdcDHzMoCpKk2WBiRmrMwX
vMQ4KtyLeNtTRkFe0FigiF5wlvIkCqKuc8370TEfkn/6D0Ph1ui1weNcKSt1eJIW
wIrIZmYsHGM1vlfijFLG+5viiGaVKCJHFVJq8IpXD0FwH8yUvqLkyAUPKGB2xHy/
VqVabjtZIz8CXU1F6szN/CvPa+kCnJgxCHXjbK9B2IwM49CqJD9SnrYfimiKeBtL
POUeGSYFZWk7BS5oLGdWwvHaajd/M5w7wdImezUNIrWyjCneZk7iEI/Viqa6ykQK
o1IX7DMQ2fYt9PDEkRW16ZjQM3EFsin7s+M02iA6LWlC8kgZx1Nqose+bX1WwpPp
omCsxSDLmjyw+hT0GFBISzR25dCSy5m/ZDSDT3OkO5dCSnPTWVYs9hiuqD1Z8/EP
TP1cq8M/LFVxQn5jR+xIgd6uc71oI9JWb7b6YGv8vtNTwad3zphhz9BjzcStOsXP
+wQeG/1cU5gZuIfkg8K4qdLVMZVuOgP1/EOF+0UtjlTClG5bG+/wZBFhb4oKggRI
/FiKOFZPAsNBDYYG+To9861JyiEsFymM928CI+DSCVhr/ObVEbBtiHXWCNShGp6m
syhJWDZkQG8jD2x/8VvhzFAFsghaoH2G0kakQiCm2bfBVAooZCkZeHSMbO/SGnWm
F4HMk0Egu8UAoD4TUZYj3A+5sHSXwe7QTWFFtOF9mztkoYwM5a/H9tX80vTTSK7p
EARLRPhn+93vwCmymioKJlO5/rMu+o487p8HhRajwabOWIVrprwv+rIPw+RcD/o7
YKqC8hrhIYYVLlv4afUk1Bm7PzwXlYyUA0NU5DYAGSyWxJCjzKwievgcQYM4WAm0
cr/Gn2YI406s/wCkN4+Y1F/+M18pN5R3RPBkhXZQfkh213tIzROhH/CJxz/GEDCE
ey3A4yNO5V/xMDMovqnY8+E95TwQfR/GCMuRq9IqNPxiDPGFCBDCTClXfXuoPhvy
igJtjolJaeokCHUK+B/PhNHEAH1trzpsjdYaZFW1p6jnVd+Ve+TCIPWOvl/raCTH
dgAsh+Ui6J76pV0f8eOg+X3PjC+XZKoSJ8NfqBVsu9IM+kn7QAimi/bHk3a7NR4a
lhG00is35+AzXNz+tW39W8LipxZruNu7YLr6z0QEFxRRM5OKTOPUqa7F2hnZupfc
Ny98BD7luvFfquk7eIkwO92yqfORp/755YcLu7fACuwlSW82LAZFEraooGjtxb4m
vK2QkT5cTjmGSldQga7RHoqfzOtzVUGCh5uLPiZqAi3F2KmzKuwaDfsMrRp//MET
20WawnLb8gqUkMgjraXY1+jOXRpBWSYtxiXY7gxk2aBjmr1eOP1jgGDodczOUkD3
teigm3rxKZjGqghuFQtPtBxXGXSF7XmI8u3oalgbgE28xWolOFDt2LMqfwNJ6XOd
CloaVp4qniM+Usxk6NcLPGCSaJ3Q28ks9wxKWfyx2f3olFtMbUQX8Wq1j+f2wFZi
Qx8pKJHtU/Jt1dZYMXZ4ad4xaqQLDNGkvV7q5vZzcyumxa31BvHNB8saIsFFCADf
9Nq6fF+E8KuYgqM2qTJ/zfB4dHesY9aPFr4rI0e8QCDZxwlU7P+cRMMQcN05uAjG
HM6fmtrlXXQcbAWkwHAvmsD31r+znTZzpZ4nUSuzzI6HJDyqrtWOmWscZhuBt2ZQ
syz3pUiPTQQiqydsAPY89kZQeNBCsKc47HERni1/xKWkB+gQKm//DlTlCCiomumy
GQVS9E84OTkuJE01kc9pq940N0VOX3wFhtcFT8Av4ykp8Yf/r+Wirz4C7knz+Ery
98ry2KfA0ml5FjJUpduvl915TX+3rap6FZiMz9Cw27MF6FgAXudewCMj6vr52msO
E1b2wNxuyfDBw3AtsG4y/LASEto9KR79iN/oSwc+Qrl6800Hc/Q3wdMm7MzoLrSg
64Ek1dfziS00qpXgZOVuvcq/akJ3yteuCVz6O1zT+lm8/2a6xKlTGcVnE6sq/npz
DBocxFcgTL4ONbznaTMnQJ+e8+oG1d2wA8hKPA1cC93CZmIAIAXHwovgiHP2kq9a
004TyAYvc+Ne/mLQ092dsHEzwaGd81ioZcXsc68xp6Idppo2U6UU6h4cFN3G+5BP
pdS/EoSrGHA6f9tqi+IgwAwzQmixy5muFskXpS6iOzS3rZ1WDxt+L7WPscTbi4Ym
wFnfMLoMgYvDUGqxaMf4IarDd6S+vVLIs22CWJb1FZggS9E7ch3w2cKp00ch1dQd
v7naaQvWfT+AA1CWzgMKce65R1MeL5or3NPSuvt6yGdU54DRxRZtJPRerTzR2tOS
0gdv90q5AwlqDcid+oo0P/YT0RjrP5twB4JKGwYJWOqNa3sBiEa8TuR0JaHDX3BY
HwkT/BbvevkMvwK1b8IdP3XhYHrgerMfHs5Y77EoUItrEJVRfL+/LVD7U6FCmJ0q
P0K6fIvmkn0C1mWz7IlEfzDLYiEkw01KvBWF1GdS8VjdqIEJ+LWQ1OIu2H0EtgJz
piGMAC7Y80RefXHwm58D2YcQWMkCjaquXXRj2VUmxVkSVm/JJsnFatc4EyhNdnyU
SOVOWGAYbC4A11mHStGc1zPpmuBTR8Gitdw0rKYLydLjTVEtU6VzBK8EKvPlDtH2
s07A4vA/PdezAkLV6XskzxlEud/rvGxpjQnkGaL2gzrgEkeTjHot1l8bHo6xifpQ
sWeMP/ApOLo81PPStPc83Or75sV1Y4P1lnyi07YsynODcov7ILwOckUJZtn8/v0Y
BeppH7PpnJBTE/g7H+k1ynNbiuFkE6TxabMhrn0N72si7sG3wcBOt0eNhIUrPybV
OrW4Xlj+Tg0iSkvFlz76XDigpPGoVfWI0zmBFMLVIxGr7baxC/8ZyRr90ayFbzWD
Fg6SwMHPSU8SJYb1X8UCv5xCVhgezQdXJwlZ5nx3QJjpfKcOxCJOH7Lcw2IYLEiy
WkYzKj50edlIzJ3jetQSFg2pmm+IF34Ir3Cgo2VqnnbSp1pJfS0WZRdhfdNyTE8k
Iev0Y5aSP5yS5ZFasfz8M4CpvRd8OwvBC86ZfKAmvq/lYW99+sIwhoSkxKZHpUDp
BBmdOlC9cVZoGU9cvZrWTjLyIBlkI6ThXlz8qAb+I4h/9+n/SGLirbT9wKnK89Iw
gJvcTasUjZZWlvRVu1+gfLL8NXYc72a/6eToA5aCv+FnfZpMJK5AO7yhCcmG1Crj
JeslvIBIFobFRBA7h3y88BNVcpr+n8qHB+k5AH6ouxqStI4w8d9h/LD+fp3V6MM+
GQhGUzhuxo1IRrLE7oG3VC7iIb44NgbRbCA75SWdZNIpiiYqxM4+H2KmcE9H3KRV
jFOsTRPCy6KRvjMVv/Vlh7AduXLy+B0q/2exsXDQ53EfyU2slcGVpuKVcqoUD9e0
+h6AyClmpGDofn99l0q2M4TA18u+gwbYpP5VcQlcWfRQDO0ZpDbt4E6QgBXapakz
jIxhViRHbdPFxLm9e0pYmSYj0u2Z9F6bfhblC7Buauv0II/QeIkKTiPr5FbUOnge
pPWR6nN9yPb9Ek/JFSd3Z3g577+rjBDO56BEckWC6FqzQ0B1dRES13gijeGU0k0u
uDBN/RQkP5jfxKNU+uiGKODKfOpp1pkqojW2Hm2M1SpWYuCBacg6dbvTTilYM2H7
MDNPvx36jEJwEyrqCQiy+93Y3WkSnuo23yaSqFH4ezXNXWyx27OlEpz/c/U3kZj2
d5rH2vBdffWzjYuLsNmPggS5waxIEa9bP1ANvo+K9lBYjFpNBwkKES9dPPdG12EK
ht0v6QVl3Gf75k3Pcp7QZzIhGQbT0rSUrvDvtuGgECJBvfaANI4GAtlF7scOHlzw
hZxBPLEP3iR3a9faFr8s/ksgRvL3/3Mz9bGxnP7VZXDT04fYz+yfousBf2NL71OE
xUjQA0pZtRmzciA+pQMf1slofTHI1YdVN9cHFI3h5eaDrKvO2xzUgQIR5vLq591q
A3WHKwhVyH16iWrt37i1zu1BydG3OFLAgoS6Z2rW4zAUC5GSpiKf/Gft5q9pA8iY
0p5FYZ0Ds5xOenHDwl+Kzt0XfaunPdTny611PibsVnOAapuQlaPCu3JwILuKyaEr
xhoVQ3GmqGrtHiTP+i7yLpzyPGuEu+b1uXw7x/4aQHpINOUIAhVrP+VsLNZsIxuj
AECeZQJzHYCyfMmJEne7JWNUArzvlGylss1DP24zoaIS3pl9LwImvnQ0iIni5kW1
WWDU5mwATWqodhWwbSOHLkVOB16gFBrwJHlafcf08dmS0OupvXYhSY1KAJPJs8IR
Mw31XgNaQwWshjm1gIwpI7wIWmG/EQssPe+/KnQc1nXm/3qB7tSQseI1MB0Mi1qy
uTiqPOeZGQ7MG4MWK9qEr0rbHeAGLkTlar47MTznPvd51SXFc8YDJhgEWRxMGIGh
2EWbr2o3p1OOzqsryL1a1Jlp9rawk2MLMxa4xoq0k+Mg5b4MS2rUse46wRdkIBHw
6BnooJVT3c9bXp3f2LUPfkPhKEsPIy9Lw35Uru7Y/W9q/+VeD+zXS9uR0a1emavG
8UiKxibG9M1BIB0n04jVCGJ3p9N2npX4QT1pwhyfTCtNJVTY3Iv6VNJRTbwZQMg5
XF81/3q7WU8akKwGka3fScEeq0oUvMXoWUyaZ8iuOUpOvDPOcx9iFgMIGj4f7F1z
CsfUoOHpdcwM+weoG2QB+Q1AKGg5aq8dOCjRaEpeVfwM4wVXxrrSggM6S2bKhN7w
z7s1WH1i4Hlz/biLIE9/SXaHONNRlCn/xC9D2YHGDXBhg7XqHlxmW9TjMlfjpYZi
HqQXf7dgxyQs5DlvqaftrEXsKhBaJuWL+4u2Ls1bmBFCxKXI09a/tbAkgugOUKfY
RD3JiVpbiBvPoRx4P0Xzu4SarwrUg5bTyYjdJhmeCh/6NToXHPeDqWdPgZKaDvbb
kVL28nd/wMreDipyw9JB/sTOk4Uy5q3/zYz1kQt4ZaXDtYWHV3SLVhHiA/NGpTty
kWjFrl8BHqM8/WCcwPJCIA==
`pragma protect end_protected
