// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
E+2L4mhpK5HMsRFnlp9BuLOwss++Zdg0lNHnTzJ6snB1pdOKdL8crsNGHfpTMMYNrlGHzMccU7MK
xr7T+8Lvpj0FQ09zY2H1OaTgDQgVvmpg9qeTaiCxE+kA+q7pDtQpHGUm5q60MiBEYWHjaa3YBQbI
pCCJEN+9jSfXXW8xAVaW5Tacqv/dhS+8aAIa9bBo6AbCTn9vpEJwRLGRSgk9mboWFx0kl1VjQDzW
5ulWFvp4PUwwTcLcM4jVWZOp6KZVtmL9gNS/imuEycFVbOys5y5kQFZfUefQa0YrmmZePYHy+B8k
qwFm8kat7/cwS4yBaLjOWA1JDNnhG1LwCJ5hYA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 18096)
mvIKtS2CBY6YMeSAqYRXOcLJn+DytcEgUdeiFMhQV+MNHRb4YBiIQjRo79BKGVQ5O4kWtzaT37X/
JJ4NU6JZipu8ch7CDJ4cHLJQTq0xoQYLqD9+5LE+McL/sI47yOPrpU71z0Shfyv/oUvIS2SAaBQT
OdHJwGdsDFbEToYLsGEnIHbOH28Po9bIYejnR1ot9rmgA8HF3LwVPd2wFXdPTkpfE01SWCx3JMp+
ONkR9CChk3YlFS9mvgHy1L8y4kZr8083uksQYevH7klonTEF4z08UGAYgctG09wjVmHF61RIYj6J
Qi0NDIgQL89LTPNIIzA/E++puYbM68c/bpO3abmMGi/LWbSoFStomItO84JDpoIYgcsoaXNhCPb9
ezP71798xAw9JXOVeLaGFI+JVGYqjyYxG826ivLRrQY4S2WFNYlDoYiwOw1aF+oqJFTqdgA8pDML
fcI2+8MLD4crEgoQ6qgwyNy5qAeaDeNobeRGphCj8A7vGDwIV6Z1gmHItJHAB6PjcdNBY3WhX7dC
GLBXgyhTiX4fpi4iPJ3dPzqvz0OC0w119fdp5odA5pXLXRs5Pbz+GmhieZFKgUcrr71TyyZXjL37
48ZjQA3F12fwEOuCPLdTiRw17zk5zrAbRTWJYR4t4ipchqAbG1AYnkTEOmmPkR72gz52e7RhXxA3
pzhyfmCzokOx7AWvxsksKRMMJ9DLRPVrc0VIYBejar7/VMVt7QXXWDJNlT1MGewbGAdXO3Hdas98
6ov3VGgVtDCNjZACn0/7AqBUDWvtlAOgPZJjCIaZ16JA49fpdygMNuJ2lQSiv8CGt0ImjtSioXQF
LfVx2a+vzNSGRFlap36HrSjbod7mfGTGDmaB2Fx1rlZoreL81KluBfx0Amf9dJ2qA20rEgeOi2rh
PQzyCnf2CWQlba+OfeUGKFr/tyZLRtzC8MGYIz4D0KKLJaIj4y7TUIzucI4MZD1GRTu97IyeliJb
YC3s1noTIkRZiGKbmiL9OrvyTr0MWbhewxyzGxpmWrKDPC4QU6eozFrtZe9nl65a0FWAMySaVrWi
80bhuxld9RumzTSPRbPFYepiNMDu+dPwVgDkDSNtIeghOnatGdEQdx+xsfJUUUHUV18FYqZDk2da
YaORA8tKqHzeT5721OJU1TIxPIh4NZwOsbCO3pc3/SBVZWwi+d+YKEknS1Ou+h8/mS+B9YnEp5H7
ZzqcYijJRKZbXdqUSGZ1Egpel4C6COU9CL9kUKU6r7W7qKT38kpZ0bxj9kIleevdRV9sMYJOHiys
VH720DvawLvpwIKp1iX+mC+doIvMmNYvIVNSuttHjVnTED2LU+27ba7nJi1qVoEGHFy11W9xPm1p
Rc/5bhPIysMnNhHIs8043UAr+VFh1Glp/K6vFBXUortJRg03hgEc5HUOFBUlKmspkxT3ZsYCiaOV
ItR96UB5b2+fXZMG8ZY/uM518VjUullwb5yf/Ioe7vCjn2MWWUjw9D0Zq5UWtYQTwuGWBlF53Qn/
PeHdOXZrTnpWptFqkqHSo1D4gfKA5HCMMtFOTs+a9MLijGCPjWoUu6t3b2jZsEfA2VOIYm8bn3+X
uw/U84bphvmsdwRvmY9EeRqvZPBmKjBL8Dc0BLnDCI6S9wYxZJFjrP2kuVt5j33Ta0Vc4vzQkwNH
j5FmH+VWGPzrCPJ7CbuhjIMUUaKiY9OQbVobVl+3xYfAaV7mDnpE69PVbMASvD3/Z0633wzTzuy3
3ZSuOPy93sWGSFwq3MQZO9v8Ol/8eN3HaAsp2OwSZ/Rz9jcLI0LNtcKuU/mOs0pNrLpo+HJcJ6GZ
IKP2uY9N4vaWnVM2wt5fWtikcNcvLWofHaK9dQVYaDSfxC0HPodDi3XRBvfMR63Mcd42ngyBxeZd
6qnzTBRkXGJwWvVmm3HEmEQIbI2UrhtH3UL7kV33n6PnZ3dndoE5/ugsXsWPf2srff9mDiU9YiNH
qJIIfHxbM+n3sPos3p9F3/i7Dpo6k0mCDKEzPlFW1BQMPLtWjP4GYeEvq4TA+SSQgYj0eT/xS6IR
wfP24mAI8ZM3MqZa5Chd3nD/MSjcVYM09NyJQ1B+RVlj2YPDhB4Wwl91TfeEfVN0AMPJFpXcskYc
ewze+cj1F5nI1AIWf7FWT+BNwMI4D392eixAIrQnrSA7rV/LeT0e7hhQVLgoZHWE8F2Dr/Gn0eFh
A2s8J0ccmbdf645xwfOQojssrdcF3MKDcIsy5AM8zwBJ9qHbRZK0Ndo/DyMCLC24nsGeFgcsn4Rd
3xRNybpPpM2ztGXC5D8J+QpOoblo7eoOiI/JIo2lGHfUqxEoA1dtnyzHJEMJ56cndx9F2D3vq9DT
E9FesWwi7QvKprRbM08jqYUwSK9FQ86Km39OITpyTxGH9mhjikSz/ul/X2LyJobgPIh5lmrY9dTU
PHuB2A6xGmsX2KTz19i15/uQ5ZHp4tWnolL5hnNHk6nhSkUaq/RJ1MzdQ8+sUBotSH0QnsbpFOxF
eEd7kh2Gz7n2hsWJ+qpt0jD0bwchYap1yRx8BGq542sWDkgUg7EZmUuPPhDOw6hM+HCQ3Ee0ZBpV
ghB4x89hjq4qpSjjfy7+QH8nOYApQIxM936OfIYTDRFmZCjQkR40apQmJF1ZmMDIAbGpw4N7lTKY
2Yrx37myEHd1+LIih0m9vvmD976gT4Iw90EkDCmH3VTGy2ygdg6/rDUZpzN1zaid3fOMeAVvFSen
tsmK0XNu5hfCr8L2A/kGlTecEOuLJBd050+3Mejt16upXQZJ9mdnMYPuFMj23iuq995nR4cGlbsv
SsJlLkgE9+6nL5cIPyWWA6H6Zvvo5LgIgsAepyEcYISjdOJ9TowPcIbOdso76rvDItNz80FJD4Tz
kwhYtkv3Ih3OnayBK1v7tSV8E0Vwo4pqcRW8eNJSofjCmSM8IFDeI5AUBC7UGvsWJz0I/+YkAIwi
J9942fBS/kF49X+XlFKZ6181PRK0csBpEN/PsmWZMMkoyfXwKIPPCLCRH/fpT7TlYzGIZJI97tka
NUp4kOPic3ZRX7jhwZFTAMy8xm129NJgZq/EfueeZX583HH0NWpfKclLFS6QxO0e/CsKBZ/G4HAe
OUfrgVwq6XzvHeMo5f88rz3O2p4zIoXk6W4FAJZa/Xt5izf8lJEZN31j8DSy9rmNE+yj/1GJ4HT/
tk4mXmsfSJgQMNjR/yRWC5FtNbvPmmyM6XnIH3il3TWHiE+hw9C6ORwb3eD3dtmrg2gdFQWFxsa4
GOOMsjv+bYK/lC0hQEYF4oE86AQBWypC52VbloWc7KPME5E1HEDb6w5fNM9u6pGeGup7vaRJgkbh
Iy9Wy/9S7bH4v5pUCCpsSsr3y7UY3GjfNEUWkCn9e9K8XgY951SV4cxxrO8X8GvkQimSBMR1fPc8
tLwoHHXZBsSYEn9QgY5ItCwOlhJaUjq51dmceGxtuYrdzpNX8z7jCdpN/YefL6Tb0fPa84wHZGcV
zyMn0wLYBnCo6D0CpC0+5N8ESljP4GDFuOcJL1PwCK2/Fc4UinA/MaRxUY5W0uZi7IU/DxXW2GJA
iYRj2U0hQcEFNm7qly+qIzsEW8IxPLZazfdysbGkgpk/W+YsTKgF84ZFHKdhQf9YD8k3vmx5SRHk
G42CI/gi0Z9X4AWiiWen/+pYa6IOgMNBHGVDjuwDv+kwCB6qd7D2g+mi8xwAknKQnbVvplU0IBKJ
Vj+dPkoENzTn2RZiUYCbQI9wsGgPWEWmmm+U8eGnFeODz30luTsn99JHaWFPVgh2ZIAuLo/BYIK4
VoqJND0hnHJsFe3P+yC1pLSR7FR+Njt41fRa7Wfs36iBty64ywOiA/cvKcedDQmhMej08w2+kpxn
agkTTVkCDMCV0VtPNqV847IZJfp3+FRAM3yOqc+X3BPtYNLsfgNqbKGq+czl0Bk4BMGv/0AnDn1V
fUkE+NfYqqtsjmRGH4xlvBylkaWapqoiNmZpd5W6tU1rXR9k+kC2EPpkE7ay6PKdHvRyqPAV9XTw
EBDdcYuCXN070Gh99kwdwbmjTTS9I8lYZX5xtD+9CKm3lae0BGJFiAPRnqXhk2bbZ9wor69cPOOg
KlSqK/SDwP62a5azel/5rjn0bXOToR6Q4LzmFX9I8RnT7Foz6ijFPwJD6Ysf3Srb/HTMCn/T8gFI
ppZWtasjmkCXPFHPnUVZPle975rblpIldp5mwNuBmeFZT3fVah4Mh9LaK/QuGNlJzUaBXOet/ena
s18iaSaldeClslFXt4CLRchbtGuT9ecpHZSHeAVPGDZrxO/pdn7MYUu0TBhxIUbUuHSP+tqVikqD
M/69K1zCxRpBomqP7tMDVfIr9a6iEqbVV2RHHo5SAFtCW3M/LLnCf41j7R2AKm1vGerGCE+BDsEo
VBJhO+41PVB9Wx7KLJ5tBpHEX9inTS0WI1bPgzrFgFVycDsqHTTZuCeRHxR4ZWPV7eVG03Inc5Cd
ek5YXETfDUIdEtLxAziN1p0E8hsQpdaCV0bFCBPKCIEZOMln/e9IkcssWnEnCluMN1g75FSScsSl
lFvQHl63J72yNfrZ+6giPCrg412SdT0IuzqbpInfAC+kw8qh/ynwZLQahEDkpdsNrx4GkobEZYUb
MY/lmDH5Lbc98mEwPLoQz63lrPc3KVfZDoQyuQ+lh2FPiiddCtXB0EutU4L4esy5QSmaxxqpBqoh
8R+BBDJrYQJIRt6Y6HS/cylvGwWQogGvnMZbkqNuCuBBkh8r977VmcqhzAOVbJSqej7kPn6KNEA6
u3PzMHbxtERCIigN37tV4+LXucj9dw5NWhJiifU/dS+FIeodPPThxJZuxR3RZ4Zm+Up5t7N5D7WO
OskA1YbXSilPVHBmdnsCUHZ2Yc4slRlDuz8nql0lg6H+DzrafRaymFF3E03iNR3AHb54l3L3+Btm
UtWKeDuhrz8fUruoKvjl/aqqENNKL4bEmpQVAZhsE6eug9FoUD10MhSrm+QPvWegpEnq3A3c4Xto
ASDyOvuSVmD/QparY7Te7G0Q9ZDlHWmWycsKDWaDWM3MghH74HtC/cWlbCswISdS79GFTFBSM2bF
qu/af5J9B1tA6UriDVizK5bCELUNt6QB6eQDbrM0FPqTlQ6SHNo1TIhtKHREb1m/2lEg9NjPk6V9
5JRvY3buS3kmfNS4f+at6nCXtVwRhYzBcdedGE+0It1TYyz0C69qM45K0APrpCK4PzWT6h3TtMGf
wNfP1prSIT/Z/zgNs0SJteuSr/XMv+0ttonk5ExHpSUgVyCcTNFUp72XC6W5EfOO1srEHXaAWTGc
I2KGDa3T3HUnIYYn9Pqyf+4Narp/4pbUm/KuwIrSyHOFC1SsGjfLdsWwGRow8PLFDPHu8otvXeXl
OS8zSbSMKxNsjkZQRSe+rRRWPmgP9YDukKgtbkyEw1Arwyv2dcnHU+VaA2tmenJOPLkMKGGsuPIp
kMH81FUSCXjSikapGXD9NKwTTEg7+zJfnf8zKWlqJq0kc7MxTGj+XWZyUWN+sUoSIzyZlDsjgUN0
1LU9tdzkij3pIbz43zcGgxT/DWBqR3GOm6ssb05hJulZgsZ8IzwQzUpfjD01Cf503L24sGh9oE2S
eXlnajjbd8BOoBtfFYzOjfW0RjAG48Md1pSHW83Hi1n1esmiGtC7V1E8STJf0xp67KbvhnBlMjvq
afFUSGRTJt1sa/gSuOeAVwRPYD2uBk02O0jWSy6WdZohVt2Fvp+n9mc7dCo51/SANcE77N0qtLmS
rcD5WjVENu015RosajXOOznEZ7c3F8Rp96xNzMYbQrHDsFi1/2NN5S++RzTXSeGri2+e6a0w7QAo
xdaehcto4rP3a108b8sujUiNyaZ16Rj/I0WOG95x1EfZaXbzV32F31ca7G9DB/FT+bbp7fiUHGYb
iXuuYimxzphnr2L6MVzs9u8AwH6V1heQeaOdc9rjksqhpQQ16UNC2UabumBLa1eRSOuE1eSjw0Ev
PGvogFNW7NYhgLx+VGiz1VjatvQK0k67mJ2sxXhHYS5jZCrqcn0m78QQgu5TQoIOEdUv6NeotaZW
F1EHiUZff/ep1Ghz8BkyQK4W8pylb2ri52NQmc5DcAA9FRb0xW96fn7EVdLiIMaOW//SnqG8VnUD
C24EqneMlK+yQFZBrNhgRfzBfvtR6N8pN7/p1ikBZ8ek5rZdLeg8nbb1j93eY2/FWrHZeSPQrrDD
vAko512+pJwdy+JGqNQSoBv9a+G5/dagwi7C8FJuPYf05cpf6rxkn/sKt36WlIR9DAXAglG9+He2
2ftIeLS4nZaRGYQZuV4wMwHUs8AD4v4P3pHQqdOvgVljQeo2dk7nUI2rjIFQN+eE7SD+cXmmSqMM
ZWjqQsV8LjlG38V52J485eQwBRUVMtrUn5a2B3f4xlpG6XxJu49r78kLpMv8n6rHjdRiK3cxZUMo
BL9O234P5ZXdi7A7r2IuRx+f8IT8T9SJ2cBwvOgXbn1hquOt8R31MNB0+oSjKwPNJsfcYNxfXPgo
Ykf/Dm2kaXRpLZGWzhvk73SFz3xBTYD4MmVKqUWrOZ3VtzN98Rxo4k8kyDs6ulcATo75zggu6jzI
laGCvlRRPxUSxgx7D4xLFcDyFC19lgC968XLF2RSIZjr8xRntsRurkK39KYzOz5eSlQ03wun/MF7
hLgiaXtDcoWKyyDVAGvo7jKqg1lLkpCwmInerKPuHYGbYZ4eCIw5qZ99kZdH9Q06utDJQmZDaIwM
+RLeH4iRfBmG7Gcm2UWNSqL2IfVhxr4PdmpvmXQF0Nu8VcMESxO1hIXEzf+fa24rIyyURV26mPR4
Mtu5uwYrdgjHnZEJlNoXMVWqyZAC8n6aQLdLJMAct1t81tDRstpLj7tnD1pVT+gqB0CZJowdJ+EE
EMDVOV3t1zHjlzJJY+xWPxzupZLsRDk8II7OZvWAT9cRokdRBz+P5AWu/VlsMEIRJ8LcEyM3Z8mG
lhaMA4e0ZX24S7KJLLVsFoFnN1eGpTmTcWXj13I7Bm9tPvXQdXBxQU91IeGw6aNi/colxS8gLr6g
oY0Tw4DyNR1XCIs8a/rhdW7DzOcI1YS7RJW+Cp1eOSrR8KgiuWFPuURtldnti8h0ekfeFnqsAe6a
NBEkBSfpr9/ZdwCxHQ0JoAT2aIaX7NYUfSomrZFGJaTN3h++mbQJjrOPLMKQBHVxrKxLjfdrSqo0
BW2H1rCgLQ+Ghc1R29zCc39s4wqvs0wMVwGEX9pWOxxSYDfin9M3GYaeGFZuzG0FOAHH1dq5nu0b
zrl+6nLmE/BZS+Mn1VKf9vPIng3pg/3Qsjq7zGZiurUm8kuK1rxIMwMM0u0lGdftlQmIgig18z6S
HxWzDBtkRt+oVc7pYfc+QDebzL6lu5fTKFDJPgvaOHEN3GARSIXizcP9vlk9GPYyyLZYUusNzyfv
cJ2otaKXBbCzFeNG17PMOlp5qilGLptADDBMV9ZuY30R8gspVm9TstBG4Kjhs054hWNwIQNRkzN7
Ag/W4nAfmjcuwE176CZwV+9pPqNZyu6jdXQdaOvoeI4eD6rPHd/+IeOkXcfe6/lt/R2JTVDAtDli
+c35JpsxyP9wGYTlGkZzPeAkEX2Df3LOuHewm0kPh+xlYMThtZBIBL7GkgbDvUQEcQtUbaIkXrgE
gDVZftG4PfIdWfVgiMEGacY50oVz1lIXBoJ+vdaH0jnAAPwyGJNBkqgdtuV/JrNtTQE2q+hlwbRU
T2KvJgiaUiqPNo9f+2InjjEeMPqS2jSnPO7rd7izUn5YDPw9zKe1qnW0UFivHQBj3IMJPL4F2O0V
QHH1up8n7uBLNgl8vG3qFTagbdrv973kXK5gpsNDWxAJ45b9GUDm+3naK4Oh6Hpep2EHxkFTYfNt
JKJsuzcgcMOcleydCPkilmT9bCxESVLOdr5uaY7qSjFVD4g60sSiIx5Aprvsv5nphKag1RaKW8KL
E61OEYiCJ6+kxMcgk1Ygry099WnnW1z4rd/kYkAOMS4GdnCACsmoZRYb413Z5yHJlKAQvp4WSrv3
+FYpNjSqgKh187a/S55S49NI3Cp7/k3w0mTwtBppbpK5AUmtesuHNLbTiSDN9vxGIvfGqyYocZVM
n0UTCQMGF05px1CXu//BS9uo8vEup4+Dcw72Q43QW47V7V5xIGQPCTkzUbrGphBUMJgN8Qpv6bNi
Nf/NKfMx1j865W/FrMH2vN2RB9VYh1gA0hdHsTmZOH9OmCKrqPlBf0jbiozG2033f71/yg+ERkyF
5l7UWVlWzmZZDNXk1/4lXDuNShfigrF08kvCjbJKYHKPuLxC1cRkFdQrzIMG5EUpaK5wjdZ7fxye
t8zv8AK+d4aQpQaBbPpOybvMA2MkCCrDjLNpxgpH3bQlEnjscDX4jvsrUJsVtcm1gRGa1QUB93as
jOXSWOz4+jDy8NyV9IlGMw02i/DxmMvxW7xgdrYx+qlnqhxwE1SlrqwhV82ySjCqiOccIe9SsH4S
T5T9o+Beq0qFHpOqiax3sE07Hkquhyn4QuqlU+2r16BKU9IWkr9PH+nBHBxPCzjlyFCBx9orhSEh
yX1bbsjFyV8AhMfgbPQgMG/0qC3L2eSiXPex5oT8bSQk0HPCzeZqSnA63c4VqgEiOy+YRnItuDU8
RsUBzt4TqHh5/dUL6hY97q18/l6A58VdISxBbzbekToye4dsjLxBaTf+OEZuWmX/Ln8XPtcwKUdw
HGU0u6GSlUE2jcv7aFl3v1LtNB3UHispcIHSfJNlpQbJ+SoLlBrCb5Or7XTErzVyVmJcZZj9+mV9
0WcgFrBd7JWyOoYXNc1wF16zMYdRu6cudjwZMAg5nwUdD+c/k99WXGr64NVniGFWoYiigTHtquRi
LEGjh1C4QH6YDK7dyrBSvDjGjC3w6evrcTST/v+rgxX+fnT3RPa6sCC2ARWXqvqyCqSTYt1aDP93
hxa/T6delSYuWwY8B9zFl7bA9zEXFC73f2U1ewg1Hird8ivISH1ke6490nDc6nFq5wAN/gs9Hqf5
rAXWdDYcjdW2I9+w/gCjujMqUaWa/5PjAqtiP9qMefkzX1PPqnTeCgSjGi3DFN18icv3YLXpccjd
omM8Ka8timDtxX6gVH7ZMImYUZ8Z3KKYoMULtbrjBGBYNrCb2rUhNFRwAmX51ofCkwjezprJrbv+
L8U1nBjHCyFgEmMJ24gqpucVaa/A/yPl+wktk4emNrAVF9oXwwZaxoycOhxaQdNY0gvQDspADUob
SAnw4yY2prfuYngL9b2dStLzChx9+BnqXQ6NugFQzmPXMmI+ZSiP0+MWLiDTjF4srSu1BwFG60XF
9Aed+kyoPZmAopfPFXWgdcH9WZfCsfLFzvBzed60d3rIXoVRKQDIEmj5HHVY7lCydIC8kzYC+Zy/
gk7a5KL9WYzks/2ehxcfFqKIgcQ4SyLz788EUgvKnz6XmDN24sJNFQo4G4Zqe0Z488NONjIH+shD
lmE4vW5BwoHFOqVEwI/tkXKxMQhCzqgQWi4+whKlOjpJiRceNxUovoPv0L1jT5ekBistVAf75fNi
sXbErQjJrlQdrbbCvKQSyA/6D3s8iPdU+6+3FG1DxRAKCowJxqTzZHdaJ/oL9TJVEt3KDAGx2E+4
R6xMwCc495x3dOlV2hHAoHPIRsu78A8eRlFEYV+JivSb0cTH51a6hiDXpQsOUdJvrknLyy4EteAj
M8w6aQLc9J/fSrLudnRD6ux7agx98Rvvv8LczZfl9Dr4rFe41GtgXIJReXaZD2kjqYZkNkK8wxNj
eSmPzZdibwN5/VvZhKBtPvLrAoF1s/NFI5zDshCndgW2LsQ/W5geR3R5FKFrYwyTPEUmr+1BGXcX
BTgkRTsbk9r1shzLsdu1igJq7QKNSvRNq59YIKBVvMh9i1WM9OmPvtQPnX6EZ2PBpJbijybMQw0U
bL7AgKiYVfAJL+sze3bKf01QrxpXkOPPY1255/JyyzMYZ8Y7O6pumUI2/JbkhkA1xVO15xdh0Wws
68N8XhxapIAb8OKnzxs3pfmb6xmzCUseB70L/vD0tgJw8z0f0mXnBWV6IuiVsdmh/xv3mXIpZ3pr
RcBl7ut1D7XG3yZhdBRbFjQHgH4kaSZLzd3dQhjT1kCtnpxwbtuxyweaN8P9D+fjrxmDncPwZlKa
yR+/BA4nEk8mLF6FLt3/sfBQlHLpCviBWJNd1pcX0OnFWHgC5kQHf44srd1XlKJSBg/Lz4C1JaEv
N1YFJdGwX3r0mDvC6j3S/2LNC3EOohR9CuQcouor5W4wLUm/FoUdXF9Z2/usn/kA3GyVBChNKsdT
qUyX5gDzYq5egVXTOk1aiohuCds7A4JUpCyT29cMJQQ8xqFfZnqbuJ4NU7M0GX/KaS9kmxMuI9oZ
jvvaDuvkmwcyG2QLViGBccG2xRoe52iUUes/FqQQumsmVzCx2dtcJUZ6z0c1BnGVRlOkkiT/8/Q9
WvXguAM2kvDOgLa+C0C5JsbusxftbP2nLAmFk9rUQX8T0Zz1lvPwPIsqkAKcpiKGpnVvSSjA3c4D
UI9NJ3wszXu3BadUpVMDLWdo+xRDUwUzanfYtlMdkTlHnQ/e6k1BVXs6q/LbeOFFpWUs32gnBUc2
CNku6491qvfT+1VbFZ3kH6CQkpSco4TBLAhKFNWDKjE1IzZyczkD4Vk+012CRGXVgCTZrMZN7qPC
59s/7IO6UhSat3dB4de68ghalnQVdknDywGpweUkDz9jsMJ3H3DBXKEHnyvx5nEbGoRYBgzQ908u
LCrCqNu0o4OX6xZnVwznfMaGL+2NrXYU0CJkzJ1UMu6Cv8aefVhyvjPs2TIaA6cI5J1KVWAS0U4L
tdBiJI7EmwtPQeNXwS5nbTE48OvvnUgyNoCYfVE30eR3hJ/HUD7Rn5xLLxsZ29XUElvLLnkUkEKk
1SVWRzcWuY9Z87VaAocH7bC6yO7ncPxvrWhFm2SUS1ugwiGDRQLnOxJVMWjTTaR4EAJiwX7HpqLf
QVWbiVDKMNHazDkWGfCZ1rW3SHbbwKTmsebu2c1B34t7TplSyvfT/jiyYwTDcpYMF+1zm12HYgMK
77gYYvVhKTgi9RdZpkDiT9h9qcRHo25oVPttjQ6/20g1ExcFZyE3f1CIDCw9IrX+bGRwYPY10fIj
myr8dQWDfsVGsZPVBJTd904yA62jQtjchcAfQRx6vDA98DjeIGFPy8NtJ5EBgnRhFAAZU5d8J45w
iWzncwteqPoP5XzJ6TZ896ByJfD/opJg0kz+j47lIm4Oe+IO4rBXejHl0qhCSOdPOXS3zxbOl3dl
voU1O7ugWkXoE2BujxArU+d3zbzc786k6UFd1VkIIOoBr0eVYIpjynR133BnHnoPU2hP3bGXP13Y
ZV9d52DdSTNL/vHnlhgqDRxIpLTPcHijFQ2u8ycYPXfzY/3kXrcTlzRkycXhcUeTPFpNORu7DENO
6Pon2eOOk4y2/hIBIJGeE7L+DY9naNtWBkNPupMH5kXv/9TcNHe9ZHFH3F4ZmX9mZMqj+4ybRJF3
s0dj2qnBdOJRiLleVGb5fkw1qT/KdPvezcfGbVpw2AXfYFzAG1c3pkyP9HQqUV+nB1SpXGeHmA7b
ZuybOaBkIW+6pr3iJJu15+lgCnxf8bpsfB11hqXg1REicqcS8sjcqiW82eGigdHUQK0NLphdpVCI
j++6Iz3pQXThcu+XWPosYHGVVSYqEamggpqkMwu7E4hHIjDtxQ13bYWZYszMXIXJhoiibyoc7lVW
LJRGE1vqKcj401rvDfNeA0LvQrbk46BmeAqR9cM9WMaxDgfDvEll+hNEpgNnsecW54Lnk8t3uplf
+qbezNHYM0T1QRE06JkJmlEBJ18IQSi20lNAfr3M12Fx3oXvCgI5djdSVbwIK7+Dj8wc8xGl1heD
978I6Q08hZAHT7bDpKzEvN48WOe5S/AnBlen8m03PmncG1V5lM7bdvZ5QAYblaje9myx7FaVRLF3
FdLrHKof3aYwMF0SlU0GpKYJGwEcfFOmYWCHlwTo5Ul2RdZjMiXx9v8aNxod31DxgWUmsi8pRuld
yzjjvo80gW80Rx0tK4w+yqOo45CB+fMQk3VqcoHnwYhnc+yzdWdVQAe4iGT2RuwZbi7NwzOPnB76
boXyYuDdGpnqiC+kLh0PQIfSf0JoM96uWFk/GV03MrVkGGWP/6ecAl5LTyY26XPARvm6PHSbqi2m
YkHQU6sjXqIIeTPqx2beMFZYGgHJZkrd5rWjg33btuAsQrF3OOoc4Z6x4fvr6cSuDUz388cfXb0z
heaY2f+t2qki/OtQKqaJGLTSfX3sFBeWD8ztUjuralVG9KlHD8uGf/GiarUPBGPBevFwuFL8ZVft
LLzEb0rsdSBsXEU/IAwl1MAnj/BtSJIOOWrPx4UFGsSabEOT/CYVOjpqfe+nhCqfRtN339hId0ot
2gImegtgiOV1onuBnKjrKroFetJRl+CsVa8wAhBiCw/QskVxlcblA1zw37SmBZywseZcIYFl+vit
2p+uXWYNmhPxsxGPt/+OnUo2A7XWbr5bAZ4UmWeXZz+1eYGq4KdUsCoaiJ5NGCubF7I5nx7ika9V
5UMTiw60XUfEtEVk5CTaBcyEABuXeI/UtgtA5piQYIXkcKSEB3zp6Kb+uZ8Ul73lsG+s8I/FjjFX
glhbXyIVqtcebTOphxWOvRNEV9IZ1YLJEC4CGTH27pzmO0yNo+g5KTv6OFbPVJXQekj0T1nZFCJ7
r8/z4w7gGcZ4DLDA6GP7pE+Gz23a3zf4/Lf03DDvZpFvD2sHVXwCqbvjyV50jMIDvjOm61Hc/tED
TSRtDql3G93+e4y8vnD/5Y8U1L4vfzQEp5esB8pwEMTbXPhLmJtXxdP8JpUhUmw1OQ17PUB1m7u1
bkLiRjfsuut9a7o8x+3TcFDBxYXQyDViiPhabYABDtfe/W43ZAvmF9A3/s8TzlATW1eSwZUVjajc
OHgay+64TdVCbqcfYOyalCrGuFKLSKxpS2lhP/JagmWatqJcrrDjXKIZJ0w7DJ7BuaFzAVkAbvtr
7SuiqFCdFEsZd9wFAmAua3+y1iR5i/lujzZOGHM8ENswYGthb6HWcSD68nO0rCP3CxQ1xtmjHTgk
+Tc51XT5tnebBOnGPDE9FGAVGyP7yQZ+7D8czdHQ2mVdbeuE4prCNn8eb/e1TtCo0fXxCSA1Ionf
EAyX7jweJ5EzlCxZp29ku4OakqDK8TgnAhJdyikYUJ+7Leu+T4uqWyDYlWamraehJ7e87+arsrJl
HYiCrYT8lJ4tdu+8oo/vjym9tCybX3KwBkyUnf0FMzw9eMdd0V5RbRytHOeqM8gQSojM476XlB+0
zb3DHbAwH0xZv3HThK7+B1hvhZqEubPcdD8ez+UmKlYT0mDMirhOLGU8dWGpo3OceGMEQNiK56is
tUeKnTUfd3iW9mUwqEX5RlYEuit66Bix61Igz2ozRFXj2ba+zSUxbQ/BLRGJFa9X29RBQwgRKYNM
Pk+xjvDGfpIDhmFgToeleslmsOIwjJgQcBukx1D6O3lTNVM3fPFBld+2QoxoGSLJShZxAUoVp7yX
gy3x0/9BC4wYNOfbxddB1usbvhhy49qeE+MEML4YdiTn7XXjWfXzBfA29vFlNYKFqKxCSaEVItYE
0DGb3LtlI/5J7AmzgW0dxpsja7dveYJoXgHOV3I4FAE/3O1Q3YWQrwPYKD2vk8gZmwyakQwwK9AC
q4oxy9ppskZv2+zlAqOKo22fKfF1n37FSf4ORTtWxEXaYYmdF/G+iZIvX3P7u+87XT0z8yD2BC9l
rQhAQbcTO1YNHv0TTMRLOb5jxL3/PmvbNWUXOpfcJnRqNBmf1CZeEeSz+3c2JtIlOZjfYG1Y/Cx8
BxReJ3RLeoi+9wW6RBpv8t3L5ZPY5IiwFbTTShmiWwG5RDrQJvmsPVZrVGQQOIjT8JO6MCeY0XKi
1qLUzt5rV6x9Y6boOPlcVsXCJHHNZEUCErRRgZlbY6x8BsjZ5tskpQvnmK/TdsNQR9it/DGOY8Fe
aPxRg/63zNyBOnDiOBxXWvNpRTzZ9rwLUHMPyxLONphYJk8nz8ET/qD4bdTF7QLscBQyYVY5AikD
+YnkNP60F4/tVseCiScZqpcavBTNnYQl6MhrmEzlBs893TZbmMQQl5XhbOuXeJPbbVkzNK/xI1qK
zPG3RWTWFPcLIqyZxb5jkEjjocMrrl9KMLyZu2MzYhg9GU0xJTV/6/iOtGpOyi7r927IVh0SIMtu
VA3CGqK3VtpKubcELFw+ukDTkMk/m/b2RiXaFPQ39w+9z8MwkcqY0nbWvkqDF0CWuxxDeLF/okYv
9Dr9ODuog6nvs5wCz6RBo78YzG8DQkaDe915fKRFIj3pW1sH+vyos5AVkhlCgLtgLYUFGKJz24Ck
XAwHoCm7zZ8TPiNYL2Cq+Mtlv+ZYPMMAiixa6aV8bYBOI9cZpkDvBjaUSTLbZ8zMUFwIktL62Nu4
V/kmYHjtVSandMNTAFNdiiU7ddZSnaNI7Q/q5Yp75ljLo0I+I7MIwIGCEF+1+jGEoQV9KIZLU0/Z
kaGu3/MKUAB/gu0hI1Wx5YtE5NofoxIOXxRdpSMZL/rMbl54vFQ68lHJXN9noFcCQFBeFtscd6/o
kuPv1QbTGxbW6kwV73H1XDEK+izAeSjxRbUW0Ergh1PTANFIM9y+ImOrsXlGpAHS7GiKmrvFyNr7
vHZ4XGfnKd6H2eELlPqLm3oomFnOQQ2/EFWnT8B/cKwK/O4MvoeF4/d62wRWpECoJ3qd55xoWCEM
XLPuX/erGCqv+jR9dLFotOY4KOQkOo6iyrfZF1o8ZTZ/LKmYwxTS0NiOSU+DwbMqGO2LTLJXYmiF
2ksITANRW61TBGH9LaQO2Er1VovmxW4NdOfZkAaDDakV8FVd1HoxknzS3Suet8gM/Qd6hg76psYh
kGutiy2Nhx7tOUNpBwN9clpASrpZ5VwyL+OgpsF26CAuiIHYgWkE8gIldhdTbFmtbRKbcJjSarUm
qpOu/fFRstzgb92HuakeUJ/EXhA70UqpZu7D9rl9Fim68PU2rgpR9eNrqGB9xX6QM8dbA3K1jfsD
H9MoSLmfGRHFhxN1DFMApq4Jw4QhGCGdvqPvjzwQHJO0B5fxeqKkxsC0HqjMac3OovJAu4NGpEgQ
iOY9IOI4CA2t/uPwt3+xbhoBIQPGXxhlH210UZ9ijrgQfvV2RBT9YFlvxl4/Uh4HTYF5Dw/M23/F
rP4IA07bDuwyVnj5OBCzK642D+OZtpnTMZqUBAi6R8Zb+7r/etJCxWcMplsE1JIMMRpDiMSSnP7l
wJR3ByuMhXBnDEUSeXBLdfoX7ZftUKjDoTNHPrvj2f5wDckovR+VMn3s8pQSpjuaBrdKT+LtiN1W
KNsREebqZaEKOU9hSW5sxkghOXiTkXu8Fnoalqc3juafSfF1dcS3kOcXzgoNxxID+/W4lV0GRlVP
Hpn7pHNZSgHxztro4vzyasAAh1d+unSVoVZMor2i2kODgdGRVXUlOMGaMPeLDnwWBpzQNYZy3cAy
SlQGFvknPYIgFIxmgx+PodC6NbaS0R0aM7WFVnccn/qhiKq2bHFcBWhtw7a2oiDD3fQ5WoNMbPZH
itPyt6jjEApB37zE/3RpVlU1sZb1DHNMtP1jjztgfNF/v/FJOoUxL3gce2kOch3ePAMOSK0wcCOp
R0CetOyo467PbgCd1vCufZzwUEe9tzDzKLwhZP5JmiccwPN8sMRbhr8l/0Tfcxb8U/qOniTZ5VEL
HJitRnTdZUq11H2uwSAzM2F3vOv6apahRaiDFkhPBTB5HlhrhW6xQHyjI25+czmZQumGf+uoJIhq
tzpLcNT8CVN/pH3kI+D2aDGkA2B2EoPqaHcwmv2FbwbaHThhP1IemDVmgLIvN36AMcpGw6Y6lKyS
pBrulWQgE1T7qOjcPUclfmKXiZEscSMQZofwWwcgtPUZJJiSpt+v4IQIPOsJZfCbWmMhB9yqaVn/
U5C3E7d8Nehrf6NE7qg3Ma+95sSm0IDyfBtN8XVDgyTaORSNqbKAS6qXeAdjDF6hKfav077oDnVJ
ojFuvC5nxOCXAMSbGaZS9l0eGRj9GF7UK9YsG7rt/IAT13OmJD19j0GWgBSwNcUufiSrgs2qD5+t
g6Hbg8F8rUAvAIz1VRmpjyCgeLFkgw75oS+UOxNG+rjaQ6wzBLFCK3m2ibCjMQ1r47fMKNf+U3Vi
AOOGTu++UYJIuleCmMz0+/HgRlxGT50DcrfG0bur4EbRzJ1I2a4eME/BjfPv0cLo0G+AtPAUeJa0
Z851Sromtz8itayU2xfh3cdQgL32nImKvIG/OovWLNk1ea8LTuvG44vWE+6dohenX2pw01N3Y6fq
CRVKFM5ix+8CsPCUkaNa/z9lIxDkfiR7KCJnIBMWavVcdJebxLHpCbN+RpcODFRwq4RcI2e8om2A
Q30VRqn+XteAj3u59eDpzNpA3DA0P3osdR9H9t6KzPFg0ZJDIPJBsyaqxEHI0sdWk1uqFsUtm1Mn
7DZB3AnzIfTAeRMoXrjRgpJlvb+kFKvOjsGJc6HKuqHKdAvhZoNE669oCQcWdj7Qd/AG6O9Ax2cb
2cr1/DYl9IXTq+XYUXm3gwXGVJn4zsoGxUELFIwZwS7jgxTySpEkVmReOCCP/qE0PUFS3iT98qLh
bvw8qHcXdb68EaG14AHU+bcq3G9cLL6S1bHrHFKMpit5XgIoNLy+04twm8o+FmrmDEhlU2IXWLQX
0hpS9Yz+vMQLlBvvBy5uvjDPFcOKAGl5TeQ0yveqIu0SGgieH4wzoLcDDsCs3+okfKLIRL8/Lc4Q
yc3swAQOgZWYczWnRGPPutKLoORmLadRUJeyZAC7meue4FxEEPh+xhBM5JAH2j4uDEgPq7hCVUTK
txbZ1gdmf/B4/A2XxzsiYyVLL0kM/wcXC+Nz2ZOKNsgSTgVK01wwQE+0zQEdHWeWr++z/C1fO1gV
KW5xTvIh7zi1tF5S+P16G+F4iB5nvW//rG/WKTtpA5qyWkjLcXZJq34i3SgdS9jFYRQYlQpHIytI
3IHfAFiaWHjMDEDjNMy3CZhy1jHQNOs3Q/ERJz5sJwslJycy43+sZgnx9J9PooE8ZokEEZA25pdL
x4Me99DNR8fioP4HVUsSBEo3YHpk7ui/EF3p6zHBWfOxMhkn8ti/98V6uXDFSQ9h95/keVj4TlS9
DO3cBMa7WdsDss0AKt4cmO/pzuAwHlqmC4JfD7zIuXTXVZowx4BIyESnCLLVp7/V4+0klR860uNA
oPx18nuTISlLQ0vTBIp/takf5sPYXYxkcN1B6QANJ8iVIWHzzjn2BUPjuTG9zxtsL3/Mo05iFrlK
VAttAzhcBLTuh1Turq5IA8KF5656g3m1MMcul4UnsRDEENQs6W7nIXoDyWHxMB8NRWKiO8nHNgUA
27cch6mWt0JkBF2J29zfWl38gFCgHxcy313TMN3P980fV/AjOFz1+TPHbsZq+5vCybQiplGZ1w7+
QmZOb7TT+dWBZoA5NFqZQT5lkUQjS0xrXoM7ZYCvrvJW4eozKQHTl1Jv8Xqst9fPdb3qvJhwYduB
LRBAc/x75RrOjo2BntI6uJFuYT8E+lyFVURAjGxW+5cYUA33MEvEuYFJzuU6LyGmG2WGSQvgCraL
aNgi+CPfGisAPT6vsasqQ5yppcdBV3Ke8eEUSEsnSBnGX+Oww95hPmE6CL49aMi7TFXlssjRPz3A
BVug4irUxXfxRO1R0tvhljrgNSmq1pO9iSvypzQ6kLoHxcLsY3cjKaoax+tpX0WQbwGkJVS2FTkb
GYzOgbk1+r+NNn4DfDQgkumfvheNsEkUL6gjrKD3K9YbXOdhERXQaYJA6WZtwJ/+ZFeHsqPSgY8P
YfMbs1ro3EdPH2wxT7GKZ4nOrZtmPa1uAIT4g7t43HPL4U6713vK3hLExQoFUCtZ+WH97JJ5m0iv
B9XfnGXIjwa2NQowJ2Dl1zLRiyAhCHpvX9sU1rbVdJU/sGzA6d5ztvA5WkQz0sWFnrcxprQYlHye
zG/ZF6Tk4G5q6VtPYkl3WqIXXIsyXdV01Z9dLCH1iPQz8qGtADZRI5QRh9jF30Czdr2h8jy0aqFl
w6c4rD23Z9fSuXHIDVISeYikHx/9nMySzDNyZPiPYDj2oYEAiC7mvs5fajeHh/2YQI54oOyLQ4a2
qywN9sBEwrdRsVrvE0JsSeQw+GKFNQMmFmYSDxIYWsC7N6ADu1FXQ7uS9ueFyn07kdX8/EmVGV1g
BI+hE/3bsBRBq2367xubFbuOLIalkj6qtlaMmO5Oth+Og1qI4vZYbI/8rg6NSJ7D10wljTFr277w
N43Nku6ND1Xmn4edzPJMoCHeAPlTk+e1c6wIF8z8nel48RosDQ5qybC++QUxtgkK3PtKl6Yj1stg
Z6qoo6LRmHrpI63J6BD1sfPLcbdMm581l/L3+yl6PKlwTXWy57PZBzP+gqMHF8CoRVm70BX+IykA
KNiTV3UIkbYoE0FvAuWlzIb457qW4LIbs5QiDRXGOOVYIXbEvQG0fGn6b9amSFgCijHfIeI8ZVAT
ZsT7Wt0HnEhCXeCb4EIfcVVFazKKusq0vl5apGD+yz01b+CcBBtwTZpRf0K/3k25GixvRABd+Pkw
REgXK/MgFqM3CM7ZhqC6XgZFp6RsnusPOC+Ag+J9fxMMURZTt7WSUWq1fG4PDepSx6vLh4oFVOuH
ne31a7Pl46uyzHSFQukuscIsJS7jXKrGkKdDLJR9qrt0hmEFfOzsJQL6uFCJZyVIzBxZ4B3vpwZh
0oGhJUmDF9N9CmMXUMI6MF5zqEA5hr6hFK3ySpUNzI0jZHnXHaikeFcFxpuDwexxcsFpnlzI+gN8
z42y3iz9A2y9Haxjeyq70ZEG8Vgcw3k35OJZzTbjJ3IH5UcxrhQMXucpbz3H4buDaokJeEELvk9F
GbQNx1tA0LLtoXDjuGl+e8kBRGJjTqm669BZIy89v7P6jg6dUW1MF/AsxYkiDX5AJbFu0xISAOJk
r/4t7vdflI5fxxQ9VNZpXTQ69uvn0r1/NwPZ5XTy1AjxI5zwHmgYkoBcYkBJFFM0BdLZ6J3hrgq2
PDvWSTNL82iHXTFbpY68+6RepK7Cq8Tn3MNTsP1dsXkB9CNTXDIrbcgin1cCk8XwG0KBroV8cie5
N5RQkPnLIs8qGr03XIiatcYcHnvF4bPsdt7HRVWEOD3wCoLg1Sto1PBqwp/iCOITw3BFPK+411j4
O96cGXqoBGiVY8OGSW4c1hz0bOeSqxbWAToWYq7z1aIo7BWHWMWJq+bfH3D0uKKByotwW26tl+bu
HbL1eHYdICB1DqIP4wq6wkUiFuTpf7X96OEiSSyYvLcTH9nrFaLuOjLvsj2VIiN5Fkphlvqk3By+
rZ58VyX1ggaySob2cDf/9NlcgsGFDRI/4UCdVf95MGVs2Dm10qiJYH7fppdgRKVsWRKa+dwzSpwb
oEF6t+O5q41Y+lxbp2SCC0Tm277yHL6a9SZ6UyH3S1tnk7ptqGjznp8+VZY3M8uY6pSRy0MjXQQf
VIzQjx6uiBdOu70D+PamXhV5dnFZz07+ZvYcZriftNwTwJQb4eqF9cFZtWzFxaD33bm5z6vcTZMh
wMusUudHPTagUeNqL1c7ERCYZt97l/KSzguT8pWHbAerUwSX/kCDDbT8t4d+YRNZpUq3HiRuff16
fTCg9ElfEYcC7R37iuEaWgsOC0Zjgxkm2BOlwwPffGXsNap7nA5Elj0KF9gBDJivl15GTwjEWag/
qH9+JaiXIiUNjEFvNZ3uFyw3nc/iQCiD/GWm8KoLkSxYWNTEZp8cnA+rXUaEjO2ToiFN/QBeYJKP
AUziD0hdw1UDDwU1MzUZSrByHsoi+LUMoEqiPCHxYYpDuIMmXgYB9/GK4bLv8ri1QWl3T4HaSKfr
OA/RwIq1p1w4MxJ98lqLdqR11aDYzOMy2lmhKDPD4dFG9pIHr78LS8lb6W+p5qGXr/XkBsYz8rQz
5FNVMSEcKguN3k55at+mYsRWxxfNAK4U+rwjqCnZy3+cj5GYIKrv4WHh+/tIwqmfIecKS0lk0xrt
tLnvKGFhITSo17uxBq3q7JqWtfd2jxifNm7VloUBGMuIUXcnr3VfQYrjDuRJPEMP/1XIKydkAyJM
2yruOkvlhhs6YcRu1sWve/4cX5GY/5oasPt/sZihRdG/m0nhxBYgz1g72YzVqzHdsaVfPj+9ta56
8jv90Xc+GQaF1R+O3tmLGNxIpRWrEYtLaQcO+pezIyb3ArQKCZ3s571HBptsoVuqGiwwkoaU04xZ
YPZXDJmdV2DGXn1aFrCZEPI6Eo1JA+GlUV2cSqK2yR5eaiUOBT1+7z7wugQaM67n9sdhk3EULpqs
27R7rYjqi8/Cv+oYKjBu3UxVtZXqWfuW/BxA/XWt76Tuvb8NjjfyWa2jyMmTwxxo9iCmZwyoa9/b
3Tm/Fh/sCHmunH0/pYbpAOYzQn3NUmy7xok0XL+38FI3EqH92OoBsOXPNXGSaGumM+1yKlWeeRqV
aNJqJ2VfGcGNKQrO4bI8+22G2jLtv+KDyyvETfxsS5aijcMEfffqQ5qNW7Eci7WscviX9U5mjPYf
zn5F71+zcaL6MSnUYq0PpH0yBHtk3Doqb9PbBomFCUqEwovl8ULTEyir0gx8slS/N0XWc9TabOUi
D7wNnWcHgpSih8VzzGhJgxCuSU3CW0UEkZr4n8UiwavS2jn01ODMWkblyuM2IsB7e6sYtOTOMIiz
ot9DgqcYmcO2BgPXjnz6f3WVpCudLw9PlUfF/djVE0IBivR+lP+FBAUi9ju0NNN9K49NyBrWZ938
Rw+Yj/ujpItKhj2AU2ZMhTIZdZL5cOw+VcH+Sk08imGxKDES1JMcUf4JKClEgv556EDswGuokEP0
jeFz+c4SFFM3Jxl8O/ZV3PGhUXj6cGd9tOmi2CmWaGBrpWgsA5f1iZ+Do8xzSLsfgWirceUcPBAG
VfTE2SbvtsIpWJdBAwYAwB7SN+4JcMLRZtv5Vn5MzJxSR5dgQNQeL+tr+zWdeF/M47Nn7k9cQv5g
cAZqYFQXBXLOq0HhQPMY/DAtkhs2U6rEspBU0QUROc8HIKnEdh0PON2pFcaG3lQ1QwZfDvfv9mB2
VR4TyyFGHwSrFG5ufm7t7qSe1oQlLlTvI5g2vklFagtmlUwfCm4VXq32QRDTXlwRdcyfy9q1VBp0
fbMgRVeBy3OSzB1GgDiv6q2N+H+jKiJ9N3u3J6Tdq88sAY83D/rKrdAe6659c+jQO7zNxlHP7XjM
do69G7ludXKdFXGGg3z769QjHIAJlAoi6ABfCeuUrgx63sTlgIzzAU3eft9oHexyjVbnftuGCqWR
e4qii89WsF8coIvoS4WMmA1dvjuAPXLkXXDl8pT6DZjbErdCArbz9RG89dpuCYiHdjfekOi9KiG9
bS7jKuIstNGlOm+ybo8ubExX5iuused4ArTf2TD324P2t+FXnf1CTFdchpbzawH1fdIiwtGlkeDr
19J3YVMUnKrq/TBf3NbPQKK397bZqXiQtprcceiy5XYmdMzWcIYpjLlr2C4Uq8RKJ5cOlyNkQbB2
ktnAI7pTQFDnV5+53e5WDu30WWzUmOmpYhIh4HZM6U7kaJ+3nhoHKGJ6A19tO8Rg0eOslo3CsWx2
fyCO62oX1wnlA+PiTPquaMSRJF1vHHDYnyK4O+RuspWiKCM+tDJuNK57iarEfqNtme/EFQFVJnol
eUN8QY+MT1lerjahXSDa8KETka1lNMFztlCpBA5XbA7ZvlwezUkvB4jz8TlqafSviZ+O4X/TWcRG
4sWKzLz0iK/R0OR7etUer4uzG5vOeWp388zCkf2VIBPwcO7R2H6877xRqlRvEkxyEuGChM7Ox8Fr
llaO+10w2HVxZoFZYzNCir4OHez9KHUDaMV+Vb//s/QzyATSNcWVzTHgEJMB57fyiw+0kk24Dyl2
DEaUPm1qwaVgpx3oRx7cq1hsx4OKeLsgBijJpePf/cZA45iOsCKCzbjaypes8tOM3mR/ha/QoPdn
6nGWZa11mffEjeRm6Gn02OVNiy7JDd2QpdKbLRcg9f0kUnVLOfqyaxrHvqZ7X5M0vytDb0a2r77j
jBgWpgZo5ImjVyjaYcb8cjVrkeOp51ziezpbOvr6s6o9dwu6m8rGx3N1VeTB8hxuFPLDFElqDKsO
21Ke8P3XwH7iXzdEph441OgRwonNe5DSi59iP+Z3a9tDlz0isvF6e0aZOsdSTa+57Spvxe4CZckJ
zug4NVFUfOPAAJynN1hMN2Gi1RwSDqBm1VxmyY+cAMyiapaWIEBWkrTeIYGyIaLphD31zL2pAiNZ
AD0NnBCH6MiL1KT5xH95QOjItsTJQB/fEZchI18Dl6NVgrwHDJbdznz+SdqDs4RZS7oON6/vTBTK
kz8mhYeDsIr5+rSPOL0jBdGHx5mdfqrFj91sTHWk9Na4e5Qc4pKp5VdUJmIYLfcz5VQjA14KEICu
7wg69MDjDkKSQC/vjNgttG6v6jkZLlsRfVlb9pcmlRQJEQfZowSOar4t4nKRaZK6AtoLzHUzEIgu
nFYJ+YP3kYiACADkXJN0hXQPukIWXP0WyC3hBsUZnZVUOymTPpjyOD0dcZoFcA9P3yMu8Wlblq7Z
bxo+yy+RzW8B7qpNo8ehEB3pkNUQbPxHPCvwlMyHnMCzzV9/UQQoE9AiYqHOxiPDnERnSMwCB6Pm
UEXd3IOGAjo0nurNOkxlks8F6gdU8DJfa216/oiBjux1Toni8y6dYAgmbdtb38UESxqB555S3X+S
pbCss76DgrdHIPeqAmZQAhlek6kTjehczSHm42jE+lwQx/5k3Kbfkp6oXkKUKg1y3q2BoV4EEi0z
kKFRqbXKvoz200VYLu1aqWoRNS+oipNXdg/wU+3hMusRJm48Zjo3ktJ4+LXkAn7r8EgDV9kIopAR
+sYFR/6qiNGAj/11obrMmaZxxWUPP0WLC5xFYKBwBSdik1TODJ36wpFzPOW28PD0Qeh9X7FW3YGs
EET/OhI0RVcJCtDFGo4ljKhVk2MYjr4ANEIfNCt6FLO6Qh5K1mnl7+xKaf+nwjLENpApmdI18Do8
bBXSzcz8awX1WyhK3K7uY9UL53uEs61dNQcEc/bLdaIvnMXFWHz0LfnMi52yZFPUoWyrQrSd/g1P
fDZ7z1Rx/lwcgjuaCUFibxORXTNvgtFrM6iLoNraL6hp9Rresmdn1f7uLqJ2CE21WYbsjZOIKyAe
G+0LEN8x/qLznz6Lcv8sIKfzJS8fkh09Jo4LSWEbpTQe6TBccOj2YlwP7kq3GJ4LL/BCA40xUTq+
Zd7GUSqUpCAipQhEHV1BSPeKVNMjKHE5DkILg4vwA7ONaiqT7omf3UPN8M9Tz+q2QU+YWM87nlP6
hGFlazP1OYLhnZQlKF9sF2irFK9ayZ+h+pBL85ZdpGuiu1wz+K+dZZuq+bzFk53SFu6g7xxdsWjT
0I2JjFVgbAamiHEPdCzZenPoOgJrLUsyY7yvJTVeR07QRZuWV+gmv08c3uM18w1IAfAWndous29y
0mzwOGkK+j/vGK/gIDlO+qU//exCsp9J8jpNE1256nKWJ0rckdkEMgoys6tt4ykfjSfBakaMd+ds
EaWsvXAs5deFmV3E8qmulvvNOmxv5a9Mt1b+NaxHd7KiUogHvY/RO4cM8GQDPB0IcVLRf7EnZ4/p
We0Jy3EWM+CVlqEe2ojqNwRznDLgrICNFT9pa7lkheT/5yWaUhb5P30W6mMsOCiIK6kAHLhNttCv
z1mnT0wqDjt4OQdDmj48WqD/EEm2mDxmp/ToDNcMnwLe6KjBZFwy0cwbSjXe97HFkJmANfk9X/r0
+dW3BMKcyCslVfoIc8P57zCiOqKVNzG61sr7E/5ZtzCTKsjHlamvlitbp2dDPoal/Nrbk2BNfMVc
DbRsLGPZQReLNnB6Mg6iEpUCAhtHEPAmN6gFd3Stt2K/EmLwd6mnaOjDm9bvHoJjkC5JQr+HB3P4
ULtk7mNBeepcpQiCIrBCSlDuqP21tokFDwhE
`pragma protect end_protected
