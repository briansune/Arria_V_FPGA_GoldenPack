// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:28 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R9vFsbjGjNPH5NYX4Ktql4da5CoFwl5VPYIpNtagqDqIah3C6hXMWpaA1GNRJ8bO
SUdqzZVr9tmpbVDRRP05BwRyOviJXVGanx9TTD1/yeR9jOQbsTWBm+4TbxAcXhYv
Y7UZdGnC4fFe3BFrwZdKo9CQw07wzxxhxp5/wegWdUw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
hUs+oWU/jWKwTGc6aG0xhqgaWyyokimgmkfSGiaUv2eho03zbnaGk8CT6pmoZv3p
8vMrNy/E+oiJ3bWu0VKRFkL7Qf11XrbITRp70Cn78U9DJIwcCb0xv/mIokM1tzK0
P8F6ThQS1kCnsiK7gy8A2MRtrmM56sp3WJ66Yf3T3YmlOXSRAfNPeRB4Ctyy9THi
zcmwi63g2dX5yZ9+6hiuovohFOQ6dmGO4UeG7SXFEbtI/Z8syhebei3Nr03qmx94
xFpM3BDHbhKwMXgaNW7ce1iyouR1hrqmaGLBx2hZPLgt7p95sHbuGqZBYq9Ool8M
5IRAGPeZSJbBh79sTZsJIcL1zRBouWyU8R1xlB8Nl3h5qhs1R0/j1EW47XKzpRr6
q2Bmd3c4KkDM9HvfMTU2DDIpzivxBVSVp5oXRxN6GbnWSRi7siHGHFOtGC+60WI1
43f+IC1idL8QhMUG6jSz8aL+od5WppI4WtRRwlreF12BBTrIG60HHrvyvxKHVnjo
BSUbPv0j7rjWqScejtUFnE/mmIXTbUjTzo0L3bxlTrqpVlLHUBnS9UVuzx4wCvNk
14i1+38nTwu8outfGoq0KovrIDG/sao/xjQMLWi23DyBrmokMzEIZwcojTLHrxc8
6vIGquaoJSe4kjP7b0mH3aV9K2pUG7blF86tIg3ETvrsfkkdDxO3Yrf3nCp9Zso1
YFX9uKzo7Z+U4G99DLZbC6JKcIsuFMh+AVDH+Ai5amI1u9/Ln32aH0HRziMf2i9v
pKXOeEFKWoXjscyu+FD2p5ScfqBOS9ygM75AJdZokQQaXmuvDxvkTYCseKRzzMuB
gZqdxvUEs/dR7RqtA5l3J3N8F7EFsIfRBhiuTn8YU1W1V32QnhvBYIw/lXy5hqCZ
qoaXkLX3YVL65HU38pI5rfKR/LwWrTO6ojvquu7Sb3sJysyqCy0gODevdzczKjo9
Envbl1ytR8IGlaPHOe5FXViz0AIs2uHaYe4BRslu6TCWkTznwHf75DpDYbJ/mEMF
IWs1EsQNfxNOxHdczC9j8zs2jvKV8VmxJepstFre0DO4kXKlbU8XfnyvLlEb1FFU
p8K3k7hlkOhXggZpkqPaaPyPcxOMM3oPNRxc3ziv/RHRNkKaGZA1Xz6jqliVP1tB
DLvhA+QOfrTKSQajo0So60bYzwMfDcNNUOkbtXODcyDyE9O/v3fN6WGbgptaPL6h
mISMEWjxvjCQmmOeRhJh8BixLP4o4PE5VslIx1r0JmEuO0ErNjgtd4AjG0I7VGOk
RfNSSmMgLiS/dKoUIXcvEs1BAxfD3ShPK1NPu5UniDp1NiXmIUfkndsglwMu8Y5v
IfJ32HsHcQfFJHzLGATBkll8N+5fQpvgtGRkT7WjT6hD6w0XLLkRq5VF5rsFjtXS
u4fdQ8GcDgXlns606OfwFtmcKUtF0atKxGzhNBDB/Sl1gNfwxj8y07sm50xTOV83
KX5o6uY21hypzvvEtqfk6khK1DPn2AhtHq3Nmv36+9ItEAUnjchmvBdsjh+qCS1e
8WqeQck6XjSLNvxcFzRX3iktQo8VoXdiUBo59RLvr5cquUIU5eaLcVpa9sWTsEes
c85Eq7K9AWKzawlw02h7bb2r8E0KLB/T6xVq70FO6WiShmHNCqmRE41ymJlBQhOn
iIHHLPVvRGJwO2J0HYTnMN+b0TuR2GPxwryJNKpweDKcn1kxXpxIzvGsE0cFOdAO
JW6zHZWhrOlqI+34gPA7hrm7Ygti5X/vCFlRqyOpOd1vdyYi2of350umkrIWuGwd
pBzdAt0jqay7T57v6tgquq+6eYk/9W6gvi1AGA9k4htWLcNN2YH91vhiT983fiIv
ugObU7zAveUecbmW4n3JBGl1+fDuIjVYG6IMpAwKBSC4y9VSOKNFNdFnoM3fRtn9
ZK1+sEMGQWHXyH0Yg+Xvax0swmcq/d+cPFpHwwT5xu2rVycoZxQMeFJH2rZcZJXB
9DOhJxqO961VJzKfoUD6f6m4MXQUwzEStEPh7rkMA1RGmihneeZx5zxa242nT4IV
ivg628ggKkLqIaDve4fS47pv1KpX5fsNWrc+J7GVT2b2rXbK0f393a+QuvRDS/nE
CzGtH4Rcsi5WgMPragdgZKCKWRNpWay6gYKdLvYwc4XLxl4lgKTHYBCalirKGJ1N
Z7WmV1Fo79tKqEvsF6XJND6KsFbgt1mu+XdbYfg3yzDc1qBGSvXP7pNQhuwPMYFJ
EZT6ca0uTacWsrPIuu4e9in2Reb3s+D03zVhKxV+Tg8+7vg3ikzCO2Z2DwOht+lF
fN03HESLOqIleXSiDmjJsT4UsJJPX/8SgV7z8acKaAANVP2rzbQAapnyPAY4P/Bl
cKnhyC94+Du8ec5LEcgFgrvda84XG5JNqvx8vt7OVBMWi0ltql6jh7qFGuGfVxYQ
NkbmEXhvKC/N2u77YyFE1x7AuXrkIqH+jiLMKSmRh1LV4TCxmZgWPqD8djlKfxkM
tnxz7c3YbdZFfdB7EghL++cJnzhHOFZ/6eJjb1I0u2n8hVEI7zSEVwQbQS8HYVMA
Q7xxQVUlq75j4Wu1j+xQDO+IbCtZgn+5+Hn0QT3Cl2+Jy0I/aT0yl6cQ7wU48Prd
r3QmRvykExXZYgF4Aed2y+0+ZNH/YuEIY6ap8XyhRKoeyq3X3CQf4vE/0yqVxGnB
PqL57YeazuZQmbe1YFFvDWrxO4xlD9VbkGKpB/4X0Mck9W9MLizD6HzWrnREfA7W
7s/zkuKGOPGAQvrqnUtmqC9ixPB6RntadX2TOJ2u0EFZYmHd7xVsTtFeHDXcO8ES
qm0heqNr+MI96auM8B5uLUvvWKcMsty0vXI0otKSbr6yGkegr4OKf21nV0jZtLeA
NYer3eunmAwq4zLXNS7JTeuTOYGgMHW0i1MJ1Yo8iebAFIXMu5n0LX/k/JEJsGKh
Ent/XGOtBcoKUdQ46ZMkRQUDnZ/frmquoY3eiwY1kFWWk2MeIXCdZglbJOBD7323
EWUa3OoI/FsL2QQnGX6LsKM08vo32SkSOS1uFd0vdt9mOUxeR8jLcrcRb3ZodKyv
nVT932JgqRFGMoRES9LxGc16birP9r7c3ft+yc42FE6uHqVoKx7aNwZ3Fwlr3qPe
7wCHrEsL+SlW+vKPAJPaQxqqHBDc5DNJ2lLfj0LI2tSX9WzhZ13KlDFiAf0oq6gS
EtN4eW4sFZyVy3wfPoX+vWtfpiEbQtsgMI+95+EHfnfhzgOofiQnr2VoUj29Oxir
jNaDVVIFj8N0mlkSYI3m0uybzPSiKJERfZG043Vej/K+8kaRKynLQBHcc7wNBxRY
6da1gmDLitO6OENxVhRR3lyiPhSGfHE7R39gsCzU2UoMG+75X3HNkXvI5hWdDB0s
7wYJL6dbPdJnk6lyO2//YouRenjrOtGZazAClsVlsGpLv5ATdRvJKDRkEwyfHhl7
uOcYuYvXzDGIFxlw0svZAI1X7JK+AurpXq5h9gYo6EB5uYZB4bB2OzDnm7o+LSgP
Zk0bWw4Of11tqQg1vnafn+5dvEvakOAs90fvMkXqwEplWQCkTPPfiDaoBkPHoSHk
FqClCRD3YWOTVuET7v9qgd/PnKyOXVIfaJKI3Wvh0DJX7IS7t9qZrIXzaRtKzAeM
VKzAiHvUMQ9i0j6V4cVYOeirVATVSW4faWZGfHfuawdNZbbqz6WAM7f1RKt/GsJc
B1jz4d/x30TuCSiAbGLmWQxtzWVaVZx/X9YTLUnO20J8fjRBfBJK5uglmr5eXo3d
vIU33vASyZOhRQABvr9t5OVsqpM37cBynrCOhC6Sfhg4furL0OYluB2ot1AWTCPL
Nover9PyhBakQUJQPBG9+C71HUd/YYPrO12oT5idTDckc1DKRZCV/JrRp7BeU4Wx
WSXtTr+eZUscGy10n1qDCRtSL3d/kgRn+z8M443g2DpTSahsx9AYb2pQoI47Cul2
bjb+0g045DVwPxX5MPPTdlHdY3cE6V/Sku0w7+v7fFrvuvVEmPPF6KjmML/VtrNz
+ScpJa5QB54dS9WMN/9Do9gh2zLd7WVAOoryBlCtG8dpaPfyODARlJ8Y2FgCsNiA
Xnt5OJPe4aNJbkmRnGqc+sqDavjWepXIgwV/p1/D+whlqZw+l+nA4BbluGQS9z6D
IaOv9hXZS8NBFXviexaVSX3Vdt1lqBCN0QK4/Z3/lBas8jDKjZR2BHRG2Dy+aDdq
E9PyXGg5dH3OM+nlr3quI8goEkCS8SwOqz+fe1nn67l+0tWddpp7U/FwCvExj9h0
ouvoFFVnq+mjVAHB3vRuWxoIEYqhCuMKkKZSKQj11Kft6evTK/olTcyOYGbgTtmp
aRwcgVbMB8B5fqUOY5HsBg==
`pragma protect end_protected
