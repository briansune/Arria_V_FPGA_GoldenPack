// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
s8e64ZLhmUA1Qicj7uOLizodbaYgMPHy+P7pN5Sk6bmm1Qn0VwuEDSTg8DqPf4gWDxmyFyl4hjm6
l8O2Xhv+6DSjFzr3Ou9wBzEA3PQsQOy49WsDJXfJbaqR7/hr3fIvUtEf2VHyQNZG62j9SXvcfOgU
Y6ZnhQ2oetmOItMcAiiL1ek9b16z4UDoLaJdCpKMrd4bIceFBW/CyBK4kvNeiC9yo+4KOkGIvmhz
y3dSftgIf07UyIXlwTFb+jQzVfP3f0NDvYInOykKoYEC8dcp6/cJ33br8H9ony4UID90JOKrd+BS
UVHaybTPa3Lxai+kAHKwBScnP5h3A76gE/IZkQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24880)
FWIJg32hRvoBr/nWmPA8h42zBHRm5mETgjIJcVOnycMX3LXMCWF7jlK/4cJxnCngBpxN0proUo0Z
PvOvVVQlTwP5hrxcklat58Ex5O/aGpsLs+Rox9DIdWjfSL3drx8dk4VnN9thBe5ol9ERC0SVHflY
ZPyWPJ8w/4s824cT6+syYDWAhvTZ1kPfxYfy2H3ooTfiAKb9pv5zrKhfKNA4oPL+nPAoVIcHne0A
vQmIOsNJE0x116gBzG8NxafOl8rtKFIvYBhmAwcBXfe8c6mnt0A/5H+aCFozjUX3vnO8XBJe10oS
v9I+JOLoQSCg8kyBWTYywe9t1WhBkQCvO+7XywUb2ACpKSrFEMxeWAcYt56upRebLl96g2zxnLDo
a701TerdKhqDKcxflFXp+TbCmU6kjz4KEwXdQWocWGdNudJoOUGvBS+E4oAo9Oyyvh/d34yje8ig
aGCqAgMA8auoSjAvxLoYag+Z5rXT/V/ZgdNVKqsBy8gk9rgUdjA7gD9L9iVGZ2kz/HiIIWF/vOuN
6Y8QuvwCQjoC83vOZQz1pey//pbFKBCeHqfuLyTo7izDcMyVtSXBLr11TKJtx3YtHx9q3JYpxxxO
ziHQfUkld3uOzHd5w7LA9oJqg6fUHJFHDP0tLWjxkKd3VzRcxwc+NTtIXgUh+bRvqsTlwVY6RoI5
nytQlvN59f4naPzxwe8BdAF2pa4s6ZscNLELLJKlJJbSYP4b/5sxhJsMqjnVnxsmQzAR3RETFcFR
Kt+wg+6IHJMQGm7Rff279FewHEf0hyXR4qFIjErgbNK+H2intCSMLrUoLmLoXio5Bdh9y2MHNgL3
Kc/wOUshahw8A51XKUlx1FAxx6W9396xfwlOvWxigzEHJ5gPaA6B4WLcjmK+frlOIB8CxqHC/k5v
noFg3DVx5rqxDz9DXURKWa/pNYEGIb9eFvccsnvd6g96qYe3lpceuyXl8mCpw1SDU9H+/gjyGyXS
OiAVYpN09/VgbRNYE53hmtOxvoQjrzSMF+B0uZOhNctmVH53IfpzvRO0wWbFKbm2UUPwLsT1MnmV
eW9/AHLPkwPqTnQqtu1aE2Sg8YYo73L0gJkyuScUq9YDLvf10K8zWsApKQ9J9t6UFhNl0u7uIhQI
mVb9sPNIwpukCP2JIEzgNHQY1w2SvZeMv6s0yY7PB1CQk3X/9oFn5tPYUBBDoW4mvJqB3D/ssQ1X
kmE/Jnp68iFxdgqTZc7/rlhGUmFqCWKUPjIbj8sEAzz2RFkZXq4cThV6kQc3fccp9CzfmVf8fqVB
inSTaEj0QJay1bs4qQYp8M9ctT24eFMX5wwLvK7ntUsiADwmR3AVfDP6IDacRR9jRNj3tJIk/uTJ
rfOy5OWH7dxyXyAS/VUGIw9HahG0k+SXYYlWIpmLRNAMkbEmZ3QqRfq+ighqs2Z1fotNF46dTSd6
dVyAJJA2VQqQw0PXJ4coFB6ppJbUy/7LbnpXjZjqHYZyeykQjjvTzO5TgWiDDveRHEG49PG+nydp
TrSFpAcJLFLHihxyilNyix7nyj1Ph/n+4yixTDRD/BWPCUvjDxPJRbo1qJX2c6MgYL+ub1QR3nTw
Q//cZDzdG9VfZtO/Dn7uED5gUfjwdSMRH5xr3NcIhu4TH5xdHKF58gCTPl0T+MTEZ0XngSzKAwoF
WAnmL6V9xLdYFlnPXmOfecAzwjjIYF02oaa4jJcSBomnIiGvzYWroxFIIuU9ZqABfowpP+PdnrOI
l1ayP0UWdu+ZxmtnkdMqr1/x6EpO4zH6vJxKoUkk/Rvj+4y1Fbo27ZEGPoOi1hbV2mduNuQQZVGb
2eaUHiUvvlx+WLr8M5E2At04E/Hg/Uppujt4c193RnVL5n3wbIM3EuSMCGfQ0JEeuXXZ0WSrZv0L
g8P/MnVbvayyJmoXYzxjsZDTRsmTrQlBeAAlSW60Bk7ty6/b7FY4Q+XlnjzDqp56O58FNapjAOOl
0FaZGTxT2PADzBuNJVf5erbIpkIQuxhG28f9Ok2yZoHZiPWgBzfuJgfbRJ97L590BbGQi4w2JJmP
8DhEenbebvVmrkB7AlkO3QxyZickTsQQkYYikHzSx+Greuv+HSiyC9lJNtvLET6ESMBwteQQet5S
1YqNGKgjH6ZMbbfcDFhkgjcADFw0WjC54+nJwNm5V9kzdJ96FlM7+kh8dZfRU2kHYHjhmvzfcVWz
nD5T1Mey/XXP+4HEXcL3b9rS05SBj9Cv5Mt31s5Oo9Le+CV+ky2fSvH6cTtYhP/4/gBTaDmpkMLb
PrmHqHnDvBTtoSZHA7EOHsAkkVKXI9bLhXhtmsRuqV991otX+VTsGfNRYMoj9V3ta0o7RPntxIqh
9SDWYw2CAC2wMz4I0p/p5LRPhvCyvTWKnt25YrUlgJSdTKLdy3ruepaKyLxpRuIzoXSew73fFnJd
nclQzn5EiMbu/J1gOSjj9g77ztGejyi2G1pWkULVnZUZKemkSWYetgacWBO9FCemqH+ZQRBpv86M
OcnCVjW+DFEIySMa2U4VjihEzlypRZZTmrKGDInvD/OlB5DnXMgalL76W/ZAiDPiDEhTuDiJsFia
EE8FD0fwiIkAU4aK2zIn69LlWBnxdcvSvlxbA21pevdoDjKwjxOPcloayW4dQd6qm7XuzSR7osS3
wlT/NR8kwFa1BemuJBPTIdDQh1ti0u2x5u28GWpIxeH12JAu8jYUFOlpqQBwfqJe6SBvH1WnHJTM
9lPKznktmZsW1PYbBUFhDk1z7FZSbgDavrj5QI5h2Kv8XXGjyrmE+rgwpAHcQzp5xMd3gZkha8+R
HuTyzI4W1jG3SycEjwWJugDCorThW6QQR8fX8tFhe5EmoKVP4TqOHsiEbLWDolkFlWSD+w47b6BK
+LJsK64yuBg0+9otkRVY9s0FYW6ezSv2wyye7Z+xKj3J+Z9pUVTSkBt2nZ9QBEPkWqdysgWG0p4+
1OXsXiLp+YwAyvrLy1DA62DbYH3HaHFmGt7sxv39jhIX7MD/3AN/ObFbkJWIcriOtkFYYLgdPWl3
V9CWrPtqDYU4GQGIE5o9zu/0wqpO5FkEsgbXU5q9U0aR9yNZbo7u8juonzjWywaJ1e+1FT8uVS65
ENJDDf1JcWvkh+D+5q/Ap+Zbd8Eq4J6W+NfdQYyER2RAhlKht//RzGkbMh7GJhTnvu4HqTrAimtz
IBUsCWCCATS6A7F1NPEVvcuMIjg8nf0Eo4b18ZEIBzGnfP1mjCM5zIshhqNWz/NIdI9E6KSQKry+
dusrWIOmFRWCBLXgiPFJpxVrQRJLWICOa0poeUL0+2BljYYDNpwyPKrpQFqOwaPr9P/5q6v94sHA
4tYqjfla2l7yvscPGKtEOoNkmhFkH4ychx29XwY7E7K+BqHbR5yo81DuCQdDP8NpEa+vNAAv01A1
lRI6x2HHvsVuRL7CZv9uzvJoHcVq51GCQVz4lwqjebAzernF+088aT9sVobQPifIrrwS9p6Cln+U
GuKdi7nQSrsTo7NR0un2jh7DyPxBXu6ZcDV+16oZVXFWpSlfMW1IxQTksB0QmFkFu0KLIrrUvJYL
JL6jYVlPhwi15nVLTHdQGCyuvvZXhsK27TX6GMS6FfXJKWQCzNbxJ5almnXRB2nEbgeu0OR/oGLB
ifkkpgv1TMeXstIvcWcmHMiodPqzt1RrtWflqEtm4ZOMGt9GglfrAJeKim2jmG1q7Gn7JDJLw2cM
CUFezXVuuRsnQUu+lrfIJQb3LWoRbsESIDrvvvEuNx4IZqA5ZfxU5YE1mDsdoN3rDItJQKD6iQFf
sKnRZYiXPfDBzZYIsw5CrKM9BAdDiVB+QEaNbaGZg/MftJFyUi/Jo6ifPtZyndA7r8QcMu6whUri
Pjhwk/lja146V14m/jWGAN8r6I9zA9doEGPuLd3QqsNM7OrxIlSO2EQwi0ItFPFctO/iUMOsYI+U
hJBNAns2PMhCKma9CIg6RXDSqoJ5Mufci2YHf8FlUrgrdjkNUpikh0kh7d8JSH8907Qu0WQrRApX
3fDIHxN97uBcXXs05adiJJg0jolcqCEPo9rrYAgBd9durfxiYwtYI1F7gX1xfB/P9+VoINTiXSY2
BTsaKQkQF6sSxQ9h2fPpyF58m3vyAnIorbzSTlu4Qd8zJb6ZQAjSHuZuMaJGWNNK8Icd7auCQkVY
a0FAaEO2LrkNg58KopWVml/GJZfPESUn6jJ9mZ6L069SbMutYNsgfRNLNDbYk0ghan+77x571eP6
hFGMDNniHZM9MKgNFi0SCObtLeiaQYkmCwd7zi5tMWx4HAhE11mzIj0nn/1qQHj70uF+le+lKPN4
CfL8bxmoA6j2jUTxGiiDY1kCxr+8lqc1+xx7n10b8QekBOIcUEL6a/3l4RWSxTzWKLwtva3mtlqT
3gNyf0VIIllzeg9ObtOMye+iNd+LpfICShl+dCLks4nBG1etwth1Qz0cwHPeegjozRoxF3iUqSUE
vYh4nIb40UFP1tijmrO3wDw8Lb+mLVIInSL6f051eYOalLYiTFx55B79AhHcH39AIpNFFDaXgYoq
m+sk18y5d/CYTe2jhBuJNAvmJ59uA5ge7aX18/uZH1SOzm0s7okS0E15mU36s6qSHKKlFAzb0qxz
IqtSqF0tUbPydK9oYV+3GuidgOre2F3TF9h57Vwvks8zaGP+a64+GS4I+cOzPnwLDqkKHQ973Uxw
pKLzyyNQWkhxrO28P2q7qQP1vJZBGd6kaO6RmFCC5SLkt1occeYb/KCKnfXUxRuBiz5BtY6Ejw+O
c1Z5ztpnsFjPmpzpK77Mooz4RmiVb2gse3ennbFQctH1vXMz7LLX/b4ve0eEMQ+WegW4PkcbW/y3
JtOnYftAHO8gD17EaQnb/GPnkylBw39cyGQqRlOGqmPocMw38U7MLCXtfmZBh3dpPeJgsvBSKX4Y
WiwZZhwHwNzT7lR6L1rl/+Zcv6NDJqwLpeU2J35MiKJfnYyi0g213+hbaUO1Fop94iuSjIo+Y5Qr
QjXH7mC97qqe/pwEQTNoY7PaXxCWTRqFnrpuQKqG8eENDgEhxsu26/lvKdOlLE/Az0xhuyMduBd7
oqz98doFU6LqKClgrK8uqPjrlrcl8teMRMWed1QAHa97NQzcM6G1ESj3teGE1Fe37IcgQG8/cMOV
Re7qihYy5jtzPatIS6v/KvyIlIoFr4jBYszquUPtGaHMcSdIWWkt5wMEbeIwSKGADuZssxk2RySu
R3STXSOjPRNMjJYFB/TVnaQrFABGnl0ycS8hFYHRcP77eyWiDqC0X+HryB5vw1UXOgJ0YxgeqS2T
DPUXM5Ijz5xiysCfYZjM2CGyWGKjG+av0BWstiLQ2tzvNUf5E8ITObZcq2zEyjR0Ql3FN/gpqR9Q
78zt22GlTA+6QGlDcJN/qhi2LTBmFJmM2ZLlYN6mP/uyYFsmKL6JH7NcWALP7jFldxTntGbnn7Bi
EqaQ0idkU2cuR81nirew0s/jMPINevBTxdd3eTULpT6dskGov4uotWRIxxiorJdMOR3oKwJEm3DH
DiSrBmPQpgfac5X3TU9CDFKxC9dsa3MYFxNmnByHr3KCfjeVWz4a5mwgluSZM+AAF7jNFgfndZ93
WnMX3keeFqP1sTkjZ59P7khgfnyHXh7fe1vzfe6wQ91ZjU1DphFKf91yzJOlWSF3WU30erStcmRN
wKZho1wuykrS14k0uTn8la81zSk+IKMA8cryXgJctGv/6Cl5iAS7EargBRtr41T2WNMnkqO6MfG1
HeRglPP1wkkjC4ZubNim1ydQ5mgTejdIfyTCCdRGIuJbEBfCay+7ohFjiE+AaP0qZFBvfxuXPjjD
Tw3YE7j6yj8NLPc/AUST+PQC7YvVyBYEUQ3sBUgU1XRTxXBnc+OuN5rtFiGAiXukqvP4/SAJdNK4
LAkaagmkeLlFGRZIUPLAh9GBe8urE9KnjvkFcaIE7s070An8WhcRDS2Yv7snF0fkwf7/GtEY3Pli
54xJ6ABnEbSYSbKoqr5vZA/BKSAl6QZQR8dNFdRASEkiy7/7h4ES0f0PMGxoLoyqstZ/0eU4YNIC
HQmCx+SyYxYVW2+P/+xj4vUAwDGjOwin718jwrTAg0echoxANpbrdRyeDdTa/UkchAbjNW4pEGnD
P/uqFBDv4mB8Mtn7XJlf6XC0pQ6g75CyDolx5o4e548sFgN9x5U5y01AnBSGDnblTMzoaP5GZjEB
wtnHT6/oqRf5XUee3iITgclWjbXRiDA/DvMWCwlwSsPSOmQWn1EdlPPtFhWTPVnRe7+HQ0EQfcq5
3zcWxnomeZQEoeZ07KUCGhXRazLNPFJAs5l0PzU/FV+qT3glgHzoJ+sYeV3ocaAcb9mwvAmlYIFv
z7hYZnQ8t9JNliNujV/3rsoSE1+Gb+p7R6nLXoNuJ0IIJfqPBHPFLG32V235NJjZB6fn5oZJ7qnA
PtHnfo9Put0YKcPzCICxIXFA+jp8gXE68Nb+jiFwa4hJ2yuOXQ045Zp7NL1V85rJ2EX1x7SWRYM8
Wup+6SnL34jE3eyIs4hPcUj85dhyke8eG18LwRfq+5AKRhW4w6ATAEyVoGUvUXQ6Pmkp6alYi3OO
KXmiacextp3TDjsx9Ms2iCUrTu25M5+sZWsXvwB3lB6x4d4ZXSpj61qtZXBHyDxFuYL3yvZE8PIw
dl4403y54fmrqy9ZJbJcobBr0X6Gdz2R11e69E2HNVwoiQmjcDBfmZcNxXYtJInR4NCEwXNVq2ss
Fh4CjfXGNsSEizCzipxV85n3E4wA1BmEijSJ7upzRI4x5ya4e9BuT6QVtAwWhOBZ1BsDuz4acrvJ
mAVpafo+QBiaDG0Jk7Jz72nd5Tjb93V5IuaWHnCw0pHvFB8x6j4xeZ8DTqlpcw/TDgeL38rhrIAl
tLxruZl3z/PcJaKf4F1Dlxc9h1ENeEiRLSGJC5Gf8k0g9JJd/2zVwkPCFbE1JZXuiwgiQ3KXXTba
uKWqUeItn1v+zx4aeUHMxxrKnFndY1O1cDf0DB8jwGYLOhM8U+zsuRUxCkArB8tbM7SDa4JNaOqH
ipc7M3SiUP6+pSiPErhL/f0z1VAgMf7SE89OsjuTGBXvkxwCbnq5ncJ/pkQbO97nTINRHRF50ChW
e/AZpANjkiUued72mxtEtsS1mJfgT4mPma5RMMF17CkyrlnnwTxs42wpraNOrxpopslF9NFJOz8N
7tAkzxtN8TJlziacVNXJfvb6ngUSplMH5W+ibnSJyOb7pKshB1ToBSQmt61kNzz1A3iL+Nu48bvt
GJ1y3/fPff49H82JO5KYgL5DK8ZTk3RR6QmzS5UUBsbzCSuxXs2WDFweHtvuDg2VjXcia1xpuzH0
CMPOXNcmGHIhJOHKU/jYYr8FCRyGKFZNz1+1HXNlJhjIVMYtIIptaZXyWwgg97uXHoEYERI6KByL
cpm4aWZhaUU1QlMQ9xc02dzHAN59uX37nA2MMano6sOp56nHNSPryEjqERzDS2emFFatDWehhyNe
JbgFSFj5Hvgr9ckUuold7JSPv8fN2lInmSpOozxIiJsZQtjfnE32mnmS+acOEMNkWkEaBQ4zhXn7
jlbY5tQivyi6jyyGKmIweDR5tiXI3s4P4xdL1+m1qsF46fnBC1saUEq08JiBfDJj25/+tcg8A5Lr
nxCk3OxvWjw3Z7SZRKoL0mp0eI12/YP8tcG6p6PESajXquBTmwKNUesTRWEOI/ZcuJGc1nZeDJ5e
NgOp4H0OEvJoDbmZch97z/zUXf3fiEoEISDDf/hEkgL72meAGHScjwR9kSgHWLIwFHVMOk5a1LIF
DQw4qh2tw8/QcAIB9dI3ZQnHC7NQb+BKiaF8xNQ9YHavik5IT7maHo8/vcWgrHp/9d7oaiPjJgGk
WduPzh2von6mIUKnS0ll41fDjQo7Km6mTwNk9voUH1aKgw8X9a0i3PAqxOFDAJiQYAjbTmNinln7
BdPNvZxNEfx34qu6Bu5jWzuhN5y+lmnJqdN7E1BJInlMFws5GBIR4wAMafUUNkA3ajyeOkl4a8jE
cxjDDi7ZPpgtYM9vB6Vz1XIf6rJIC3FEsKo7br69XIDPNXLgJiMGv+lL+SSHtnTxnV1+rpDiSiYk
z9dxsx6CeIiIvvvZwue20pwY5c1tFCQAoUHK6jLHxOW7egjAAjek7zNzOqVOQy6j9zyRfEmf2oXl
bRLJpLtI6QHJp/HdA1NOoP3ErVAjzPdC+yqIVyTcTt4nLiCrTLfSh0pUUd1MP/Wa/hyzkbAwQQSI
wnyo4wZXSwXJ6T+DPZx+o4YBk0JHHgm7dCs3EGF8XLJoktJ9z8XE6mSlDylHeNxnHMZhHP9xTmRB
OjvSBC5ldt6rzw8oZVCkohz8tb3KYe7ccjG7EixXLcKSQVZPcIjuRcIYUOgBkPjpO6RGuG+udEi8
CctJmZxMT3asMEc44LTYu9cybsJnPU6KgNfF862JIJX8h+0eWTifX5Egf5Caa3OUwdQ/3Z5YUBTX
j0UM8wP3K8722QY45A5PAXasPn2PJHHNDGL81dWVsoxTIqr9i6H8OnD1W6VvwWGBJ9zYnw1ecQEv
6tRGBEXNyp9gghuBC74XUjZJoxKyBi46Rbz8Fnwa8RJroSr7L9S9QK2J0i6c/uvrtIIXzEWgk5GA
Llddgy1rTU8zZ48tdKsgxuQKvtkPYvcN+iIwhwwsoQ6cSQws1ZKzEhy+Dml/HtW5gTjGWaDahlfF
JTgjU0IC2txYYIKTx1M+Pw1F68v9P05ilEJgneOEgUfeP7Puo/b7G+UkAZuUR/ewB7UFXjV9NWf9
wbDt0+h2jHRNMFMr5z1L35+/SqroD3ovQG+l8o3onUlbXs549K3p/OAS3GRN6GdWxPwUyXY+QFxi
4edU76rFoqvHDNPQZprX9kMMwOdczOWeM/Ge1JBfbtJAU6SYAPCkFM+2pcUjsXxdquZc+zDZy5ql
nAcqkkgM9N5owTwNXTi9aek09hIEeIqi7Uc/Olv7uhSNM2ndF4rlDTmrjb4eeG8PQURfFfefC49g
x8FwP094W5xSaHwhUNCpp5tTyifPDvXGya8onxZZ8URC9Xqv/ZyElVgMWk5Fbkf3+oI40iL2iqdk
pflBRZMYLl7zY+rlceoMJwbooZkGshdTNiqNzbu3PbPzP0YnOInEXaun//oZmV5clKWq1LxhSO0F
0ygbbJcq8sWl9fvOfOln51SLJuRmwLZp3PH4KGZgf+cWno1pw8AsNwd4iOawhjlVieEJ5sgJNnFi
jtnw7p+nBf6SA75kYyDeBdE78D7VReOPi3UC2G8ROCibbWRg3xve/Z5Oc/G+/vFsHnmhcsYE6KDa
z3YUF1mipv57bYv2a+OVv6R6d+s3SmCZxbIBe7FN7M/DmtubkU853zKuaYyCEoqoNRG18p2DjeP1
K9Cj4LRiuGBBPF5JTcnYam7sc8jWBPIpWpcpB77IJxKTFSVXWVQ6bo+I93raIZdpEqY+kfUxTGMK
fBoU0OM83I7LBSjhCD0FrGP4WhX6X3nmLjwboYJsZf4uK00Rf2EYnjQl+EuInvdTpeF3wCygSgr+
4WkZMWkNDsRONOhDPDQYXoYI72FcZwP79W1018Ea947LLHLOYDDZDvXk2wfhaNEDb7zQu0hnO4S/
kU0g9X7pk5nrog/RFWWrF0syDQjrL0Ch7QS4tWo8Bc58t5wJ4b5OS4yh0y3Ur8By+aJyfz+NNSTH
gPGPtuSQWsP2XikRO2X8GPupfMTAJkuWApvcAnLYu2wcwrTRKFu3QmpQvtkq1+wqIfXkXJUVZlZZ
Q3XsmvZryflVIazIldoWNDzrIlYC9gv1WthqyVb40zRKyuVO6SrReLbE/xd7pUgIHMRn0q77j6Kn
qwcsQ5uAV1TZnLenszFmX6UK2s6AcRwd5vCDzRxnCw8k+AThDxaOZwd4NSoshU9zEQgJ2EuxUw4n
3XdAj+ALpcSor+r4uQPknAfEen5k38Zu1g6511BfMuD8L1bpUcCtaqvjTt4I4A8Wd9clUYX566eE
6mM2vffmztpLPnuapHl1Mh3p81X8PoHNLuPUzC92nyhCpiZTcmzafRsxKhzxi1vaMLHlCUfJllts
cxqjM7FGjJijAYkM+zdkIKn7by1h+4TZ68t5JT5jpu/ugOg1mXyQ/CziDuf9I2KevOF5BFHBV/oY
tinAm/q4/jLVKKSHBc7ORxBYbrvCW5EIPqhy6HtyJLH/jB1QI8iXGJOnK0x5BJR4MpLr0k01gUAF
tZsrzVdHzliF56zyMpPjd2pxNjooaB2RXVjC0Yjy63rOv6VEju0eLGEuRcyDOaXzLGnDuOlLC6Vf
0tEazS9x7SlYEsDwjrST+GfF7zYzGxCYSZ0urmAoViaz6GcHY5ZWl4/BP4y6VYnub0QwReyfkhoh
zwD8jl/fgMRKvsmPgin8X++X8FwPj/zV4UZMG+B2s0RO9e5v+T/z+nq5jrIULytxBRGfAMc5BfdW
3mR6YWe8cgaDD93xP/JUCi6P9SKI2nLloZEeeV3BMTEBtZ49pz4V96m6Jc1+D4FN8CJ2rBl+R46/
QNfF7EjUyYWzH37WdRIrRSxB5SBxmY5Ty/ASxMuM+zC13BJDpV9zsH3OfGSrmso4k1+dAZX2zR5A
FYuYA9zPxVN5vFU5qvthOH9LspcqNHQs80SJxqsUDul9fLirmqT/djPAE1lA3lLKaZo1rh/pqExc
5iHtKKBLbnc68Rv7ajqeJRKDwERD34zfvj29bzpPuFKeH5b5VW8tSe+ARLRhOfvStqLbSQ0nA1Nq
3sRFvGdywXgbTfdjl5Fc+Wa11ZhvpLVwKPRfLwtAI4JJq6NVoItQ7Fuhm00fJ3KTsSx0mwcZ0Ls1
Fdj0iJtzHG+s8JcFnwB7FJMsQVaY3Th7o+v95FKdNDe8gdZa+NORXJGmX/N7J/Owsb0pcqu7VKoO
fm0VkJ3PiKO6hqCzuTwhRL8qxKnvCdx7g4NQw4/a0Z3wWpIgde5wztJugA5LOjn+ImoUTfciSL8x
i93bN8LArH4IWmZHzXCyh/scFmseC4aR3b2B8N1v+3dcqh7ENp5fnzGFS91vd3WxdgSM+RWyR3JR
9hyGVW7qaFidffTTk/vhku0+jBLUxlWtEdBOzIXiorZQprVknR6EYXwvgjoAGxDjHxF5hXYfZtng
KtWTjLhETOuD3Wt0h7wvCVaUd7MtVGgHRKij6EkqHFZTehOAoTjhgGLfhXgnsE43Bavyl3KGs16s
Fsc6oFRQqyLkJhNMuzIprOEppnK3GN/ig5ZyuhenUxrCOyPIfuK8aWjZ3m3ao3RklXXNMqDg0CmM
Nr+ySFQTbA+kiTdKIgPrl7PM5T5SyPOEfdm81w30AOrzByOmr2vyEBnft0U5S5atQ1Oc3YSKUNCw
iQ3hNX4r7eIKHik+QyNkPM9Itw8Z1DHbssYp8vtHOMYRDaBi2l3ObQgZvF0ssYM9+gurzWmpCaP8
upYNpRUirXIVezPG+IwVJuRpl/7gTs20jcHG2nUg8H2y4/89NYyrM76zmiRuYwBMqxl4awh1Wk0h
qu9GRa50Irhbm8LELa7cVp12paEVBjZgifr619sSFYjSmK0Nm1KDBPlWeCqEiDHfKygizHiykBOu
iZuvDnUtcXJzIxZzhu3DARwMjg8PhP2J0xfltwnsIn+9Fm3zo6x4Uir/veK/7YxPfBxIRti3uvcd
O7ZizhZUGiqwOVlVm7w6Kki+csYN4OnDJei4dWqTFGys3dg62dki9wzW5KVNvajhITUVUwPTMiEs
eYDlAsnb96lwQPtylTO2cZ+uaH7N8OX4lZ851jYjqx1v7M0LLjroMzBbMoZbB4eL3GwXStsDQ8r5
My1d3NUcStO+wtfnOp0ntVt+x73GHUIp4q8fVuEUmWF7XaEUz5peVxzyh+PrsBqtyPtEa9MbH5LT
IOKlGQhk8fAKAR9XUWGgUwH6Wh0bazs63PWmTqpKSOrr9hHPigLSpVwPg9Qj1YLQWiGYuoLbD1yt
UinS0n+nYlU+3fxVkfyqSL1EQnMIy2kyJYfVskx5t6Ul7IWTfS5Ujv2fgfBg2TvaZqDuaeFqfkN4
0GjYpTk8eDMsYTlENHmLWhHW3pWe3wDEwyCFcYPLN6/NWHuP6KCC1zK/xeItBD9VIfJA0GnnyBcj
aSOQxcsfxGoYdkT6ssj/cKvNYtqveDuDPE1AvxssrFzaU9rPeq5AyuyMu32Q1kjJpC4HAZcjp4XZ
DxuukeeFWfiaJX5/OTBf4XDe9YHr0n1G2YJSQcraF8uUdadbtKXxKy8N1dIADpXHyl1S0RSdP6Qc
5HAEA7TwWFooPpszspSMoNwOvHjAfUyENYnhgbNdWXEdBE8ESKd8VKksC4DzE3FwJF41PZAwjbtf
PLpp7n8kvpnI7PYaF8OxeFGqucjS6VY+wexpdnozHXI8nlV58QI/aeAlowC3YuqzFIRBBGmRq7Gs
oCDSObkXf+uNSzAyL4rr8jR5jzda2lqfE/qleyT5n5O1n1xRuyH2fFscs8/BuLxjFBJuFpoGJvq/
2GGriRl0DeC1/KlNNhpRLkfzU8JEPynkQAUOTw6RW9Fjgj1TtGZOGbM1RmjWLNYv2wnaTmH3N5Gc
hpd79ttsYMwLYTiHNOGgqBUmPlE8vB1DoWcAKizLHp6CfWcRG5oUWC9f2a8b4UvK1/OkfUtw+lwt
yFbLfJCoTi4mfc/hOqJEuHZO+IB5EOJ5l+smPUkCd+Yz7TPHrELra3HAP2BZLEcnFNXy0jZWSL7x
KC/9I8UZuvK8KzgF0uLM6OygQj8e5U+m1kzsvDnBJkpTOacWYXRNPd17G6324pPhdnQ3Hzehrz9P
zP1sYShxGTNMxZwqCmLlHsBSBpsCXD4YzUsu16gSaXPq1SeuHDAVQXv/fT76Sn33AWx69zcFYaRA
YmVhQOWcf6PwCp7noi7Jnr9Hpcj34Jo/JL3k0y82s+KnmdEggh5FcymygExwG+Z3hzKak28ctv6M
9wuSMv+u+sgOak4kV9hNMKOrba0ukk3Egz9wXzgeDkBzBOKhxEudRuO6a7/4lMJzkXsE9e2rORow
7MSP0tjGryhRAKQw7qjffUnC/kMlsVTYxi0+G+guv+bOCDrHP8QoQu/m3csANYlMJ45vJtDuu+ha
opzEr305TLk1EKqUIVHWc6e18ZV14FxPufoD20+jEU07jE7vQ7B6E7DaP6tx156Mhg1ll0RIdBDn
jDOIGnlHc7JOM3fOh3KsPU8AZnxBmYHmdNgzDH86N0cyI5oPN0zwkc1foVomP4JQ7kTGwDnMCHbu
11Zd4Sy1vSLv6FDCAzdfkMyPY/yO+hfW1FwlZQuHV1rS/0HHFa95Lxlf6bIxE0tzMzbnosKvT/yc
iONpqddctuIB4gLL6ejgWEHIiHagu/wJHTY6ukmaZtb6pS4rgRfcYLdmlKgoUhNDt5TEHG9bowms
faXxtiia+JZ+cqQ0/veo6GfCuhCoLGOYr9GGkHETdSw9LvcR1Zv6u6R1BoiqWyhVkDtD0m+sq9Zl
/JpEVGwKIYLLGBHVHGaeDJvOOQ6b9SZ/LcS4lAYLAkP65Eky4RUyoKzEN+o8Wb9v9sT2ZaeowiCN
XpjV+ufIyOkis0EdTw79em1UGKWS9z2+kLa3fhJBLPR+vjS0Fn4a7qZJSPtZVTvtVO9OrJFEI4Vi
QOkZR87/pRmrBUqNnmK2BvhbjyStGEivC84qTEpjPclH8HmoLD1n8sjzpVWewr2AdTSqzNNgbxrA
W+LYTehCtduCYwZdrDEmuSa98j5/zMaJ2+CxDwc4TKR3m0W5DOMlfG9UFHIOzx7ZngykSwoZIiiU
FGBBp1BkW1l2DEki0OxIPace1nKh55EeKCqrfWu+3D/7U7YSdHCUR7Ei+BOVt2tBEU+OdHRVw6Ul
HhQ/lP48moBMEJNrb5+NRNp8s23htdTHg6/HIuBXoNg0w/3Viquvl+hYIs+R+S+pAKTJN6klU3T8
ENhYqpzZCybZNvem3DT3n2A0gEM1gmnyLAtOvdgOMr8mAxoinD51WVmhjV7Ga8PHceDdnP56r0Yv
HV0yon2bLUm952U+9zxM5MMlRvIJcHTli1LFNGbvzPNJhuRj59yPRSyc8qs5kqi5adncPVo5FOiL
UuF2Ron8VCE3BxWHyEZ0DPAJPu0hmhnw7u9PLWdkmHc19qznUEDguK8n/p5OwvvjGmx0urzKCo6u
0djzXE8RtBWfIlz6i7SzvJ+jR1Gh/pk0bBB2mmUGiR/JATfDpERLy+VFdhIDRMKgplV+o7+KdbDE
zZs0BU5++uVCUIFOx6pG022D1qBJsbBbxUuZvtlw2GN0ezcgDyyBos4kq7yjYAZggC8V4ZAQ0AHZ
mhm7ew9r5Kl13rN5DB/hC9QlWhBXz75UIC5I0bQymYatxNCtOZdRqn4FbaHgRlhXpb4YvHduvrcf
cFv8wB51Kj/gh8glBuzP7AyVhNzwb4usIHRX8gJh9vbltrgzORCItuET0rSqg/OtwyH2WCKeTwnI
4ehZd2CAwMpSkk9oCTUmAKkUYqPp/Lxq1ZqsnxfauMHhYXG74Sj903bsxTHWx2bJPDDrWsd2tmLR
HAR14bbrpzno/hdByG9VENGnqnGDMyERP2N0JkSab+++sM9vDO8MRVZIX16CQP2P8y5gzouMcHC/
JljTtvOJdS1Xm7jcB8bDTyEwxWiCxTI4t/Avnq+KZKWDCgn2ny/XiHoyMPJLtGBF+B2g7AL3D3m2
sEG8WjRbGPU8fBL82WyGF8G8MG3qIgfuwQoZ+tbmA/PPTMRFqGmzNTZtIQvnGL5EliLEy+tVjhPu
kwo+w4CsMiYNHBLctLWVmF1sRbvUFOKElHJ3+ULgtz3ShNFbJ2Zm+VAosv7nB4tANoORzSlc5btp
CG+HWYC1Z8pjKf/9UTYXLrdVrT+AunJjsEjgtqtwAXlZUjUJYHEim7fRz8cGNFwo8oaAeiNsZpwk
Yaf/DS1yRczNuESWE+yBmuiSbIf2afDrQxL8CqXzkZRYc6CZJjoipxKP7Bc/w7UBj5Qp7XjWHGhD
pQM0lGnkgebmDjijHaVymuAvNulXR5nXWxEK0ejuheh4N3l8WowxJrtMVVRCYJCeBSb+IbYml1q4
bbhkgfRR5w7Niw+o/6lxCfp7dBUAHqqsfGzsWxDNEofnFdegs993ARvUuHJp2EL8TuYri6XwwqUv
ZHbFUf87ImLeyV2NgkdDWw0MKZU1CP0v7oLZQ14nbFtip0oK7bCl7tiADhciLyNanPgr41Egbzxe
qspN1rHAg4REqUk3J2Nvg05fUOY3ZPOdiPrYokHvgnFekJKg9LQA1IKSGn5Czn9LC3eTnfE/pSq1
VZhxhrxyX8QCxoySZAdtS6z5dz6pOEW8zbUFeuF6qab1IZ41ZFYxQbWoqgfTy1OYUphyxGF14BX9
JS8b7y4GngxUGtx8QzUH5S4NK2W5MHYNA6oOaCuEdFhLQ3KyyW5sR54KuJcyv344pC9yiruLV0pP
p2XN3vqbLuMHhi2vKl6mr57CRd/nMBY1lF6edWRAA2tguOeL2KSK0hJhsq7v563AY/wsclmeGb7T
sCf0qU6RdTZh7ygh+A/q5U5bQzH2mnvnKJz//Klz+nsqTq9jTGIuLpDNA91KzrR0KkQQPlb0bDUs
GIltRag5unTPkpioPLSIl5GT6x6z12UdclDVwwUnrmrgBIeLGsjBFDnhDTYj2OnCUF7jzB5ZeyDc
jfaiKkssh+gTFr3ilb3IAk1dLch+MohMY6v93VgMf/i+5mnjBgh0PqqaeI9Yu7YoKRwVciHf/692
QNWZwhUXMRCrqYYPh0hHho+/pYU2vXUjdVA8a3p8GOy42kh4CWBF66kzA1bT8aUpq854oGamm2IW
lpDeiYBA859CAawK2ByaAmWupdMD6x8Y2yTUJ6G8+lRpNUwkQBM0R997U8OioxpcbVPc13VelXp8
Dhv0Z2Pcn7tjD7AN+wVZ/1fUDpTi/n2Cp2ccQb06heh7qoa5VOnbTW2slh8chAb54z54rnWk3uB/
WEVbLq3vOsphffNwZ4/iuIhqA72QfeUeXVAyPiMHB1iPsXVETrmNI5Ko51iSg7b/rXtTxIXmeLsY
7AiuOVAES0koS12aLFOeYaNlxhgiAVlInfEw1NYIWaszsqu3PVqaSmqkVGflvYc/4quNxYHOYSWa
53uZPEgn7BNjOyo4T4jVpF0vRyhuDro3zy1/Czcyv+4Hawu1jNxsD/UVKLMjggCwwJ+tLX0PqUx6
YhorizFyG0LhP47oMKPs/26sY06bbmjUg+aq7b4C3Hm19W2TCrfnPKHLQy1725+sQne/r7YgYGfh
AXsKKpLG7UfMvIsNjuHn8Kqygxzc6izzNBrsj/EZ8Y72vYgZQV0qbENsUmCB+/noYxpLxwExk/Wx
c8IBiY9+bB+BM0smz5N092qO69Yl6otdc1xHDL5VUdWSsan+JWXRpgQEOG0gIQQAcs1iNiRMSh5s
jluARMSI04eQx8Gj2oCnQMBQsWntaSLd8QMkvmUB46KlidpJlhpE4fXVSDN5lxGYoRlZR6fycyVt
E8JeGly+P3+DQf5RAQ4ih/CpCGq+izH9DVPI8+pTmJzAtkhxHsCKNwIg5VGaz1/heZkXI6F9R8m+
3pWXhPEv4gzr4O5ZOTYkf5/DrR7aGLGfneFj6QgmZHaJKmYtlsBuEGb/PYNxFnUMoZ1sbEi3qqjt
l+pxefImi4eydgTtJsPYJvUQBU71VA1Dq5+nayYmDfJusGRHvs/W2KmoWGE/qspi8XYTHljXa3RH
xddkS36n8vC21o1mjGibXyj5XeiBxwi+m20U5jzk7ojtEMaj+yRw5N1BVhb5t/fUduQM66Q6Pt1p
qkjszg7F/ezyBA4pQu/VwJCTx+jHnlAdUey6F1j+YsK3bzZd9WgJ8lOIJ3Ud50vupSBlLHDvLv+j
plRi3LPz8sURyNksmRSkENE8knpVMHnPlur4aVXHDwsRIGVCo74fzdBY08OlbeLBcF1rl338DxWp
TExtra/AR+OpfqgDUe24McOoYpQQp2MMJ898Kx+YDuJnvWapzNL0QTSQFUcUcvwmXSFVPpxgfdZs
GdRNWqaMylUu6M4Oy1kGReNuExR6U2V1Od967wz8nfG/NIpsG60zjQ94R/flUzaNaRvFyjAkCiNs
M9fxLwnd/cCROWUnvhM0AtKr/8Vq00jGaqxM0vTVeztJ2JVIwh6z9ihMvG7XURGL5LVCLWKfW68I
gWSxThopemcgfsFJNV6mB/QrFdX6PqiTGxMFY18+XhOEBCjF6AnUebR5u0J8kQFnYXxZGDokqu7i
MPQKfwdqtvF1zPRVN4AXHDaxi2QFS8YpZyLiVN439sNT2sWQUBfCwuAaanP0pbwyfr8PhzvdLTVp
IXFpNbRMJ5Wpsk6zBscOMbQBuNqAo2nq4sr7k+EvxJ7uSiuK18WWVViy122BJzUNzSpjdEOvGBpB
lIun6UcYVJhYsSaDCCH4cnCiM8sYPj274Ov7V/wFp5p3ioxbptS5RrZCjk/wCDI0nFCkaxySr8xU
0rNFOgcarMUsywRUdiWaFzOJA5+9QU4v7fcHP5cVUsYgsLeTiaa2uPm1nHvdauo7McqNZYD1ANFV
6djMFvLXdR7NUyTMB4diICi9TlIS2oNKEZNy5Xit0bTIeQCVGhKjTIW68Y9V1A/HiyDhNwt9tyMV
8BHJ/XqK8T/gnu3GtcSuxBteDXjGRrDjQry7K+3vrUnnbDNfo+mflc2IoRbBmVAf3O1v57pd+J6Q
y2ZtWj1vnBVOvaoorPhcM9ymfCtI20sVF6YkfyAAvY+yDzEcIKJRqU2kV8pbVOI6JLYDokUaFCUe
3Lr6q/ZxMl85iEBjaiRYPbpueFRmy+N9sBByBawTSkj4TFkL1+A7gD9OvASNBG6TI1rVXH2mxR71
k6XReW5eDgwEcrdVqoe02bF+0FBcsqyprxlnD+9Hv94tPfu32OMwQIbViH8eEyeb2e7QLv6KM3gX
xYmapcQkoSzer7Kkvgf/tKWIsX3IQsScNdoSy3Byw5hITdViMX5x9W7nfsJlmqKJbjkeIV1HrnOf
eYvp0IkPjA4mW+xvo7+umv4H46wFXEvy6b/pc0TXNrHZ0hyZEhac9lMEMi8iAqn4kSdxTq9H5et0
PDIUJzWd1mys0IuIYvZ0Xs3K8SA/1LOZujiPSjUVf1e0UN/t4j3rlt4EphPlZTJrYhCX4BPRSZ4T
ImBAmlPyeVQpnzOOKFGvdV/cpdO3Q2RxT89XDS6iI+iSLFmBE8wiDm/MCjVlSLFq/2NbhOFYs0lE
f0eeh+wGyjCiUZHyNNAiQPnar0dPsqtl8HbX9FJ3aqunc1TGHRFcHqTG9w54gsNSGjq9FMmyy6jb
N6gWiARZecAWbotYksoqeO0n8GffiDGhJi/yMC2BdO2H113K5TN5v3ly41mXsV8IvGXhz1B5wFrw
9yBbTJ+InKzR46XcLWBp61deTDqgBDd05LqI7MWKEDukF+CG6OLfN4+j3nkDRjKpoDx3OE4jt48K
ISDW2bHbPz2Y/z/Zco61i5lNyQ3G8pJHWiNYqRsUuW1Xo8fmN+oWVo50poolbrX35wT5ne146UWc
nF6sZhR4EBZyE0OBA2cT/WGSmR+yWlr5Tj5J3nd8nO+wJtHoaAJhSbNeEzNKfrDbDqDPrOwLaU6t
E1WpLJaKJSXFOvBwmOrsAVeodaNfJ1zOBR4Z3Fk0LunrjwXOxtCZY8FclyIGLHZzIY7WLXgHNiwH
EEpi/k1iJexPv/Z1QONyY2vVviekDaSfKhCsZECDXL0yMCu4lkYjqxuxU62wlc8txGltTR9+dG9F
Z7XuvR8J3NEqoD5L01lzRicbX5yTj50mbooZhDvrymGCTrFnv1V6doP1PmhPDHKcKsnV8DaRiCmn
+dyRV7DSduKX5yyqD3bBsWlRxJlWVIaboew+xfv8071WxtEr2u4h2G00SByagEf7qYtlyz1LsXdr
/cHBz5zyrE6wgEyh2HPLXSV87dr+gF0MlzhKgZ07nUVoYMhMEeDTR492ICkere/BxT8m3BLI1z6m
Kxq8VoKc0k2qSb3WM7v9K6Gipux4C3EXzeGNL2nJujC1Wm+gGghkyov1AHyE8FbBbOTb9f+HN0Wu
fs84ev00etwa++Acn93CHnmWrqj2paF4yTqA/es+ySK81HJl5AVZQdckdBhd4QJGMY8TD6DxKgU8
AOFibWVxX6l0vQPvk+6djGLOgoA25oMaF6aqzi+tQazIBNRzJ+dZUKL5/GtsPcNR7i008YCOlM1h
xuXzgaHDqJrLxR3aozWWbaiFIHCOgRQXOM+873RA8MCcok4o2thLnuQw0niSKSudeNFBTsMocdNR
Y9WLQsQoyJKSb78OJgN8/OtXbrxBpRXrrzlp3M1hJuQ70yfsibX5wg/Id8UJjxjvvKF9Y4ux/pJ8
KHZRSubNlJXcZWws9rxDxvB4k7/32EcPga0zqlbOYlH2ztvAHoDYrHKBclD74sb9dZpHkP+jKipX
BL54obYsSIWuo9AYQGS8YvD7q+SLL8aqZIXutMw6E+TC/y0gxDk2fsdjecUqnSWLC5nr17pR10QN
tOofnEutzya/gvS61zfThznbRB7YwfhrCtDlzRDBUGqnQpdZi3sbnRxLzZRn+E6kq/xj+9d0FLxE
5P/f4kKXcFIVvkVw/AghtMbnxZhlkC+jDfDVhaurvQfxeEO9VHg7Wb0RuXOVIZ3XRb6Ro3RILS/2
LTRdEI3fvu8po0lkCoTNyzZThnchYQpQVbibh39OHVqc850TsO8KsoIfEZWnWdbHGbDKoFy76/jT
ZoyHyy3PB2ccz8MUYDFmAr6xjkjzcdS8KPOo4iARyZzcy0d9ErHC5RfH5LoFTWeLdsr8XzqlODWU
qGQE6tb4OUBAAQrzwOis/wG5qcQbU8YLc2q/Mueui6/8on6hJ8bZzApqSDbZfpTk5jpYq301EKz3
I8veqmT8ks+qiFsThmzZqOybA08oSXT+lEBivzptABDP5f1FMy78/wi/ZMJpDh46nFyaxPukRcqe
HacphxeQksVPni1Wz+lutO05atH20xO+mxzkDA8ndwywClKkb9Do2f8jytk1Cigv+BiGyd4UslLw
jEZqaoCZq9+XyAI2UaRQCu0GnYrd3UzioZZVyCoHJYioeuUE4T40P57rlCpWdd4ceC2xl1VoGxiW
uwZWiLe+RnDVGLj4R3HbC7xqhMNmB8qGUgxtOhGfONvzegcIfH7+dXTva2faUV/HEnzA0HIOl/w7
OWBApQdUrBoQIxArg+7Y8vGxzTaJh1CZrAQxb6B2hM4mR5refiZ208x1ccS0qLU/IPzaYEQtYKTV
JFcTrczWwkxrP694KrILi1ge46I7BZOK+gfmHiGU0yAbZyD+pzIPVTQjvSwuUEoPrPHEWeIP2zYG
LlH/ZZq5nbJuCWOyW1GQpd6D01XQmOWg/KMV9TCeHdXTW1v+j6awUO9qig4h2AK4QuC5L+uT9vfj
X/qLrtDDrmj5CKsJSz5iL54dMhQHivbktMkj3/JxzWEVXa01v1xIIVU4pY8O50Tgy4GSdsFUc5ck
BUX4MqTO2c0x6vQcT2vrf+V6yzCqhEor5uXglwcgizE3/wmrDvCgr7kjPQ+NTctLJhaPI49UQB5p
jF07tTyj4aNA40DeBqX3gqbtw1mt3yocgNNEuz16M2UCAcZiu/EhrGgxUMzxLRYYJN0Tx3NiGs37
tlFNRETJ/uygYSwonpvLUlNeyRpmMDrjPs+ktmer99b6zLxv9bOV+sHZSl+s6RgrwlBr8HFf2AW9
iq28/jq1/oaU2Sh+It+AuWio7z5LNHlDMvpeLBC2+l8L4uggdllpmCj28xQAmFf3kRJULuWCJMM7
lKI2ZcqquEJGK6IwflydS8v0hDMSFpjJQPr1MV1VIaGWF+Mzb9PZ5eqA+oCPwtgEzNuqjFcOkhHA
maxTzxbz6QL76Hv1bqqr4eyS3YQItqdhBqfjcFsfdGfg6X8x8gjcGtfLAjvT8UJICneqgfXPr+Po
osOw0dmhV9MbcISqLVIhmJUEeteiBxmADhHybnrOFrRqiMJRyAlEeC7WEmvu3ZuJ5GWWwdoH1/r5
NyJslVXSR6crq4lWzaP0X8cbKRtb4eUVXgy0xgyBrEGbYAY/+COgYK4+w7V798aSfvywtLX+sz9s
T+64fNPSpAjRNfjX/0av6c/R/JRNJGT8Y775qlh73PiHkVgXyJCoTrzsmAGWM1Y8oh3s1xnqK9Gt
6h1FWBdDRiQtIEoGRsz+dkq5IkvIERDFTPUgWJTBza2hXPPjYDxPzfxg2OcnKpQTqQT9PulXeQW+
moFrnFDkxKvrQTJDc3PbMMl23luud4G9V5e5gdWANmSmMwFAJRWMlHYqaDL26+CexqzSafUIYoRR
XNz51KXQbgWudLNTvZxTf3gshPt6MyCMoe8bY6xdsMPobShEZdjZHE6qchUtAs+axCr+jmFR12sV
eiRUf8pvnjHZjzc5znhRruUm5iGTZWiApQs5lEXhMk501iwyEkqHa5crcrbI2hlKJfryvT4n8Msx
bneQyuhTuu2P5k8Vz+QU5rwAok91jgS4vn3PxMhsi58cncfMVTSPo8DN5T+jS4bMGt+IDmUlOj0m
CqhmR4C23OcTdnQbHblGt55og1r+Bt1W2jUG6RPTvo6nAZnhkg0ZZG2XHSLu7AK/Kln9u3wYVrv3
d9VcPCdQ8Z4D9S1uSzrKw+A9ttKGL9HdJtMGglJ9f3N2gsz25XnQyBZQdxvTYDr2HKvFwvN/9itO
OyoZWolrYIoid4zKc4X3oxm8GFwu42XdCR9OncOzkntZQWwkrL3NDlufHwHxIvvsGIeUbtduM4AE
VPFcNpnsuUBuclbWpAlHKJwFOaNFwCsu76ySW3gUIyVkva9IBO5H5ZRTpkpo7k4tWbJJ6AgRKl7y
vb+BHADpTatdnX/QBnCzd+LDpQL0Vt+FlMxDSCf/KOn8MxkX212FXLJybdsoQzQpKJYVmtjjdH3H
K7N2ljtH7JTDxC4fodAUEvfmypptHQzOvQ676OiVc4n1S4a1WhKfGYhP6BTn6XNq7SNRtoPJg/p1
W9/wFmF1jvmAN1n8xLGqbU8IECAQ7RG0R3cVGvDpBTmQADIfewvC7LqAnUW8Nku3KtaQSOvVbnf6
fmXHvCScdMLEzhg1fGlHBDuZfVk3WSEGpn/VgPNWLPx5nVFYpMtISdfh8lARfJzoDq+pctWIwZWV
34BSEZmX6ImcRI+3bXtTNAt7Gs1XStl7XLjUtbVTHi6e556ucvrZta5ulqgEJ80Yv3PihViiYVRv
8BlJZdMW8nCcoFJ+pr83j52pt3F1U88qxhYxAcxkMwTrfnavdfp1EvZXiL1TyfqN78zSu1SEpGsk
WmjLytr3207G47PEVUrByMdO3N4UePC/qzcKQoTU/79REhoOwWnadvKX3X1s/4q2qZQF8FizxprP
TUObg+xkIEtRD5qciDkLSa0DpHdPnuU5RmMD0ePO/RXsa8mD4xzo0uFEJ0Ta5B1QQpWF1F+P15S4
C5fTybPQUuLkj80bclgPhYpjAJUcc1uSoHfxScCEGpKxj+JGcYJMwazJK36Pm1Vz9f+65rcOy0tH
o1yJg69Xcm8PDxErjHGciINpYnd3dCfYefD9JGjmQc/NHz33HrENxyDL/W9ywOx+/dgZ01tnzpv5
qUrR0rKrtBPEi3thBXFFzBI3ffA4TKvm2hhsPgoya/RjqcrenT6AHu/izvdWpT+62aTF+WRoJUhr
eJaAYAdpozW2nZjjep1mmmNq4guxTu11qWnY/3l57YkCMtkN2ny7h925X1JHAtvY0BbLMFCUPLdb
YeFusmxmrkJlbr/HOF+OMRpnc4sFiv/pQM7jI5wxnd/K6BUEm78Dc5kXzCSsP0uSmvmHuTaeVnMD
ce2nNoSCvVdIpyTL5oP8IpLfTrxJp2gBhTMVkZTZyDe/R3Y1zd2bGMijkqar99QrElZicDYoqoVw
M+4oIA6oXPJ1M1Fqk91Xur/jukG1pyO0ZoEKXmtIVKTfk3U7sWbFReZIid6BTgRN7fGNhCG9jU6R
apCIwUEmFPQRPrm14wyOpnQpPWnIuQi9zRJY6myrNTOL0MbeiDRA6gulRV1xAMyTqMGX1MtWos2d
tMaQAreKXx2jhKrgvtcBc3kSqb7NcgxPpOvW65YGNsnsDHg8HrwowNex6zyRC2MytneLRbR4wpPL
R0tjDYC9RHo3Crobz2fOeKDYOPqizmU4CzAz7GnIdu2Ul8JCqxi1bnNbAzD2U9DyBYZ2igbxstoL
L3v9603BXgIobMRE4h2V7RUjXYkr1BEsdlxIgMYi8dzgCgeRtdcgSbqeHwpyqNzMhB0laQMHz8Sw
4fI5JozbWWqjchgU46VAk3LXpd0+PS/7qnjYQtNqYqb+57QmZksf0WiNto37nJKFNULloCYum58I
qPgGaw3xQGz9onKS0FSbJLpSICEgkMQORUufy73+5Xk8B2dCupX5LhnWpXLDCvUHtV2rAalTemyf
O4nVD6CR8mykoCX5TFdLtaVx7Y9UQ6Ae1zvBXTlMAqvIFXMuUgzbFqaU81ANKk8WBGzVXkR9JjRq
amGxYIvR9zaQup1x1C/qM6FQTeSGRsd63PYN6276jdIdg2CXzPyj5EH8KOR/SWDJUtLJe83JYSDM
8pr4N40sNR7rWtB86Bu79kZlpMm4bEx9PH3ZhliL+YOXJLTzsoHZVHVsweXDBICE/J7CTwEbusG/
UH385B05VFdqld9EOW9M4+5d2Cp1KIbcZiRbSyIlGl3byjC/2H6wCc0gXpDtPfNps8ngNG44PiSv
U3FQgvwPC48ClEBu4TXZh/3tTIpU31Al3HE8Ji4KFZ38CNuzANAyePzvZI2+WSiSSbS87BNP/I0j
ZQ1x6mrE3f1bPht6ffhCsveYW8PZGDt/uVXuUs2IKEMjm48EeBlE4a7PyLkhg4SPKa7j/PDU1IuC
A1PWYjhHm+zqPASYFQxcMmCNdAgg2N5wF9oMUTYMZAb1DZww2lFiOBeqFS3JyATbfECSEbXadJsj
k8jeZxu/fSkHedDjRgA0lQbMuI7VYtfd8jUlmRSRU4unA7eMlYh7dGxnysDhLSTuvNpv3Vy63IKo
NRMlFmUyEKVbye8lek0yyBTJbrmUgnR+nuQDSDFJqFAdsP8YYceOtgQwnxQa/P4lM0cHUbEASwN7
2LgMdLfOLvS552yo6lu5b9NoF9cluvYCK2qz8YFuiw/qVCmOnhFqMy7iEbWv2y9r+osDLojylnPi
lcJroI9hu25mq+4O8oT8o7LvFTXpKlBYu3dbmROB8EMdHiufOd1ZfIlYDFGoBiNt6pYVxO2f9hjO
oKX9Mq86hZgj29eu4YkZ41TOpbWlB6FvE7y0kmPsH2YM1Tza6p7HvR7tGMCBGs/1xXb1CcfdD4+X
vRznfiCFYUYFFNyl/kjdH5zfTYpvxsLAlf/dJa2v/qSBF3qNO0JNp3CSqwYM/x84ulFUgJTHUE66
7d8QwA1tFNtoKD+NKMrhZDcZq/OAF2rOJ7St5WBviaFqlhfmzm/4sK/QswS5GSA44Gloe63JwYyA
L77LwngD7zZtJ7Nw9Wx2QCv6yAFgQJl8UfRKusK0mN5MxoieAvk5Gb1KsA3O2juj0r/DeKdUMLTK
kav+x31i7TYDJmZlEtv4y3h068uDPV9tftBTjeb4YjtBySt5De47ZslKhAXOMhhRgitF1xEEtauO
9tko7QqO0DsV7JhbctZpqJIjQurw5lrd7rvLk0Qy649N3GpNfe6CsKs70GJTqf0v8VZGHQ8KVBFP
2GYuE4OfdNqvE1eaeJ89jTxhAQUDjX5UqnGs+t6888XqfIoNvgsqC1xmixvRG86jD/IGLrRQuN9U
fn+okqb8kmDiR22hbPb1DNysG8HXo/HrwgwGeeq2E+e4da9suRvDyMPx77ckQIomLYcGGbAUWRP0
wCs7f/OZDxNQJzoyukpabM9zPh0CuxHTwG7mymRztTfEBRgqEKCrOkQEdz4slqryKLv9kmIyLAn+
6C8WK10zQ4owoOKn+In0HxSoAzYFoddjUiPRCIbskjjRtCv6M81TN8I/PrRxCcpYX+iGNuuzGwp9
IeG7qauJ5ulDzw3W42hRy+0hN8AlncjhHolXp6JY5vdlZ0q4YMeGd4kEpyLyEYFMMsvWYfQZQyxE
qU+2Xcq8LcwjanacvbPUSCinMViuyOHCgle1YpGSCAOPVNmACMOnGHGATc9/bvii1AXe0VOu8e6i
6XJ+h6SfcKuHUgYg6RgfmmQb397PqGMr6KnlOfk9EJqRwLWUgTuSIvRf1oFGgIJr3Q2s5M6OT/H2
A6TiUlBEbka0uX6qvYaU8Fv8B7bL0goLpSKVC6sWow/NDNXOiJycVX+Bv7Bv2ec+77afD6ibWnEf
za9Q/5WKR8ci9osHaA8pdWSv/vPuiLZNp51YtUQNR5eoJhbc01KxMqiqUb/oTdSO7NsPxvBtezdd
GIuQvbZVS1MgtkH8OMVY1MbfSilNcV0PjPwgzUNiYmq3qzrtYsYw2FuKvZbvvJEGf908i6hOiaMv
cSFj6xxl7YIxx2ACzSQPKJSDzayEmy7fo0CWrBj5OhOWBamczVI4OQ1nmWnGEtFASMq6Mkr47bVp
tsiSrD3YUwrsDN9OSzz5iQpJXJ5rvrloVz7r9Sfnct8KE3TjJrsaEjtPxc8702VB2Tgulmd2+XCb
szwHS2aiATgo6vahvsUQ+1AOL1afAKpq9qmdMAgOF56qlMNgjIDpXIhkAWtQ+X5q8BllRLDe29s2
eN7w2bgSoM77imN9pd5Efj7fWdpKlrtBAfJT6H4CWWCH88AkCSAjLobLUG47X1UrhCFvd+y3XK9N
p4Ifh+4+7BBf4Wgjkp34JNhaB4pGAoJCetc7BncpcsVxvLPDR+o2twYjSf2uBle4AvzoPWHAltjf
c3JmgAZJTR58euCGIIsgzpXnybEerTMRV19l0NXw6qpXFVpBdRV4u72aCCs+J7IPHiqT6KW86d7a
sSS4/vu48wvgW07ZYht69dNunjMYOa9wS1gBe1rhaQpz8SDvlApZdeyVZhRD2+6DIVufX7Ht545+
KlCKXmlhtoAmF+2mVaSlhk0ApYxCDy4mxDm4V4SBnZbX/rgtXu8qXUuj2o4zcq60A27qCbdcHh+8
MKoyYNIRqdYP14Q9hOqFyZMFl3HPPq42dVSTOXHB3Gef0vtf9qKZnG5GYw+yPNOxR7++WINkDckC
+BamoVXfn1X2DQH/eFy1racyEZmRy7+PNk7rcwWY5HpBaEYejgMYoiVl8MJz1vMwzSgL1dCIzT+9
FqkNDO7hEYV0sgsAuSDLVMvox216SqYlG8RB25I8I3QF9EXbeJ2cM8Veh3l8++1/UBKhVjVz+CgW
fGHnZxyKTjNdov48GNWV1oykF1rKJiHYcq4abEKdlLqqUNJZWY3ib4otoxy5n1xdcUrKsSjk1mBZ
SLmqtq0pGP+jMChZq47yWc4Xx6lWrnXUFaJAn2QAMbjonh46YEltPmddKz48LopakuHKeAVM6pol
hIkFT/NxN1853dNkhJqAlwqtSO0KYE3DF9/sMzpGKdE0/rAtGK3VjQaFiTWNOwR4dB8aEZ6ZHuJa
B+VLfpnUoBtjcdODWK5+yawDjECvFBRaaMZqTwV+Ewi9n+uPPdi46qSmk0d1MlDnAjTGpKXQOwxy
ewzJqWogD8oZst/awmDNRFDGGPR4dasNf6yGjq8LFhgcGJasVLRXtjX22BAIw3zIhqAqL/ZWrKoD
ffp5CndBYpS1qvWBzAnJgWuBrSTGEDwcbYMp6wshme43sAAaR9clnChuz/j/y6A7XRQnA4KuufpO
NgQvulzlydQNCp1MaGsdVIHk9OZhLJkk6VUYS+MRLwofxfZle+Q6tF3k9r2Z5uHHzqcn9H2pyqLR
Rrch6XH5eTzg4WM4vZ5f+mNHMlee/222X7+T/KgPFpyEwNE6LJ8kCiht7MUxb1adygacH/VDEHR4
jS/oMVzriRT2rjfaOh+evGPXNAYG59hQlV7rziWIHbUY9yzW9FQRq2+yMhV0Qg74V74EDHtgW8t8
MJ6sLP48H8PWB/cbAQBEY8SRXTR4+b/WrmhQNxUKV5CoVMuvETyt6ZK710IPTrK476vkxT1vZ1YU
utdKp80BMfVqSoTwwlE1eTCICcE25S0jntIsHPpkG9827siR4COGMAdYrMyqSYgXTbnScyPdVeRh
0yF7j2Hs4SG5/CvsblspLS/ThN5sP8IEi6xTlhl6yFWxC2olQOAsjU0iYuFTvB7ubVjZI5nzGZh1
XhWYqwZhNnMK7HEKroGM/AarUOVIOY1/dPxXRVKoTjrw28ly8RWtOzYDspsp2g924FRQOIIWWHtm
rkIC8vsw/BO9npeL/Y+uy47M6wRr2YqRz5pDsRthGJn9NhC/1tK9w+nz+zffoXZHuzC1Ox7LQSXs
9dZ6HZW+i5nMVVH1O9712Ztzvhmcht6bbJ1MO27S5rwwkj7yDwFvx4FBMnOydBijZ68UQDuexyfk
g3cydCyK7FPg8pD2cCyFmUrpvRNq7OpzrSRyquuP7PwoPVWTiQ0mox+M9PlQTkXnMJWVsR34ye7m
JOiOVLNyZmcuE7DptvPAq5mTf9vl1ZbqRlQ2xDXlqAWAJ7fOMm0cgErogAr9/BB1a3uNmUMiGve9
bbcV5Z2asBgO3t6WxrMX5FCVoL2TioPqhR7271EYp2Mx5mv7Ps3eOMTsiAP/9MDL0JV7hs5C2W0F
/2MEpeJfp5LyDpXgTCGhTnqg2p/TJk4lKW5O5By+VIOCEIRtF7IUntBUPDZoXMs3OFtp2E4rqdZU
SFalGnvIixgpNCXY+0wL6VLlH895ytsrA9UOn/6dirb0e4UuV18W6RIaFj+yRFgnt983YDrcimNT
mb6O9jYBBfRdmKTAlsADeHmpPyOlhiJabuQdYkCQzQjfuBt/rA0JbylV2nzpUFqQzBUrdw1hEgd5
cmPG/8C39rqwikoXkiT/LC37AIvnDoHOqoKTojkeKpgQQZxh4mkj9awcOc7R/8EGz4UJnCR+Lp1b
8/E15NsStwWp92J5yMgv94sqCrqhafsk6iGwlCC/+0uWP/B9OWueVgdyCegieii5DTQBeWerDn12
G2ccZaNCurjb/L5560nkPoXm7J3mXht2gdWB/NQUNl+j0nH57oGkk1ODWXqoXT78uJjPBg1DZI4G
RAteNKo4CARrzCr+yuKElLGECpcRguhsQ9G/QHsMHi9KlDnYRhkCxrJDAAy0CrDfohUrq0GNhlSZ
fipIF5ds5u/E28vMsxMqB/Rk7ceaQZBxDb8cG0LsMKSGNHrlCZjGDn2N6l0DwyU1suF6cIvaaxdi
scSkgBppdclbUOJ9JAPpy0Ms4Hid+9umPEKsM7DNIWdNPdYfpL30R20/E6EdOZbhS2a0u/TWPfkB
reEJAKq5eGGOCRE8QQr6gx6inpRz4nkRpTcBv9ckM7ULmsqOj/LwcyrKPv5rj9eU+dyT8XWLmozW
J7MQXYllv7BcfN04rPWsyrOk9hZ4qh3BdDMYE8oZC0Bt7EXwTtEFsybgBP4KlSH0GtnFo9ouEsD0
hMLYl7+DOut5ptqo0q/Mcs3z1P8xo/JD1O2LrCgGJfx4EolFwGtjURbpj0VFp6Ck8swzq9USORUQ
/wnwftgGnd+0hHZVew6fKOXAy3rd1JOrfhN1qdJFJXylog4kUAtd38EWZtqwEzI2UO4qulVgjZng
fj7szpDk48uzNyLKRkqQEYnyQ9M49T6lyjm6Nc6mYN6brrByOu+g7e5GrHvxykQ7WpitGUBxsXje
InfvcXlG2QPjnEd9bcGHh6HrDJTsVtlpI741GFFmqjViX46KDhEAw4ksa8XDShq3tBcIY9jLfm23
A0v8RHCauiTc31x+c0Vv6schDCm4HJ9Gcgzow89QAsym+eOPreH6nLyttzcWfIFtpp6Mtj6qO+aq
m407Qo8t68bOP0V49l5w5RB1GT1Niyi3Ewwjn9dBIt3bV9vVUnu0AdYOwu/vaTY+6gXp6PvnyihT
2rkgn+hpi0l2XwsXZyZvaKBgbLXWOBRwP7NTbcMdnrxrhLJVBp/gSI48FYk0DNsDH4gEGkjB1xa9
q1S2hKaBcWQctBwzi4hxBhC9bse5fs89FBL+nh1OP66IX1IYcKUknajut6RU0Z7Z3w6GZ9A0SpNu
o8mL2DKcS3xly+529rUbKYG9C1SYbBj3Whh3qq/8QYvcIoCr42mzyc/VvAtsbGQH0ibjW1z0doWr
3R1GX+b3UVu4tXn/Lw7eKgCijbXg1b+nzOOVrIVYtcHR2KbTfPHgTkR2lGsujxNl8dJIxQAW2wVr
IdMoixe0qq/9P3PskHIWHNQO0fiTYYkW1AemcKANTENf94pVKPHMB4wj4/79pbYXDdXSSkDWK9GI
eS5ilxkosla9Ff7+p4gdF/OfWSoSlJFEjaBN2ZhV5jnwG6yoRuSFoqNxy+rpu9P00pzQvhlllrCV
0nHZ14z84pqX10a7HIJOqw7Wh6Il6l29ZjF4PJ5NENZe0xNuLgppLArHoFQEIx/j6V7iy/p+saU+
14CV9f632LbFor5AvFNwB5g7FZSROeo8TtZJBwNVdB2e9IHXqw+3mv6IgDwYrB4kN4w1idkgBq7l
vZ5Phrvf4zuIKINJUd6ReZhwZ+972WIY2QoxOfHLNkgE1xtLxG4magbvNzInHytKi4ucTFYppTks
6An0DYleuhgVtoYmk+V61ID+r3/0y9hTBuG+oN9OVzv7pQjt720OaKgmywU+dGkHDo7M1XejVkKS
pfnqpEJCOrscdmMW1RMq7V62ZQ7292e2vc9/XoN1NQTkpo+NFGC5emIx9hTtsxWxEys9rQj8DINR
GLohoH1Sg3mqRn4ZmmVwKqTObV9dxZ6ff/K8vXQolkTsn3/hrSzSYEYUG8szBNIBh0hxGavs+r6t
aQqYd8xIzvjecDBhHVuaumY/sCRqftMMy24zjOIsuu5L3ufgcUUPJ3A4lbcuYRN21u4LypioHSRJ
kByp4yrysWTW7uBBwDj/vZ47mebRqyK/4HryvWncBpHrsn8C9kwis5I4P6GpPFVwlfQxoD+jvuyG
T/tc/hEcAknASggQSZXetwcIRLAfHqn9jj3BccfOcB+cgF2m4kTzhXapoAdbhrWZzZqGsLG5ZVh+
upntxJpmCIgtmNApQzoPlFObMv5fmlFg37v10bnAfJs7i6CeMYyMTXCWFowjXEicJ+PBOoHr+5R/
TAB9z9mZaIvP6THgajC4ifmfwgJrHgQC75l2YIs0DC8uydbI10g+w2wmmt0c9Ark392zJwaajt8m
bQaym1oPvNdJ99N1FmHiCWPAChAPwD5x0HBeiccupkC+l0hIY/MiPY2KmU23NwHyd9oVjoBu9ENf
B6FmW8wY4cAK4CRwut6H5A3LVxZe9hq7hKdFQLHYn8kPwyJjVdBwcAmIRnUgPgjwJkM6UJjy71Vf
9s9Cont4tjXCuFeGVfTW+KsGBYxG0pZdGjZFc3FxNbCXF6iGOLgPMra/ZdqOXrjNQnezqnSABmv3
0b6/QGO/ZSIV3vM7zl2Q7rfNhAeeaELyF8GBPUoWa/DBP1QIR7RkPKCCxFdYCbIDK1Y8O2OrWBpC
Tror6dklotpDCcX8k9Y6zi7VNrofqhRH/d02ZU04B3QxMWwEFj4Ay4p3C34QOPPzL23hQik2sC2B
EfQrtaCkD+sYnldTbtktbXQUztevy9SVlRpPAm9K/kr1ym3ob1i47Br/AaNahjWnwzAr1zuJ0Ktc
4OCcjgX3DmZ7LPu+5ftARl2u9mYmegPi9LnaTOMAlPTqLU85RwhC06SsaNj98kAfHBylg3oTNeAo
v40swToSN2QyFBIIyYmq3n6I4boyCuJi2CDatED697116ZSkaTejk1MX9jF8EMmdvLkXsPZ4HFnd
itA475DRZs3Gz7OXoHTBvSZAVfSNbrewfr/09NkIDhF+wtqMxyWeU93FsUBqZBY6k/mcBUzobBvf
sQaj/QohcWZx3q6ve70gugDJQvzvq072nT2OO/TJ7XXtIGYt4zVFmH18Wbp2bQiZVutPEChNzGrH
iq5l1Yc5y5I3sJnnZRiZQRBe43qDWoOITqLjHNLl3R12auVecgOFemF+LrrfhdKeGNJ4LB2NMq4C
pg0EFH02zfFj3a2uqfTb1RZ/WrRZiW+zg4CcOfnVel3XuthSbwZTt7UPmDpx4MxMa5OO8AnG1DLN
xZ89rdOkVVOf2lstueIC3yNydLJg2Lc9VncgobbVC4xpSQ4JrMmlL9zyaDiQHvwxsehSndaJwQmW
i+GvA7Cf6GgDPT7uOz6uLkYX/oOtbuta2hNDTIlFYv46PBplshh65aRSxlKsj+ajGdYOho3Uv/Sm
7nHZE79RItopX12lacqGsJ6NoJDT8bJ+j7mHcYl6EHcGMEso3wu5fXUHlbD+mmznBhid6hBD+x0/
68d4DaNL+ia5Pyztuu+Y2bSCumbVmCe72H8UIogZy41PTFiZkugxmhw5LqUq5I6wyUyqq0n2cOdW
CItjGIgn4X9olE+/coLIpnxtGEDiCA7WG9DIWymZ78YfhGWQ8wyjXCZUPH2VBN64g09B8fGseGFh
Z9QiQK6Zg4Z2gAuSKo1Imp70xFfQNiItwIYTOPUv/t26NvktLKBRwUo4My5kfAAx7EmmKiYACQO7
8WEgg3/wzBUEZ4xf/LGytUb+MNxfLkommfN5HFZgfgAogcw19vuXUM6ck1trl2btHY5gD88L2juG
tQYmJPqg80+5MFMEN+WzDMtvCfAAu5bWFcmPqpXWV2s1rOpdisK8dAWBIe3bqE0ioF0VGZmVueh1
S2GB+4z5QthVp1FXLW9VYGA4WpW13izA+Y+DnhIaeProAzngvIvtFUjBfpvqciIKh2MrWcfEovGh
qfUEN1Wbloxj/soobdC0DtNlkPCe1zt91c2qz89OmXTS7Y81LTWXnn9u3j2WDWkaxe578BXC/d/W
6miOOtdsOrxEQzyVzoysa62V6BMYgly63yMGs+xHfyt7/iQR0NY7VQbIPBJxfQHPfmDaJE7XSfPX
Oc8XEolTByWepWuG7YTGLGBSD5vIc+FhmR/tFg5JEx0UIWejaJtX0n7Dn9luLm7AkjUrWkuVzS3J
aa1+ZfgABhJsvglP/S3sK2mhFUCgNkj/U8n+VRa6bQZ8Dpbsf+NgYF6JKbx45YUKUZ4m/NpQtmo8
nxz4jx7SvWGBTOwFaRsLEPpThvdPs9Pex+GUZNAvtG3w2qjV6TjfBlu4Bu8dDwqAsHi595z4JmwQ
VVu8PsS+KT1Ge2EoYcizVbCIFIiVXBsG2Qz+z0fKlWTiLrjHHK3ttnNFhLXG9/A699ROrIfOLfOT
X5MVCINIrTcUwm97s0v/RoT+v0ZfZ7l4qhi5VQM23VKuyd0EHspXm3vORLatTNVylgMNO19eIeAk
bXwDzYa5EtiZKpMJ2LhBxxOfJ3OU5Cr6W8FVafZa4kOad62gr7NOmAf6YTBi20aH+gWJ8ZN/vZGJ
jxQBx56J7HW6MDcCl4RoypnoN0/kZFst7B/mZA2ZSUMfG02vaGXHD9Q1uiJ51VH2vI/ZyQ1H4Llt
yHRL26bUumO5dhLCR6sv3JEc3Jwes+QU6gtZ3LXd6/ZjvAA7HnG1XDf0yI9EfpWigoItcoCVraOs
NHtYO3yPgZ4sw1AC1PMY177GL4v7her3sNl/erIcY2xpdQjs1zhj0eDHlOwRwiMHwTeaB80dhLbK
A1MgFigMXWhIo2ZT3OjR6JrZZMTyOjnSZ+AFw0pVNR0kKxMijJUjYfONsx0wA7IWMkPPnQsPzoR+
op3JlOqYGgFC+bfy0ay3gCdudp13MW39uRd4ia8MA1ElguI3KVxYxeHkzTDM4d+VXH+NxU4+OITV
OyV7ToXzV+AqSiwkQgEQwHxDYWmZ+jYZb+4ERlud/yeXq0OTNLK+5WuiVnUX3J0ZB44M27r5ml95
bX5qDuZiqPc5U23RPhu0/7wCy0fVmkTGpeqpNKOmCA7ZNy5HP4UUIMImj0A+dKwkiyzRiZo/QAGu
E6CCE6slM/jnHpXPjnQKp286wBvWln478YzQlA==
`pragma protect end_protected
