// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:27:11 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XaSbWoQcSgrDfMff3irgvfkaK/0p/sl2gKHrSPjwa32U+F8TX7y0IsBvbaphMjXy
KyNEslxpeBx8MHDFtJk/Y3X9+Gx0t26ItqCq5n3/tnk8MH0icmloCHHhlgZxwKTa
I+pzefV5UtsYp27NNT2D19YqAUwHxoku8AfF0ONMKws=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5520)
+iow7dMsUwDf/4PIR3QvCwwGZKhOb2b7bPaqdQA+TahfvlNr4Xg1aJ3rPFSILyf5
Jfm65L2fv/9xcSOoZCCHYE8i5JR0aOykfpANJeKKKXF3reBGan7WahrT9SU1cP+R
uiBIVKHwUPQIblnIjQKqOhYQzg4WtgXjfNe6uO+8g12XaSQzt+GJIjJqwYHuksIr
sSVLX9NYYsTiaW+ElLfHg3T1lSWebLMe/ODjKAUAXLTLuhVl1Qy58a6h7lhXeOPo
dE9J/oxI0sw8HlWmWuAbEgfe6Y5N8nKL99x3jrU1CixUS7iu3DdcQmWRyVLZAXvV
tfI3DXbzFiSm5yx3lDxaCwgtthsq1DiOMk6jfEQQ4THV0oIlwLD+ekbVMIndDYma
05CgI/bpy3z5bApO04Zoekc6UVtS5yBtiG0z6pXTuD9fkfdtNzfMrPZkT8aoHhjs
mPJSGohWBCGU1IipJRIcArg4weWl3mm3wmsneTYHripfFq7cdOOgegvhHKV57olo
Av92hG3eYceLcX2ec5mYIK9WHwoYK+qXM/SWMxYvW9O5Bqm3f8VRShtxNCSxuhEK
xC75yarCMS16CPESeAiTbyI+YDBADNRfSvKaC8iITSH7YndZ+ghiTWxlikoP08FY
l22VhOPkadGHclv1OVOkRuTL/Shiegcj9U3RBnlNYjfYkkV54ss2hFFxGRfJV/jf
/yvKqEC1rne5RthCBEoMUbLi4lGi/4vuwZVgMtDyiL8VZyGK4wZIQeswOB7Llzbp
W35pZxJBhOULHnRDhKkoyifgVAR8otumD6rTINjgyCKMLHPhT1/ZhxCjYovUiPQ0
hyMaZZ3N3fVPIz07x/wovLwvbfezoDBRLwTSiqPvvoAx9GzHlbEPj6Hf7jg6RLKn
FMehlunxHTHXMEFkYTCWjzsb+HPLKL2dPxwH0HLN+j4l6aI990Po/5M/oFOdZKY7
Akr+26LfGuSq8GtOlJ22XjXzEXb0XWLvzhP7HiXlGRlnf2U3wBmOw710o6IkzbpH
oinDjarF1FBp4nCjak6+kjDIaTUnHqT0q/nEZlATcUMKhwP12tDzsDvWm6J4GADv
UDpxVWwbeZsdBWwUfzMhiaxzHZh2Bb+CHgv59Hy5btqc2/WJ2t+vW+H/7lJoVzMi
m1a0Ks7YrGtIZTF9ZYkWQd/668Hqk4CU7081Kmo7q5kt2FgNefAIZo8mSXnZmErD
zuHns4XqtJ9rTS8Bv+bvUCv23ij4KPD+q1YQJXFmqjYxnnJgF8Fnrqm6hw0ukw8T
9Du4BxFt6Qy0xoKtOWST+A65zfqZXHCLIxrZX9OtOLeXUiHiIymdS/fKB3uZZSLb
USAc8W2lhIkER7o7NrIe30U3RUX9J++en1bbcYQkdE78munP2m63p1Wf25Ms2gb1
W1zeN7wSJiP0nEdR/g5Ksu5NN397i+6s575CBvZtTlZ70mqWZmzmtmKBfnb4h4Et
0+qU/OgiY33C2HfOOo0bhN/BhyJXVhp2D7s6FUErLDgPcLELB0SzIQ84nJctoQ/W
WC1hNXT1XpyYBhlP2//Jxemz+ONykIbjAFhUUD9Ra0pijkZ0N+1orr7r3JaxPxa0
1aMvvU97Ry20vuH04YTiNmV448/uvrTt/AFNkG7crUQUxFNcrxv/fjn5aWzxSTyF
ogL868/VvsWCPk9ET15UyaAGhOuyKxHHY9StM5l3KPGrDqYdolBo4AHHpGUSbXpj
UNopDdIgcguP5pZi6fR/GjYMewrw453srpnHJSTBSQegqjFMvSGxi1GAOYPLLWak
wwKN2Ld1a5o2Bwyl+TSpz0kQIiBwARD8vrRL96rQDPKNA1Wlcy+Pw1kksakOK4+6
iLnwIuE9+LJfKRJP0cma8swJ0Y+F5KnRl30QYR8uTbwMH9erW6679FWpl81GebCr
1B0rHWsOBwJ64U74ET2kUnJAYMR2CzrRmlSepcxddTA7BGba7CtiwP1tA+ruxwex
YH2cDcu9t0LDZH0uHdjHI2soA4Ilt8SOApWpaDcto6Wxs34eAjujMaS9Ze7YYSjb
3hnY9ho1THN6fttbHty57Pb/Ez17TL9nUaA6mwKGsAvExU9jPRYxsd3G7X9fhs8h
uC4cPZE7eu9CamQMLo0L6D6SrvnDP6uneg9AI9/kYo7s1jIwe59KWLcLP19WQiyJ
ZxNo2uqphKnKfOY8IA453ew9FN0fif1pgwdL0fdiyufuznJwmZkJnh799Ffm7n2R
0CDaLJxREuHXkwxNUBsbMhAo9LAEQY21Cjpa3VvOYIG3sNoyWSZrGEMaJExvQ/lb
akZnc/vLG+k8ddao3I5NPzQguuurpaf1KPpZDdoaBaJZcZY0yyUFQOliQ8E9Usg2
XWZdC6D0mrmdeb7TR0d5FI7rMeld1dgZHpXQktiMk0LszUagY0rgiXPYbPDUjLIt
vxa3a1mSqSsG3RWojWQDlyKKE7dB/h+XX7IjM5c62OPpnOqol/LmOjqWWpTO3SEX
GRrw4zFrP+R+Wb1RmYsTEMcpn1evqMzh9hiYrq1hNoSLOnd1q7+8dX5/PD3Y3UEW
F3XimSRVcQxforHGfkFVDcykFMEL5qoUZjorU6WqkElakXfMkbYxUN6F5pMI16uT
+zCU1iGe/I9WD5/xM3L7MegIT5khwGto029LGEFOrVLzKA74ffd2vv8HcJHv1qd9
YwKU6+LuBzoLxcVXWLHAAMKruik74nIN41z+awbwpiUAbSOWmCJmusxgnS7YEUJi
czgRGTRzZl3UQh9e4ECx6vXgaKBU6AgYpRbwAYeInK2KOjXAYRGpXncHQc5Mytk3
H+C+QrfJPurfyqE/iWe3ZAsqcMeP1kOdS1YfL7JNvHCC68CwnrP3ulXinE3Lb9pj
E60u+BKZchCN2XCil2DXxWmrrRUXJ+0BaZumtF3nm+Omb2KQ7dxrFWLzvv/NdIAi
ICdErR+4YkdJDPC3566zGye1J9MxDwU1FzXYhxWqx3qbgFK+2jku1sm2F3bhH/d7
yFcTv97MyEO1lH8fjQFOByVKTsn2PfJgae+ZjRSVDog/6xlt4Bavi/py5Z7zNOch
y6NVDgbH6mMkiYYLPWmTrgbWlIYh5TaWlgRWZr/5oXFKAwzoHYq3k8cSw9UNKsyU
cg64I2pUJdLf29jJpgLqe2j3gyXFjFCTsc+U+LTCixWrsQ4EGhMpKosu/1LB7/eN
G1E+McsFXZzfSaigvNZk+E9sBJzERlzLzscYaUd/FaPS6WjH/DhJ7e+2evBu/u/7
Ki7W9fsjyobFkC9QZl3+25031jdjoirTm8YsN75Uybvaf7nih9zF/lWiH+71007z
oNRgPbcwAdZgdh58ewUHxwzvE38/JGQ1psM0M9ebKArgC8hiSCbfAlNgkmPz0KIa
p8fCzdeKPlbguMuad9Rn4WYv5ZevSBMAFvKLI6MmNYZ9JvePRrzMyHE07A7JAGa6
1AxA3IBNfVfK7WoQzK0XhthdmZ/68+K9uxlIUotBc/g2yN+GvgcjyfDeAuQHddh0
1FRc4EgiG/U8Y7ansiO1bgxWDSkGA6zajm40PdeSbYQcqgwgVanhDl8UV/hGevUH
ZF0VlU1zxQ0lielys+iJM+OR1spscYagUiAMohfmJUilu6IA4uEhSBPGlwCbqA9H
ACZt2sU/FFL6GICLr0CfdPA1dbLA4iSKyroBgj7gdMmMClYE4axw6Omc2/11rO0F
vGtO+JmEF0dolc0inm9vokY4mOP6R6Ga+tocY2UN/RiCqRQSFDJa9QoGLD0U8/3d
NpCZxWoDXJd4TTLF/XUB1M4TlOvfIeeC+tF1FLHfqABj/E+v06D0jmJB1gPgyM4D
jOgJ61RGf7FF+zAs8ThM8imqe9AwfuQUbHyChz7X0ntVv08+bAcfkrcGrGGdV371
c1Ca7WJd8n3DgHWS6ECBEUiG6+YROnUaMZBpUX8l3XhcExSBRChbSKtS9OasfSgF
dDg4EmW2NPxyPGzhiNycv6WobwiF1u1cNf8Al7acGgCZQ464KLLJKxaS33l/AOPM
Gzf3xW1gK5lXvjM4uZygZPKXb4rAFv70oFMH7L3RRyZI74aRAB+T9ARwCx6yRl5b
il4PJajCWThFfqcbW72YmXSHuov0ubaXt80Hd/DYoWuQEDomXQw+dBAjDEqMPyoQ
tEgpGqzkYyTz9dr49urPP3H1OYlaU5CZE6dtwiWxticePDzRD7pY817bhkUiLuMX
EBCPHOaPmxlFC4OMMjmu++lFvV5DjBGBNK/y5JZckPgEvjOti/j8xYMwVxbmdD3L
6z/J2EJeEirL2gOTi6RnVJWjHBCBsZVtEsmg3CpAUaFp7SJD51eFLHbaHGGMkTzI
SG67Zs56TzCjrXkmg8p5GCqOBfOo3xiNFNdJ00Jl9A+B1PrkX9YmX9OJhmt4wVO8
rMa4fsswX5H50eJ9RT0yUGnn+QxLpplae6EM+aJobIs4sC7Xeoe2YOoZecKK+rlv
0xbErDjjwkS/wEkG70Ehduqe/p4J1sAORSZ1cr9VRqzd0RqgyQYkxA89ekglFuF9
TnmbMuYMQBYJlf5evLqAXEu9c/pheBDZjBMH3QMCVzkah5RlJME2yN/IUYA/yDo8
hgYRWbn5TBXbLbhkxt0RQubPrm1XvbKdV0DLvLd+IocV6g3UwkvDh/z152axt4DN
CY1u6WZPH5gPO2oJv/nNOVYi/U99Y3DNkTAoeyo4N++RbpAxfu0Z4eGWo30iNHge
FdihLTBDCuKOHvHAMt3Kpiy8epzFdoAz9PXRekFznbTRFANQfUgjVPO46oxYsMcw
QHTv8QNtisU8SZbRmKk1wq77+cBmCZ8epBYubYaWXOYm/hDLJfKQhIOi1Uek0Jly
qczIWgyS9SrSeP4E0AWXBpmiqjSgGT8MKZMTpohYcLD1+cROSYBoJpDsqHRXzvpn
4Xug4YNEcQ2i0IBQMe8lTx/oaxWjY3Fg/SoCazoOlBk0PwUjr6INDRuAZBhYnRjQ
BjZZHT/h4BhUWdY+CNKfowPhYljw5ZGW/4TiJHxklTFBKp771U6HdWahYsSWb0h/
HAn87bCW8eDJsoEfV8RNoc0pYesKe4O7AHScIUAGtgbXswUGUQMvq6KkvcUczLRF
pRNKZUIXzTv8YFOAZPwth/rh1QGQNPya2/sUB/DRF3WFOThxl2XXAiJk1iI7Y+5F
r6X4sl4XTwNh8M7kTSjKlTQiaIV2z9e2lavGTaWanViOmw2sb+gF1gEVc0DAwlow
y2f7lx/1FUsQK6qBsR+MPXXQ8FftujeYDG/5Ev0jzUut0y3t0OgjYmcK3WMH1kV/
JMolE96gSZNbeXdxK0mmr38grm1ADsp+nMalbnTsyyMIvHn6eQ6y/8bzOEfnLc1a
ypf+oichf6asYWIfjYvaukDnDwjG2SiNXIoQLtOSVZ2rtN1JpUVkOHdiY48nkmRQ
PCSsk8cNTnQw9mNfg4pY+v4pOVfcrNUIXcL7kDbEp5k48IaBxikLOAR0dHBXaC+9
CaZ5MhJmPsGD7Yg9OTKe7wI6KILb3h2zYakcCao9/sb+ntAdqcEBAfAzLCj9Nic3
6g1pY5CsqE+GVLmEcdKZkq9fXCopM4jWeyvKov1yQKVwAx/YdKMFp5scXz6VZP/g
WLtyypdUpDBC7hUAX4bT1ECne9tPBkYUCvVjJgdC1QZF5SWwGHZeAvVjbetHGz8g
v2SbVsnlS7cd2elr4fsfDqISL3b24LNZXkBojB0ryK9krSQ5KJuT+8kjH0NeBQKm
5vKQPQNiabE66C4GM/pIDgq4YBeYVhjRgpHEnP+2klt9lSkY0mQRyiH/8oaF7twx
+a+3RcDwniH2IhOEwXvlOThVotMmGaw6Wc+XsTH8HXijdSBxoX5VUkJs8heZxDHD
f09+26O6Vi113YIkxjhPVh/D43cbrf0iiHKGSMeaZA65o/rLLmOmi1i1XTkw2ZF7
8rufwYcTQbeCwIDafGebR4UTw55iOXwmYhvim6ib7OBuow+9RARsKkOejXFDeLlv
0q9/6U3SG79u5s20Fz4hPYV6vey0wD6J/OdNlpHUq4NOUIhpHtqRkmQZEF14p7cf
n/Uk0gnsB/d6fItktz6GFIbij1Oi+N7Q3HfftNWor8SK4WhKx9mlHm04nyTnBZWa
1KJnAqPwGy/5X345nM/6Sakscf6tj8cbep6RS3Qk95qOl5mqdFcgbThItfSBaahU
6xv9R/blDqw4lYZMoxpVOtJyBEgwiq7AcNv2AMoY5OYvSB8e8PUY2LIhR99Mjdlb
scJPI5I7msSOvfKTg6g/ZIR5oM/NZzT0WMpbVSA46iyYEX/y5i1cJAYtPxkagQr4
4S7R8ypU+bw8UsESUL9zZwKag/iznWaKhsbUlUMZ5WFaMHz8X36akp095NxAUrW1
LiyYkNgCdgOe4c2j8u2GEpOgIOd1f+ndpfVUwEPdfIb2fHCkFO2iQnpS1xmYL5/8
OToee37BvDmLVU/0CVKz0kM67SpGNDHfSQ7NFP76LKAaZ+ibAbTAH2u5I8s04UKs
Bo8hORdixLS9iieD17xxCX6ak4xAU02+gi45dJMc6gDPt8YmlOfkhw7G+J5NA22D
LfhRrOLCYs/TrIiZnD4peu7hNnGOgHZVGXh3hxlYFNNx0KxlcC51OLaP9XbNBi2+
M5WnV36vyiDSPTImxYyGGO/ZMtzPKESmT9E/eFkjSEAd5/GDyDEuuntqczohGKmh
HG1lkNooL5WYxgpf53z5r/GEM4K0JxkD91946j9d7T94Lxcr3zwbXt1LLcX0uisT
P5meyi+wPUn3UOG32xxAMgjVZNN8cs1prudxOu5sPDVRwv/rRCm4RTymXyT9zwMF
eQOdHwbYdJsHL2j2aa/VXJC2BPjvCbwKpSJg/ZcYzbL3tUZLqBmzFv+KPqEh9r02
YJ//NgmMziGgDNPDrEznXAIKkThqZ21lShE+9Cmmhq952LotwSLhTqJP61K41FgS
FjxTlgj2cXtFGTCIy0vggp+yEO1Y60DBxTJ9lKlPkwVyLxIoA+avNsQFKmUMB4k7
y+BYBetfYrD3M1xnZVHn/Z3EQcxJ1kkTXMbIlM47S6UVYbamecU9Vovosm9jKRoy
nFGqSYnLt/GyGqlRk2cKqRfvWHvQYXc851mI+EbVDMr6B8ocC8HAiSrsmPtmy1OF
JUfB8yNDCaXn6hScVZAKoE/Ub+usG0oqEL6QAzhDaJyqROrm/DxOfWKt0+IV3wPq
TRlZbODJ73oBGZ4+40yHcnQHcpiepKDr6k0XMU4YFMwj8huc4Zqzk/reTqXbEckQ
5WTlbkC3iVrFGKTVYoSaP4xD+gly47asQTz7g77VgGuc1cpclgf1N62NGcK68aMu
`pragma protect end_protected
