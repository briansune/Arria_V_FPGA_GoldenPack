// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:22 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PM16YX0XE0oQB0EWGKmI2tfmCkk4ofthP6wjJFjSqOGxIUURv6h9kfjFdAE/AAD0
Mk8syuUHwQQ8niKHN/Fyw8zTGaj2S4MU2yFaIqhiIkrDN4bsTAsP+Vdi4n5rkT/b
35ku3ksKFHGQOmyZ3SlDXEXC89vPC+TFM37yJxeTJFI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33696)
MquBlh1TcYjfHBR5FD17qExzqSuk4iKlgVDDYUgE7VgpucJGvvjuazLNFFBVmCOp
sRv9m61hkw7/Xr3o7/a6Q3VbF78avtsEb1fngBo3+Bbimz55Tvsokt33La2a7GSv
SUrRAWrVOY+FhG8q5qOgVbtuTXoHPqP3F2A8CQsy4wXvudeAv1JdwG8DgYnF7gpz
2GCRarREWhX2uB1oBcDM4dSzScwjp1KIEGMLAK4GWbcuImq4lAbvdlNqrpPj01oI
dWPvE2Ft494v6c08G3ytPm54qX+Ez+QSfD9BQ5Y8Cli/F5KD+lpKKjcVwVmoemqy
POFzTnDG/4y8ABpqdpHroFSFy6By0rLq/nUTRHHz4sEombxmjmdN8zLOwdX5rurT
fxu0MkFQlXgPZqSoXCg66QcbU6zyNRws3jkULTALY/XZMQcjdE0iH6U21qSyurXC
IrT3XqOyff5aXwftq1P/dYu7NYGqQDhAFf0DTXPFFsdoheFUIcxtqjxEp6+7wjXd
8eZG73yzlsWbm32tqIarmUY4sZH/JwneK0ahKz6LUfIuyJ/cg5IMjuHQntXkJq6y
aQXZmRKrs5pEplTmx7q25QOWRVrbUur5LLbLHGPEYWMXdMK101e7ed4RH2DNVh1I
nIScmsay1dvHE5Y/tSmxUL748yIRPU+ae2nEj9f513pDAiwP59/W03yNA7/UYYMY
YbCNgoj0TwSqOtfXb+5xp6oyHUWROKfzmqA2NWiENaa0Qgr80LBgrDiq5oTdy6Is
FBjLHwynt7wsC/IhPx6WuSPIYAcDrG/GLYOjtXbSPc4123WipO42PcS/oz7VT1zH
ywHU0Ayc1vkZFAVsnrKSlNwk1WXN5VZYUwgfht8Wuv+WAUsqTV8sViTUkCM36VCb
gJF1cNfxgNRhrS5UFWjtxXAxRTyl0HZI4VQ+hvxnFrgWYGZQt4FDJP2Mt1mF6LZ+
nsjLZ3ONaGQrMdpjwkKuOX0DKrJK89OFb79IofN/buTNMV5adS9r3Gt/JPjbU7KP
LYbjHopu8mA6LFsGB6h6RjuDIX1t/lGBgb8nwlMfW1WzQH63EKuqfLe7VLnLF3Xf
R8katHkcKQ3Opphv6ppK/1V3412LRmqAa6kGh2tuPnXUKEwvdxyI1JmY6FtUmAY1
7eiHkFCW3/2VttwOaUWabA3n2rHnQaoTSbtNLk2p+Uzhx8/lALJT7ZbTkjTArMCj
5h9KyzJEIuDZDaPmPE8wnYJBdhhjlB/QX6gUXLrRpVrv7cfqjY9FIcT5Ev9PRPS0
Gobrm9V29uSlZlCrLs0bpzFxj5le6kD3VpeRGPOfJ1nRqsqH/7ctxsRAa00LFB8J
EtvznXzPsp2/5EV1rjphMTNCl6rHitWeJS0HRVS+r1Vmg9EeuJ+QSrW9wOMQxtuV
7ofGUwB4e8W1R3MzP8bZng9IQW7GRC2IZKTk6A/8+Z5dpUsHBB0kp4cpEYxbWZgy
9+4GqBjsrn7SorGevcRRiET5aMCOPivgizjan1INQasEs5OXuMrT9g7Tort9LwLN
idnQUKn3CtM7wLTw7ddWxsKSBRHKv2djk7oSk1DS/AvZoipJagE29SlZjcfN/oyA
G67LQkCbROjUwkgbkLnXLFvO9ARmBFSiJfPWpx4zUlL4gzgrCPKinS5HHCfFfbgj
SSL/j5flWJPiIXa7F4Gjf8ezxxJ9Yg2tia/Aljx2U289oW1V1ny167dEXbHwAWj5
Gwx8I+dkT7wKHEl8nENxwIOH5Kf699bYz4mhNAHA5ty1AjYS2XzrIAwg7K6L2UjJ
YLYCcvZNFprXHbUhkf7aNG05KIpaIuE91dimHyjSyYeJvhJMOb1q50nSIv+x2ZPo
QpXG8mIULTNofGXhuLGv8JM8oo8wqKQMcqT2Gx0yZcRAtSAIrHOWpg2cOIx4lZlP
4BeK/q7cSHD+1zhraMwy6MogQtqLUaJ5M0VJjPZjuWAFCja6ip6nHW4qFbULiY1o
6sUMFb2Lmmof7WiDvlRQaYyvDM+ZRgkrqUTgqrR9+1MdQoTsnhYhNw/BXyfqKjb+
G3RuC0u/CW8Nazh9/jTTNenTNzlO3w9UNQbjQgq/Fqxhb0uJxdnTg5FELuINlgGa
IJi99WUS/d31UV09bGXKCJz+wjrxey85HuNPtbNv2YFsNcl9WitMNYRWvHzuc9Ed
3Eu9LVyf7Krr129VWBoGG0oSmu36SmHApFliexXpnTNCArVpBye/szhsfKjCWNlA
bve0Yp5HvW3RKsaJ82AyNNcKWf5tm8X6xpRsLAyrL+W0RtUWdC2p1pOFWykyFGqi
vBMTZJDz4TMbAhKPWWIOVWL63VgNaZxvVU3O2lwaTPOCPYCjthtyhJIhHo/pKBTl
dYm2Gya82+1ZSXtoeshAUAe7vB4hfkg9LfhdeAwDstsvpKbC3iQDJg8vG8LrDCL1
w6K4M4V8aLes32Npx4pmtwZXs/UG4bPoNHIefmpyMZnoLVuTx7jNd9MKX+KEySRw
jDGD667HMz8T9EDwsIpj2k3lgvRRzm9t2bzLL5siKmbAsHmn+t0O+xEOK+Y417Ql
2h1GOYb1UDyyLfLBxTSp5w0SXoS/vP8WyvOsEVs0fm81Qo0qFzmmRk62R4YRWjtL
/+pL76kmdyWflJ79RGYypOrfWIUKUFshYv/SVAsTDDj3DJhpNuZ3a9XR7lsLF+Kr
a7gHxIIHupxVdKTCFAE7KPFyBVbwQqEKTyn6gOVQ85ULI5Wsx0mAfXObB9Dd3wql
j1vtji8cv/wKon/zf6fTEC9XgfLxtc/Ea+Kt/qXOOzAjvMQiCV+gkUBBj3gvuVUw
VWF948T74CLFfAp5k1RJVS9inPx5sDdeCQuwJNOYeRVlipIO2XjkIlQ6pfFqHgA0
3tSkwckCGKPkWCte7gaxBroFWfnVzw+IOpcJaIFurwbRxKG3eq/rqLZOC7GQF/M+
KGO08jyr2RUNI3Q5tThEHfQVz+v8fuf3hqe8BUGB4dnGOr65WIfK7t0uHnF61wet
iFuSeHKaDEQOmkISizKIwST3YvV4lmF5nBEG3f1/WHnaOsXXH3KiuW4nLK0r9vAH
DrIc0nVWvyePdoHSGSgT1akYjAC1zQDZILGEYoArwbZ4G0dkfA8OF3jxXAtMpbFi
0RWA0Lfuug2KP4Nhh88tLrYq8gP1kEb4DBv3qwFEWkWHy62hMofJ+weKrH2kFXW0
qy+IlW2h2sqzi3lJAKotc5rjT6HP2lNjAAZQYQzRbYb/QTUYxCV4yvybOlNpwRU9
iqkDKS2Uk704V3ejdGqQk+k9RFSXzcd/95bBjO+qm7RZJoyHvHRez9GlvFjifLje
E9f8QyTg8elR7YrslDO9yj734+Tacl0ny72BkzKwDqq0claDXbNprtUtYnug9gDK
VtkKaGv18ApZMT2OVEgUGt71//xreCAmdXV13KcFRPoxVXIoCLvo7WtgBEAKl8Uf
RyTTfcZItUTqRkoXHN7gDDrjwl7WVrr69j5ZZHg+O5W1QA4bd6ingRGc3S5B/Vkn
IdKUmtUFH3epzn6Mn2eFGEpTBComVd7QiUz0jVcEHyeIh23gLJOQHT3VzkaLJe0u
anVSuVYNJ7LmlskpnTDkw3vOElUFDAAPQ9z+XFwCh34Orh4ClwWiCIHyg6IHCRdf
0eIh3pk40T4DQ4MNabZNBGQAa/VL4AP72e/JM4DQN+rMw6pcnGxLxuzpVhl+ObvR
wLcDWxE7PyHtkU+ESH3mtCSxdtAXdhP2e0wV1pVrlzThHERojr6MfowfdGuMziHs
nBbp8hkIm+K83JvDcye4z4tYkDPxwDuC5K/7KxNtb3k6V83nS0lemdAAHNxIrtIv
yzW0fO3zlRvfg1wkfnDmIDIDrUcNBAxPJshpOhb15U3jEF/0p6TiMVUURYgKhb6Z
Dr4mS7GV34AkjcwJ+McWcUtQEGOs/cjwKNZmy6OQICXYSiK73QGPhRjObi0rDMdg
M1DO+mFxoLUaW9tdl8ZsuNhqsrGbKf9fS6uDM7yxvXhqdBDibPFJjmhKq7zV6BEb
7M5sohy1moE7NNhVDanC+49jTSW+YCOcaMRbrAJ6J+YNhVSREiCswdU6/jCa8RRd
yAigDNa7QrDTjdtLGbKGV+Ej1JvKXINEOJveQD6zrh/Geti3/EydPlPn8nOlVSH/
RgW4EeBJT57yC/AOT26vZBXCSNS9SJQF5tV6eSBxvY9mVaRR+AiuAR1K3rwCpQ+g
9R1glumWYiLQh7carB1KJMbYfA1atoMTftkGJ+ubpI/S6usugx6wTWdPtjvXj1am
vuKe/ebmiIuvyY0snOAJkVgTpy0Z41UIgFb6hNERzlgBvRUfohY6UIf873MAsID+
f3YWR2HuNH66RNVlmgvjBhxoi8Wj7KqY8OpZZlCKHkLFYUdMTnTE51EGlsMD6zwP
fHdAqYd1d5Mn59M7Dfdm261nCkPTHc7htgjRHPlWzVKZrXs4Qopz6ks3DzIy1sHl
Dz4EHkGLKsi3q3e96HR4hWeqbNKE2VVffq8HPzujjWq2csU9c/aBdHbcMAh3pJCk
tFA2IBNf6gMesdJAINsVO+YYLHvO56RgjrJSaH8H+1OJWWy326QtLJwwtnDm+g0H
qkCjPSthdsHwOezpP4FevklBaQWG4ljJlLEZOFGj3LcsTA5soxuDInUHVXBiGMLi
kojp4kk8hqKO/yFKr6pmiybleqzll0hwK0UkrajyDU0w6BuNnQJN/55T2At3Ajwl
GfOp3TRiwLmQrpgoejET6kLnA5p5riMAc3+knDJytzB1gpeqjaOl389GmX1zxD9R
CMuJNax3qZzh/h4bOHK0fkdhzmiemiHWVo0ekzt7UHC64M84rveQ3ahXvluYs3vj
EZLplG4GuVTyF9vu3rOnl3TkI7Hk2pP4YqPXMH9wjEemfyGTrTkwLLfEN3jgu609
aRbtJoFoFsh6s7DgveP2QlV8vc6gImvVaRzrn6gkAiL/PDT1gBzcfLxyQmh6mqLE
rLCNVyz4mDxyFHYCU0y7kitdvRUlHiYArxJuGqGO6uAiTVr4/k0r2hXY+O1i93d6
zbYGVlZgDl1maZe7hEYxcgYCHRam4acdIUyBlgvT9dY1gqJ19qij9xEgDJx9ac8m
NccaBRHOXmgDnYnHP1QZY0YKGuZNfi/msg98dNno7UM8VBTqVSilcTXH06q79Nao
H0UhzM8FBVjnzoktncOfX9w4WIDDhqeM8edTk7vFzJm2cCNU0796PpCT2gyptOoY
8ttKDzBx+6ZwShzo6rkNZlKLtKU51QHnyZMKmHJr0h7U1hXD6les5RmRj5z/F+ZD
4p4GmAqDXvprVBOdQ77a5lqnW3PUUxvjPGET5KMXY7XE8Moy0vzWX7/DMzSyL47R
IEUpSyOR9ay3otNG8Nqec1ITcnSZaszY/2DnEm0dq3m7lW8NfCgguSbwzbk/hfBA
ElxucHWBuM9RVW0bzHdRtPNLeHF8lYgPzjjgiKnYofQa2SDHwG9N06oBO3skB+KC
IGsG/1mqfGdstw9TIQXZHJ2CcLNmzjvt8igYcyptipsJEeV3Uuu9ULRs/37cMmfp
myPb3ZIioQbyvq/kaGUuX+Cfnz3AMINvBDiHlt/UOW6diS7hAVBrX+iH8RXVW8vw
AudihqBVptaQijj8Il5EfHIjnEjsxkO6Jo51eTDVkhXVOlggR/032lHsZqe7k8ka
PdJOGNwwKou9ctpDdhCeim8uf3mkbtwuyeqWCTATOMcDgjaaAFBQMMD79BbtPAf9
Sdiu5E2tknIFNyisvipbAV8uOC1hMz3YuWBxRLWqNOgujqSo9wyzSI1VhjEbxNm2
PNTN+mqvxRIAntKKeAfZkSs4yqFjh2esex01tK3KOnBCw/oYEIRwNGrxGgl0NKEq
0u09dPpUr47smLHqPM5Y6VZYHmKB2nfYY0O1Uw5gtuMp//UI7UVYxb+O4FWAwram
tmXQLz7AfSvbGbpbo5vRP0oy6OYrRsX47Lwa1wuB6Nq638TO3TPmO0154+wMc8kz
nujbCuhAOGSIMcUsctrc1J+l2db0YXlxXR72uwTiJis918CoNtrxQD68UUYPYgHE
u7v5SAFdSmhSZIVhcE07rHWfn8kwm75WLWnqc0y+oHnDfkbX9WhZEvDA7fuMupqt
hs09Idh2jdRGxc5CkW0R5oaD6EDIIZpUxJATF5/GFR9iWi9p7J0Dd1QD262sx/CP
G5oRBaOjXkFPkXQ6sXlsQmJK93diUgiQbtwIJw4SJ7Ze5CsAQad+UAo+Dr9fQNsy
wECAaSsuAsy7EuTDCmAS65ADSXvCaAjDTiXHmIzpMrfgkA8JLjn0yZ3kyWq/VA46
zqC8fqMgQumiNw7N4yhL9qSMloHJ9pzbaZoe7Yt3HdQ5uMFH3nIkBPnT5iPLbemB
nlelot4SAyRzq9vVUoi1VHBvIh2z4WKtFDk6/gD1uxdgJw6m1ouvXlhlxFYOEOYO
rUdsMhidy4LZudyTW4goFqfzc/7s2XKmfCxOy6KtzQrgXson21H65hySjD3V3JGW
LzjyGjyYwZwsU1M//tIx0JEnB5rHsULHaosQqVYMhnTTSnZ0BmZFJPlw4pAoYKtH
Lkbv5QBJGes4Ev0c9ttFbh270AP4CK8oAcC01yegE0g0wk/46kjp7MrwnkRbphFn
qQ8ooSXuUOX88Q9RmFGz2pXuES0Q5AnTlkMejCXbdCszUti+WCvszs4nDThG5j8D
VzBmEtuQh+6DG5wLBFwPn4KBqsXzmVnAb4puRkpHfQ1bPUDtu0MVI3jv9nrPMGYF
96K/g/JVVDcFDhyiUJJNNb9386Eeamyl+i9kCvImW6NTF81T35P5Tqh7jsIFz13W
7BdQPkll6RxH/ho0jXt4NI2CB6o7ZXohgGw1zO9Jd6bMxYppuqCsemEecEl4X0FH
usWDYikx4ETIzTtwKXKQGTTY3C5lKAkjXf0XW5Muh14FhP6oli7lSWtlxOH/Ut1i
l5K4VYbhsimhgRfG0J0dH3ah7cgJxNwDsoHK8nxBkQbt6ZahmmJFeKwMoDJ8kN2t
HSSiIx3VJoXUqieeMOwm00t+8kmFZv1us3GeIDwhNgvbocFogs7cdhAG7jMgRdnz
s7M4ObcvvIJ4Y6NdOEnN1Q9WvlcnT7V+zW/L6/f9g9VzMjVncH8iCLc2ZiHq68kd
2BpPqvq7FFijvIQO5Bo+hLkByjRlJbBLvwUrnEkWvrECiVpNi7t1n/UfDHT7Qb0V
buGsrkIwdW14r9fEPNM/wRV2PKx1l7ZC5SyAELBJLaM3f8ucA7fPaBo5Ate9Nfu4
qYl5pLL5/sqYtPcmGHdrt8JdoiXIB84hiUieZoUVVyq4GamlgdZaKxhjatc9YApu
f3VAF56PdSLFmmhurIaUK58nIBafk1Gaa7Lwg6Nah5kzIMOH2k1247DtvUUE0c60
CFOtXrp3lpd8MasRx00Ikf5bCP85m5pIdGeyIuWG7/iEF5Taqo+dPvYB+SXn6R2m
JwpenfR+qDqSDP2F7spO/pmQDKBnBbGdQeFbcqfoVPbcVF0sFaRCd+a8dU4FBVYa
vIbTOXzuKAUMCzM1LLGViIPesb7OUD5OiV2A6WutIAkdo26Ti/T2KGCTYFv7cmy1
YVmklHZUFOh59LC9bNaYBgRzHkHuiNXkwU3zJR5xCFpGdvCfs+S+IfPM0x1ipQh6
gFdWuL1IFBaqudq+PHJ7PD66/ad0xEkb8XUmEkILnXmPyrMg6w1N9ljGtb47Hvpi
tpye1hHI1Kh5ipJKuC1GDutvAHyfWtxBsCl/R+JtMqgyOUTOX/kkQF0frT1ww0uT
KgYZbUwHLkzx5d50GpaLXwSLThwlbZ9HVepwYDmfulxcDPnSEpTYqdKX9PP9fU0k
OINdIeEfZ7Jti68qddLn4nIKiUImGMTtAuw0T3LxqxklFB4ltcdmVvAPWmUSzqpZ
uFIXMkotjEQTwhhJchqaWtNK7aedPDr0TQOEhR45QtQmCKJmgzaN5JnhEfsqgy62
Z64t9XRH6kTYVF3AwBXpniQ2AqWvH19WstdS0iQHd8RjvYyV1XLmlCWmjh5xmz1h
+UtNJe/dO0E6kwM2Cbd8MDsB+OKrOUJFpDSNMoqbm6F7Os9EVufphmhXpre87ijQ
kdTrm62hTsHnH6kEsanAy7aIOUosOamj1cuwUSnDEiJ4vQXudr1OTXZ7IA0tSmSy
9KUQEKdM1uJZ32DaOxMNWbEg19pON0XtcRFJLR2pC/6AgK529nKsxjJRXX7NyUI3
PAtgOMdTXCZr3yIYmlW7UFj7cuzLTX1zxr0bi1+gZ5tnovXVt0TT3TVCpKeoIgJw
mxGP7cmfW+W0eJg0kWz91AzMwjs+tdDGJ07hCqiErnNw8JyQPMvKjew/BOvYAIB1
kk0DT8TkCNsBLwImPgf/J1f+0BPHGAflydDH0W9o/zKyz3tQJBc7kyL8rHu5NqUJ
v5wjkjmnLW6Z/APIkxKMh+56ucKtdQ8Q2b3ICTwOXsSGTVFNxX17ZAcyL4VSkiYw
pXCVxnnv2xWnzWENaHS+LF7dLJ3cglbKRPu0fLrShcS3TUFCxHIKx7htBkUYraT6
TIzUUN1oPHbSduJgcR4Vxm9Fx8TyChSw9TMsxPWhK1je4RBvo7goKOJtC+wgji0M
Az5+dyzx9icWTPd1wJucobavtJ1IctgYipvLdWFr5dOYgghn1hu/IFm/U+DQ7zBk
MJgnXzNHgCOvqDxHoAjOlXrZE4ODon4pof76t67tL6/YdkqBwGyeSHWNwx8CnoaJ
7SNE+9Yk0wghwVlU8WAfG7lVEnr6iNjdi4rh3q+UKkE3Taimsh12FmqdAIUfK2gF
ecFZCm82vdxWBdwEFtUdCTPqdT8k8L6oD295kLCSY733A3DKRS0Y8gJaWvNL2CeH
CChADKquIXhHtuhnLv4mGqF6E75ANsVCcLfhOPLc3AN+kq5WwBvDyuYjcaakEVQK
m9CU/hUZ0roVuiqIuZg0vQhaI69IPbWvqn57VWPZGD3ecEpcuuvWucJt00RWPyCF
kaZnu398ukFAwQ0hOfBSc5/4D5GHRHMFtKKL1y+oR/CV3uPjzLSf71nOaLBYeaYY
hIHkbYfTDgOQOhcszDyVjHPbEih6wCo5tcJNZ7Ypj3XtnucIuSjL5+9gr/HwiK3w
E2K4nOWcIxE626di6LsLzn4z47Csg2Z3Dno+FjvzpVfEUuYPaZZVCwBTmKCWx5PA
wGYhmL3rjuVlpScLS1sV9wwTQuRpNXq35/immNdL5e3jUbmaXrgzCg9H19Mq9xjG
F6I0/mbgDSyY8XzA5XRtVf8hz9klgGJhx9XjV6/T7rmK/E0r48qAYu2tpz0VVoZA
H87sHCUx10kdSTOV5N6fEYyzLflZ0pa9z+vQBKbr35A6/zZYY66EKQ/mx5fQV+Ae
m/o0Nzxv1ipy6p3JD23u59KO0vaZrEkHmYlwVzqCCUJl2WFzBYzZswIpqHDEDsOP
z/4pLjBQycnh21r7Me3tsScwMA8VGHBPkl3aCvOfBOl8lWaRmOpSVTNhDr9q0iUd
xrWhl7Z3HXnB2VVvT8WRJFYQD9R2CRjNbsgzttFabsy5YCv7dEzVr4PRe7so+HTo
ixazgEjpWzZWI21xm+W2xQPN/2OpyU+sI4fEq2lLe25u4RZlL1y6w2N5yo0mN5f7
3dhX1QKBbQU0sMPXCz2CWVkEXrp3n/t3KFq6+kAnYtY+Ume9KKouJu44OOYa87LY
6IF8tU94gkWgKtZns0zsHWK0KfWJG2PTHOTzm7SVg4QtJQYuj0ZR1TfgvRVCR5KX
guuw93fohaTITnTvSz5DZtIxo3Cern9MoWHR/gPpDWmkcKncZLM4oyE7fziHJ7cG
jhsi6+oymTbox8k+L5ogl6OuJ8DhQwYV6+KM5Q778/vOjljqbmvWRsL4jv2d5zSS
vKmprrOEYbPQFV8v+dSgl0TdgOScIl1mMP4neQQl12UYMApfevoUshgrHmqiqoCC
5CEQT65ee+ZkwYwg5Ox6+MuT6u2c88lrz9WDg/0Q0RT8pM8qFMLRcTnR4T/Md4nM
tGm+bF2C9UsLEP/JO8RqF4UPj3cpQ3MvIKkaFu8/ooFfHCwBku8UGPjBT27jZ/SF
RbrEiaMm++ZqX3jIOmPsoX56U7RbOHLVh33pqwgNtFzYsvLvrxAWcoZITJA7VzvE
ekysM1Wcb/tW3b1uBbov43rljmzDRRoZW8ZbamL/XOHm3Kg/aPjXjEquG0OLmrPT
uVo/gOgUGvjfl83+a76D5gKiyVB5nDY4L++l2ZdSG2rslIAlqOSVxmBCraCsxoQs
WKCYTAtbmCJkRipPFs5+gOUPH+um6HxqlCeBUSj0/J25YMdTqMmXhMUuJZAtBOEi
EMFDrAaXCzmqatNVNeg6wUsffk7u6qB8b9vovOuwqlVGY35v1yUa5ePA9KRdfwHc
L+C3O/WE/USrdLgBRlm6M9bRCzuj/FGzI/afpZkUJq//5PB73keXzgmMbMhvvRQ4
cj8jnrrvYMCVP6ba8b0ZWnuGibp0zfvTZB3eFduSGVh+R17DX1Ppg2P0nZsexvAD
d3oUmHLGMgR45W8vEJdUkgQ/dF+fM2IHc1Dum2O/kCZZHRRrMT540XmoE6OGEb9X
zG4fhElnzzIOxQf0apVg15H+hl/dw5RR++Csq4R8LeEByszcqXiGgj60/it6JNME
Ak6ig8D2KydSxUX2VzNMAwneGySPR7diFNi0PGwrFHubOVaUlU9EYUaGqh993MO2
xMqQb6xzaZT2rwfSeqtyVG0ggBvmnvGn5iVOnmkxoRkg2b9do+oOeJQmI5KmQ6Bx
k138z0ARycb9/+eebCpu1EK20uZptVtJiP9oSR8CQG/DgMCx/ni/iIJJtiQWoK7r
DXUay7isocm7BQYZ5Q4n8VQgqp1S9J0VbHbI8emrOmfn81Vt+/VjYoM0Y4H6hTwY
kodoeyoHhOxKISCMLUmW5d9ns3ua2CFpvQCz5AlPBqWvQLT8JHR4aHiPNGGPuNB8
nqer2REarDr2hbBd973FSQoKusjLAyMGU19Ygh40NNXWqYBV1kvAOYyZEgG0tqRY
vFRwfVkhLJFyifiGNZho7bmaYWAh2yAIjgiHtHYykyzGQygTqrTVg9PHk5mhQT+5
nG6iuMDvP0pJv1SjZLWDAZspxW6oHbLXuwy/2bpo5t/ahhjjQqWXMelM/D0egJ1f
qxyGhGpAf07NMIWlMWSdk8IYCRvjqPyhRJIbKAtJC7JXo2Ib6vlhY3B2bXEwvBPz
pHH6EPmh8scm2xkPXPwBcMoyZU4Xcfufws2+3JEn3VIMyAe1Cmn5Qo+u0sJFr3lb
t2ITCqkdQyWlyUuiyFG5HxrQVolSkWcRZsVNF+Z9BCKxvrbbCddqmZGWJ8DbrNoL
ctM4AaYjNPhajvv7rNjC/5+FpwRpjMl2CXRTXcQ9vJqRgIWF4fFDm/7yCQuFWGSB
UHxwCahJjBXQIf5SvrMk0ohwgreEsnSdd2Zrx6qsLkH22kUbveg/MbgZ6swlzLRk
ZlzQypwrr8b3sPxgPkshWWhqq4Pl4/HyPg9Bw/a/8Dzvn8ar2h2aEFT1ut4ljl0h
6ZVi63ouhb/TZwHCmKIPDi+dGK+zsFWjdUkFgSy5aGkoac8GAR6YbzGPauscXtXt
p+qKu2259SpevExAsFbNTAzSD1vPCUFKClazpt6Wms7yH7tUFjCZNqOZosh3Eo2A
W7rxkInqoVF65pQ5Fn/A/0FJAtKSMUPCoOXGpnwbXhH3d5bY8YDAQYDiIhLxsrKN
2/ysm5FtT5MYbUjhY1+MbqVlwz8Zq7ATY1IHrb+DAQNchUVS0By/L4XW1DRxSU3V
ohHfaGb/xQlzlv0DSwnXozaxQVAD7oDZoc5xVOGoyUyEGeWU0nvNKUHyv+oIPfAt
jx0yJyXRSgDWbGfPdXQzVLg+3Q/A8ONrxEL806ah18d0xjG2T/aOX9kIreT2ndIp
ewAQEEpY/VNzGZfch7xcMHgrl21Fx5cKP69wt/eZXpbzScitPebkGo9p1YtWR/p9
UgVUF8sLT7UOx1K+bqNYjgkHrIhoNr/bjMspgYkQRiaVtMp4xjfMY/QDbrMgsqFa
LUVVcVtCvA8fGA2hkKLTyG0/2l7BFolzsqC0vh3ujeNHSZAceFro1Omv7pKGBbn3
rP5rIKAP2mn2lfy6F3fIJ/0oqiJjMsDBNU+HHb2+HhWNLOgbmhNnrCJ7hTAAQBhp
+Ap5c7DRJ7qTz+z3Ywm9jznHGKmzXj7VZfNuxHTPbNSfH8GP2Qi8rbn872RYVwFL
I+UWqzFX6+R6FMX5gaQcd3zgSrb0ZNPzK6Q+y4NSwGoDO3dr5QJg6wgPl4uXKOoj
S05TRMKcpGVrq0tL1onRU00jdsanKOzLrvBERB04Y2bC1PWgtCnnD2buHhJ8XXUQ
G4njF+1sKIxKltwiSuUn3liU9GVnZeBW7cgp/2iAS9TQi4q7wJruamDeB54B0RlS
0TWF4N/VnD9EvmUmuXx4oQ33HjLIMqnMChuUJ4Ka1CSQFdY+OcxgY6jj/MdKMgSz
7tLjguisOLrNEBm8og6KL4VTW226gMDNDxwCIxuhB/zj44XEat/A5NtuQR0j3pjh
IZXR1aPMma78uYuW7+x84fILwf3zGGSarBogVTv2kkJ+lAXmBWXEoFFBx+IMyi8w
5iXIKkyZjVUN6WkJjOFPOhI+toPGHqivSIEcKgyb0+4KAii/yCx9uNlIn6iKaY4E
WvDytjGKdE0E+VX0Ex+xFMGADn0gDSd6UtzxcQbRxQ2q06AB475Gfbm97A4qE9r+
uEq/jkmWyDqx4t2Zs7GXeKI/U1z9miQ7p9Wo36BDBDyX3C2S+PFvSihNwUhZzvn5
slZGmHotzZKCSsJ+KaT8a/4oZW2fg+p7junkE3N+4io9JGqwMeQOXDqSzu76Vs6q
WSpAvKuRuXkW7hD8c2dLKGnKtzKCLmJLxZLhz5GBVALpg3vQ8Zzk33BaBDw6Qi7S
6K2G+cumKRz+/MGDGXfB/hbNBiE+TzKdt3F3YBGkwVG4G2HRLhVY5MAmtGdTYeDY
kAb56gYabH47gxFauowF0Sks4M/S0nj87Xpw//3hG8EMQqSbDVzEbPXb04Nyc5gS
geUU3wMIUdw+B7CmKnAPCunwI2acjINFYlqZZT5GowqcTTwAJVs3Vhg7l0Z7oeR3
yZyIiCXBxQ9wgDsWAxRwModQeza5ReoxamBvNdZLKv9tqhBk2tBucDr6FklxoFYt
Ngq6uE78XQB8xDgQXlCeKKfkD2rvrfbNkvYsoXjP8QSZKFSAl+2M6fSK6z+INm0E
11l/ucIVZuWew4aIlBmQL7P3raUMQSEoHW35lEpgjYaB+TldzINxe/FPYED7R0Yi
yNXcDroVXTvu0KoH+fivp0Qhvst/kmJRVUtSn83MI/6ZSZyntSn3OI/tJGExb9e/
tl2wBfoqtQblB3RAzziBTMnQYfnS2oZyJkiaGH4ealKsLbPJPy7UOaH1aN/oVTO+
rcuBR7Ld332/HzlbKQ+V/dSa8ZF8GkI5YWARtHdIjuNuKjyKUuP7auV9fpraotXo
L126TYUasEI0QxfDQlQnz6cR1KJea7b/i0nZg41CjVnjpoJR/pO78DpLpZHIRRJM
1ERvSzgyyzzCvzfD9JkSW/cR/a0SmnXxUoy2hISz3LBiF7aM0NKBC6GLrFq981JY
rdU+NHms0N0YYF42VeCnZwyEHB8UpBhZB3v3NXcwNS8CkdvsPUMl0ov2iDeE7K8Z
GZchySERHxUT5aDxgetOrPmfaAKgo8h48Sp6GYSxb+DG3CDbNeOKzssHeq86VvSz
DQbWoKEXqiNKjAOXlwCfOXCYmCPSpI3cOzVY09t6GyohhfV0YpRsjoq6rht2oAdZ
1Rznjia89exjpKvfr5oLX5C6OMlaHbn14QazCeJ+Qcrj9XlmriHq65Pg1ww1SfCu
AEPhC0bfQJoyOOaP7Y630bBmoCr0EEFKvwMFiCHnFUcz7hCiyD2NxsC63I7UQWPh
CKaoOdUOZE1hg+SWnqpYnFr4op884AY47xh7m13Ggfbh2zuW3jYztYEPi6XfWwqv
KDmvVK454uA+xL7fALEKPjmD2AbZenH2Qcmm/5448NGtf2ByJmAv/EDGtBnOiDtH
tHYTS1FcJs5uRGuefFzPoR0/dmdPGucfYDzc+Azy7AT7CT+HPwxfvAIzI87079jF
glD4C7/ppNNEDl/RNcB3/2I55zvQmEv0+OenLb4pddWqRYcIt5FUlUudLL07D8wU
BoPP1IhkhhYTf59g2RJ/7F2xn85N/9AYjrLBsSxXyiwZz+yZuarHDOIRoRi/a3Th
QXbqJ6GDa71ltNenozrZnkjirL1GlChhYam19dCgfxOQc05bOwcOImDP0+smK3O1
N53z4ioDkA+5oP51H3AUt418LXXubVpnQyhMYEsvG9/j6+qGLGuNoTWnKjYPHH0x
aiZue//1ceOMBkoXUKRE1bW+rONWCCC0+6OI6bS572lX1BTSDeqojffRQFb2BcyP
+8IS7V2r1EG2jmQXwPuYghM5oFuiJO2/35Wnm0tRDu3bV+VphxXhpPyyUmF6hgRr
dEO3fZDFvqp8BAYTgJ8XKTiuk2fz6RXnpBSmuBmeopxEISDdvSiZhjEB5ogkGfq0
IDrVeqyMU0/VJzj/4zmbxFFAZoU9RajyocTSIcqAkBeLJfrvGqIctk5CAEz+tXen
Mt3NAEh1OZoeJ/0YjibrxTfg83i1VkgN8hJS4g0qEkJDKKC20W9th/Neg1lUCmD2
DkaneoTvu9UB0boPKl034cWoZBHC1JO6+E7fEpEIwqLrupAp1/uhTIuBSM49cYkr
rGxBKto9HzaUeY0JDE+RIYMKac2CVj0zCoY4ciZONE/SlS9hLkMrk8HzePEInXsi
qD2HIuxbhCYQEpSF8OF+G4L8tZnt3TIv9D7hVV2WRDi51+D2DjgNW7IMASs4BYox
KbT6XUNfNaM6tCrQxNb4FwuhbePh0ICDH41Zkc9yYGMadPYRMi7zuZ8/COYdulyC
vAOjHpGJDdFMOMZzynbPQadMAqYlBIq7qxXhvKKiJ2kQlBSL0NXog6UDTPwnK1JP
T36Q8viuQPpLnqhrkvoJRejysD7Js0NE6umDvUMiqv+TpeI/vDjpXoOItgeYzVaF
e+EGdOp9sptJ20QA+rm8qIDWtoaHYA+m5s3WoRYAYT+mr11trZ8cjd5swFDl06E/
NqNpJPPa9Rojt1P1n4O4yGf4BLlxEm1aPSZkZPHJFDmJnoewI5wjAvXzh1Oc1ze2
SlZobJ9qo9jjFBxWFPf2A5zaakpsROou1nmYP51dKDdXHdp391NJurnl46pJwUqV
WUQu/AcF+GUZxDG8W5HvuwWADYQYw0WPYOc9eTSVnMQ8W8vupeLfrCqb1gDN/kKx
zkSM6KoR3a+dwLeQ9VV/M5YHfs7x+Nf9MmCowMRaqqnPmquu3b/5SLRL09sN0+Lc
dsNM/DnT/AAdsHUx17D+g1QHo5rcz5tty+23+kpHA5G20IptPB4dSuitmUq/6UAa
rnzOaU/Px4A53b746+/uX/qvbIvhnb3rsh2ogLB3+4o58zf18U4GurZJ6IIchBME
LX45TRb55ctgK/fPrWFX34QfGiQlTN4/seX0SyQAIMXrHnkxazSSZLSvm67DQjJh
5mEPuTHGOUuxRdV7TklBJmiLLJzfXT75pte3tdxF8nYWd6lyYpheQvZmuEDedwUM
iW1ATSpzgGtImz6oydHRHv81YCI50nL7VPy/VmchHi7Owf1Cyu1FGk6OYRF3XlrW
xmcc69ctQs+cZMi/eV/qL/MYzzEgMKpYvdiCy23hEiKuek0X06V2ZS+wyd1Q0FjB
wfY49+MthZfkowRqHjp3Ok1a/i2OQIG48Rg5v9PXL/ZHovsJyA5xC2n9ayjUiTCa
z1VnUlIBzfcjZLoK+3sq7iKgbbjdlAiEGjgtiqx/xyHMYU0dTd7Bm994K48gVxTl
rTwhmltj0t1l3V7/Lp92NUw7BPaJtoJXZm83cPSNKS/lzrrQGwoIpiJjB2t8nXmm
lnAYYWs4A9V6/NCg0oDLlB043SPAK0PAXq5mwEE/qS/ohr0xwWX0xHFUX4q6XHgm
cmDma1PNM2Y6JqeUBrLE/KBHsmkTdtGkzLJJRo2ipDkCC2CaeK9fCu/PpUz+JpBF
ub6NhXaUOXzy9JgvYGNGxAVc4Ox22fDcXGrj7F0GhIVWqQA0IblYbZouthX3kYqn
eN+7OsUyROvnKAJ+pqtvbTmPo2NpbJv7wV2HP38uHtEs6JhZEaZW/Tg0ibiJJZNh
ZeduR42OpkeQ/hl2X5twq8Crskq3fn3XiCeTjgEFW7TpQglV3LG8NjyPfh0IN42E
dKD/6Re6MBPotnB1Eg3X76nVQR3tEl52avDUzJmTI/UM7oOjcq8GhCf3Mg1FetVi
trYJ73yxUEd3OWNYyD67QrpDX2hVbYKVex9ggeYT3Xrw9bhIl664+LeOe3a7jF37
dfSlgPoGUajOAl0UgtIhlrugTUBMSoEHf5AzCLWzo5VevnwY+goBb9yrJiBtRqyg
VCaa0SE0tGJFHq23KtgB75BZrXzks9nMNxwnMjh+0afImXnC3ii4r/kMdGOxiNfC
9Ly5x8DZ28hEfJzL+A2qBRYxKMlRwY+EI3bPVaSGIFLLN4NyH7XAILlyCQzAr3p2
AaoqL6wT8qXH5nI5PqpAAt0rpBzYnX34cAEuAs4Vx1N4b3D4RrzRLGv0citLMA9s
xCw2LbI0H1mi1nW54W7WkovUWNC1SFjM3/G0sGCSEHSiIUxpD/9QoLiA83kBLpZB
aXCIoXkb/ylwsqzHAg+c56TvPyaelg5u4NNNs4QpNRVFj2plQowVNHndic3saQ/Q
ir7GmKCVhHN6QS9wwHOfK3wMuUuUnvqQMxcFe+EuQbiPAibrIPOY9bjVtfq2xRBo
WEOApy88IlVt1VOgnEDz7/wWVFaPXu7fxlbvqQxdTwoH/GDOv50fVrwCRlPyC1Wf
v/5QXWEHSait372JEbhlVLjErMce9/1hYLuf3o/mD34LcGca9c29++Ck0VkaAwa/
SuSUCXl2ak7Ek0NyEgh6mD7MnlZJw7TTUVYgER/cXQ2F8Dc2U7YSsP0jTtr0uZW8
AQ/ZM7AHjyJbUFK0QzeXbuc9ZMlYJrIWzSOTHpWMKAqgGW8lkefg6nX1jc6xvmMN
ivxgudOM1Cn41yj+x0z0/81+4roxK9CMZ8jOr9BpAyIFOuyS/bGCnBuhARBP6B44
zG6AViWt8Ll/NvDSjKoA1FOgBQGOaTzugq0LwIHF4XScF6g2EReKtxLeHonXmGPb
NnT2r4e5T9FByVHGxWvtVApLj+R5ItsIsm3kqD40WmPzpsMBKspzJ8kMf4W5ryD2
E4LZmN7ryVOtjPwCiSXoPrCvmPVapLQ5MGKkeRqIcomlHOyidw532HFsMTtpp3cv
avdy21mdAwqzh9uVx85amtMUc79go0v71ecyQ4NgdyBCs4igZCyaQGNAOmUcoi46
V5pHJQaVn6YzjfbfpKt++Xxy47G0oZv9ZWiZEngyDI/ix5q82FwNAJNFKkzV5OLP
oAfaAd3VpP1eNamLvdU/ox/4Sn91hqceeM+O6IWojHIcVtYFzyHugxtc6CEAMr/4
tubrwVxY7I2iKjAxvoxi6HV3jY+rkdO3r2ZfWG223UNTtFbXuXoKtVzOgSzkiig/
7Qycob/kdULUpdnVwSAstRW7BH6sWhJsnXrNzlI0IYpsKJLqjvytOaNZDDlsNRn0
qnU5IQjEux5a8p9fmBPVd2QgWoxnVR47q7rMrJk/EuN64X6ecISF5mRsYKG/P4Qp
Wxi1e77nKvHSOpMGSe81KaezSyQmZd44J22gAQywHc70gF0L0zKGwlBWVZ0eGRu9
m00afJlJd8uXYL1nrduQ8BBFlaVyNM7uKZVZ7pBBDFH+lYkpB/VNYFkb9tJM6jxT
HSIijFUKeVGVeTsTUV2I0mir8C4gYfm8jn2m3or52Y65T0qKX8svH2mchH/8VVe/
A7pkAJpxLI/G5zA20gwA495nXajbhUq5IanrhIKRGwHOqjnIz4lBpPQcOvn9mFqW
Ay+gLKNCSMVicIunXTIAsMvOtINNmIZ3SzNQYMBYgVkQaq/Ttw0EuX+4iuPMqc0l
Pv9Z2DIWis2e0jw3o9a27cyWAmi6WYK/QWmZRRa4fiCAZGacKjfQ4GOttIlvTtsC
4Fk7F9dHL9AWnl5blXXMOAXisz2NsyISzErRwVFIXcPicukwjIULcPsRTnSob0hI
Ja4fhElyicVBpf3o4bDmye/gTG21VEaaEyFP7VOKezAnzy8O3K9i3Bz7i1/I5KNB
KHOkLTHET39MWObmZIN1XYSSzaCWKKogZGdu0HTu3iHBzZIsVxQWUuF6wRSkayS3
35Vv4N+OAV3n0tQ2PUtGAHpGFcFDCebK2lZEt4YnPYsvywTxWStmFL20ldeZ+K98
/KXHwILZAeNQM/noEhDdIuuAZhklitaqCpBhMQUQQrBLXw3PYMAgMbNb7tQPP95F
ve2326k1fNFEHKwb4bML3Z+CJl5DsTZA9Wb067BPFvZGHJs5u4YCONCeppbN+JCo
JauDOxAsZFfXxVK6fatmlAatdgJyx1k2wYaDV+iyZW61vaCS2cEIAK1Ki3iSLJZ5
V2LkTN60r5HASz51ad8EI9bmPEQYtccw++KeHZX2wSGHxjxWKz+sSApnBl7ygKsC
Yuq4SGXL83aD59ctAZWsvoWgh7YfDSVsawBCN0w+kfza0ilNUmTUDFh6VVy6Sf2g
849qJwnHjXrLDi8amXZwZkkhSMy++jjbswbUQWIF5iLRQhnmvb7WdinMtMVn2hO0
SkNyO/CeKRL4uW6byROxSmY/AavadaMyBPVsac2bZUTqpfMO0YQCAp3vakl96L1a
2uOr0gpLAD+snB8bhxomLwp2g1KaKw7/oCNmUD+LW1PxP45OoLy0Kc59B3fB4TYK
5vQqRuiBqukPHzin7PTDHixnlpqoz8B4TC8Is2sharwb4tBZfrLWstkzIANW51y1
XJlWdIGRB1AcSfBq52DIUitIO5kt8EXIWJLGL0WqQhK7wAaUwem3+hF7DUBZho+V
thmLr2GXzyPkK1CHe8q+K9QFdJgML8a3Ix+uQop6ngt9Zpvrou5YqOuIsNr1dp/J
NUgo3s47wgEl7A8xHxvBOJ1Z09yVGL7+6a1TQYnlJkEMMVGhqRKz1ikoQQCgRmtK
VrJI5Sdnlcx4m7ODA4eOVLVUcwyfmB+PPC9kDpNSPV9iXMajffXoviQS/Qq5ZQB9
G2EBkmJzcBaIYgZVYxWNuscMX8bpt6SSK+cfbHV2qx+TQL5U/Y0qKLF4o72zM1Mn
eUS+1zzYgtYF6H+BfqdweRGMxki7SOblzDpFFvd3iFgFhS6HFZCgjMW9rpi3VU2A
SKz7MZbQV80OzjmkaO/sb6c+/qevYNgRNa81GmxR3JaCkb/Tyqy8GEzU2EGVCYM4
g+VxiZuTLUvF6z4yE5ehzh28Sg9skZIEdgBTwN66jdEGFsTtPoZ+k2M2PE3edyES
oVf27IqI3rap/VUicqDaGrm3D+GMR3WKN9lhBja+AxVqjEF1C2/iEF9dMExTSWwa
VSeH88jexl1z1Za6gsofCMDQAvLWO6dc44q/hUe/KXMsRWpE+W0JuH74caGcW/rq
jKiFyTVRd0EGVqHYWbbtcDDNHuloGfGgS69XruQzyYpknTC3nRbtTzJFK8grKA30
DoZDUsGklgHThhm9bJyideXhvW/OrDBXa0lxFt222d13z25xsvWOuKARLiths6AJ
ZWJ690JH8pUNSWHhNSHVYTViGfBqw6GfBKc1f+g3lXkxoSROJlNpisbBV0JrXEKA
MtS2kfvvX2pbKmGzyBNWLZTzi82nn+rHBay+ZFd7dT+osZL8yvmJEJ/g26GwJ8ug
8uoBEZeruR8nFtKM1f8p1+eiwUCkGxt3gELWVcnHFCDaZvmBENKBBHuEfeXUPF+4
gMZCsopPsL4S6rEk6kNhR9H0t6cBNjrS1iQ3mavv9Bdd++P0hNcJP/jrZZASoC6q
Q4O0My+OgDtSreAw9s67Xe4bFVa9jGylmazGiKYL5m5vh42xsyqBFKLTMf8nOcGa
PjC7jjtBLDmQKYnpos3jG0EBGEA3UgpKCIvPdOcfw9Dw8zvfpuCOwflQ+ThbAuU7
Q+81fl6eFAU+v8ECl3jR8vTd7ImklyT+LDuNL1M0y8gz2GaD7jOPKj624e1oHzvP
uePZm7U9WFxaMY8qoecu9ANA+kD2OGkk95Pm4lADJwCpoUQDZnmhqf2+o65M/qCX
6TEM52yJVJqdiySQkERKTYqe3+3QYtK/EbRcTeQyr3IJVMlka7Wro9hIv44DirZK
7ASUkEcqtiz+cqDQ5UI1QSolnQyZd83++UpwbTk5BtbkW7WOGZ0ZwnvDao/DirkM
baKTJ9HpP1/v4MZ3YqZYZGB25Po27z0dJXcGZ9XbZOHgDoUbfzwWzN9uLYulif4t
sv9u+u7h67iqk74y8PH2xQ/Da1x6B/u/Ak9VwbadvuE1IXM80zfpfUzJHomDlJpf
coPbvxpGSSUk8K+j8ZYSbpWQMS0J6Qyc3FBpFU2/yVoF+CD2lMzoqugC5l+4fy+O
S22HmzaLdvJkQFf0FsbtAXHYsB8AEq/As+rhKP8rLZJOplHfLZUq1IrVc3BOOZRC
wOve5IrNoAn+8sYpygAs1Yy6/JhxMZ7g0Y7oudDm+XxJ7kYJ+5dtB/AgLHQ9nNmE
GO7oVWNRQYdI8akS2MV0M3yjcdR9Tpi4NPqCm7J004fV4nG89+CA58rC1iC9kjIl
oasMHvEYPoTTDevXLzzV4jzP17EB0SlTu8NBQzq6drcBIEsibf2OjtYCEb21Yp87
wjJKApD+xeqOF8bagKxEhcFeorkUrnapBfyU95C1Aucu7tGlX/nm3j1WywH2wVaj
bAWJVur449KipM+6zoLvXLRSzf1hwQVUXt3INn29vQlq+pkQ5MP8rouk2c6O8iWW
1vKuRFK/4hfxbWr4O4Kfrh3y/S68m+ttHAFSdotC5sSU5mmNOnpBL+EI8sQ7vsAF
jC+MkF8IKefH2+ZPDV/Atts+NvyxXDrc5N06r6ojsqDpmfOyCXfNf4wBE/TKpAIi
KiU7kKm1Q4+B+LmwpcaCVdu1MFJznfB6vMACohATbbzaI7YH6nwXnVK5L+Iv2rIX
ChvUTUq/YSq8D6PntcsIx9pvX+JzIOjHnFrNVbft4jsjHgeFEickkfvKLCvzahAe
2cvlC8ifKXVpVpbOxo8+OcUNUsNkyL0JybIMoW3HHSwUCRYmWo96bo7R0RmL1qHj
oBr6S7bXO6cQ3cO+veFDQfI6eegVzSHuIeVr1qfADNq1DWhxNH30lI7nvGE4xsYZ
xTD3xOIh7R8u7Ry0YctZ/Kcz/1xd+vI3CXsjzsxnz4TN5qEzQsryKPHRtyIkbE6X
jmw3D39QNzUpNqC3aEOE6G9CH99TFOaO7X3lvwRB7PyaNJfMUXlsIHiNqWTnGcRZ
iGqQoWA/JMgv0C1HNmLlR1THq9Wqz9qwNUEHN6wVRhSCPl2WkABK0BteuxV1pbNB
6TYqC1IWIs4jxu1NbYSyCzHZfMydUTa95AwSHgebnu7Ee1+oB2U4Q1wj4fxXhzKX
mif+w+3yYftekmum18G2gxXJ02CbCu0vvxrbdOJtqFYOe0gnGHV+9CnzE9mcc2Y2
mNDK54uUh20cpq2cIT61gt6Ep/CbB8WJF8/PK24lMhrHvaW2/lIBl/8SVUX/7Hf/
nheaB574ZLQUquME1Fha9v2RkAKBBPA0Tl23tlW/77MSPcrZCKko7TkJo9fn8D9H
TfVWFcw+r+oW7PG4tdD3d3Q4lKEeOAtBHBLj4GJ1M8sNKtsPtnkBB2+hfTYRMTBk
D5m0NsRVlLgJSXcnfS+kQBc3B7wfGa+/dfhHR3lolBbIjn3QrJsthm2rTqV/UtG9
ksLFd2xrTLzEKV6iCHUCZMcWhj9ecIUAejhRrkGyHhxd0vQauQTpizr7paNcR2Tg
bXCxk+QtiSx6qJTWaPE5SwMMABiCJDWCKKcw6xULMbd1Cvee2y39FXdLEipmpnhc
tsCmgYjb92AaKIqBrZCCnAucQnSB+NDS2PXZyhrWzMoIW/EdHGZdhJxALIoRkLs/
84yyqElg3DbQFlNFS59eN/Tri9VrTYMhPirIC2AgL+oeP1Ssrj3ZhlhbNw3FDbRt
DbKm2iezMsXlqpC6wISanzxqWP8occi+y884G/8f3N4GmbJ7zTULpa8QYvYkdq7U
k3Zemv8f/67Tda0pfA1Jr+pI+TTMnneD616ZqC5tJqRRzmSrIRlzINxi5cm7KtT3
+68ZpLn3M9uttZaF02/FSYTRjQW/vBrgxJ47qmzvg1xpiV6aXyFIxrQ9r96kZgLc
jd1Hf0cihdZub87X0C3TE+VwAtUHImgt7XoXsrEpWFhB74/Gac4UGi3YzkQziYmh
Fm8/8+EwWNeNheIoTFtoAfF9WFbA0G67rU5FRUkO84QYt901Y5HabGn+7uPy1P1D
aOivDT2jIzRVQh87SbNhmlC4eMqisbSGukcPFHim35yieKzVWeJHawqVmKEa4fq4
mjtMrQw+8MdlUbujogd78rD9+LFXskXdi9AYnZN3QL8s8DEit4gmuZCgP+AEH5Cf
tLBPgZX3i73acN5tbYZXlr7WUsJV3KZn5YBy2vHCjjMb71Nrtqn6RQj/aIQmlA+W
r0KfIYz2iR8CW8PBNp56WbSXsQU4TZ9dA29rqoMmI3A4ojWD3Iir/AhDNQS1ONlS
UULy50BMC/fGuzLhmkpyY4Czk1uitlquBi7BS5IsIMSSq1gtNhLoj9mecn7wD5Fz
5GyEHrlqWM59fWIYq5j1Ce7xH39lb4mqV58yQ0P2MIZIHddqphwJMR+jzt+9B8+t
0HgHsee/lNldvcvg6TTxDy2q23oNu+1Khxmc8u2hzd+lEI8dZ1GJhk1/IQ54oDEk
M/PmdBAoYRgg080ei7yjY17gwlFq5z0Az6ToiwepoNv4xjWFvmi3NUBaHo/thUU9
dc7RvYMls+HognYxVt6IjZTSBPUsk7nJrNge3JV8Dde6TpsYNMkMzXrGm8C13gOL
FbSM1K93gwYLGa89dQy2e36f2jEdHo0urZq3gkadqMSc1ajx2lydao+fX4uLx5tp
kr/Wnooz8nnibG+5+/UKjnJWLa+3aJANacwggZKyEDjofd8nCdd+3kz+N6bQl+m+
Fi1nJJTUhJlhdks4PO8SZVA1p1OYKbh+uqsTI/QQ4s3QXvq3pnO2BYCEdukuPRBG
DC6B+951/SC4ugLbogxk/NfMtyMJunYtzuMBojLvKYEqRPZ9ztBUrw8X/7QFflBo
1Gt6P+knHa5UVghxmpyQ81H49f7AUyvjQ72BR4bG1LDixJptc9lxGlkXkD813d/C
HrzVF7M8ghfOQVIxrqkK/fuN/02TlYitDJPniJLp72sptbusVsG5w72JP4UCQ5fr
Qu1+eIBQO2cmh7Ij7oq8uivntM/7YxJ+xXAWXUnHiY43XWhGHC5qYM/HvargrnE8
rwM5hT5+pistuwuneEOilDJtGmh4sYgHPeL+n0N2BdY41w9xfb1Z6JgQ3/EZGkgj
dGsT0VZ9un5lUjO3UToUciTVXPeeiWcpEGuIECBOMRvrq+6x73WvMe8VHLQzp9/z
+GXPzB7QAk+ntqz8D1GpbkOwFWO4vl53ySTZNgwkZQmJJM/YYhbT5fppaoGMDBfz
Z4asb1JRao3GNSpF2ya6rh2mVpEv+vDKucLffbu0yp6QZttKthLwMrjERH+FvcFZ
k9ZkkR9gBRiYiotFlAIY3BFapxUBysm0u2MzgrwNDrZnrDvIZllyhKwfVwKk0vY9
hMxDisClwARAidKxhb7XKTYbLAV+SUb28z0TOA540v1c0usnV5PC6TKgY7CQJ+7R
AlpH4L2kk5pYyuVv4/6BpA8JH6CtNR95xjmI4A/73O169sJzSAL3nt9VIxUBT8hw
WTAeu0ItRWop8aulKaBD2GBh0Yq2D1vayuP3n9fVPcTn+ADTQT9DS282u+go2tHK
I3w0yJetZL72PzHgn7X+pNgnyrtFlQSmgklY1tCBUDCrLOS0kONtd0phjhglYNgZ
gmAR02ZcZaOym3eLKmtrUkXmhpg4zm80HKw86cZEQd5AAKqIUJPJnuJXD6zPotdp
Y2BqKonsc/7y2drg/6/HAnxLFzxFO6TnF+EN4xFxCgOmmk5kRiiZAZLNl33T2pbG
C7AriDb8NSWKZk67VsXSJlpEqcmhTrz595LU4qOAeD5Qdt36PrcllGxsylbP6Fcz
qaH0MlBUvAIrv0xWrrsljqLIsVrWj5QzOVYGzBvPYAGk3A+FI5yG39DV9ti/UmmK
hFymIZqN9EYCRdyUxfi7u+NJDQX8PVRqoFulIvo8wHRShExHixBddlCD973cZMHs
8K0SnxGkMa2svSPn0QUSjZ5BGuToYk8WFxF0IpDypG/PtIB9p0j1OlDhXrdOPqam
VM/1L1bAG+Q6pDKlUDv0As4RDiBcOQA31k5OldtgXcwPydqsheGQXPYVdkyb8MWT
n2dfySGNHeQCZRBszlvquAQbKL45L8NO/xTRcuBFhJdRSCT1ZbnsOcbObWg2t4TN
+iVLlxtWwIeNC1ojQoHOVbKGKLlvlX7170UyMTLiijW+QZ5PTrAJqTCDCTaoJhYW
KhumuLkDGPjGlWFiWZoFYGf7cuuzDCO/Xyj7ysaEERmGyDXt8N+47onQOATfA0/u
4c6GlNJMowGngbgih4kjZ1PWWkp6D69v7IrHkFZGChBpYEEdC3tt7y8MbiL/RaLR
33mCL/ETr1nXusG+WOTxaqHNN3Yao+dkkN5bOg3YPAU6YNYCtWcosXNTlHX9KcOU
hEyyIIoCv4Sz3mRHO31ihmdbnudApI4YX9e/szn/1Kwt/x1Y5QIYoxuTCnRTncjV
2ABmNIQTt8Ig3b20MvmOemMa+MtNZY5YyR5tCh6SWRqCXQOFYH7aJR8pOxqwO/xE
ApfviI9hDYNnbY45YU3ZrsigJkPFaf2Vrn1MIWNRasJ4SRKqslEcGz7L99t+4mGz
x5YhoK8bDSiamUD0Ny9Bs2hudL08Mpphmp3OTyNmLHNyyEIkHqhPlD/4tJ+d/Z7n
N0tDVR4nL13H1qulgFa/ARBwFeFDWrN2fzSL8OW7krFURfSZw3aNU9WhQWvBGwA4
8OFWYjOUZPoNSkQIHpuHcrVLhec2IkQDRM80yZgocbsV748imqeRcIsek0SEUjlz
C1SW4Cm5k/TonUVe8Gp+2oqkSHIHA+RtEe2Vn9tHI6JkQQIhboIEX6pMHSg3KJRW
Y/QaW1oD6jM7BznyJ9P5M0t1zytwkNXJqBkYvszr2+eTWRgQbAwuAGNDod5k+/HY
d4SNVMDU6PLJQR7TVXuM/4Dx+Y+LfDmrvSmT85S+8NZCjOwu2dVcmQ/ABHthUguO
xvCXTfAlvxeAf7V43ROVER9AIUKY9xGHiyTjuidYQ9KYTgzXK2q+/srklcNhqPx3
9+G5B+//O7PX7TgJsxeHInZMjo4ckJGq5Gjxk1eLvC7Ib3lX6yFSm0eSue+OGt9J
LUHhcmEVbyiLWHWelUNT1OyO2eHpRhs08bH+L2pYB+sHLP9HJ9cH5liYx1Y5o+f4
hWWZyxuEXVk1RGWjXZdWdzsf0ijLbYH2h++4X6imVjrtHcb9c43SXI7Msk2NgFCo
qAVtgNW3Nn/T7fYfnVUjtbkBr05VK+FqpqFB1fH7YZdSjIv5pGwep0Yds8x+Sgqg
YCe6ZlwmlcObazlwWLMCkJlHiS+kEqlxrbou2whlOo/I7eSSA5AS6XSLWO7pEk14
2Poh7vzD/T9xiq7Xy4nBOggJ+pvhSQKqE+kwRiAR+FBgtk/HUEBGNYctuybKWOOY
sZpg2Tw112gKlFDtlkE8/nM7SJg05CvG3Qs2QlsmozFThzePq1/1vrYrHp4ff+wg
js+bixR5POBSH4fCmtk+F+8WPJ1gBvXEv+yV7R9lPZmshwPpaAFfvghmF/A6tWK6
lc4UuSL7b2mS5HXxPe21VWGJmt3AhQpsjRdZ79Q+4adRVxB/p8pzpK0a4DLL8qEO
Objn472atM6vz8EwefUF9KWvE4F7+bvfmQky/P11r9y8cfoGiJk0p1fPXv5tIape
vvrcftp97Jg2lc0qwDp2pOrD1Wn1wIVKRtEFOP/dk7vR1L9K+Gzsqol5tC0kSdYQ
4njScnzkd06CKC90+r3RJi/JCMJmuw8q8xXnmYKMIr1d+CneNYo4BaH4GuN9jHeY
InGZa4Zx24lO+59VNHpkqR+SWmhHmyTBdqqy+LeiYDKPxgU6zZFfLMQfk+K4cuXx
B+l3xXJPFIddLr/tFBdi1buKw2+N2QJ15xB64sMje5qasXOXn5HhO3xxXfCZjkv7
uiknAKZ7rTgqWtuYtJMubAGpdcb0Ow3tt4P4+FQFLNEF+uaQJRLkXR5CKPxmPRBL
ZT8Gng4yUk1IrVYABwCaMJ0Fs3zGcM7vcLBDi5hXodByzhKvfkFboSZkqRmg5+BI
pBgyoPZKLnT8eSmoqxdH9S7z6BvSpM9a/1cgtNn5k0gs4bSld2QVNnao46KkSwjJ
Lhik1KxKh8WEt5khxP5IfvHeRXkdW5KdPXmbMX4qQvQ3e62Lc37/sBJ2Yva0pcty
rmZ71QDkSPBPL11sX2mBdrciz9TsC8DbNVlcEu3LMo+ctesFYC9qxdYXTT9QyS4c
iGIaFF+fSQK+04azasplGyUKOXz6SBjvlxgD7Y4DYoLImme2A2WNGXrPQV6CE8qp
tCi2DgfSx3iOux87DDkFAPdtywBj9rpZ4cBPFIu89zzs/aVhysBc3JloTyrmc9VM
i7Qo47C99/wumTkAmtNigPGWAT3giQOrNYYx3VJ+O3c30kalBc/MJxS5OVyusYUZ
E8O0jcpWB1KnVxLKjbxcDti4+Y15Igj9wgflJxu12XIZ+y+sOqQHQt1zbxiVFOdw
I7GZcfV4S+d8j9VUv+tLIbM1vRAbOw+PSmVq4BW2UKOztfmxT7sTlqCow+uheXuX
yB/IEwZ7pEDA2TjcHKQQfrEiN7OTvuJ/6jfMPkdYdttobm42DeN7DXg2JdSLZHmc
bn0mj3Ttj341kqTrbYXByRz7Y/6q1c3TlnLIE9BA/SsZ/ZHp8GwDJFDQ0h74XXaV
1QEQyAz72EgF990ZvRH9hCRw/pS5QLDlYOmkTZvJ4NKRwFqSn3L9Vh+IlzRonmkb
jTmD64w9Ku/VgyiHcuurKvIV7kwC24AbqZnDrE4lVP5P756Fx25x9J3TtP0L7NAw
oU1yTam3GkyeTLmqio0f2QqlAxqiqlvPeQfZBBXEOEHLSsARxa8akIdRZbPRhAp8
ekqdYVY/EiZLIP4Gt/HhPCxJMt1Tr+TYZJSH6fGV6tDMz70u0NQcZbQcwXTztKoC
HLirrDQiZ6bJg8Gs/SxhQMTm0ojcu+MyOSxm35HWI1xPf5g6mg4x/eaPcc0QuK8g
dCjeKSOhSwyUPy+np9TpNDOGxQB5fzO+TBfkzMQ/cMR3OIQaJQpOil2a4ECFDyxB
vvCcLwTKBT5Yoc01hTv47FSR2iGADNJOSvm8mQ+LfD8idpWNOQTerox7wFY0kiex
vMsjMgbijW2kSOfgu6pYtKxace/Ve9/Hs+ixI9Jq33ObFxnMHEoSRlTc1k/cVT+s
JG4gMlYbSTv0ZMBjm2UazD5PyxziH5UA6/V3iflE7Fg51NFyed55MXT+VnEYSBza
uP/Ke9B4sTymuAgnoP/EFfrgwIMJIf9UqJpqf4BIKtU8/GBO8RGlIt7JGMz/KPFQ
FYakZdyqL++CZjPa1uOqjAzbe9HyDelXeNnrnl+DUhnFJoKYY90FUkSDlpENfr2t
iRPSeCN18NfpgUL/569ytPJRkQ8RmegEbw+Rp7atCs+T62tXw1HGqlPKyEYGO9QQ
diVVogKR2NhnxlBA5RD5Z3alC+4owDQoKI5OteCGpkOPl/pIU25gBh+Gn1ke1o4K
Wa2wweMLIGD0tNdrzbJjCcQ9Gm5xgnuIRKG/CRyNiEXoa9/4gmYYxaiPs+quOzxN
vjAlUSCLqf0blbZWJ79MaNVoOyrHGqmIA4L2tH1pxuirFNxzLmli8wBE8Jhfa600
MpJ5mP+MEBp9SGcX65oN92bFEbXL6CycSERWQMEXNDfE1YmEa9TTPz/iLqKk6osz
YusV9zbffzv0H+/QBD8JGKHV3Rh21m3y0UYQUqTv95t/ojoXF5hvBzjZgCxR2swF
P0bWHTlu2apc0jfAux+TgaJCD+EeBXjF/ZJomWT500OGoWIcq2lv6Y3ru0iN2ICl
5MzHEOS2d6rAZpnHZYoWDxGHbdevQsttvlW5KElj6G0IvqTJQaW1vATcDP7r65gQ
6TUC+cwApQFoRIOJteCHFGbfzOCWS1Ms7vmoRedJQVHts7r0CtwaYAGHv1Bc1I8g
yzPB8gAyUIh2Nsa6g0zeIxKNu3ORBlSyHUZKZz0mHRCFvy6sm0U49zEguNZI+R0j
qIh6iQwpySTevo+6Nc4QqMvOUhov9kQqq82V/x+nbfeJxA7mCma6WdDfiZxk3mD9
zZXiavyU9dlMorGFQHOvHqU9W0i02y5ovgQtGNFmi3w9yEmRQt+DOCtfPUvCHyvF
VllufpmNnocsLuzAsH+vtCFDQcOrIiabt/Wnq8yrO2ZlOL60IUz/TLOvGPHWQCB9
tEbpv84c15S6en+2LPnqPOXOM9L4pGW0IpGXrIScUkZwbB1wjPxIngYCJlAV/Xxg
Xtmpw3DclqYVIYmUwN6rZK+7uwfs97024QqScap1ll8oJsxQ7UzwbZ6ihnuMwO7a
W9+hiewrBFjau1P+D6vAvVG8krYCe/BcN1C/cX1FJWbke/5M8lA7AKyBKpFSc2DP
vinz90+UjnVeHCTi1OEFCHI6GKBLlQq7xdHYll/zgtq9Mxq+TCZmF7e4t+aeEYte
GTUSI5PYqtxn/x/pLe4qOSkZtNWTHjtxYtsyf9AZb1EZ1z4FPw0Ndrcy8+rhJV0X
m/pp5Kgb456sdnY6WpQo4HlmgA0YrKbJV1ZsZC2M4pDXvgy+WaDMA+4MtU3QAEq8
i4tyrZEgvehBTHFQ9+o4yHYvBDEJTVb3/29ArWaiHKxcNnQa8SVCLLIq3QLz4VMn
5tTtR9jvTtGsGpCze5+qDUsk+1Rm8NwLt9NhV9grp3x8Jjf1eSB8tALWzznL3KBG
0hV//xza5UIXwfIODywkIQMWVX4wQ3S2s01kkXZ0IRydUE6uB+9DAm/l3NHUyHZ2
yxCE71VEkirP+r2GvFABCBqtYmuzHdNdi7oRz2Dah0NOqUtF04xNPBrA5AsaCizB
xJVdN75/xIZbUnoJUzegLNer380VKDmp1OW22bgDvy742TcQVNhbCQS2WUPlO2Md
hcRLJrtO7MuzZhnAjFGM8jd3JB0qUkcnhk0h/HY1dae3JMhbngFurntzrYqrdvTR
EQV/RBGZh0Pgo+vxRjJF0MlaT8Q5sPPXwuGS0K3joyvKJjUnuKjjK4F4AbpRR/xR
yxDrv+7uUvGCGoRX4CJPvqAzlp1OlkKWK2NTFmYHlIJxLpqQ7GzF3c1s0RWUsXUh
W3nqF9rtFLoktUbhSd4zZ7LRpJSsG9jPLLQXjZT+aXVWHHA7m33tPhz4PoDQKTTA
XQhOOLv1CpJi7Huk3N1gJpG2JaTrr8xl+MnwzUXpNhJwFwXaEWfHdKzOmLeyzkjs
bDxgaYsRMEZizZJYzN4x3ep/EC6eVh9JonHkYnAfxRI12C3nCa43sMTWkMnfZCOJ
Tf+YYD6+1honf6/w/BsvsruHa+0Ylp812fMZrukcYmuua3DM7XRgjtirGsgmGClr
DEj77wvMSmsgMnNSRzLAdMcwfFOco6fVe5UiK4959sbkNoV+FpH6Por3bgFGjJUc
dIEJA9iCUWiwvsYXVYTv5Zm2gvn1IdI5aMeNs2VYEM4Y5O5ZYJpYIuh6dBTc4EwJ
3eDnE0UrCP9fHYnm9ECMtJgMWGp/kosRv61i8ZMPjwZTZELvjEW8m+zhW+782L7S
TBP+TrSBx2qC+zMCpy5PBQLYMJeQRTay5ZoGlEdSkTfHVld3R/WuUOqqljJ+utAB
uoEOufV9dgmwS9wXGyGF5LzNfSMcy3o1EjwzFl62z6i8YJsfBWEMQ7ecgSXTOWZU
pquhQqIscW2ot6Fm3k37xDMkOeLtSi1Pw+TNTM71OuBZxBwZyC2g+MnDEKNiDxGW
JxHJQN+tS4XoYJpJEkXt5mpB1PM9rb0LK7517Jwr6NuXbk4Tim3FiS2jSSCrgm9Q
Dx5hDWT5VmjnBdjFhXVrtSVrhWrpxWd3evKBbSW8+YHA6zFW8BAjZqm68BKgIH80
e38bDmHebWZbEbleiTRWEXu8zhiNH1A5BggBHiGgrbwTFefBJoiEIhlFelUJ2/Y9
ZwFMWPvztT7H/kBmyjBxwydiGQxiDbUrJvrznxymP/nPUaj1fGfpNTqHPRiWAL+1
96TCB4jvhUTq1POVRkzpDQIrQZ0D1vipo1CtYB+vmYHYQNNGzu2CVg0JHpJPBicu
p5aed5HKn+I54YQ2sNR8kx0zwXL1IEZmxe9CsGG3iZPcyhVYgaCwlI7SmZn4M3dU
ucViNJh7AtY1zxY0Clun+0//YEKEe7sTKmRNi4PG4P9Q3nP1yQKvmb1eQtkDqcIJ
F79ftButRynCMDivUpJsIyEzAgoTzrXQ0b5RZLrrJWWfLirdxJ+j/kxRvadhJ287
YPSbxfoZcTvlS5/+EnZ/NRyUIG34gcHSkjCKj//9TV2H6jucfMrHePivwq1aSE9p
EcSn84XTUNmidym9+oAhsZ2rRObYcww+6rVAj5MIqNS4b6Ny3C4NZB0sxnz7Se75
kOMj5aHj7TXrpiGIZviFdEFDTQLxozI2cT/7mkNhkyBkNs17N3fUD8I9jnEy4dBk
mFBkTAYgCAIGGIY8tzu03xc338g5EqZEJqsLzOxEglQYmPyyMx4e/EZlLOIXtLF3
4VyQcnoYK+QgoiUVcKSHDv/o+QdfZazeyAzgEwFf3g2LGnTeEONqzjqQJ6G3fFBB
ExWRPDORo/i3/BgsHLH7JXSr7LbXb+XSNY4q9kg05hXYCNBqzFf9ub2DXgviflLd
ExpPt9m5TMlLa/lEwHyJ+ptxx5MtgvhkH7njvnekHtNYYsVRgBPoc6u5fmpyoXS3
dPvZgR+2VXCCub+EJZkfeVWVp73YB0MIuA0aGNDuZ0ZQTjLHOyuMWTmD1EZnwTCK
w5NTOH5TR5uSYTczuQMLXg+SKDhoNNgLzx9uD5cE65sczQ8u9hfphlnHtenpWCwJ
59sGPu+xxsvzW4D7GCHX9zpedZecfzPzIP3KpTlMIJZOQeiiicd24fzKoRosEfbx
zuxJ+WfPTvw3fBOMBJhDWE81Ui8HS5jklV/HwmaC8PcKTIeZMDBTR8LBeOsiIEut
QfLjgwfFOLFScxy/qbTT64IWfhb71+gERCYK5Ds5eeg2kLY3S8J0qSQIB2nfq3Pk
aAAAsHWKpv4jupfsTmbr3ZsQqEVl6g1DH2guBCVD4F5Q9J06y4FLWladoy0NE1rs
I/fimtFrV7QBYj0Js/Cc/07hbbagpnvhWTTTADwVX2+6BAIUl8/LUvBcDoa3eOtC
pH8Quk1Ir53jlrb5S5hr3fHsc7p/V0Auvy1qBZS4K9HKNB/I6qj0OHgnk/5dws/h
EGi3jblCnjtGmirOIdrcJuMlRHMLEmFy+E1R2Bm2u/i4svB0ymThYaNl+85Os+Qp
JqJr2Jiw7VdyNSKkgOSP18Gj4aW4YRtBBKz+h5C7cRsHQ/Ctgtbl93eGK6Erm9kg
/v0PlppEKMjdUyfl9BGFhOyjwSHABTgnMvKRCmrOvfBquv1ZQgc2gVOYU820A1Gu
ljvbVrdjRVInUJWYLR0mzMmOqPW/n1o3q0YhAwx9hkc37NGjToNAfSJSRE0+Xa4b
GOQdF3E0loHfgwZtbCma9fur1UfkA2HGsWhDrrFgCAh8LZWPhQFDM4o8vvAp1gIb
IhYNTT44avPDUf1lGcXkEEoKE3h7tizl8mAfhghQ9809wSHBavFu6zg+V4UnqqVX
exmBqY86VyBjarflgcXeeZV8Ov04ipZdc6vtqSP8Rx/SP6HLXfrU82GFQUzz4k+p
rPYUryX5/2raZnFhUzZg4wCBtCTLWSWa8+43rCW70DuvtH1Qpv867Hll/3Dg1x6Y
j4B+fu0zod5YZ6nOCHh5wTRdMkQ4DucxRms1SfuTcC15BloHcTLvJG0BNuFTebo2
dPzDkGz/7w1vr0Q/FhIbIHZamk5ebn74x/zTDRV9zeV0wLwGPZw+c0qwehlerIsO
Iprig0SlFER1yVh9owzq+IKOpg3Kql8cVafm1gqiTvh6peasGHnc1+0Pjqp3666t
mHX6b5PtEsVb5zdzKyHNqMynLsp/c+wIELqOIuk2CUm7nrdoRYRyAnng7cW8Xlju
xdhawMAEjrlXa1keeSdLFRNt8ioxoVwlS+27sC8K+SephY6U3pKQDNNhPoA15kOi
/7fBHNcoTc9QYm6HMYRsI7wbCM38R8sjHFtbg5cKxm4FUKDXMatOM81uW8HWkL5Q
GV99ZWIWQ+BGfiXRHKMKtb74aghKRugLlSZpUaM0P80vWxv9KBDYz/CtesZgdlGa
R2HKnFeeej4m87GOzOv5d+MtsSCB2Ltof/YdyhUFbPL1PK/tSbYJt7DawhBr07LP
OsBdzHU0APAYCJFu/PYBlfK1Dy6pHjDu8+xZ/415VylnLRRLcENQG/M6O/zJy1nB
3ZkxKKxcfV6peO1+HsFz48fwY440eJ1FuFX1+eUaHIJQF709nrVJ/zMZ2MMyHfFY
2ks/Jr9KjmoErnF7zDA+F2ip5JYmrPPin0gOgA+/bukLePhvG9j8jUU8fds9Tw7I
KVb4R2tjwINH5yiiUmBiGp2pvMJKnaup5OwgZheyYMxQB7F03TV32+/G1V0AUYdH
XWzI6TX6UAW0xoFtfambcVvcCU5ZtqUM8F57mJ3JoctbmmctpWV9sRHWq1fCMQQe
HRsYxtrLyqR+/wkyksObqobSCnV0t41Df9pdfBgUYDerBF0gM4znYmcpKpzEK2ud
fXKvUchlQ0/UCPY/Dy35Hp5mrk4L4TrQbkJve876mxzfpQttvHm+qxbZvJG4hzjQ
+4PbLQBViidhjCrnkrh6J4cSLTAVPh9EunlfLfDuDM4MOhB4yHJOSH7ZHr5GkRoz
6PNaaDkV3c0Zv4hdXtuJMSx5oYcoZQjX0eWBvt0qP1TrSiBhAo9y2lg4s9GKpEjX
R9FlhgpsTzTFZnurlTpMczjjifwak7wUoE4cJedUK4iOBgWmfjQlzcwE0i4r/+F9
EvfODG1sss+BrCryKvrGsBWgeCTfpM6bHYH8I3y8qdMfojUlpAs0y3Cd9qBCaPPP
itWE7UvyXpn9J3kzqRqnBI9ijUjqWOB2YK6J/7u5yFMhbF6CXzAJSzonXCL4ITkN
BJeEt7OzANe/uiVp07d0wM+QGIbjJqxk1pi6+zpOR+8dwRMrAFR8FY7cUWjwMHvZ
V+NUrND+3O+oRiy3q+V766rXTk4TI5epicbBCw1hgqz79TIYdmq6nsFYXvmz+Piu
oa30V1AO2XSxXeZmo9H3uYTxQoZGsKxGnPUfwFbTDMp4q/GT7hXJ1WSpLjoy1N2s
OvuQIa3nu1clQm4roPbxnhJ19r8njJR6mScWom36CN86txkHY1s8RzhylMx0v3iA
a9skhHFMxLJhepQdj40dMOLML575WOEmtfiFRl+I84pxMIM+/sLo/pV0fG/eUv+O
0DmyXSG3XLE8ykJwwCZSFy3AqnblC0QHucyd3StBOyDKdwG3EryKLx8l59kcEfts
8NShqwUgIa30Sk87HC4tq3hAcgBokkeSHHlKb74IKfWslz6iUX1t1uYFnh9511b4
ShHURFUA/h6o6vDqjmb/ojZa+mH6qfoVKDJTdZjQ3Mda3Kalxlb3osvj48JokZXM
/v5bQHc9wv6myWBW1ylGqUP1IyMZqoq4OaKK9xXHFrQ2+/DDtNTOzNPHi38+B6m5
tiPMrNmXXY//iKS0KvtF/UjIyIK99NMyVGQBJxkawqbiLEty2+UXR9gdjWKefo9T
gs1OzPBxTmuX/eu3bjL0dCh9Z5JxKP95W57ePe2Bbr6/KhRmCTfegm1POVn3eX6g
2wgeuRwI4ByGzQOs33GDV/rGZoro/2SpAkTI5mbii6zW+QerZXgSjt9KIftkoO9Q
zwgOy3rt1aatut37j2nfr9lEtwCC0h72FhFuncqu/299AImRMCXYw5xRBJjGYTG4
DzlnVoUQiZbR6gBsyymEg+UcteYUDrTYd2Y2OTi2fZx5jSq2ZLolerfThokU+2Ka
LnYQPyUSqTVZVZPP/Ss3RGuTTrfux7jxNMVMekk2DtQCV55EJbMPcV7NJA/WYfKN
xRUlET1J3qxm4TeU0rM1NV4BAqkdGQE7uvFQ9reww/Q0/GScHe3WptHgm7AUXtf0
vu/Mf9YPRv1I9W1u/KWcQaGDlm8wGKz7WZu/VjMl404fff3byER76qjQxlrTGiYo
3ogn2R3ClpuJ8Ji2h8FRVTqDgWPpRQMvS1IfS0Y2kA9bw2F4R4ADdyh1Tf+3L0uF
YNMHXV/BqWLLcZlcpcEyIvKd+l/NBtGpzaofrQLla7ZYdSRSR27PaAzTuPqhcwqR
vUhf+1JFD9RDVWIGkfaqGq7G1F66//Cn/m3AXegtbhu7r0qX+vdzWsnsL7vvDlvx
4491fM9t6tI9TaVR5pwF/l+ttVBfByi9ch4W33viTaxtafuRWnHyyS6MS/j2q+FK
6H6tBGuuV9xh9Rh3te64Tn6yCwFLaYN62EXTPXmIdxUhlosj2mpaoCE5wAwI/SqE
lR7rkdCiQWCkPFe/BQ6EvE/A5yNicsNu1r0a/J9uMKyfhGiKvQcAqfLziV+ZCSM1
pGoeEbsR5INkOzkCVZKry8aehQ19vhadqBE8xQk3qiK93kQTNUCxJwMO6h0R5zls
ibTtpk7U3em2OEHzoYPgPQrG7QGNHmsdm6ivvFAMjmRcdsdvbPzRoBvO7xjGyKr6
88QNKenaJGzClAA3Pla3XF9GIk2pUDq2Nd7oYHt4ix2+s6oTnnSkRRyAGMuE4uga
BMcQ4XeMVCN9VwLATQMYMIQbbblCdSG1omYRoC1uKEhGKmZASnqJ2+9Lu6WIwkwh
i6AgiNTtohB0cgJPYplnXH94piDt43pajUzrGNMUyKJE2sBrx1P7ye9kiAatYmic
Zaca3iy5sKiTnqzwKwPMuaVNxrqJozm/EAKJjMrxFNBo2b3BFt7DG6LnidWwLc9+
DsN9dhhz8efAS22UZ1k+idWKJf11G9KhiCtXpbFVk3ezt/xfx/iB9hj0/QcDDB4F
TGp5W5jVIr33ApxHyI5IIkVUDdH1pxWdGKV5aQf38puLK82WDqDPimPP2b7Q4jjx
O5dNwrMofbfkH7ulBA5J3vAtOF6GTfu0Lkms95pNi5pP1T+1zZIP0gGIcQ3Y2wAC
f9AYOJ5hszPnzSbiurYmB8VS4VFlIv/npiDG2DZICFFb7de2r/W2PcxYMaN2xLfw
XsZjc/UIaB+37hYUV5zLpPb3SJD0II3dORgTk81AnVOP5FzXAUZghqBxQQR2HtXb
vs3d3Pvh8YiKNwlAGVUtW1eq0A2RH4jnZVXH5GVNNemVjIdOEgn1F4b0z29BOGm2
Xyg8CiSjueP3JatLos88fpxaWvIMKleVuf7HkUU2mj0Uc3bjZHDWSwWbHaZy9gTU
eiRIjnWzn0R4MC/ATHYDJxx5HTo9ewPKS8pvgvTwdBuO7QHtb5AXnojb1ALnMijD
q07n6mcpcatKTnfy/OeJwFTifI0neOWQeOocT9r12MlXtwUxqyAVQ0tQf7lSrW23
xIPN/eH1hWzjYM7t71aVYw9UlTzLUXnNQOHdbeyLibu8twtCmaUm0VlE67rs8AG4
qIluX4aHJ3NAMWmxcDid+AoioB6K4/X2llWr9TPaD9NCOGnbO1+gyT/B7SoBWSOi
ZhkE0otSnRWG24ZDPmlnDrLtmhQ1KHPN1unpdVygXQbl7zTBY7j6eAhq5l/n+7OJ
OYjA+iTCHLG+fsNaXUQ4eiMvyW/6X8Y6UZbhPr7grmq+OLLnTOhUjnZmj+npfdJI
OmKa5Qp2qFWnzygrU31diHbMh1DLy69/gE8voW/xRruP+IDDMsw5VBfOzrYBZHXx
ttRsYnrs1rZ5HM6/UhgH7bYN6HTqXUsqZdqGcq16Q/5YTZPCfHCwahI3Jk0ssEG/
2vyv4Utla7FM7vOKJtT9lepasKlUH58EJlvz7FXcYsH4O4aLYicIVEEa89qqWrkh
84wblW1UAr6hVqD5eroqQsURRuRUcxtCTt2bOowlRSPyFJg6mK/H55JisPaKo0Y/
b6O5xg9TTrXV8ziwZcjN3Am2vBKMazafy/N8uP+hc85CKlPRaFkwj5LxlzSaZ/rY
U0zaHdXmYKY1VYSk+09F+DDDZFRk0wOW79HeSdSRqws3Ikosg4KFEF1wgOAxJKUd
OlWLTc3lRzxiDe49utKUEWYoEtbG/p2EdIbNnw3vJZx3Gf1sMdCLN2bS1DNaeV7L
ibp5nLDdoM+FssR4VyfZd79FLEgdECpdfrM8uxo7Ogt6hZfRveZ29+pdjHMY07Cr
Op8CVSqCPxlLZ+Wof6+EGh7ESOP4o9ZVjJMNV4BMS/tGH4aSVH9jzo6hnNVAWvvh
xfNWBg2CV7FSRjYhCehc1jF8sqXstZ1mC6SY1/Ot9jsloBkhj5kwXkebj7DK1lcz
O2O6MhFqHFz1lw5bRWAr0IKH17Sh0vnSYXAj7ruRFF6SuVLWYfoiBLYWpuXAQjHe
JwyNKE5aDdz4wVEopjGcEdVnEqfeSkiF/EwoaUf3fMA5PIZmMLi/3X1VrElSSuXU
bGM0mTDGgoWTyI2MZ/r1VIe/rwIIFHEFRsaWcUhBr4jRUz1qcCvuTb1Ujp38SAOu
oATdVYKWWvskvGzNtgrKluextnjZ4M2tsrdmWWVutwvS100ZZNWDnBdU9v9x8vM9
BaUtT+61oCZ0WdvcAfo6HXrFunprCCTaf2QdUowgiu5MG34Bo0sWzSWLy+77Cytk
HIwRONIlHEfMRrPNHQQfBYV6YMbKXKVhhoWkq62Ug+APlBDTx4OHPdqQiJLqS7jF
sQKsS8GokBzrHkwuwjFqQc/0m0TsM+fvp150j46lRfeJZO6myDpUZU0PiQS324t3
vBJHhct/d3Bfyy5k8ZIJoA3v/pFWDncY0oYCY67zbbML3irxvnrCIf3wcldyoPZs
yfzkK/yhd4XoP+WRgFaNMRwqq58kwMuBCN/iKVnjCCkmZwLPOFHdpqD0c9U8FMnM
SpsbERkPQimZBDvSuiNhfBaIsDPdC61Q2eXq3Lz4AMUim28O2kcJQqC1Ef/riAuW
JXAP4vGhqz0wvMRCqzupgR5eGxVybGzRz+gWjRn80U+3GPsWXnLPcIs8e4wogode
H5lexCbhyimgTbSmOEj4rVRv2R1twqinXX1MFuTzpHAu3gYcAxxitkMlQXbEsgRp
JzXalvvsxJdH2vERRCfs91/VOK910nCT+FOFuyzohVV5ao9xJjbGxJrzvDEymJJg
TyMOxv4XDRvD3DHHvfmTJtArRNT4VMMrgOdlPgdMZBGQuX8GkUHrtesWVYdLOaV1
uxkiBnMSA4Y8XzukqjtLUMgY3JSM87NX0qagJz5yp7uXSWgCEo1WU8/d9uJhvlY8
zjDBI94xfYyTpSeZufPoX+2VfsmH+St8rd0+sITNRpraa1qufDXsge03tF99cZUJ
otLIZTnn1jvRfoc3EjBTGJvCWaST43WvApqA0oWEvvmFd2X0N+SB6J/lJMvThoit
BAcL0TLd+ymg2ogDmEBJQKht8vaJek1eNSyki9cPQ+JpJw34nf2oIlTy/6H8ZKzN
4qM9uqX7CLzhY+L0mPj2so7GM65C2a3t1LkbUTsCviMPjLzXQmoVD2QsCn/qG5x8
2T253m92zSJgJYuyYI7GHCE0VNVC03osKgzXoY9fqPG/FpgcSeSO7zGfMX5gHP+i
xA5VQsXwMuKNpbj8JjQHqZZHtPdAriqy+VCQPuW2yWtlGQicmL7IXNPM5szlAqsz
VFhHEVPLrD5dRRL2+QuFY5bnOSNFiR2lstPQvGlqIaUyV9J/bly7WqqoC8XWYiI4
8xpPmB0l3gnqE5/3sQJTnlVfZdv7KD0O5hkCfc5uq94bAM7IMTkXEvqXWCn01h0J
VPlaM94lgKD4A5G2puVAEaIeIu+CQO5nyM90XoR8Qd4ttxK90bB+cGmsrB4ac4R3
FMsB3SFA3yjzFhMyKtlX5P86GOoDIKQN/rpLS1K0yhH9M/jgbd9+sjP8wkGKyQkX
c1h5KHvEJGa+qHcIH+yC8ZvFpjSjdBCBlYQLyhKfC8CKv2+f91d+CqaqmiMTX49M
xQmf3esDuBguN6mrYTM9iT9C7cmuXjtUiuMo0116DmEjUvGQsTLmjrbDvsdWu3Dn
CybIqXCi+tpouDsSqfL6dOSwc0Vgy27uB2rNvUAJdrrjDEct246agw3OTkE5GUGP
o9xNyb9AKh0RIaO6tn+cukcxZ4HHA2TiVXD8qZg0L5S5gGLDahtzy8wgxc4wbNIq
kqzlK3SUoHZZkPzsVFLfkYQU2wE3KuWDul/lKJ3C54q9jgaobvZIjz6PD/mqMII1
8BGO4MCXKNemUK/2AffNrg1K2DiKesX0gHYBTXIczeTawEo3Z4bpkyppvFIGz6xt
Nb7bpKKUYMqyIfXjk46AwTeKOlcp3OYjf6N3Q6aIFLLyqOiEpFpzGryryrOI8ywI
vDctc7pdWf75qZTVSaO8Fb3hAmjQe2ht8y+4IEacCz4/eDHmgMuDQV15Etm3tRhK
p3a+ftfDz78Ot/YntQfP27i1cwuDu/wv+2DyJJwn4i6WcJ4KKhZXEme/ZZFXuL14
U/Ip/CSJNBDBz7BDIxUkJFukF1AxBZoxYgJdvMralvQc4j4EudyfWzCS698mXK/S
n0rbaNRcSXEbViu+WBU0OhIKBu8jGcUyLrBBd7ExXAq43UlxAPEscIel/gDV+06S
bxCtDIg0yQ6ySsB+QxI5rKDSBxgmTYLe56utcc4RxtyvNcqxGUbq/HPZGSMdYbnd
QxNLxMdFb8Mvs3Zdqdxmi9lBBsAb1LFF8sTyjBgvWJ5nG4Gmif9dMSnVcM6U4xld
bWe6uUxvW04Wuh2dzHPo035R6Kz8vi3PrY/1wZ3b9huDwzdbIQmTdq7dTwDFIn26
myIVzsrQwZVAKDy0kXFEBoWLTb+VDeQAalju5r/rysKC+gKL3HwFeh1KZGy3K/N0
LdRW1zoDIAnA3rvdijTxfgHH+Xgkn2vRTHjS3wuT/5niuAFOWNwwO/pAA1X/wXy/
bN9WFMF/u6niwJ0r8ovFB5063Ia4IhLtFk4UJvGQ8S+t6zk6n4d3Cd27dfDncDiQ
8wNnFAD06lU0nETHlgINFyWlkDYWXO7Pe1phY/3Y9X1bJpYcp7Kaa8ILkvtiG86p
cHBQxzChFsC/xmAiD9u69vZSQxL+72nzE9YtzziBDEzFS/T4jxn0uy43+vvtRuUs
kObOJ9Bd7RfEdmfiTLBruytW3wo24ScDvUtH+IfAxlcrILjotqT+IySgqS5KUX0V
GNw2bb+Kc8f2/PJiRPiR/42GkqunvewuUQic8ISKgb0e67Bgt32Ogh6ZAY+Q+K0P
CI44BUDITIUuyMw9H/UoNrztswKnTdVV68MftYuMDTlK4H5V3YnzWpcI1JO72E/2
Xd6q+KwZtr417jDakx6XpljpsIGx5d/NTNQDFdC0kTifV1xSmGHQ8UTcMhU+O1Ab
37m8WcgBOSqZKEhlw8Tgffb5YoQYn/lOxJTJtuGRuH2E7VitN2n6NAR4ue8sAIIh
jZPsoMLRG3gsSjuWwivQD5eKGjXUVveK294vJenNhfU3ziGmvuoXNP1EYtP+Txzh
cDYUI5SfU44Mz2FQlpSZA4WY7Bl8nVgsVtwrpCyrIRHYJX9yOjHIHB0UZkeZ+vb+
2pea77BRe4o6qpisYxzLzBAGg2DoGikK9eYHsTZdP4aRCkJf4limSwDaclouQHAp
LdEiy7NqHkeoJLtMp5Srk6lnwDG6UKfb7UlV8hXw+L/BFe7XrmWpd04Ojg8bJpcY
uOjJPTGq6CwSn3JR4+B9QOSskm79a0eByIWwFWfGg//wkjZQPwmpE57GRnUel6ej
spjaTNnzSN/WH/6H484SuE3yzrQ/dp2IMyInpYhlVVINq0xakseE4lSe6DzRckS4
85WwRDLThhOvvERK5yueJOTNJpjPG61Bm5R35dkY9ZmVG7WqzjKjmJJdIitP3SlU
jaGHmjU6nQL83eisRbxWKi0ADi5yG3xoKww2I0ImWU1jtiSjd7uSbTAw8nI7vwba
MnEuKM7jgkT2VLIU3V7Pgwb9eHac2ewSjGfJj/kgGSpHrJXXytrwZA71FYKWRjdK
xVKVJhIEKlHuP/AScsmPNI9Vsj2unmuCb+EgCkMXOArGFPE38cqvnerTINdKFyH4
bYLcSWeWTml1TGeF+qPlRsIaN+c6Bpl8gU4+/NtHANKPRSz5/u/AOxwgINlQEU/o
kI52/JlI0khhWrSWpKVRRm2eRJb9iuVCsP6czLUK/YaPgrUzqToCeHtQvTz16FSw
qoJ8D0BTNdwdrrS9Qmbe7wczgifwzG9+tswBhT/olFR+GJ28IGM/9hcyY7ePmjLm
3V+qiMOcvn2mR1ByqnbkxcKRNrVZdO2OMcchoM7oncD/wDj4mkTjVylCg9d9GBx9
YUZ/fc7efEAJMTeMk+PWvu/cawO/pERhZz0Eq8N40Q8oXqWggEpy0YWNwJMEWnUo
39GzNImGGd5TyX1r3mVKqSGCROwqqptG/KyY8KSZkDO+mEKuMBpnBlNXGI36NcJ8
REyQwEjTBGxd1/bizOOxNKNS9qNuA5t0fYSw6ZI4xZasLOToL4ow5vSVsbu7Jmxk
aoPqs6hG7GzB3ViKRMn3itT/rEPQIJT4b6NXk6ZAWhfWxHkS8CUpO6TV/yZZVdD+
kSwShGyhxfRH3+Eo7kh3v6muBrxuo+4wOKP2eFZVEt/yJ+fMAFNYHsVQxKktbgOp
Ngu7bpX+VoB16oCgUolshvmQFZ8XLbCHtKUGzlbmpaadXF4wXCnK2pTMoTNIDxis
c0nZiueAwztbGGqxaTy5Hr/zqnYLK3TXgq/5bFgMh3TN9AEnoAHuZxlbI3yawjWv
1biM89Mm7HRHdQCbLxW/jhS3Of7c8Y8lOUWZWa5R5J5/76DplN7jmLV3Xr6dRQ3f
62anzueeexcN77xsNXsPWfslCNcmsF/ISlRpeLc92zA8dR9vkKiFgOIyzfF1vcEg
tF3O+aaUBJNtvGTD7Pocn4jLbtNAiMmlwgXKvcWu6Gu6DsmQijk9D3ZvGCKBp/DU
nxDNmwAV0vadD7uFoJ+WtxyBpa+x+kzdSGvwWbWwX0bIsd5yks+9cuaMHthrZiX7
Bz3YTx7okfL/FoINTKAYnRc+Cis7jKKGh/WbhMkqmuzzFebEVg64hpZA7bCZcHPU
GQq0NOLg8E03/Qz5hX2PUfBsmMN/zhqdFf3dsMzC7bf6LaBJ7RrP7VO3/Jwd4VMx
BkktBxNskfdEqIlDV6QnJMKFLv69cWrPlPW8bQoTem60MtRUKOpTpxyVPLXA3Ndq
kuqi0aA46NonzTXc6plGTcQymcx0O/qmQ0zMf5LhNBtF2sn0puO9oCcRH09+hbzj
5lWQoMAH+RP27FJjZknapKJBp3DITrS4sCmVT6W73KSE5pnlu3WaBCbq0oxQX/Dm
g50cY4BjJkFrnziPEs2JAJZeuXG/2pKRuYFOYrkm2BNAGfqg+I8uAb5KAZkwveuf
eiO4w+8Kvn4VU7hhFgPIKHLYBlegAWGmZVpHJghohAc73hlIBR3OhTEjCS49ZsVw
SAoeLdP1/GmsyYxDeYCwXspQJlPxJ8/pLxt1GW/5vmwDWFl/5RSM4Oo/oy5q8Fdh
4j1qlzOJUpe5FksG1BFMrKLXA1/UIw0JiX77f8rvJPPAYtXA0KH90qkxFlk/B5j/
VCTySdEUIP/wB//gDGJSYuLyGUJP3xggV70fo5v7FyVW3vUDtdZnVAIfAqNny957
2jPyFffmbQsUkXWQA1J0pmc0IDuedmZSyf5Mh5F0cKn+HjXpjnRnZiMi6LFDZfHD
OMzYtkyuLOzX3hJd+hgMEJVLpeIhEh7bwm+B5fd6av63LyrD8bENMSp/InPyuoTR
+6tznxkIyjEQeZjin9LrpDMmHp5kBsxigNH1Dz2/ONDaeVlJHnuwySLy21wfyAE8
EbXh9v79rNqLYYz4+wa99xXXjQRmZsEj6WpJwZepy0kdW8zRhX8Tn5Vjm3wDBDiE
TVTM96y/m7ByNmo6TOL7mq0BrMEeuLCE1IblvEXpbNFqcDQNJf4yQ5C02g8LhuR1
+4N22xlAC5Dq3LIuHPHy4fQTmcUseY5idU8NL1wBqwbmD5AJfCBPrGiISCJX5Fdc
vX6rntc+vGpl8YQtYodZ8Gn0r2/xwveUk6rL/1xp60K5TdrMW6PR+w6AiopszxDa
eELboZ/8e/T9JLH3dXOJMJhwC772J3YLIZu1Hjva9fRUKPkURue+VSCGeFhqf2TY
chH+SozcbDDsSF4z8/2cNLEiCAgrLgVUGdjQeyyNap1kzrevouA4Kk1m9IFAaSfk
3z/HM74G9ffsP7uXVgcOl7qS+CSeZKHX4mzIffiW/j+16Kr1ENqZ0M7XFzebOj9T
ktibTBkGnBCf4Gw/I0vS6O+5X3BNahEmB6DeIZGPVy0w2LOQPLcGWTDhzDoLTz06
qlFzGdZq0rhgAxfJfghoynePakds5dWlbBNItBna/AgG9rBpCV9ZgcjAsiJLNlYv
5osTzJOsaBPHmtSoGH46X8O5ZOqwxzKEl9G1GR1fMrkUy7GvKr67K8DrXovXIQsm
NfjNPKj8a8kbs8o8wK4U0vTXle9NVTCOmjb2t7UZrxzF5xe4T0PAQAHcBnFWdPzA
bCrEpf77sn6QTM2lgiTK4KV2SUXCboQgfnA3DfFP6Kn/CMEu7yz9NFeRt14XlKnx
yJ/H7Ikm9knMnMBnCe/zLXqesdM2/ZaIkbdfdi9bWbpd934uwFXvxrQCXS3BH2AQ
wlrpbd2p2704UL8+YYsMa0GPlq7NdbH/UGEPmM2qAHxQn1TdJVvfahpumvdylAy5
rz99z2oKKYa1naYhEB5pzDbtYiDu04/rsDpvAjb7CxB5Jlv3p8TXGliIGGkMcfSe
bJhDpiyMXn96+mjp7+HcPaqUknrXhMIDbsh8qC1kMmMRwOX1rMXsZkSOtKWtF2tS
icN5V+M2EQe/vLYMEmgVjfoO754Mu+UL/5Z8id+9TcDGm+dEWNvg1ltmsweBSRLu
Zt0XpIzmmeGeDcQmAycx7WJkFxY0V30pcaA+W3M5A+UClalEnY0tlgkvwMBWF4jb
3kUD7WGPtwsKSO+YmWYccg+nR67V5+FcRKLzbT05mDod1vmVLjpfyJ/FeG8ANUqe
8RpLpnVOWtZ+TMzArJ0lZTWcpEZZrcPPhyh1o0NyWM3mEG/67VLbjioSmwxpRSGX
sQmJcbUEP30Xs/DFoXhkEoxg2q77W+XBOmRSjy51gN12ezepaoiZH7kKG65wT13U
sYn3JLAh7kohB8ZhVguxb6rL262dMnyb+WS/OTBfxliMq7vYZ6Az08WikH2WBr75
cNQZFmVGYLX4echrC+bxr4OpfWIonGdTPqLPoLOY5o9n81bTmvSaFFYlMbJD+VSk
07iFxwNeDkNZgDzoEbmrySgOu3Q7tuqzm16bOv+PNxMTECpPWRJBzrhZCSJYSF/J
XB9XfCTKjO4WfrjLOzPATTuAjh6fHLim4cPZKnw6f83TaSMSzdbY2bgoRrC9ldFn
PbsEUP6pBM1ptaQL+P2cDkWCxXwYSMgFhlYVvcNuxtG9MhE61nOnaACKHpVG3sK0
lQj5vPXZwJBLXpNPvqkaXXDPn/zTrg57w7t/JoQoXKpnq1RxRy7/C81vbdJZR6Uc
rJIb8zgt7WZxIVfWLDyZ9KHiUWeO7CGwY31h4AjrSBZ1Ke+DLR3C0R2clQGCsrUU
1tExVnSpU6K+5zqxj9vLphaxM15QpYuQH7E5z35qw7CzUqnW4C1khklb7Lyj8gRH
lQ+f8GRT1oabzpFHObx6VaSDatp/474l54Yv8po1iNKmZPUHLYARVSseyq4WwYRN
akYt6fk+0QNneOZVFOpMZDxgFGcb3+9kZ99dX25BdHuIiwJ4XrhL1haVK11jo8YL
NA0Fguj9zCMeolS1qBhSmJ+AXJ2054ao/aPSIyhe/BG3EkMIQEkwDBc6shFNaJSd
Qh9r/r6v/v+wL6ZwIrtXAyCl6buAF4x4FirPK6PNS8bc9Xa7KqcU97bYxVmuYPg1
Eb0jfQ4isLJ3gXm6UKD1iI58C3uOq8SLO6YCBMOu4C7e34sJDzjLXP6Cd3npPJpc
82uFMbdEkx/uOOpiEkwDwyv60s5Ui8qRB9E2YmHB/AGiT78h3DMSE0hmtuYaPme3
jflN6yN3VrP22IcB7NfGao9B5FPOBEqIYxDU96qLGsk9v1nXHh/K9GDOI7+TSpZz
bPi1Yd0msrHMOgO5Q14RBRu+KaXVpQEKgaky0+E7X/zGWBBFpwStFRK4i2oabnrW
H1jUfBvMosbsqzljdAh4kgt6wdFTFhBFpPC4IAuEcc24i7GL5xbsYNvyl0tnGASz
`pragma protect end_protected
