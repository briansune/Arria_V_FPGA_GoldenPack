// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:29 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B5BxK1jMVXKX6mO/Sa63m7knjtTPoBBYe1AqqUavTDpFfvG8d6Jf143cJtqCMO+D
/meczSpHPzEVJic1lRfnXgwRt9RWVfbaJfq9P9EjMh4Y1N8MCbY0GURY64MhJcIw
ByObsZC2+IepihR4kX7xWPqjlNY3Aa34Zpid34G6CJI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
UWGK1a2JfE9v1agzHpsibBbUGJ8CVYfH8NS7EXtiDk0B+VRWhBJbjlJWqShH/AId
9iUGay6EMebri+NOvi0kCghzDN7sqLImRS0Abg0gNI76/0F/ZlRHgvDxXESJAiKj
6dtrYPzXpZTvKJY8B2R9iOQ7ABKDDAzTOCoVuN98olODEWoSXwmrNHWuj39kbsJu
KARRBZQ8RXkjAB7MgcitxlBSHnGN+33S6BPSht2sk31gwmrDbTbmGxc4xB+D97mW
EeIF7A/RyAYrAm/ZAO9NBCNHUEv8uQdRjQzQfcvd7cI7CYMtCcrDGR6X/M6gW4cN
t4jDFwCFDMwVDxlwWUqx1qqcnQzdXULgVkUxI8okvXm1IGG71lcuV5C1GxCzV6q2
+TXEMIMFTuFnZVWfRXuifsK6cbnN0M6HMYkg24zvCpMWaKGoUQSmMSmZ0npArxQ+
xC0fQoFuapKSWxpmPMRlKDwYPL+8BJtFf+Ngf59PJdEe9wHZjQCOmJapctPPlIMB
7QWj6k0LPxlpgUbmBuUhx/zNScL8cII8dYyVKYfX6UAesONSqjI//D0O3wRrEzpa
jdBkvsWIgl8RwCEjK/gi35D7HNf3mjZZMRX27SBKhFMGrZv1S8vl2N08zN8p/KOp
lBy9zdkM0LwuPq73wi/2VDS6RvbPawdMcvNwJIUN6iqNS7aEjaZaPnPMUhHjHRok
N2o/NnTz1qo0xfaujncBszSMha1uvBHRJDbnFkO/2DjHOpCnWbaQRc21oEKZ+T0I
UXqvzSKg66ih9t8dIt6DplccBzvWzNWfhVpXil+RWKJpfZ0jdMjruGOUMy4ItMqH
c9x/zQl3MBR/JEZnPdRxjNIZEf7Z/PBl7plbqrsmNWa6/9d+P1OU0u1aSKfPi8rC
Gt9XgCQ6LRzo/kCvnqF+gLr5OqLVRwWhFZ0udv0Xe11jUbOPTZ4kd7xdcJ6n4xwf
07G13Gyo0rdooo2hQaQa2fTQiT3vE0IOBxx7dQFQdc0KlE4aD5Cjg3w4wKLiz+st
ZeCpLgQ1+ue+hArsPB1FvekmmTKmOHL87/xBPEQ9nobvxHh0e8M7s1LVlMlhzurz
ZEzeBsp6TkiNix965pNDtS+YU/lZ43x1kflXpD+IokoxzXV0OVZekGCNs1RRg3f8
9g9mUb2lQEVG0QzUm+OuQ0pXmW1cuIueisiNHExbbAkDU/RXGSAH0A9VYcm92T0Y
z58iagzcy+CCc8eFqcn3rxMiGs9csQYEB4FzLtRehpx3ZtFmMyp2kyzuXXNj2H7V
TwyLmJUq8eLmIhkvMOjSsMwTLR1Mu5/1VZjrfsoYPSpoN8CRg/VWQJEcWZ2ni3zv
2hKvfrbjY4cFjRCouif/Z4zWqxNyrnZDcMAAPI33ZiIXUawQOk66cNtOEu8nXtXW
95TapkCMDvy+ODKw5Q+rAz6UnoDdl9Uc9VXTKgqdEG1DXPZ/LVCmD+E1BuyGkqB3
wUVQ+SgjVWirDeMPSDiMiVrrmPbtoP4OUPLHu5NojkvKW+k3qyLTymszZfLB+REf
NeP+HPFMC0bPLel5RxHhVO6r2+v7H9lMiC/1cZz0s2dHxjw8ZICiQvVRD+tpqtXa
BN2eGDQZ1PP15Jsd0KpZPvlCMOh26VYRuhkWJiMdxiFZRDcChti5HSN7yiMV5GeV
9SN5Hv2alUg5AHvzN+oYsjCojGkVB1wzYW4iIQeR6umiypyk40o7D1krs5t4hqDb
DBwhWbBYLwyFl6p3T6cxJtUX0qbrp3ZnL30y0gBNWIFpmem0aD4EoB8rMBaaFhL0
H3C7My3W/3JyG7jEbnoRCF97niyOfxNI7jc0mkrP3pvyxr7GPLMEnih2dOD31vYh
dQy49ngTu1BGvPUoVGMqWicVkda6tLcVmaJQcQeVcy5xJE6BdXL52favENmjYDVg
RneaBSCdQ84SuwWdaKpo1SRI+9NDjm9MEkMC1TQQRpBmY4LYQudR1bEAp9DzXZX4
NIB0rHUidmdVPwgVZ/XCD7hKD9xfBMYyLNUOkk/uUMyaz4603mKuS7Ai3bmAwN7J
V5aN/y11hUAk+OEaDHPLCZLWro8rrAOhShO2LbeMALTfzyE8t4AkFqKXO7Vj4tr6
uPa888zWjqNA8J0yBouzOtpZioBz48RXaIYWNUGERo3V9I6EJHx2tdv4fjXb9DE9
hdGI6/5pugTpe9976448eLgQL6I5KLVdN1lU/6qW3v5TLF5G6otIn/8v3dFJ2Qo5
AVutwJnw+l34r5wHcFRu6S4KanKDXl/YAGeR9dWOYFvWaacE4R7mLAGUjoNG1Mfz
ZcAamRvzm7Wc+XfSBa0CfQDnkGFtB1QLppx/Z2eouTWxWoBswLaSlbzeOkQjIQSC
zQ5g+HhwIlP2lI9ZVNEyMPVeONGHWVy8u/ahYzCt1QvemRYOuTvoqglPiYaHslvo
Goj/EHmQ3SokF58FUQ731BI+ciMVzkJqQskXO25ZqW6a8mordtwArZyL5vXOAPi4
1IrWwTPPDN/9dy8ooyImZLor74Bza2z8JIjzwtU+U5NfKOlkbD0Ynn0PzgyHnhPV
nVulPw/IPc2jXZuxeLTtTKLOIJKcX2A2bkELKU7GQolumHWUy7NligBbS1ShD4VN
0kBakSzdb50cLjhMMTiicN8QgF2/EOg7LuSOrQWLcVrf12F4kuYTDpGG6kjTzPkz
AB+IZAVir4HlrDc5wPz7e3xYmohB2PhUrgKsN7mRjzup4ucm2qzJolktVUfS9AOW
c/gNcX4C1J/jwK+fG9x4qJF7M6IDsVI5weh6ZV1Kpjrc7FSAk7vVu8Q9CbFTCrQT
Wj7ba19vvGR2gG0xZJCDYd5cVFPoseZNWjD/9IeMofUcD2EbYoJ/5DJN5+Y4suyk
ohBCyp5tNnCRiaHbOQU65dIZVOco2C1f0rtm7w3jSDiEtemHannnQtLFmxI8ukcd
uDmo6MR9pD7Ua7HdFMDBX3RMh5TqMHh+/9/LCCzPAoFX7YsLyuOSCPcd6dcLjKzs
TIWr167Cm3Ozh4eLOh1B7ccgzLVM1863203eqYPhJL9Szg2MDNSBeLF7JMjFOBXo
2kD6BmI962eAwee5UC6tvkMvkHr0krbN8lyISJ0DMNmr/0u0mV7ZKPEKzesGNFFS
`pragma protect end_protected
