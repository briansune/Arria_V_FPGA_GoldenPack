// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:23 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VkQ0yC4OGH1tvkMM6KPgyonp8Vp4WtcAV1Suii0wVQ40mtA25/IHt0ZX2192JaSs
euZyDJdmAIYcZMQ6JYmomSIJ7dIV/RHYjvdHYNqbi81lfr9THkPIEz0UmbGXFmvD
sG93SgSP+whpj3dmv5YLiH7w9e0/iMbQOV+ivWyk9R0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6528)
wHGAipp5L+CW03wNeOWKPyUVpfkmMZ0gNby0JhhGI7lLLhEmfqWYO17nci+SVK6n
zJMxi0VplWmuWrUHGogP5ugo6ejZURUheYFel2TKvtqCWk+Vbr1UDnB1MpIxHpIj
+8Bbr9c26DEXC6MM3AYZhBGqDvM8cpWZSsb4acoP6RPZzEjSAj3Xd408EoAXEROx
0cWYfnFUw72JRYdvS9C//6ajL6i5byouQHhprjE6R+JqkBEiDsbf2OSR806Nnaf6
ZaR2OvsguGZyvBG8fFdaBJoaa0M8sk4Bpu3klmpgWOuhAW1TAVCnbxU0UOiv5Ze6
/f2qBPCHHxF48SXAKj8rzH+oWV2+zCWqztoNnVcqy4i83hf6fZgKQHuJSnvy4lRX
LFMgcRUgIiN4cIrklwNkxcvRpSCZ1HPyvv4H1J6VEJiCrWOUwEbKHzySA+UG23dm
JRJSj4Shkd9KlCFIw62u7qJ3O476PurCWExXCX4G9ZfLMMoeBcTxazCcJQEZlhh6
wfkiTJ81gRdS+d9WSHCuC5IpTP8WInw8xNg6ZnavnxLFgl/wFbkAN1HCy5K6nam3
Blb/qO0Lxwux0voMpFw7jal+45F9UE8BJfF/jMN12qLmW/gao0TM1n41pLFt9aZN
K2pHPXXvavJq1QHWq4yUUzt2BNbQfP3cVi8Ov9Idgew64MZbxsE9QeCSSubvI0kc
nWYwgwkwhnsTQcf76dGCiQfF+A4aNWxKegqABgOz+SdmgxISHROWDLl7TV5KL2Vz
gCRIJU3msczDrQWYDorc15xgwM8uiaD8hPM/HBImyOwxS6gjTuUz1BmRJnoBAvmY
ii+2xlltbZaMpO/MSoIDtFoh+B6N9Feah1Grok7iRcfFTK5p9rFoYv4fKt/it0We
qTOCkjeNGxx5RZEWMevxTIEzPsLOZDkpOIawnhStaNI27BxdQ5eJnGatd6RUcdtm
iEYM1Ns85dIOL6eJ9cvlzk/Ni+xe9Y45nwmPTcB6CbnnY/YEQT5ZVunTw81nJwLG
rEQGT1iH8Hdr94BnOdQs+sjI3MwoITt2xMhdkGfRFbW+Q5PKY5VqCARxsm6nfEVE
6tTPXTf/JG9fe1TBvMW83bTZHMF8oHdYxES6EQj2VlHNRHHI6ww/aI1nDSttbxv+
nram/Ek/vjn2rDX97KwbiB9nCiqrW3MBgXhpqejafGD/7Wxl1EULxuFR7W/s35EB
pkiOBg4r8eRMpVZTjmoTpHi+tCUK0HoSoMNSZKXGWhHdQVrin8NepCNOwiS8j7PQ
DveC5lMeXyoa6GRgYxQRZDpOpUHEJdj4UgUUJpxRPkd18XmahSLiNduX/eTLo6KN
uBvJD3G0hYKh9dy5l4nL4bUk7NmjpDFsWzuoQgi8c98VjJNA/zoH7YMMLnkC7Ilp
bEQNG19oz/ZNtE92wM2vqWMfDjvkk19UOvdLs/SeCgttQiYKW5tco3KzaNAw2vFG
+Lloemie1MAJ1raWYJkk83KHYM8Q1u/MMor45xhdwasF7n+QM6XWEMmBpPfSMnge
LMcqyrjzzUmsy/U0Ke0k5EVC0XDXicGcyde0uozBt5kDehk6gxrZBg4zogJtaJZB
VPV8FcGZUmZenI9fM9L8dYjRHe4LIseYyWPEmcMTSejq41ogNAXQiVQrz7s49Rox
n/BOB2he42Z0O9KwqbaUmvwmv6hT6/U27JzS0c756zwyajpoqKLaR5qyuHhCjyWG
P1N/ttS2GewOEe0Pt4hVWTP4KIczfbwE7usN10rvisDRwyYFSrh2F/qPHgYBfAVo
YqOK5Voe2tM2ejee1JAPaCzyHsQCoZ08zKpcD4LyLrqsi0bUVOK2E1VCKaBwfBgy
/MFy6Uh4R/h8PMI8CwnhUlBPPXuHo154UUHm43Ci9Cmrc/SgV8m3vzxGT1gG+1Rb
VnmEGkdsaldKSgEPByGZkiryhDei9xgUsXyyaIDXTJb5PzcBplDBQcEdbSBiKu3q
EvJXXqFcDau+/HIOV+vUKGiycR80Qc6oX9qJCN+Fy8goeNWeEPewd8Rghnq2wdVr
7VOE5V42bWrFlsU1tpftqEI4dHQlZt9igI2+TLrQ+r8FDoUucjftp6OS4zVED7nk
g7uyzIGUnu0NxzmoRoFD0hadthcwJ8rD4CDXGSY/4+8NYtsiIls7/hzVpbPxZkzi
iz+Z6uXUcDSBHRx7TP0DWnRAhrwC5sMY5tt1rmxMG5M87q54G9JCcdsHmtOSa0mN
9xJafnbjBtYH2GeyE8zdEZ2uRlMhWJuayd6KAxv2ei82I0ErN/7qmzev+JC9QG/E
TzNr+D586y62vb9XO4l9V4m5SaFNRhdq/36f4hmtJx8TZ+elh16zKUKY8DTMGwrV
+vpKwOwNGAVASGgMlK0bRtq9/JWzn2DrUfsU0zTai+3S1OaopZAtP9YhizbP5k5f
waB2WtklZ6x0hhiPqt5WIxLK85/ZNdxPiw21wPmzY+BqBAuy6QqIutraIMJkSbgT
yP/Tc17lmtmZxGaokB0T40krqmuHWnuoNl66w64HpaZyiP/ChCavAnMaVcjPW6Iu
xm7kKepM9WLGssA3lcf6BQKgwPcNS1oKOuBfG7TTysydy9H2TmRGNwKm8Dn+zC/5
GS2R5DmqsjlzK1Xou5/2duhKqsHlJA7pT8cfBh0T0hRGsK95xgJYc4rP9SyvRgo7
Hbr9JCiDhY8v1dBcqmqvzTSrEZZnYaLaZ4F+Vxd1K1ZWjB/dDdzJBjs0s2ODaGtL
/19CRb2Mwiz41veAMNK1INL1UicO7LZEd6VzHsgEgQFljQJahtxYVfgLuXxgKEaw
i5KrI/9VOnjIzceDEajoOg9kBP5wiECcR8B1Xsycv6XMgWO6RtGvmYSLVdK0z018
ZbKjwamvByb1i5AuCbUCKZadiN47AVUtjBOLeuq6UYxGDOC/dF7EuUHvRM9pR/n+
Ut+ZgARyZ4l5PZGHMIUJDd+8zwQ1urQKOTmAEtT0Cf9hd3ZwZh0E1cEUDcS8lvV8
G1osO2hodcONfInNGblrywlzepubnsmsNOoZyEBzUOss3OYMM0jeIUtLjdxK7ImQ
e8GWZZ3EHgkmN8Fdql52DQGNFp/H4hFqtaR67aNkoyELbGheOXmVa9HAFuMZnCbl
CTgIbkCJSAE25V+yDY4RJmoc0Lzv16+rA9k9LCgVOk92kaTNXpjF5R8a/BxuAxhs
xRmMkluiLHCCZS8AmYG4lyxqyutDtnHnZcEX0Y0wkjXv4hjGML0D5m1NZePJBooU
BPOwkGxB+RQFvR5nMrUn9P/EH6nDR3fX7pHMKWkR7BxjLnS0IJyp2W6Xp9I/Lhb9
YA6EbUYOeMWrxZm6lx/ZCwtf7RCCXd2aqGfinfbVupPrsbhBQmmJNN2RL0HfkQVp
nM1IkjKm2L4Z8YrzJakHCIXTHAu5d5auXhcRbOAoDNniyKv3XuGBM6ph4dVCGVBD
RmM7a4RdnD3D7m4mIasox+muVnafvNRcm1xuRFHn/gAWP6aikIqmfUURsyv2VAq9
S+vxIo4ZsWHW/ZygOXETdJBYnWUdYKSahVnCxyezHu9jXSuJ3kDbz5fi4RmG0sOw
YD/rfAeD9CDMnis+nqxSDhd8BbUTu3Cb8+Ao1aklp7YhZhDEI/iD44QuVLocGOVF
mEtQ19id0gj8xP9KNiD5BQC+9JIRXoRCbhA9ejuOo8HFuY3ZCmc9I6tyItcms0Nf
EyAmB25ZR3c6Eypk+cvYdsxl/iNQQ+pNazolftCnWmFqVppyRiPAufjh9MuQqJ8j
jqrYeR/q5fGVFWu0iy6OyxcHe6SD6fDn1OPwpSFHpr8gL/KYSjVi7K0Z+yL5OISy
/Fc80Nl3y32h6j5zhWS4VB9nC6LFf01EzH9qgJbzA6lIhdNVhqpKpDvPrmrPx5Pk
xwZeVlwp4lUpVzDX88BwyqWVPnLxfCs/pfSIWkGQ/4yozHgux8q2/djeiPrdyJS9
29bgrI6KJLx8Iz0gNRsikxDHoUBMBosexdSx+qSlPv9xZhabpYZZ7+Ustiu8kSmi
VfyKIpTYBQCxEm3niQwSKWYIaMXYwi01oYcTzCC1WncQ5A8Kp85YBv0V1b9AFgGE
uV2dBrnsl3sLwLorK7G5wKrXzKG6zFfq66zEI5ZI8jkb4WomNuDSqofMUsHkDZQO
g5ObRYQ+j4/g4XPIVhG2s4p6UzCpPluYUZxyWLgCzLbFZhLY6epBBaZZwruXP9Rv
pPGYBJKTuv5YCv7ariyzlLGEXr/l+/LFlHNevYHk9JY9gNcTfDqRUxxb9S2G9kyL
WC+g45b0l2LA+JK857YLTpu71bRqxjODS2SqEYibxea5V5ck5JqvvWZbIKxNbks1
SwLgvYGGLPIRy24LbNPqSm07Z1cj3qLqWXxXGyMxrAOc6S+ChZxRWa1Hb4IRhwFl
2N5+o++cXdRn44Hr0QxMIldQbnabfY0qzON4+PBEy7QxWcZMPuPWrCGkP01Zv/SE
WNnsGk8mYfpIo4FvHRNFxMxWtz16H9ZU4i2LBXUMV2d2ux/H9NlxNEy/6Q/l7zio
vVnL3E7E3XDGi/K4aIx2Pd94/QjlxztGXrhtdm55IatdjXts4SQ4HmzDi6LbuaLw
l2KG0PCJa/qrXTdLpm5O0CnzpniwTnvV1UmXfEkt6tkwXi4mPoGahotS0U8xf/fX
YKKQ6ZuU6PHU7pp/lt2mWZnNVacJN6oej8DUpf730MDmwJqO7Ms50swHaDNeID6M
xmxAspdpqTyzWlNH2y1XYC3bMVRd0IQn62KSPZnXYbyIi+Nfrr2+y7E4fsxTYueD
KaKVJCdqR85Kw5eJRfA9FhYdEULmHXHTfAYpk2EqecvaD8Oih+Da8XKJYJmjBdmy
PtGjuD9uikFkOrSsZQek9ScX5f/KEBA+w2tiJAqVljz12wDAuGRumQ3lpPYS7HLp
5+oAu0yU1fSTIHrwCIyGmTLciv7rXS2/23h4oSN25VMQwRzbuzrlBYF18pTTGhrX
S5DBYa1modA1pC2gyqEUcK7RmiIlD4rlnBSzuc5otHV6rvtam9CF62ZHl28jmAwE
u+I0WMF5vN1NIhkdaYNEzDLvieh4FIZOIC7p7I0HlnYVftELXiP1d6Krhk/n9IgT
4DkaxzC3CxUvte+8XBXdOaUClBGetwK7Cnko76QwAdIwLEI3mOrqm/QRIsWU0iGy
PyOT7AEuZnr9DyWI0awSto0JkB51fkDGv1IWnlEVdFj/5uzHJIL48TO9l49wqmou
Q5LW7xlSV4/4kalmhAm193F57xuzLl163Om9XmkXuLlKD0u6OId3vW1CmAjwNCKP
nX1+FkTAZt/AsYMrPPR+AnICUV58eP6fvU5QdQ6vZjhEJ3zD299qOMVvzKEc1oOd
DqJtfIXGm7vUyAD1kwpr8QM0RJAyPU1PWHjNPZTaXep8ZnWwTTwQ7wGE3meQU5iE
gd7p0oSOvfzpMvtvMQr9wMwX35FW6DWFnBP1hhLoicqczJWFootBnwiVtoPKjii+
XAQZdsLITMeQg0q+rzbe5UWYs7IQSZbvjGlcsxzN4MqLIq4tHDqRu8PiMs5BFnhl
TKtiAefUKveInrSHrYkRWkKjwxNqS0DQtVCFd8uUkAlzPdEwpGlvtGquVMnnD2hK
w36qwZZH7nAIqd5pCjpl6thqcqYiJ6ZkItsp95jcc0RdVXkSQZsATQB//UdvaZFc
Qe4g8vPN5VAn08u3RT6O1tF+4JvT+Qf2rg0FCvzoA5CDcsi1q6Z+f+BxnIHVJNGo
IHzM7mC4Db+KBEHBiuIe6TCqnyjbOtMpBoBzXYwegPi06z/wGAez31bDWvNAhOKt
YX2Thy3WjDy4Pu6K3TFqg5I+bYhs5fkkIZhHAQfV+ZcKwjgVyGuURnuDyDgyyazJ
SvGDSEb+j/ZlUIJfs84nL9gCGJLgwE5p1H0AHPjeQ0LwTvImd2J0p6xVRu4/1EkD
/bCT4d0sSkEkBPclzsOeOqPAHWJz4BHpBMEyLca0qjqrHlGD2u6vCpmRndhiOnWR
c1JntEhryNnbmQ4kE2xGKLoUh/L10gXmNeiQ+wpuvqGJQ7Gdiyrf8LRdUvCa/ej7
/Wr2SHXV9fdL2xk5xfw1iuY/qz9JBZErJnug6r4+QWwicYZ+l8/FxqAYBAwEnC2P
8KwuWfEij9/rEp9Tnv9vLQkzlxoltzU1sYSYPBNs/zkuUJAyq9is3EXYUb6d2NDV
YBG/OjXSSu9wsQAScHGKWsPaNvTcgCDyWbaJok178TlbYkjIeKNvR1XstB/uaLOh
438nLoyCHyn2bxcwWn4GlucQSpb50KdNn0H9u+6EmRhyokgzgfnkly3jLYSc9rvt
lrCrPUCMrb1h4AIkQtyX3ykydbq5jCz/7pp0CaMV1PZX2nUyzr3rH2OEgDzg/j49
hZygllKLeXAWwKusg3Ccvv0Kowz7ES2OKM6VdGxz8hg/3iq8gWoxKg8OCU8PE2ld
VOQhCg0mzft5JehCQRGc8WyY+pfTW3/6LOzZ6hM7f7ZNaTbgUUNSkOgDQk/iCQie
IddsAHDODQdnMmyRE49SjnhR7yG0G3Y3Lf9/Yd0TPmKJ7FtR5jI7b6c9fl9Nkut+
GqzSHtQmESiA8eVpqgxhdAJGS0LpkAaV10wnRa2EqcWAI7CQVWqIusthdWbP0j+A
svPS7lvZ2zNEG1kWRYhFiFklcaBwIM4neFZZrs2iMkP1DyFhVdEU5bIl1JO3k3fR
VhgPTz7Ki3ljrO6Cp7yey1oj55D/vU675YPShzK+EruZVTlA1dY80VTmiHESfOZ0
cXS1wA9aS9ZL10Jf1hggactCyQogMRK2SJ26ExoUIBAKRDKkqHRsZk7Jap59bsYg
rFoZlsaA7+6X+n/7ul/zQL15S2nDiuvCSfoKTqv1CJN8suQ31W5i+u8hYwiLKgfM
4pO9OZwFXsGlOQLMrXOANsoIrazJgnZjBqiDq+LofHrsgAX1ybkrNE9Qb4XQn3z8
9E3U63rlpQSYKRIE2hg3Z0SJcSxVzWQ+pTEzeIlNqJ8BHmtxSsobUu7kMOqpleDA
PhZB957LOYr4xpnEQZlKJzdR6uUBE/RhuBvEPkoCEOlxEr/3Fh/qx6pxIakDRtss
4/38wvVGwI32/v+eshJs3p+MMVDRAMkfNkf3bkDkEKQCw+LG9XYcgHOJmOG8MDgc
SRJzjjvRcWG/PWHhyJQWt5VNSx+qIpcSrOoLTB0PrgT1EgIlGe9aazt0+vJmlvmK
RWKOhG2g/gkb1icUt57ZqOCl+J0QJyX47P9FmPIw+8kvpLT4TALrtZIVLJHKU8/K
Ujm1nUcZzd01u1AOwMuPYbpxnRI97HlmxlLQWYANwsLN2VRo5n8T2w3tF/aC2dFj
xk/9YPcYwA4U80AJTP5hbWrWcbd7q+jZzyl5oaTjBtGas8480m3N+BuRRRo8dKDG
xlpobHgjKFI9Bhxa23/I/rvKjBleAfhZ8jlhLhZOALYUnECOkJ1tjSNoISc8/eyV
qzT6iiIPQP7zwGkGQmju46VOvK9xHfsf08+rFCvDGnvGAr+ySlOety0N0vbjjGMv
n9QM6JcdmQcfNYI6mbD5q2rzPA5YRn89NlU3XC0pdKnpffp3VQAtddzv/AhnZGtQ
ZdY/rSoHt2yVOSl74C0BsOy02LfiAFPj7TtCuXSa6ePyZqJQVduOfHQ0KTWNOc2n
3K8/RZ+CUkNpavEBWJ3lRkIWNLaz53Z8Rip9Xhnoy8bSV4JRlDn4Fsj4bDDsM4Ca
QPm2iX4iPmhrcfQhXNT2gd+3Y+UzktD+AHsO3hHhtlL2aNx5zxgEjQl2cQ75UomA
8nlAQVAWxQ3MLWw2qmkRb7sd6Ra7LF7sU73DY3E61IB9RqPclv8XwBGiZVA1EdTI
zAE/jntaUH4CiuiRu/Fphpx+cqe9xP1AmxqffDym/LR2kW/1GuZeep+sQdUQtfV0
h8tgNt4SEQ6BpAFw0IFjgQ2iMcAgJNC7zBf6gvHzHGGCKexWQ0EN0UFBkgjPnCJR
eg1yrhR3a6VT2Ik37PORfKaFvJupBZfO4RmqlCADYcJLihzYhfDUWSVu856JnjA+
U/g1o95jz/XC6AatMYmGMQlDkeP4n5eHq6Rsk7+J12fGtI2ofCpu0P97Qp82ebdH
M2omUeM53ZtqauB/mJ5UtAxKE0G48AOApTum9w1s669sfiGRMMbXZBASyEJAH64m
KEeKN1lhzPO5MoEXNBXoUO12Oyz1wSGZ6f2rcbB0pyLuOBRnyO9NWW7/SbJA5HnJ
T8MmJ/FkUQK9yxf2/f9hZeMKCxLqGyfKtrOF4qOH93KpBxSenw9PBSuH4viGWRc3
Fdutj8C59AVG90giVK8EvSfrcGd+kSTBI6or3y7SUKtue9aL0c8QOVE10Vg86eVZ
uj2TClytDuBVwUV9n1UfPTj262Ilj6nlnPC/Tc0zRERsd2sroPCNPPumIjUhi2ul
jER7lIIsJ87it/amkhVw0+OapgTDthw8N/fZ30whDwvxa8pkwsFINmLP58qfzm7Q
m9tekpdC4/nxkd0ZuNJXnOnnx+Yiw3dL1Htqegrfo1PcImnV96c/kHdzEYXY3hdc
l83Y5di8iGNlIqIvp2z+KHlltHGSn+x8nAnAeGwzRaM/27mtpGOAjgCI+N2lZago
arcZsNSWksZlcnXH3GA5BYOaKOMOIHJARB5wc1cm9okDxLcfJ2p1C6U2HV0kEVyZ
`pragma protect end_protected
