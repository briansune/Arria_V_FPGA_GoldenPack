// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:27 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Quog40zmoYeKyiXOC3aZAj/l6TWcmRynqM7pmF+ZN1D5wInd1f9BHfNdVmg4v3u4
viTOUmw3HRFOIQ8V4KVnXXlcS7KGIX4LDdZz88yxAGZotQI63pk9uqBfZePw8jUI
OJOhm+VNWr7xT5ZdQ7NPYqN1cNbGdT21zdG/Z51Lx9w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
GNLWLiIqT8L4N3z2yR06XqdGFU06175EcYP8Gt3GCw+RygMbW+GfNdhEkfvLiGyr
T2Wkcl13HYXdfiHuQtp9wdXEPpZ/8/dNBEuy5zfLkQJz89Oh8Rcq4Q1enpwv/7ws
AB8j3p48TZwqzCReky9IR+z+F6c3+gSBbhTeCC1EgJIp9BmCLbJqwdzBcr4cmN3D
BlSP6X8pP41ZOLubFzKQbKObPztwkR7ZkPKmcQdOz6ArFVbnfjVm49Tf9ZyAqCkm
JjwMY59BoVIwbVKGLnD8Zc/omoLG45rKpJv1BAfHzvML3XoPqQAQpSpkJ/PYD/He
4abl9tlttrFMPyFwMV2hRD94KhZ+z7meXhkjJB9Dme8j3KqWajSB4mHeujKIww4s
17tSzLPkyVwSBasXSIzQ7xOisNYx8ji+aRSvKMG2sQyAcyCIrZxcALWncqpDSXZA
13OneB/xlDMwjTQ9yWKnuvL6h/SlTYCnm+C8IODrlAMzAld/U6Qa7EYylaPdWxT6
QEWyqT+eYkYY4Nt1I5ovMqDWoIuleSsmyhnkOptTyHW+dju1TrgJkrUuczGtowXn
GoVnyarmwhscVSiGSW4RPuYuuZWp17hYDHIZVs7ghh4ocFcYnE+OGICNX0cVAuHo
+SuiS2QjSoqg/Voad9DHOIyjCL2H1ISH9qc27Zg9Ov8bo23gb6g583JFWebGyz/R
cXW8H6JO88t6UXORQpbD0z2JhfmU5EokUaxE2LLqiYZY005C9GVn7cGsT04LvEpb
bz7fClLi1WlCfkrDDTS3uJaAJKquh1N0Xc1r/BNuYtH3Y4nrcZ/61L6rMDuJnLiq
UuM20dU37aznkB8CjUlfoSxP+z408vHBjnJmFUDOy/I+krvLFxWpvz6+kxyaBwR8
yt51YBB1Q91r+KjqxmphuwRtN5MSn/XPm2t4YMAFjeAsgIIjrwKDMeOmty+gBztV
5brJ3A+NrT8MuvwMEaB+hCdeqyYvzTtX9+oHeNVmdexLLOaQAN7OhBn9Lb92+kSR
782vpGd36UcAGY+kHCehCAoe06k34dlO4CWurZ32DKPah2bnQ3/hZSrQKpjR7npW
7TS7CVWkJ0N+ZXRWTzfhZVAi/br0bkNdulfNKMcG1BR/IyLev7DFOyFYpTCNKlf1
6WMvTNjUFAlAQ5/Q+elViW3NBL8WDnvLNkEolLYBBK/OlyfjftrrpRHiGvhmW3jD
CD46UpriwFa3fP99sVuAFy3otGPLhWlLLyKSYMZOiB8R1+YsJ9N8DvhpBVWuAHJp
+ZK2LaBdyUTn1QMH6REyxDIAglZHWBDAGquUgwsqF1PFuybpI2/ntIFBi6dYspqV
uAx4owMiWx9pYVoNTMiwbbRdxVQaPctgvM3TWfsvwqRIEB/AOvw2CHKjlidXIBhJ
s44ir1b406080E3V1ozYzZFJcrM0olodCFA4p6mkUZSr3fxlwOXSnuusKpfE5b3s
FGc4lQt3HIAlHCqt2mCVaMjICA9Y6Eko9UeBiVp+xzOhjvGNPCSaIvwB3AUQMlVK
fzW/iJrlepTBVQ4pSO97GsOZK8smt/pq0Kw3LPwWZNvBDSs6zhoZ6CUIbGGr3Ijz
X8TtiSBxSiRA95OEHdr0W99GN03VLScP+d8ZErU4xm/01oxzSbxB8EOX+b+0HWL4
NV2SBDR/VYBc2/1f26W955c8bg77AyHzZLRGvirOgJ33e1bRryDssj56KGb0kTSP
kJXVNWTrrahHvfc2ZaOB8x6KFwVqNrjw0V7Dll4CwTy73lj2s8SzOBW+mSGMfk8O
/EtGC7pCoX9Z6oCWjWXMHUrGnZNXdCpaENHXAVgnuiiETCuHRB1Woa0NUSKuM7C8
wxPrHZ92Uh+HDoclKz7fpjh6s8akg9ywh3qrPm2aCocNg3iD0Us+o5LBT2u/td51
FU+rWC9r+2chnSc7EkWeMCrod0aQYViNnL602/cM7VAqw5u9emWEyN6wfNEvX84t
uvtsDDDGYeyuVHjxVqDIiO7KbBZgD98YqOgjv+v8l9fgM0sxM3FYhV84h5SwExpM
XrfQP2taKmi6tsoSIxecQ8Ts84mohMOggmSAwqRg+Zr+CjBZYnG/5KZ7rgf6xLrG
kwZIztGo6DzAy7P5xb+ASR5YyOxHPS+mY1Zy3827QY0dS5ASUnjYupWb+I+S8u9h
+32+uYNi6zUArTlTI6JP926/DXQDZ05PLbINDDNJAbhXTC9gRRTnYiwMtk/e99tS
g+sC8nMQSBbfTFnuDShRr7fC4Fiyqo4ukQpvD8Sgbe9j44ysuumLRYGv2ncV3nwf
Zged+76UKtz9PRgBmCgbRE4MYJ4smBvCXMWfTEMg6xo5A98aubI8/zuf07sA+yDD
1O6PuHtPi1lBQXfQZDfeaRDOg2kapTyhBu3TOLa5oa80V26Am0FDautlr2VNK7aw
dA844hjcycBJf7CIzqp9ePUMQg1JvfQ65/qP9quNAdsdOKu0OWKpCAhKJjOgHcHw
pqS7n0PtLjxNlCGUw3E/0Jat1rmWlIKHeBWKWoHHP8zXGfXt8QXfwcdCO56U8Qnj
Yaood6eJwyJFSbVbiyjpnONU/a/hKQRm07pA9uzhgR+dtTRMtvRY26ZniuI7xNAa
R6JFNwK8QioqBw0c+k+B9eoXpI0UHvLbGgQWcf4sfvltCKDf3qOvN8fEDjdW+60P
eXl1F3avlY+DsHJtzUynuHUMVPRVZ8D79WP379jzXwvtplNIlMDZuL+pI5CmC+E7
RUACatnB0tLg5gUGgaASnKDaKCixxSZ5gquOR8Hc1bUkAnHPcgHPVBmPMfFaj0mR
hlBT/dB2sPpsJZIsFOPPF6BRgmWppWgMKjPlrs+FJzdylLgHAcMvLbhAxD44156T
BQiuVHuFPTROg+AuqcUcYxQg6dxmbQm9luXSsM5gLaQlliIxXGRbR/t0ZXyPVINP
S79ckiU+R9PgAO+zMStr8fnun/jKCuL/O//dlx04QxHOs04nZCdzQWJFb0Qmb9vK
n/wiE/eQbMBIXavmIu2pHpZ41FRQwH9irzt981oejSG6ZnMoPfmJYV5YKX4TcbmF
iC6BKIawC5foqrJsNgQBYMFK70OUbqultY2vkLlL8Pfqm4QytYp2FqlPk9wPQ0Vh
ErpINZq1k5nKGkEVMkGUAGueYroxN1qDse3oQ/PWmp84LVVeK/GzXB0SefxirK8P
1gOJ66tgqb4FQiCBXpq5rf+Qri2XyTeU8AmVEloG5W6Dic+j2uV8Sx8Vy1CN4h/F
Ra4es3ghDw0yoWSrWEZMPudA0LJS/TbDK45EKwgXkZAG9wBQM8PISGiMSHEpic5Q
N2O/VLCgrvJO5jSMuValD8UwdZbfce3SoJRiLyfhnISSYICiV57ZhkWMHV48NRJk
SUQRHS+zUBHQ68PG7bRj5cDwk9ZQUL2xV305x0gYxOH4QrKcwVy6S0U8cX24HbjK
CVP2iSjNCkPwlzZAl2AEZV8uVij7QS8wT3IHdHV468f6xhFnM/csBcRxWBDPtyr7
/Yb0rJMmr0fLeAcWk9eKtIpbXTQ7nEQTudlNSpQ/yPsbvqHACThI/V/R6e5Be7WO
6NUk90ruyBUvj7N145aaEEwwQf0dWxqRmF15ezB+vJxvXmOynoKGE2IyyxKle9KH
HFO04DuriAzrnhrnM/xjiUA9pV3Af3TwNHSQXX3BPlDZOfg7gms1PU0dIIsaETYE
e9i8D8szIVfa9Li7Eq1G52dA9kRRmOvTtmMrw4rDRBNsCM70L5u42WWYbeUppvpb
q2jp4Z0EcneXP/UsJlbXf+BdklnDhMcd9aqbSnRrGnbQx/Z5onGbuzFtF861EOJo
pLt+AsRElj+hFwCfpFlbhxvsSWFZE5Z48mnFvDqPag61cIrH7xYPr6fr1MlODZfN
5HRZdD1lMR6LVgcte9R+siMjVzuwUslreF8jLGl/BLUy+rYH3ViWBfSgxMJbfbBP
SoKo8tvcRFexUiqoX6qR6Db4Oj8JT6CaEUa4kleLTtZ+j4+BvEbpps/BisVUHESp
PYNYKPF4znmzC0juUZCzeue6GlqiHUsfcBif4CnIXMAAI+zIIeJZRmdbAsEJ3yzb
bmwJXWITipk5NgWoDeYD5A8BdPI+0Hvrsa7cLMZaNcA5ZsX9YdjUziLgmEc/T4nV
16tsTAP65wD0wC9uKL55Mjxe/QP5vaRsi0uMu1GYeooJdLYxwy9U3OLVCjYk4QaY
Akh918PjpcjBsgd+Q317/DTBFxpwegb4rJiiVg0sR1Hbu2JguKLcoQ/gPQd/NWQC
TFBYMX4gZJN+eBHBEhBSiPH/+5Op85jb4XPKNWgYNsxVxu5945Il/HWIDG4souDd
VUB6FYo4aaK/sJ+i5yGHz1znerlFyyLsl/Qab3RrPIFRaJYPckqb7TDPDCtMOf7e
/fKYNBWxrfpvZ9aN/yY3lZqRF5Xc7qQHcLCYfRPzxuke+iHw6zICqladbjHGwD2J
IZSuunW+QxgUm0ijcKjmmFtRMXipBWh1k4N0jH/w6mry6Zb1nVF9BgSYokpNSxd8
TZPhasfDjNq63MMDVecJAFxODbe4oBkY9JTARvsXHmLEaByztJqcHZLSzliaRHgM
RPdggol+AxCOMAEmqnB6zPmMJL7Vne5DOjA9Zc3GJ80XgoMOcqMrV+bdMIAOk2eX
rzmlGZrUUPZ1KAO5NO0VpgKnW7KdmZxvRNY7gtoXKbiiBiPixd5vW73KGw6DXEPJ
SRYYrl1R0xt3sCQnI4/kkUyUX2Jd14FSLp12jO+PFqD+xTKE6QwHRJMP+uru7Rxm
3VIMjRTSd9NzUSuJhcQqUX1FknT8Ue914IOkhm/Plhg4Zrw3Nn69JPPzRLJNb9d9
1hQma1mkGOhE5MFHMHBhcGbHpxzUGnYAhK649AlznwHKOUqKLTCNHiC7sAa/P06y
Ix3SL2gbeNvGBpAVdTaEqkEEk24XY6vDuDTNo92piuobMcqH9GZ1qkMp8V5QXN52
h3SkeCZ/PJiyae36d/r/3ACKKeiMIzB9cm2g0j8E1gDdxETLWPZvt+4F0Tkym0NL
ILcOJB3+rsZEiONtCsmHmowoHglOQr7lgWUAFzeG5mqOnPJJMOfdzfAHrpfwvH0B
WadWw0FJUXRbND4DbV0oQE1P40tRTxwKhKSGcRhW2IoCTkoe3ZtQegy4d9Wh+D4x
Fzjp5eibtXfofbMDWQmNNY4ZNKqKU6jUTDrN9VG6aoBAhH317vLwF3fzKfCIJbYS
UyfxFyePoIeT3ipZuO2YaJd2n+OOvE3gBOcsNvsi+yAYyjsDH1uKsO5r5ct/DzEg
Ks1zVR//xsXDSvavPdIJkPjhndnQNTQT5ijfRuvnRDj94vbNZWIKwimu9nMi0als
hUdvlhh4/7sNwZF39WOeZSZ3B6Tiu8+yn0r1midf9WdaroCbmYcJgi9zkXFjBsu7
MBiMpzQIqsnY81VJDj5FZDvICqBSE1z+UrK3RqMQla2aKulIMouBG8v77I2JUf/g
k1dpbcldar7YTc3clJcd3aB1Wv9TQPQxC562/maJ+i4NCxVPduA1FKA9nFKZPvg7
SqlPuI6or1GQvU6nN9wRnsqj71+ZD7CObDfUM3IhciKPknDl90M6gmc0RHppzS1w
0vr1OMXwe6tTPF1t0YACcG48NEjIIHqfJyHXGDpzZKtp5k5Rh2OXaav21HXsc7ki
xyxMrjzMN8D4FCEU9b52wtE1oHDVumGlbk5rTBmDxfFvke4q1Hv7+P9HwP5EfB3s
NbNBVeXV8Mk0fTe8QvEK9Dh71rPFmdwy6k7T9SKJCJjb8aZJxR3qS756dQPNRr02
Zr8qbx64QUsrPYluCzVUzSiH8Rv0tKS0n2Xa6znVJ06zGGr39i2k4wnHyjPZopbX
ntsmN/lMdJj0kUhb9lanLocY4F+EFt3m7SSfEQ/IH0LV1xtXgl9pcC3zkTQM3PDF
2Xz8HJ0VqcRXBX2n6mOKfvK4f77e9OrhFyj0Om743WpFcnE9bqHMjV3LfoGGMEoV
6yK1k+qpPzqYqo9t5vnAQ/+FzkRHQiiB32QklJCZH3GoL83JkoTP/NjkwSeAWrio
qlCh7lHzzoEGoYCK5eK3Qh/12mkYAjxqY6MylRCWdNe4kPtv6BVNcR5o3/1fFHAd
a3gIt9RKt1oWCPXUG6ukli354BMMRcPnk/qlzGbQGGmtyO3m0CdzywJdqb6FJc9R
/ks3FWqSM3JfknnLIuQv/eE6WyGTmhGpWH1FBQNiaz8FUSMwnfUAJG4d92UYDfIb
3NB6wIbSo7QijXCul9sFbbWNKRUzozMMEd/5L3i0TC6OEVqPQS9X2pOy57kzP11i
z3FeZG3WDLdFAoo8r/KcbAuxRV689vtRNq9WpLMangkGr8Oh2wjRr8rbPUxtcqpQ
utYOfal+6mQ15bwOkSOUXrSsJqAy37nDtKy0vesYhzh17gfGPsvm0l7OTZxefgaS
6XnXcp+wdvMEX0KWs2V1bd+VVV/G9MsC9lAYNciBv/E5v7xuOR2Ckdcx9q/ByANM
+i6XWYR9g1GlUNcOepEEqkhs07m1zjl9LKADqXWKhnCeDzymXE6jXd99Z67tt8Om
LXNRE0oqzo8Q3XxrRbmd/FQ8qCqYrs5cxfNFTU6+2E7wEjXEnTQUGu3IcQ4u7u5Q
PhHHhfCTdYXavanffsmTTwUWq5larbIR4n/6JE+3Pfg6Uyw+wmxdYkwdmJDonl5U
vRVgcTsRhX3kU4UcaTCyjljjjYuX7GTJioAuJuOttaKIi6drdXqABTlu3Yf3SUSg
IpWH+rFXdtJ93DsYhF8/thO7P4w+W8ABkBZDONkg+4hoipvb8NWSAtCtyzTJD9gF
7L70ZwwFP7vfxyKHWdIWxfQ6LftF4LnWboydAyTPNaMiMON5U6aOG3CuG+QZiOje
NiA1rf+qDXuo0MPx95AoXiZdIIPSmFgdZlXYJDGqhtzoLAw0PNb664qE8RAYtnTa
z1osidFhmBhBTeYOXkkua4PNjMBhF9NWnTsxbVHL50R3tNwUAkUBK+POrZ/Hohx/
qneQSfDdNVJUXij7iLb1iq7qTdqOJ0nYw4MdJGL+5W/o4NYgxnuPF342zFryp0qo
y2NIdbzPO1Ja+qSuHvwGj7pUlK8JQCniGmd4q+Y2Ga5zgS2r/Suy1VxXRMG3sCc+
hdT5RLvktttQVqZqOH6ymTd0Q5faA/jlyqoCofwd5pSQCfad4U7vDh8d7hOibOs1
DnKrtFEX5ueHwDKUqIwc4+TFj2ZIFtuSTrVf0D3QrGgkmowZpbD9RSOFXmpudCLi
la4UXDDCZ6AYz6Vfg+dtymMii7Gr58OnS6bveRlpKeMxg/VscRomtF5D4q8Pr6OV
+IStonrdxQ0va8s9XqPULdwIXMEMTMOffCGOhQvuJv8fnBNji7mxvHaj2mzAcCQ+
9a7rwmQL+lNUXKB7Udso3aEpTZItF/np2GU+9DGxxfr2BfNBZdp/brGrMc47DEj6
5Zn74gT4u2P0hbWFjEMixK+ytJ6vLto1iXpzHGee/cxaw3nxBL+UFLZ8dvG2IPqU
MQKUZNvpNb/hGxZ3ygyTu4dwOikbe/jWbj2O/eM+IQFeQ/igOmA4OYWdscoJ0Ag5
u9oZ977p4XjlV1EiQDZRtGckFYuVPT5BjzCqzFhMKfoUKvSjlMp7mHfcBqO7lGIg
gHhn8jL3udZV3fvEP0jhK+tBlAmQtLBokwosQYbRPz4LPah7EkYhLdkGiZ+bqtJ/
tQfuni/7euySr2RcuRrxzHX3gFKGxNgh7YQO39QzfjvScU+RB0VVuSVSS7ZsQC6Q
Df+1zYl1XBtoTAhy/YgPYh6hihqJ1XiGB7P3YZKLg3PmZW+XgXl4UXRKJv80SFqr
x+NXP/PN/yk52YU+ElU+IkCYjANLGIvFb9oZ21xdb5P9XG3OOgQ8U+eZRwAkxUor
EKpu40hdhEO157TwQlAIfb+ihMmjKAji5TLkRygzO5lojBqvGASQ+r2/r20RcoEE
lCstghXcA7cjlCRzw2somyY4kXxSNNHULMqbjsxjsOLhgbLLoCsH94qk1GKAu/SW
M9eNbKhdY9r/li/h9BTGGffMVhZgJEh06aJ5iRjU9/MWuzyNzwNA4pX7EoD+A8oz
QVGYFx4XCN9zN6//kcQULqP8MEhbllWDNhr/7pCcQStlVUR59bZtGJ9vkMl8Hf5K
WyX4Kx7kERHcYSctOa83XU+fgfOeRh7Cl3QR2bCKaTs/ZzG+aN5xQ77ZSrez7Qq+
nE90L57zKPAWEdExCUywneNem0NXF7rVi7tyJklSvEz3VlKxT+SR3E7gEUTCgQuy
XLtr2ypBc7P+VdGeSOwx/v1znIn2wWX8WNHmt5pHX+tQ7skmsklcJ1tdrPTsxZKS
QJfgDBbbvjoZL+WBsvHkOBqsvAJk8syhFcOHCWcCaZMeaXbrDfss0OVUF40PsuZ3
WaHZF9KhweIOM1KHKUwgoaOhF1HYV5Wc/Ny9DMoTh5xvQbi5SwZL5RBFsTLnAOTa
b1VAO4QneW+t4a39eIWrG2pwwdUR2Sffi3cbCSD1SPus/AH5Y4hVT30fnXv613rZ
f4tfH5bZAN9WwIkl6UMaiMxNEOhUPV8btl+iQTQQLqwtlniUGrR3iEYXnk3ZVJqh
rVQiS+mUzrKCTs9I3Y9HmqaaAqww6hneaqNWMzSp3u3HKH1v1lMtDQvTUN0PyJI0
TxC0jStiSa8zeIFB9AXaljouiyqg9MV/h6KHRg68A9DYkmHxL8DNtqqshOZ8X2y5
OHWMj2u777fCvlI6lNmgulwb5bX2JIqKRf2QQ+MA7ehOD6VrF/1dfXpW8votd/ui
HLLeFUmwMVL+bwTwwrEgL//n9Mz7ZWTA+3voniItKlz/6uDvAmmutJlkd8VqXSLY
Il1Toka/bCR6k7KGCOTjv6MxFG+P9FX44wUCZ1srwzVGfchXsZRRP8MVI1j1lKON
Px4cxNEYf3AvA2RWLwe5o16ONdRAa3mZTu5XPgcruOPkgqkUVkGQIdXtNRvMhpDf
MrC4dAT/ce6+bnRKnF80hYxeLbJSKBoMd10yVjvzW1V1nzJoUeb0IR0wzxsQyZgy
ZgGrSn8N2irx5mIiLNf1oGH88n423BC/i1D3jAYi5Ob8iFp5gzPY7Te9/b9HLyFv
EcWajixvVOjXx8FINy4YtrIwL48jvRzXKCLBT7Z1F760M85IUqsKBLC4KbVjH1TH
ob/VjyGM6L9g0gEpGFf2kYiGjbsxe19XUav1FtuSmfkTU4MbMGfWCzwB8X4XxCZ3
DdCqCq1+gEUAZ7gMQO3RvxveGkiMhFBvVP1pZ40fk+wHHuZ2ENcf/gOnkf95QMsS
+ODqLaAuYJWLSOWQm58kY5Qo+UK377yYkL5KO58qd7FO5kPon45b46dCz69wQXrI
/hU/SEvt/ndagCPD574zt7VZmACVd/B7Klat8LtDYpzQHj9Kr2ljI2stycw9GTcy
iuOEaNNN8mc4OkkQOuVupogGRqlUlwFGMl3H9mzVLrOsL3H3wAvYHchf+SNgn4QB
nHz7CYbKfXaIaKdPai3QahF610gMwkiWvXow0tFOhDACNzji6nNUhqY6B1Gsyi7h
BR4vY9lA8lzgYeQFOBLk8pDWr8C7dpoGS6n979QQaT5ledR/7aS0rSv7zgdcPmel
P1QrN7jHTzR8zPn/SpZuqNnRhbmfFp32lX4KWoIh2Mr2+NB5k8hjfdzu+zhTzroy
YA9Vxg/MgmTd2PvcaJLwXTUog6gcEulvNbzv0PWBjso0nsDt5aRXUMbduryAMuEO
/Kt0nBg5egzh3dRskuwR7gw30cuypRQsoZmGn38pjSmwg9wQfrzRg6QME9/yeo0S
3HSwAvaVY+nVC6/hixw67lIsNr5R246IXbmKCtA79w0bdkkEeQxFTK1UbSrprMIU
uss2oh6m2b6bqAo+MN7caN/U3iZIIbEXjdntBVhJ4/Ag7xvlXM877awAiB/KeJOb
ft46UBCl/pPcAqsdIWiKebGO7FIJl+6YgFoml0Bs1ha6I8c4DMr/fcxFKhmM43PG
w0Ez4eG2lKmZH/9cdvR1BoHCGi/XgKABDVGzEQ37k0T1aZAhuSWS8hqSxKOOJcHx
sbtC9ZddbRkZ/LNTFtgFBD1geVsjGJTB8qF7NbqW9DUuPmlT+azHq38c+8XM5fSe
6mOA6S5YAQtVFL2TEFAET5OiXzYIpB0heKb7xoPcBUBD9OFkHqeTaySZvDYEYAX7
68rXByLOnSmh5aYFnwuU6iT7Ii97xvOmg3dYRSf3lqdngI5jhXdfreuIROGhmTmC
D6XIIi2bj24YlCmagibzSvUh7CB5f9SNXEG+GM9zWkoubIyDlj0qi6EhAmFkv+Uz
FJw7iGMswRKdatKcImh/R181mbPkvuMtf9xOZ5mxxsX48u4lVdOgDkBhiuLWqjN+
05QVbk5wSJa1dwiD393V6+vrDTIQou8xCengXPc9kSC8c1QCzZy8B5rU4r0wy7yt
rpl7OWowjQXYBElphIHdUGDf5GR5XiUJzxPimAEnt+1i8VBunp5HtRMDPx+3gbKS
w2KA3YqzZPw5LkxFujcCFcADYt19bcYd4+0hi12zU6JbhOYn58d0fQeGzGalIITm
3ISPYsC+tIphS5l+fgR/vSdjsO/LPZai4hzclfALEp5OMkg6Rb2ZEU1xZkcv/FQN
Cs8+ht6RsvJRUay+/VQpPPfmvonITCAzCLTzaftoyOTv3YXLJDSb0WS3uFD8bWUp
VbpJF1X+Cg1TuzsaKhFluCBRSzPLrYfBzEiSeyKil0pMXzopFBl/SRxRwksgeenM
RvowtiDWzv/enJJODjl1nuDZSeYHWJgMqxwLM6VRW0B9GUY646jMHfHeGmpFeW+I
OJazX8fB3Fhuw4DSBisqHmhdx8geSXyW9v0WsMS6GcEMfgMgBkCUXFsgL9ewUdsL
KFiCDEnEpUpcjm+qeN17DaUxASHtWQVIO3zi3A5q+uKXXzDDWeYAmfFUrmS+YTUR
E0qr+kfsHh2UmW1vLSqehVF/R94uKQs5Vo2RO5XS0R/Vf3bLEQmOxFRx8JDGjgy+
tHayCU7r2/oX2asigq0vVMxu2Gp8KyHGUAHGKRBiYMFFhY7ZdVdViJBKLag5zi6R
mHlpmHtVslvdqSAiBTwRu97Bkx8SSiF+8QCvNveaplxJb7+w8xcNIVlKQFGTTkSs
RApJGw5ddtlbhkin1K2adHC6D1sbFZ2AKf+UCI2fFlaXf8/LA8s9YZdx7o90vZkY
Ak+33BiINrEccGtqpmPNcwnW6JbV5X7FpccAN6jmyvpJaNqnsUtwgDzjUNzFYb3Z
pjBe/PYg3k/Q3/J8OWsMfkinILb6BgGeNTjrYizX/ehK1UasBCyIGsaNiXaDEq0q
SySTZzsdmOa98BeG/FIvtCTYcLvONCp2Ke+WF1EWJZQYoWhIZk1mHXI+ZDZbgQD+
xgGtYKru4rguK0BMXOQ7IaPIKyAnPz/f3dYLlNoDPhSheEU8kTDTSnbVJp5liTDp
Y4Zq6yLLkIuw8VyR1cf0ukRF0W7afpdxw11tLwybxPUhRsjVk+/d9QDGs+1+xN7l
TYCJtEnkq44akVfP8MBbWC/YLH21hW33A/CWhLu+8tSG7UJHc+p2tgjuGGCLWTIu
vHgWoSpM/mN2btlx1/AHmz9YIEmh9dgeDQTpEusdul/zkDF+3W+4ljH7E0FiYvmh
2Qtxmzz1peeZSILRNuN/k20OBCr/a/z/BlZkxFq1T3cxGSEXQhRxXmoJSNfMcAcn
DMhR6YopSSFseEZnkIfE9Ekh1HmmVgYl26BfECCZCDzYq+uVdhCp0NW9gFPOJss7
j3rzTdPXEl2FVTDeI/l3MmoDSHsE5iVZNKD0y8leAHoHjHYyxOWFMbhQgss/8oUL
3MZnOBFVz9HQ7IT1eqoZgkfoY2aWKUjz0t/jTsp8MudPds5ZHqkmU3xTT8jAjZ0T
+sUq1VkJBW3EdnU17rFbE+TKpHUajcDwPHU14Ied7UecwXBcCbN2JQXhVuILu3Ps
EBSIkwWgbk48Xt3wCuywtQmoTxzluum/4oVs63GaXbAU0Ah9Q+EDU4hp2KANJ2Up
hkgekCnnQaM2ryMKfBDGbFDshBiiD/ItqSfsQ5ax+coECXogJcfTtEJquoycRpQz
NdwHbHisXN65vJE+7SMVoRGaYftZgR0MYG7UX0W8lYjy0KSHXwLUhPaAh5ze3aUO
Q+026Ri8jz+kpd3k9D5J1hrPl2QWGvVZ96ky35/rP5htZhOWikGrQ1LLXdIMlZHx
5f/xlJoityLCZm9BDNjSseA6MlZirVpn0ycLOMvrPvhZBdLgN96v4HKzHHffeLQ8
qNS9Zu0Slm5WbklnpgN1VewpblGIK/StOCp0apcM7M1tnUm0dZbi+5ZQ6mzfnFij
Qd2XTiqVwjyKQYkXTWu2je36g9e2n9E/LGPHKJ4k264njtv0gqZKupJIZcH5VoWd
r6kijBGG2eH8TRQ1ZdCwoBFVNJjHoj6xhE3FK2yz4AQavATb/Fbgl2l+WMAT+6lh
3NqygGbwmLMRIYK40iYmTdJf1F5e3La4ZCyM17ch5C9RDBidr0vovcmHHO8930nj
isVXYJ1XTo3XV1jR1jpTM8arQG6H1hJI2GOIHAI/MPw3GHB2dURxbgAz3DWGvw6H
XzRAdha0Qg7VYdfS9ELkjAI9DnXWiFTu1wqlnwhGIOUDtR6VW/mayX+sDZrAZahw
wg0ZUc8/2WAYF6Q5OBmndazLE1VIIKQ/dPLtfUpYcZGlAtSGzI0PKrm2LyH2tXa2
XuOZRVcSQHRmfh5GGL19Fr+aE+Hb+GtwcYbChlRQ64GxCDmD/ElqOu1dCqEXxnSF
X2bJyMpU5ezTNM1z/eGOuY/aA/PrAQkryogAihAtMvhxhl4PQNF4pJhV9c2htYUj
3CdnZWta+tRsVBQUGxYfzxOvs7JrkxkE2QsOnUuiLFf752bFIyAEXWebZUGrcCen
B5+Hx944+2eE0d2PytuyJjTtrtxd7WeXGbRb1yKR+1a1Dc6XMhIOgfDaXeqGyKn1
mya2020iLzdb5e93C82XsS+UqgBtCC+Uo7Ct39eZq6VjF5cqGx68B2yhmju+ywzW
WMVoQZDma3R4BtfF28o+OsKsC45x0VKuEnT+M9pyCkQYuw+S6hE7Oxm7RSTkALO6
s/e5s0tdID2jvDOTmitUBCn3WQUFbvFDFMXUeOPVGvutBieYW3vK/2EkRZghwiQU
/j6WQu1yFVvFC3cSSNK38mkEODkbyoJGmeZ8st3buEW7TolKoh+o0tU9gsCd7ckb
R1NfDXcQfsejVGZsiOSv9DRi1rDqws/gqnane0fE3W5pp184lsxC24M93CMbW+Gw
PUjj/OXa7r+CH3AeI8H+dx5Xc/avpa9EZoS8wuA7g7roya5s22mHePA5Pf9Ob1Xj
Ck8xZdeWnzO65jt8Yvg4B3YmC9PP1FFr0f05WywwG4Sn/1nX2ELVLVqfKnbJcC67
ZN80new9hxY+XsDyEDhIdiT/QVrb8uNQCzbi0tl01aoEwGWGH53O1l70kWfFlTww
YDi+I0gE9ZJKx5AKMZyJd08vermV3/eA6UH5ONKj++E/MQIKGcFvM0QAOdtfMLGv
40ZwMSlzAwuHF3llcdJPC2sRoERQhp+9danVpeQDcME4J3juOroEGFm1vLRe7Rs9
s60jNzfp6E23GRNYwoMjWjEWkjujqACl89T72Z6tEqyVUZWPGAuqxuWtUI4XxKZF
FzZHCv6Bjg+KQpANVSRkY1PVRqxj1gJZjd+Fq3ghahpzccGovbymNyd/Bxg8hHya
I4+02+GeALeHIVJbWG/j+UzQKfKHL3u12wrBBIRgFLto36P+ID8k2kZXl3e9MURg
o/MgCX614dwE73LMq1zNEmmXFMOznxqWEB1G2UTtMEIG3rNQ0kjpiLkYkH49K7e7
I9d7uc/3SBpbl7MUo9opqVe6pLz0Asfn6p029eVkj+SlLJCdPMmSBc2IN/zDiPEC
P2yapGPEHgxtxylz2LUn+XFkA+Jb63OTWkBhYoYyBse1KB/dDQnm0dMKyxXjfYEA
wcbX4bR7/M5rmw6zDWJDXTnZszO4PtWgsBVH8MUM99BxBF8SM9QHVyH5X8qd7R7T
4kj7L/QqD2jK2WF8Z1hIT7nNtWTJdY7mwf5h6Yf0bQJ+UiJGY77knlDwiJfOAf1g
zja8pXF4z7YskUjZnkA1/DSZoLF/t9gmuPBKCCEcsM+cXYZpKIMKta0c0FUzdwdB
ZimNWdRjE5lbt+RFNnw0B+G1qO1J+NQtB2EwIODMUmZisWgO4q5jVMMI/18c3+8t
rZ8jpQ8+RkrsRy2Hp2R+VPaXlO3mi74IS51SzovYxdO/G7wTRHCdyELifLmCckCe
lZBhCdKVCQEIvP2pXWFXsFMKr9onk5QA513vkScACJLQJAPhCvP1I4N0+4t2IpKJ
7l6ugvHdD1tOQMIzDG6oXZ+TR5Ty/Eat0yij4tZVe8cApKRgYzbXCTECS8b9mYk1
3Jbz7lCqurhFlTDha4hg0TaS5L784nuYObUzvamnL2jaiMQWVoN41iHePL+Zi/UC
X4DXuBooi6TDnCOPLUq+huaBN2XK2w3/VDVTG4omRlDCcVftFS1BRilBnj9MRPbi
iarNBfsTiIUJ+EgBnzjktOaE98UY3sqID0yBog7WhntACNSkT8RlbU11Y7KpVygE
p3DfczM1OgjlnVYZHXO/8n5HKGofkVh150P5/fbaT/P+q31jw3LtldQcAf5BoRQ8
uGy2A8S0y0+gHHO7gkvSepUufkYVrmcM4qQfOVOiNTqivDshL+awUBzwU3BFNEn9
ZlPlSk7tBACqPvfvGbfoSu0OxSozZCHv82nTwqHKEOTJb5YHf/UwXsPN+Rn6dJwB
qHNoUKjDv/hM6OEMVbXfhls8tnNySb/Yvj1RywtmPVyo3kaNez2a02GaJVQnimyi
a/McLTKqnLDUl1NB2Etro5bMdN3tmGXpE13xP+4YKbPoTnTyMFUknCZ2Bbc/BvzG
7YKrQGTKU7DW7AEFBSeGnGtWRxq9gh3L+Ns1WG3369yylE32fiHKLQsCMi4s2k4B
fHoFUUyhbRBmYVO5zUTtxWtKZu5s+KHFY1JXy8Iq6LPzoWSGzg5uN5aS0BXENKk3
dDm7fVTwb1E2cAKpbNKOoRoZLjISrH8YgWnuyTSzEneInrK5aS5GLuVH6lqJbL2s
4aVYL1wclVI/FExPnlJ+MONhItMDsC/eeOD2U+GNloacAgc2lSat0tLX76lHyvKF
JD4QVwvXzM0v3pm6PXXmhq17B+QUNegh/5JPwoS8XAYnhDAO9vadvkHsd+PTf5GD
CGmD46Eyyd1W9mrB55bpQXCd4OED73IblhNh4IhCnDzoRWh9ojXPg5nydaLMGS3g
DiY0HJ2n1+jrivd/sWgVnAvfI2G9Tn/fnHNezHILfoQ6/ff5+dEVQnYnXIUoZYfh
bfT7SDOr+PwKNSkM4zFOYKrVjkDLdCXEKBYD0yVkFUngOBndTpF30wYXEX6zttkA
yPDgvsqn9yp74ae/yyDA89jUac/swhv7zMU/CNHJlXbB7KhLUrHPQro6QqyS+YUC
8g/AqN6LH9HpCD3lG7LrumpiiymtyALxtqWOc9TYd/ClQ004dPLZqctJJphCb6gP
1H+c9QsgCvAXDw5lu47WYF74lVZxsWbSP42ygiAnxHNnMZ503rcJf/7VUVS78nEH
2rYxb23JoI6n/a7cJQuXQI6ln9d0pXegGD0fhbEmgJUwz/mItX8AY5R/bd7HQRnu
vA5qlpsd5b3htJOyVExTOn4gcZMt7xePt3KVz5P7fZGgaMOamIS2QvhljqhXqhJt
DMRaBwP+71EX0yIZmtF++xiQ7g46yj3xHXiEZm4hkCSh5AbvUdAmF8t9Wr3O5Qvu
uw9FQIscdysIZ3tD0TnOlNaieDeDYlf1O9K4/8rGVQA2xcadvEQ7K4aK2sKBR8zV
EBURmCNlSePKkv6ceDZSCYxqP9Jnlsn79mtLPt4BvlDmPJ0opnmohgdY7Uw8FBKd
w7sRoj66pkCzRcNqI+1vEpGz//T4GS0otG7ZfOKIMbZWV8OvzPDBP4UVjWhZPFKf
DX2q6AiaVoeu/sa7INViNdqnRxQsOCJSpfVbtRoGlROevKXWbz9jSRDVKpyAQlJh
p6ANJWf4QvLaExE+cj2syjBoVnUu6iJzDtnbUrOl9sC4iwVbsnzk4nqWQrIkSYhb
mRI6WCimpdz61wxK42/bOGwPIJfwVOqcYn2i8e6BA8lrpj+CD0/Xq8fqw1zXPJRS
Od2UzFZJj7ZSD6nG1LKENKnM6hCgzIOgPIED+/4vGrkn14kjDUcGy60OX1stfXaa
jUPmgy/99RjWDcuLMvZN3hDLJRY1jocattLiWykI9bt/NZ0/2qXwzPBqASKOzjiI
/Ejk6v8J4RHQmblT+K5E2NED5zJHWka9G0df4suU3k1ej5sgcMNXHGNX8yKmNGsj
0TvXixmAmOCFSxUFbLQUp1mct3caYeSNDNJj8GXVg0gI4rThO0ann1AFLPM2QXR4
XfV8qw5fhX3izLuVDHKOmKpzjxCTN4R1MuqTiGLDfelt6jnZkvLWHAvQT2HnIe7v
6SGuO5eSXzU+pBYjd2aNBRSzvbbfx5DHkLpWj734mEYGGtl8MzvKpLxAinKHJSSY
7uG/Q4K9EN80u/9pdgQr3g6tyHxFcXcEu8DzeHqp3XvYzFiuF5s86rHrTqmflvmR
W4/AqkzMn5b4FeIWrZWcAmOdCd34gpSWKK9jMs+NYA/9cW6UjR7IMx53UHF0jQDQ
d+AtC16ZSjixJnR4KyDkKA+IltHG9UyE+GjImQyHGny+Tsn5FXdxbtSx80sX5kXC
OxqsBAeKkcV1MPWjaJXP/QuVVBcxE/wemFuQ5U/ybKXQOIsGwD8SC2/o0ogE1OGC
ALgFdTwc/N92k/UpjUmz2ImFfjHQUGsIJ8L9dLydhhQi6NJH6zigb5ZmaDU9PLv6
RkMDhFQPG4kfTssUIXU9pLR6HS15kj1AmkRZQUT2LAiPEC6wkmatJGIz3CoSjpTW
eEbWNAE1/LW91wnj0ojaHY9n3fevgg+jqxMNGmQysBw6eISW1GVO6394qHuvfjKb
/ufEfD57JeL2vMadYgV6hXeOCEQaAxg4aT0qWRSLXRylni7IUKWaYkD4ttOacKYo
sKeE9D6HL3Brpci6lKBXVECY/F7ixu9xb+w/UJOUSxWAn33Yqbl8oFLe8/e5bvmk
JagOd7zcY3V856oqaV6VWH+4ubQy+YbE+zcxFFN4ihlWOYDc0OUP+bvN9jHsi2rl
iyx2pMpd6wwlIeQhYn+Psy2MaIzt4hgkNmkHqVGaB5iLZj2e/WyQpb76aZL8yken
us4ZBvQ83QZLCh6xEMH7xBt/RD3LcJNrMTs2PrgqEDeQPB93OFSns76vq/Ie/BqU
9jJb9JZZI7klBHlb8/31M1syKqvrqbBuXpYFkx3CHzbeeesWCArJVwO0uK34ZcoK
gVnHdzeJSUC9ibYCsHVnZ5RQT+s7t+NX9XPCvdzC8rAXZzVHwEc/AFKrawa6hN8W
7rCRdFHSPmf7x1IC8PhvKrqRIFyre+EiF4bcAuQO3QdwhFz6LSNvjY+tJH1+7pN5
leKb6zZBG6jxjqJ+GdGGnuc4/4GGfxpjnG0aB31vA+bNkFwPDJ4RxTEgLwOJoE/1
beANJMmis/p1CxlW8bLMoAHbjmfyH7aOjnlHq9qupjgzv/s+ket2fqoLXaHbBYzW
FFfqNP1/KLLPecdse5eqvGxFPYEYh0wTDBePxlpuuGz+sJ0GxlOM/qM1t2aVHktC
s20sG2L62vmlbuEP30vqLs03oJoDvf6ak6rvrZ5aEyD9KhrnFG2M6oyAMsPUTsdv
dzzrzmo+LQflexMO6+k+h0cyl0SmjZoO6LbsR5Mo03ShJImPQCZcuJRpqropc8vb
i6ZU8QW8ZBzMLokY6/pwv75xCC3xPxkhTL0wX9RN5PrdiufqPk6NewkexkQDfhyJ
fSso2ITuj7gS+Znt/TmTUz5FDLgHqv7005MiPxSHb4EdxQy87+XWFZme9JzDLA1j
kUvLSSxVWOKCbnnIjG0bb5lwQwSPwJSbEdM3eUV82jFSIjrkpkQcJu7Qg/jH/lb9
wAWjAA5hAAN6KoRX2yHOEOPRGP9S+ceHVzGbbOBdxqR4jpo2AhvenYqjLpaLZpWo
jAxkKVg0ZjCs5Z+X7G4Scvx3F36fALxQk0i8P556mrSwo7b0yZk4DdSivg0Y3Ybt
2U8KGD0HZY5r7W1zdQ2UCxwcZg/rjKtZspK3Op4ftafhrZ4vNbU9h7sxjsKFfiuX
c4ka/C5AveXgm6nwuSe21hHshKp3ZBOuREevvUrXdEdc893mLaBoFfy2M0lmgJ4e
Li+fVZ6NMnd+lI7WmXAO67hNs/FiDhPZkBoWlmyjJ9u/u4dQNFSihabTSkPIgegw
1iydo487NnmrQAEJE6FS2h7C7D5VjCcE4x7gPo+TO65+3TftIKSW/OxSR3Wh3mwU
tPLEHSvkuhBn0BXFDIXI4dQ2G1VRJEd2HorrK7argWKZpKavCmjT7jsm+IGeqUHH
wrLvktpsVmY5kg4c7DP9SOQSxY8jcYQrsV3fySLpkWum/wjBHGVl7BgSXfqrN/bu
DNUdNi/q26TgUgEoUO0mHCXvswh+m2Y4msrFduVPoBkGNgjP461uEDGwUGbImQBV
oGPYN3VJl0CR0flZXG/4WtIujFuUrneAFuDkfV/7qsrwyvfudBD4Z36+WrnnGOIx
vOfVz5nxhhoHThpZuOyrmciPmA7FHv5tWmp7Uoyc2H8zla8E2B64mFmgfLtfdea+
j9kixtcRxnZC6JFSfHqQazRT8nF74BRvPudjqil+duXj9tryMWg+RfKXGhgSThmB
WqZhiqE+bW9AN4upRdgYH8Qo09ov4/mTAaJQd80xKsVg3f70fDtvsqAFhR+qv0up
9sGr4Q5DcpY2CWtu1WnlIfO5voFoQmr+90B+HIdslT/KhaPGrJlECWcoAsRDGnuE
OtD+GXbiVoZQMM4kO4c7ZKzNA3R3MpkgJeFcIdOFTLmKI44eVIrMeavdiUz+/lzj
ng6qZBHU5PKBxmoJgYsp7mFCjHkfnSjJHViOf/K4QZ42MhRDrUjM4YwdG8FAMq1y
35X9PjxlmVgiQ7ukipJNVQPKEhPqVMNED6UBTM3mg5y6HCf5VgHRd6Og9qSpNmsf
9cXMxY4oSSiNUYXl+pZEg1744fCgc27KS69d0VdZ5fNiWiD6QhGH72h4XLnf7dY7
wuxTmQs8qnYrP0x13qPce8ngln4qfI9hs7N+O5UUywxkuZBNKSaY0EbJ7v6UYFdB
xbP5Ntr3HnZcQAV/yVVS+cCcxq5+DWWC5J4bykVI/qLJY/AYbl8RP0M6nSUhllo+
xfjSIKGSBcuwiALc3RtbhFaoBY82a1iaFrN4D0c1nY3NL22k5BkzVOUfiJMSUJ1E
iXINdKm/vremarPSeTG86ov36PDDApHEB99UsZSANlLX2w6R8deqooLnQdF3DpKq
PxmZ8VhpIJSO4E3VOOdEWGsuz36YJYQ08O73361UEb0yfE0rXBsJHPi+j/cCNqbD
JKMaqKBeLmPsrG3lL+YgeD19HIyoCySGdQ1Vfo1SQkCrZXjiho7dkcxpZY0te7Ej
m7IJhjiBT4/UXM6muhMLgfs03xPwpDPn+nRU+4MVrUjaIPzF9uuC6CNRdLxmoGJc
TYOoEhqJhXSdfp9uCcxrritYmvQfb7rlK9XggiTbq7wn4IB3QzYozF5Flmr6xI3q
qNTv6O5UxseReSGud63dSqMIpHKVhb3AAD2Dpoai8yDjKaK4A2Sc6qimysEuYs97
ahEOfJw8dGZoqdwlx62E2INO4yv485K0CZvFys0FP1czDAMOlLVAvIqlM3toXdxJ
aNLdYURyq4rX01zXN82QjOGWGW1sW/6kd1tM2lHTi5dObGq6Af0PBXUz8R2cdcsp
yA2gQhXL7viGTSs5QlxmBU2Jm6Q0Eu0ID90Yr4FAeLZgjNv0V/U6Gye7HG6InrWg
Q5vdz9rLHlGlM+Q1WfUG+/E6e7DvkDC2GamYxzq713ELA++erZ7kMMu1qVs9bzKe
HW9hCnlJggORpfBWBwwJbdak8nApTXvNQW4PwEE2NGOrY9BNKqwQxdQES5fr4jjh
hyzDrCKjTYgSVTTcFPTJAh7/RW5rpn6eXuv8xRvlVdOH4yxzdCwbR6FC24th49xu
ONeD9y3eX7xChQgo3RpodJqmxeQmSVg8pocG4mSFrVIOezsSuhWkKhYrVPktp+dh
fT/8aPtU/gFnceh5ZJW3VCqkdbCJhE8gyoQ/C0ElRd8A6rDI/u1etBIo9Yn2WwP6
73RLuIbOeYUf4bFlhy3zXNFJJVcGOSQ3yeTs9nNzFN/FbTQqmc2no/Tj/T7+noT3
nMnsI5piIvm7BS/gQcRD0cji0ZUmF+MODEppF6aNauYXxmg0yTWOyI+TrvuNkQTP
OrB2kxsFhoUnmsNZmLu53ekhlRpMa+K9KireKu0J9dhklAm/jbJPuWx2MAQY/oPa
+cxVtP6ObSZJM6wfhoXJxrghIjBb7Mg6mKBlkUIpClNwEdDzZQ9x3q4kV7vTwI7U
VUU3lfVy7CNlsxgh0fcqVW5wdbzuEEcVcnAD+cogNTMwUISnsnpyMkpi9wxOOzRz
XIPk18SYVeX3oUYoFzuSp4WvsshLLdMVqCDJ/41OwRSeBMaN6IJ6en/kbYECdLGO
rYDZvUQWk4jEIA1ZJimniAUaIe0e+0kvj9slxTHkFXHX/mXNN1plUs2+oVByZhA2
KO61WqzWC407VNOeu4Np4MWcNfIQyCgUiuZiEP7oEy88kl+gk8lgbPS7BVM4KX7+
xDHIvwenDn2UI3CBHvmMMYdYDPSwaLXCfHykv/c/5yOgzap18ftEZV0HK/Ylu4pg
LFhtfRYDK97spUnBrflu1O9UCmSkTjgydhC9brZC3hW+vYhXtNKG6vdPjIHeH6qX
c5cP7G4efkzN+4UN6ZNjWbd/kYRyCP60fxZ826VHhP9C+h18OS+tAocFv/WF6odg
uzn2Qliz5IPENekk2QollpZmm1TlLaxL/xUcGKD6+hPuBJM3OmfH+vo28QvWeiUQ
79WyxiU95ClDoMfFXLG4RahDUmsqFpnFF6h/nn+16eiXYH511lBfR5uJwF4rWkqu
WlD6uYrh8yRzp85DPVGi6y7w2HJL2gdS7acmWYYoKPtV9P+AKIa/4Qy2S3bnaA3F
l6j34obHSoIxX/mWpzk5hMx/MIKMZPkg/FoqDOLIzMlWH/Ml/pRAz3+ghgVSatrF
d7Zg2Rtigqk+1PDHI69BR2ZIE5qKwi2TggeIo3hahPQhwIsrr+mv+9UmwjkzvybH
ygOTbM9ScXipWznfCmsv1GwoJipnKpT6d0ywPVw+TmKEtShOe63cRaIrzi26hPc1
Vas7V6SnlPuAW4wIxXMCyXExjko5hk9hP0U6IylEpb3ynAuxtG87MrkMH9UXN2PL
wbdjAayn1bGldihN26FUGYYhsRNe3iBTQn4foyu1AVvX3UzDWs8rHjUVkaAKKH7H
7X/BpZFBNEqqFaCb5qMF0fwjmwodyA47lr/MagSGMzTJGJyyAvd4k1mJy12M2Q28
NmIVkX+cNIfZVzggjFehU47IzAZOa3caVbNt0tiGRHk5X4VLM23FM7aXJ9WrnSpo
pJwW6y6dF+KUmkMxENk5LivhVRJeTi1/NsP2ACyPIjPimVh4f/5CtlR9IqSS+31N
a+38amK2GekkEiA8McSSdewaQmK4ZfxoRhaHaBMda8DzSx1I8qDVEpk4/T2dUPsc
3u0pPEDS0Y7Qh+XKYZnEkM+UGXh28I6Zfpc6SeR+gah5BxkpbrTmjuyo5lcasGm8
EaxALML11sqc8Vl2WmIjI+V3uy6BqaUV72cq/VsKK69xn6nmIwf2++7hUG5TN4o2
wTUJOms6I2MSnenL4WiRvUvocIZL81+iT/x+d2BKDidcvIcNZSGfRaLgiLrPLPJY
OuFrAPjXUj0t0DMw/O+e4g5Wdwc7VtXIQWlWt2wIFGf0CN4ogm7c/Og0BBjM6ISl
wMA45mf/uSWAtrpI6LIpIskEo1FZoSyGOE0FeaBMHQ/23ygDsYu1Z5315FaLkVSN
ZXtFs0ON853AcVUTY9IC61aD0MHaHERMdTuEAwclIM5tb29viCQQmwUGJEzkGE/d
1CnwCIbh128Kr7I3SmufiH6tAZtWADxY/SElr4i+8fXHKWawVM2hzQyBxxAATrgw
RLV+tD1MPQqtsK3A8Rk9yNUQf7eDu4tenrDlnzonfQ7MH2MFho4nCt49tO61mcC3
PAFfEkqaDClLnZm4jE4xYgD9yMYYZlN0LshldCcdwLyl4/3JezkOr2ADpDx1PuCN
ZLKdVkREtWehY1dS9OKwVuKSl3s9H1CCoM2aCaunaq9Jpw4g4OBVb12UgfuR3NyW
m1bwY8Ff29D/mBksVNG+yBUgaBuzD0g7MjsGHOGHnIpMpas3JqFlxob+xtx8KspQ
LWw5njfWxfUHUkCZPj2XVVzKjzirSRywx6BgQrK9h+ORpSz9CsUrK+R09VCzYZd6
8ibHSICMS3a89WtvO3+uIilfC0mt8muQY0t5WcAgmIhd9og6PSoZeZL1UR4TjI9N
/7ojLAmxP2SyaqxNUd0Qgw0EO3g5DNdO09NJVm/kNiL0BTB1Qsn+m025IJRq04wC
sLr6ACtQE1uB/IRGtn9OGU5AKtioD5IsJsOkTRB3wMpUmpM48bqlZ08EewXKd8l2
iXR5aqysAnGvkAz1L3sM92s7bgV59KSV2b4EcUkW3IuOuSHkLCvmQyymoQi9yL1+
hj5RZMjK734Y07lAwd24h/I/+aRNuuKjIygSsmjxGc4RoETzbTfr5fM2SBH/J1EZ
tiNW+whxYcSC+7KIK/cWy+9BwWGqWVRq4jMX0N4YHfnt+JEKIUSicYZqBfRX5Uxo
UrNHp43JS2BbR/6PmS4SkN9WKrX/CLOGyrlflBVSUfbbGGTjCj9bHAT9EyFXjMKW
KYvfzUUK7qmVVwUdx3cLiPmgrKfVp4L15dYKEctt+0u3gFqyv+tTxi8W4ukCQokM
Ugo54jSJHI4/WL26fsEE7x1Vwd22uhbjIxNdQAgHYHS1rzB/f5hwx1cHby/4UBSZ
dQDcQUCYUBZXKn2oU/XMxEOwTf/e6u8sCdsIsAjzd2RAoBOZYn2L9MT/SwnXny11
YgNPW5BtGeX3d+P88AQDQDqOUMPopaqmZQkFNSoK7A4IlVjyfCaVS7tm5grpXdLa
SfPfa7VXaCYc77g5h98KJWgz70jPJg6n8hSk4HnqYzLqWvrVZBm7rokAvuBPCsN+
OX9wty27HYEnEKiT4KBjFOCXN7XR0Dedj9vM4TTp2sprrhGaCSTuahw/VyEa4Tk1
vkdt7ZB7lg0HEITfUwUaaTgxYXivJZj2ZbPJPQ/1RthWSsvAXQWJpYR58aTK/IEV
XvF9yNv8g2a4KXPQC/Ksjuek+BWWM6AcvcfqI2rFpY0LJuuO7OMsQ61ecM0vfm7U
3MlG0T8DtSTTthNW8bg7Z3uFpjSE7PMzTXtiRus7O0cDFkIUz8s7zamjekzdmJj1
KKhyuz5TrFIwRDcvLn7WzkynLjtscwoG8TbauHNJGAKosgsv3B3de69hSKblSuaz
MsFZBZKy5czjo9c0yX0ZNhFh5K/luF1U4PA33dZm2s0mbnB9/gmYwZVnKJWnkSFG
Ru1hPsNAlhLdrFu8VsAYwlAwTboXqRf/3g0/aVfD4g7+Dp2XACFW25xuxgepqIZL
vmuqxgapL0AE01HKhma3LAenEgPJk2Y8zUlM+8IwcYaObKJFtVVTEHILqa/p8mNr
D8obSvhO/MlX5IRRXFE0aa7E4bALIaARP4URPLUEiQNQDn3yMS5XNKPKFbGTBnlW
/F/gpwuO3s/ybFIu+mNtXEhCmOFYDhxotPNuPDIvq5DG1U713KlkAOX+YvuLK8EY
Sa0MxYS0V1ckTj/MvhMiMc45qDFe10C8L3Pg5XaRaeOfTCJZ2Crzx1h5ix6u52km
BR8AAG0GRnqZisELfh8AgGiGYhyMeGZta2O6hj96UsfWduiTtlMs2sAq5nPfE3cm
pyLIdUsrL6/pA8+2xK2Xl3CGaprxiBRUq6hP64PkWKlG/3qwpiMrNNX+vQY8eGmU
hmXEWwwB/biAiBov48rxX8dDGgzqE7bbIngBjXrOrHLmmVeIToXxp3eBu/ZZK+AS
1bm1pUeSZLqf/dwfjirqL/9oQalKuXshtP+F87lN2UFfYFyK2eIPDOMgAFtvQ/8B
lPMsqU6gj7NS+t9/4BBSll9/F1nshBEA/FkhykgNxFCrG4WfmAycg/y1rsJlKKnv
4ahNuHbuZxI+UaG89+dubhTeB8b27x/pEbXWeDq+ZWmexY7FhO1TeaPwc3X4QGoP
P6lyRPNVcfebNLxZsGtsipZt4YykKMSguRoxnFEmKPPZeNaB4QsmOWtuSYHLk0xo
vgAgney7gtsaPQ35LTTs9Rq2WLxVTboF2RVtjeOVGLPgITfoIp5HvnwR0zY5/X2f
lR0gC27hg+Ix8JDKetCKBsHYlbWlQKL8pdwTU/3NQOZGg6+7F+KKQvdZBtStQDLL
IOSowzeGhAkvyoopo3AInaoHIzSWROWvHZcV5kdpPj8pPIr5hAEX9HEta0TcpG8N
67hP51VgRimeaG0yNDMFvYS1ml7wBov4k3iFXLYXK6o1OKhohZ8ouUrKm/wu/HE0
gALLanPI6zSksor2zaM2vfX7OrPvPSyPFUU9Vj6Ov1H4GrTSbE0NqhwFtNrzTvzS
fFj7P0aKES5aCZ+H7D5UJjKIvZ/B4UvwU8o57g+NEIhm0tAi+RQJ2ritwS5yEM/L
4hE/XmmZZfMes9ipvw9sgKfbanKDtxui+HuSuIWKrJfqTberSwnFl3fDX8JrUAzF
kFK5bCBdRSO/2tNN3qXHiuQu433EdfuNkrVe6m7/Vme+9jTUUAEZmy878I3XG+AX
r5YF1FRT0KdzOMRYylHQ8+o8pbdUK9XUi7Q1plM/arL0Z/So7lhMKUbVkb0OS/WI
K8pIavKBin9HPK03LnmqXH8bfru/JDJ0uZev0VT5O5zk0wYe/82BNUYMoJdCJkB5
2HDmQKfnaHjeTVF5s52wEV8K4IDSdMVROmFRBotgFcqLSxx0tGb8938ayBXCOAjI
+cvAr3rTSxCfXztO4wZ46XT7bUj6HGeI/Dhkpw2ZytTvCzbs4ZZ9qDvHf8HnLdKy
dqjjvzNRnfUNt47E8uro5yOnAcnuuf2L3xrIzJyYW1vVlec01mt4/PepuXFaTNQV
/cqzzfkFGkE9EiAgCCbB/pmwntZXJUACwwB0I3VF/4zn5LrTe3FNHzljhYBjqH4M
sFOpSiSHatQ8miz/6MBc2uJHP1rftd+s+fmFnWC9R7FqWFoYOSyi0+8Wq0XIu4aI
AgylBHRlWSX5QhEdjbbbTP2jAU9oQATaBu0IalLLIq1Nt/nkFTnMU+IBtRt9c4/L
VCipoCdZLW4zXA3StXySnAvRWzIgzrWdK/YpY8FQjyqsFfSKk0EY9kWurrsUGC2u
pGRek3YTm8a1W1guqJQltUzxcMaAoZSj9rXssYCsi9tv7ZQnlIz0LT2ebmxswthy
fZV6cF68AWyOAhxulBKT/rq2OFz1PN0wmnjmgvFrnxPGwZ9GCVAfeZqprMWPRSAH
JfmOx1LssmVduy1hoF1vE2YIJ4HAw9ktf+dGG/BrNCpU7I5e3c3ueSp0e5BsLHyv
yf6lwLklPuA+RWn2jCUGYCg9BxadzNhnFAMRaVvq1GJvq7gSXuuorsFfuH0WTYSF
QEVtHYIpOayefDCA+CqlkcwiTNXYxxruuFu+KsjKLbOmBhVS6dqxMJTcsIq7l/MB
6gEruhht/7aw5zZg5MkCyTcH6T6UAUuOhQOe4U5B+nbeHsowSLZklp0nJvuIjD0f
FtM3nVIpumAJ1z7joEdrfW6Lrvs3ePVpyalxAhJWEa7ngz5sn3a8IJKSQbd6FcCM
fUmE19ryvbfY7sfSlxOT9VdFeFnqcQkkjoO1MIhDVNOJz8dYnAl/m8yeQnUfeh7V
PV1ylNHUvXYJN9cfj+fpQCuP/waNqLy0heVVHBkqULlAczaQZ1le6Z7xHwovuw9H
lw3s4sf6K05fyKlqWFhfUoWqrTfBjjVWYUswxdpzu1H+m81vzLLKm1JLNeAGP7VI
FO59QbEZ8oJfheOxBjgQMnIKfl5A6WDEBO4F62zgDYwYShX6PEsnLsGHyLxL5693
1cUf9kk6FeZuBdzwTfZhq5F7HrYbWEg93Cq4oLLkiqEbI7TiS9jY5AoH0qT2o21e
YxklJTWgtSrVPgGv5d58bWBPqftEiUyam4657p3IsmElzpbRd4rvL6zehHZf21i1
kR2wYfuaYUFhPF12/WX8mz6rpfXaP5UOEeTVRh0ay+WvgDFLi885FVY0QSW17FDJ
IymMNL2ZZQRPVqBEO9glYyHyvr/k5ety69JwmRXAUxjtBhb163osMGsq0TVdtR+2
+Yg0s6exPaLd5YBzHF3HEqfGhrU14E+EWdOHXV1asQRwzkYoMmIgL4d/JtoMaSnk
7uEVDNZczhVUHaKzodtKMWNDB77nSuHcSR20fS1j5uC36aMnC7P1LEkPXutBpIi3
lnv1XqT/K2m+tCW98Q+PS/r/yz8roz11Scm49rjROivGamdWfEMvw7YPFo4JHpaU
DWLez82/2J/tU0bYg1OGBKzwbSGztOblYaBojw9HhSlvOOc1p7jqj8fBhNWmv8Ew
Q4+vh9KJuv2jJAfMfm4IfTC8H+pePB966EVahi7PS/5fSsdMYCpYQIenIZtxYbLx
rkVmfb8dQ8/uHMKfdfx4GwPE8Wh2iOW5hJjr/eR/mwcTAbgvlqpHcHLEDD1fTmfc
CGZyvoK5GshQPJ0tG4SlHEjM8cRDuvZIfN+eH+QvDA99gkI1Vkbe5gXdws6cLtmz
xRG9wQ5Ht7NdnSkErjBFOau2ojBuJgZ33PjQACu1zTDQAsiqViGUKDD/1kpry6XI
jVsUNy5BRi2WXJtDCbu1VDXisN97KZ7Mj8urtwHQoYttOAB1hRUlTL9ES3TTq9xq
TZeF86ClDIvBcQcy1hHQgkreFv7XUf01MRZVjUBxdOFlR+a7RxyC7Sh3mRFXwgAb
msrziR6L1aJbZpNAx4e/I0pLcaRVpXJG4QL0QoXOLUyqrdtnlsEF7lxfJScvr2K1
njA7mVrn0ubFKBz4HfeCATOfOHTdpuDA5PxT8Fv8jhx797+zANtQLIK/7GURf2sy
ujGT8KjvgBvnx26s0Esi9VQm1N/LiOFmWEHUx+eEndBgc1pcUeD/5H8mVSO5g+wV
7ay0Jj3rOluEHNwFW4zmzXMF9FX3/YdsRHW8O21GO6voUwG4QBmv9RT95bYTvOWs
TivBsaMRoJym3OfzTQ6JRuJI/R1Z+Hz0cEeo/sCcDTIHwXDJG32vv7DBEkhbn+B4
+EcVwDgPkLaBAR2wFwCLxiJSL4XJRoMuoD/995hwFdfAHK49+gCT/RaJi6Y/1qSB
kPM2qUtwm105oO+wV7y6ct4Rup6EhP09oaiqzMaLFJOQ6eOnkBlQgiAXJLfa/xYE
uciTu5MqKONLea6nfc5uwQ0DQaPseVD21ikYt/4L5llaLEwx9jOIJrisR6PDJ0SS
YCKCKtWvSVH8n0/mqts5/C1eEQgAiu0tob5yu2WzYAhfoTsZXQtu8zdoeuL3RUdO
Gy0wtF3Y6Trrhe1KT/NJp/jYIow4bGGdTz+R0/aY4NJ6bc13kcO3nXFD30NbW1Yq
1KoycrS49YRUgRYFwFfXvfOEzZxvbx5nbJ1i4S0Guqw5bNDfmI926Xa3BtI3hhQ1
55DdBpBY7HVtCTSGbJrwNibCB8KmkQtMxH5pIV0QCHKEp5VVBRAg3BhVIH7rG15v
hhY/ZwJ0XqCjDfM5bgAFmETdTeYU1JmVc4n6L6wRyjXiz30tsKfkbGpDsw0l5SeP
8R2+nCYGvyBbqQvDhJnLYPxbUTnx+P5hLEGeNt9E/EdZ4MYYNTCU35xpceOu4Z2p
1GnOHdtznSV7tdkRpwGG2U7nf6H58mCmz0meUl1dbAeGXHxDsL67HB2IpktH3civ
1uxgSchuPe+qvdZ9ezJXAk9bnKTlgzgGCewROzPm9pcPw/38wKD88BpHGl7AuEym
cWIQMws5KB1B28OSUxhRJXF142ndvn2FWY2Pfhr71imzG1oAre7Z3NDLIZn+5lzH
zLyeqt1nnZnMDSwzN+lcZgLhKy+N7QU7+gedtxXvpoC/s/ThpZr7NYL3kv6S17y/
9kd1JrjOhkwrEvsZcM4zWsV+aO0ieF1f6xnoBu9BGa1BAQrbo2lquXaF5ACyfqee
KGg0ApUpUnaCWTPe8tTJcI/QlgsVhRNFHaXVuRrVU5IxdxYQH3XDqUHSaOLc0dP8
q7RBSPfibzSP/N8Sljc7vQGH/ZYIIcF3V+YtqtYBs5RYDalTBlCGvaBv9BV4JJsa
8/FOGfVc3giM5L4siDOZoNT/7jUnrRJd3YJ3NLGlvbm7AuSBZZkrLlHQhbGkuzHv
ejuNaivRMDjZJkgRGLqDD/Fsq1moTxg+xYKPa57d+3UxWo0M7Wo5wT32OMf+hhCU
uTS2prU2kf+AucFSVWStwDYHsVlA0TH+vmCgmeh1uopDg7uWx31S1YjBs7UenvAK
aTfWOGPCk/9P0x45CenF7yhxWCx1mfunu9yHDAaAnH+/bqyyFTLusrxSgjaPoMq5
0U0lwbZQcKcYiUNNA+Y3H77Pa+eEzxPWLgtYRPM71oVAaXvoDqzjAu1Ju3iVpoCN
5NhyG6fUm6jOz8RBQTRTt8yAuNgXfsLZ0eds+/8Y5eZuaKwJYFb7DjRHNNOOR2We
ME2XO2wb6bd3DRjTulN7b5mi1SnaUmAHJMGJWHEYb26iGj56Cu0gdwgUK79RaT0z
Cecx8zGKx/NBOR+3tAIoxt3jSHe4WIFgl6wKYpzasqrcYAqbelPpcmFYwE7+anf+
8Vt9nz3wikkZhmK64ikxmnFjkB3Py3rL7f8SDlD+WxStixaXEYX6YfHJjaHEzIPF
KvHT/br88jAI/eJRasqdKpHSTpPln98AG677s1A3fNOBWXLiP0ScDRZH54BD6cip
kYdqoMlS1Q6g1fD1MrRstRfWGn6+ZfLzZ4tcebA2dScPw/VrSw3VQHwhOHoZQetd
nmy2gwpdoA/eGgx4cxPJSheYPcqhfWgwRvP1TBbwh7J1wU60+ByDOfae0Qq+QKPU
9LCCNBRlJj0pqQ7s8nv+NWSzqQCAXspHLkNQ9nQyBNwiGNpW+izyUxE3kCZNyY11
NcRp05BZH/85YCOFnEZQmuIDAFDQGspoWF299auflHaHiz1Bd+Uz0WGA60ux5Bo7
JXaoiYH5VESFxL2FaKxqB11JBpgulKSGGRxhPEd9ohe0d4yG8Pajvl9mtKGUUWAN
LNwvwAW4lXSPynKuTek2duZ4nXSQW/zNPvENCX1rQEwWTn9bkcpRgykc7mDMQOOG
2BEprgWmzJCwQ/LjeIFUMpeN8c/7pOPORvT6UrHZ82QP18aVGuz5aJ44BfZAsrJL
xEtF7OjhkPghlAt3AKf2iNq0aqNW3G3gmLkwg6rGj45xZ6LLFxJPWqC7IniCD7bq
Lsn7HIkAt+O3xfRos4btkuBad9xJ5lAIrB5gxATzp9xtnQfyF4QRup51dLHbaGU/
MPHXwjprgr0CRNseFnhPI50fnQMBkngCT8Qp05j3Jj50Debb+qDjGfZ6BV63D5BL
o5A1aTTva+L+AupaHlukvCpMrKfFjwgDrETkitliChl4POZEGVxOiJI8hTHvrc4J
p5P3m3ve71JTSytM8BaobjPhhJtZVRajnIUPMATg70z1AB0Evwb4Q97NZaRyYDDJ
0eq/d08YodeDiog8edxtekKE1+9z4iUX9VBn1QqHp0OlxeydBYD2hs403vJLP3bc
0JkfHt/Kl0SIXtCC8ge5j4ItqmoffxVmtngUvAwqBAvMiGxqNJE26KvYVizhCiFJ
75Wvkzusv2LyAK2bRgcv3Nf4HupiEyD/DuKgYKoAs/QmIayyf4hdr2KBrgIvnodi
QRDeKITCxFkg7uWt+r15xLW4RN6S/lZUuSjNqDxYQZkPmyYJ4fDreYw6zzz6MZ7W
6R4ScTN6yYB88XGWULmwk2A7sbfdSfg7ACizPETNVzqbMTacq/awtzKAlVMwmBzc
+wSzgVgzYOnI7hZ2bvOJHM9JmcdlZu17wZ3InM6SD3DOO9GukPOxwldHPA6yT2Yd
G4+2KcYojHiN1VOoo9u/rbKGsxymUWsbxNwvedyc+b7C198Y2HRsKsqBbLa+qSSi
Ubv02VV9W9Ck54kkEtKQ3RROsWg6t4L4oV7UpQ5kU+IlBKh+HowcXSsGCwr2V1Yu
j5ASl8YlAnqnhgNhKUW9gXGpj7d96K3aAwEG2/8lVDbkrYoEZ+FytlC3OQybzXP3
R2WEK+f+C/VxQkScH53gaei83c/Hpsj/q9oVtryseKeXUKXmhktyO0LYnM5DY5QG
RkBzgDsY6monmPViXXDZ9PIvU0+i11iCTPtLE9I2yNc1EFzO/vyGWNhAf4YNHFc2
pTYH/V5a9skdxLRSjP+1gA3JwlIns9LMmyWmpYfaxr92j4kT6uslsiXQtVOJPAEc
iXMeo2uHxq9L4ru9nbThNqBhzk6yxqrtasEHs7LcwZ7VoRT2x3Z9lgumqJCJndiq
sltzKfn/f9/iXaRP2DE8byjA0ASEUenmBSiA+v1DgCqC1KG4B61CJW599jlY7XJi
6b/yKn0vnafE3U1bs1gYgLsxjIysn5pxvKMTh4Y2bonblk9lXUSDKhYcfQD4kO6w
oZAQlNlfIjFFeGfN/QkeCJsIoB1D+QE3eLUC+gS4k3hFUu1Vv5+9VSmbfIWh7J7T
Hj3OMf60fw0mpmPG6j07Sm7Nuj6UBVcjmQ9e5kinUNRA0yQzRM32NRWaXVWboQ/Q
5FNf8D9Uth1mx+71VRPrlG7MOGa+SU5Tnj3t/yjM361zLuuwiroluIJisWi4UYTm
bwqHTWbWoHtE8Zq6rLYdlBWfcTDZLK7rC3sSTSMPLlUsSFb0r4gvv8J0UrDA/0Uj
h528rc0ta7KuBYDfGrbU5IJXpyASlaSTTMTIHl5pe6OFcvQ/bKs2Fb0uPu1JpgdE
Q4rgDZQ7tbWPPfvQWAcKYj2Ks3Z/wXaZuMakRMfcY3pJFAaqGpiHtWOu4SPwYjDr
UcGSHiq52kX1IUMw+8jCis+lwk6VLfupiyhvjwPqcX5Q0WGXzNLq8XTKd1pXZTy/
ClQIVRHL12GuCzwPvr+Np0TJEAPe73kXuP30zFWvyHZKy+fTQSGzPRNF/uXf4oYc
QJW8wjRvN7ClwHvgbyIzoZctBljLNaPYfWhiI/l92j0BIo1SuXATivqscv7sf1v7
CkstwfcMM/Jbyk4ncRMPQ/x3EhL8bA74B+002VGlfvEIQhDmrJFFbqOGL/ZM7oOx
b4bnwCR2quJ/1J/3Fk1um6gTnKgocbpwGZ7ObkHn6KCoK5wUA0zGpIN+5InGaIaQ
WqTBAmqWgeyZwV2En9v61BcJQljTXKA0kWY55ukgG0RGoeMKkciOrwxAoPkE/9Ou
uPiDYryjeOvpWHzNMxcl4CWm/WIgs1pRzCUQuBhPljClU+1Icdwzx9a1erbtxHoG
0sJej7BEjE09esD/nzefHRjdzQMkQq8XCAUew8OnbsFO560yzZf86ko2alNgk0WT
xZCg1Z3oVeGdPSStSJylhfCOnPN+0JqnfDuCMx0oESEFIhQCqAYEa+U8Jw1jQ3j6
ykUf7DG1lAmpIs73rwcFsgHm+pwexRN3OaEzHXyP9y6JQ6BTrb935xK4falB21Tv
3TodJrgN+fWSeINoEG7S0iwAl6aistMH58Fk3ISZW37EV+rZvZUCs2WWEeRA6Whd
0LofO4XTYMBwZdJIqvBifmeoMV4vpQ5pML3fMoup4uzrHuzhqTtiTJ5XV15SgsBv
/1p0xmM+ZvfUmWvxkiRgmgBk6fQ+jnDndAHuwbu6IbpfR58JKvueDBlfkwnFixR7
kscXsMkjNaX3XbwB3BkU1vq0lsUghlBIrqExh7uY0KWwGZhy9tIOj2SOXPoHnWF/
YGsMMqew6U9F9LATE84Vf387g6mYrVF2BKrrpML6eAyr5mP9KaMQTDJ6W+uYzY4a
mvNkL/o2yTUXNOeT2igUWC586JsZhBIIhhgQ2pjwwXzHhDZKDGtiQzyDopn+63zj
zOwXIVlBIqxoyEFB/rq2POfCnwdPc+KeOhgGUf6VlSMaDFuVmcTFcXkmi0drvByp
NS4JCEJlFjQbM8UXdl1ol2RWDqRBCuAmu8gzXvRjSvEzwX/mMIDM+4jebjW+/8kn
aAIPEDQy/Z92y6Cu2RIcQy2eqER4kB94hLvP2WoNybzyqyHVgMSsetw/dPEJxHH5
TnBKzU5a5oUGsj6JZw9SJb+f/W3IUnTcmpDJRW8Y4l1txKsChFMRPKAIXEu+Cm3n
LJ8GJXDB6a1OCgPfzwddj23zJI+1aLrFuM31jWfEhGT5I/LhJFSMZE9SDA4GLQwP
JbRM9L1ygMbw1J1kik6A8eCHugbO/ZhvCiZpNJwY0Zqc38cMF8RX82+GNebVX0+3
ifq0cQweOeMhyngrN+wuXq40TCml5W8medsohHnYDv9Kl95XE0SBDAttE8P1o8Uh
gYRqvzwAbQaINI29P3eupAJhzWxBieSGM3k39dnde2zdVaiI1Wcq/1dTLl3kb9dg
Mrk6jWCLfZT0gW1NOzhobZVtjwiQhDU7LD4mezEBKZctt6V6GeG4dtYAKIoNZWgK
t6He3gOOGCMPQpHBLNlR7W3qmPHwbfy/T1PxLy++vjXwlwuMe6nT1TTaqV/ou1jQ
rC2MavTSGMSJGyy58x+81TERPsGXAfeLPqpeAoLkKr7m/VaBAqyw/7eKHkxGtQr6
gON11zL06Hnr9fAm0jgVW5qz2vtFloi9nWspCsMvGK+Cs+wlmR/0phcoa8FzeatW
1UAcKYeZw6AOiRIoq/18mh2+VGpkouFPLOlYhK7mB4pbWmFbRY8TiOSykgTRAhIW
gH4Ydnd51UzDdCNPNWHpyozXANfJ0i0yQmxCEXfXUcqexZ3l7gkQHt0K+pHy4hmL
zUv3uXcYYnZ8vHffBs+FRhOK0RwtAVZ756aqEQUDwneCrG2JXv60tTuU40TAYwFf
dahB2ikQ7u4HzVZEYRKAfOU0TRP8sM3I4ir5e7uS8tM6tNSU/AtnAo6ZGzWKbJ/Y
5YYGcxE9M9497Wq/Z+i1DkeCa2oZzympRqilDaNlJsZC+fEd6bfsvfcHKNpI2mpY
muW7C6i3ojoQ3fVfIIPOjCy1DmHbXZheooLLZPxL0hxWAwq06EiUNNrzJx+arQsG
bRFMs8n0uCZGpfZHgGavtlPYD8dnGGR06fSrHHEo3FJyxSoWREiHf4kXD1EBz9WP
yu5T2Vv8g6HP1d0oDWdb3tWolNQW3h0Uos0nK0oDL+w44XqNWKvvEolcCRkAsoLF
en2tS4MF9UirZnpGOea3cGInxzC9mQUO7cEWjFKjWi2F81V+YKfQINig2QBgYG8V
8Om+GI8pACuj5xsQZ/j55Buak0o8injCSjCJn29rcFPEsDXsg/5IRqTwR002BuVn
rmc6dmWsV1iiJZtEicnbRxhAEzmRAFqdWy+XF4aNhvyFzlu6UDb9gZSUg6FtvqYL
UUNJEkcsh8XPzq0U70elNuyql0AwCIusF806yilY32FdPmA8k+97aAbBDL1wxrkt
9nX2ghsPQ7vxyTer5vSCwqFLbVXsMDZLBLGy8lTUsRgCCSzappbgusJMsR/MVafG
uDjs+IREPNIj3o9wvs4AOHPl6NpApjFWG2d3TyrOyxnWKGtuEOzXy1/jUNpZ0w+3
/xiAAxlfZ2wlQTTaBh2ObIViyIoeqU4bSLDlTZQ6woEIcLAGLzT2Cqw6XKT8GGSz
Jl9jBSrlC02JZB8KF59tlu8JtLz/wF33POlcWie9p9C1bbUDT6gdph0thN7EUV1i
NSzKDztKa0UzHejzfy+GxZeS2xccVhAhHZOPsWA0G2Tzs+OpqgGVIKRLo9GhqyUP
mHV4JePWFNJhAUvxCbNqq1izxkuaIvBhkfJEo3FzxXXnRoQ4RI8rEAdW88uZDVHl
eKorioxMOu/Up6zYuWJFfwCP5/5qwqBDDSz0eojiUrS+6hnSUhAltpzHE7qT9163
/DBbjG5GJ8ZF90F01dsR8fPUhOwNdEN9PkrPEr5Q2Le0D3FXLfD7OcDA+NfdJ8ac
N0h9r5XmOZUOJw/O0ACGWLGn0BReOoft4p6Op02q9tWbP30wX5BbMCGK9RoTiu6z
sniJE7jBSNk0QyL9job8K4r27quMoGh29+QTXrbtct03+NutIrpyW2dBr+5iuiPQ
d21BAvsXsFEsJrIfmTVG6a3A11V3FmUcQX7iUTIAQBb9gsUx39YF+CBRfaNvCFgV
Tj6vHP/xFKPAtYYn1tmE4bLffnnAVV0LfXWIjyTFbX6Kv3bgWxJJI5ddgWeWQqh3
KrHf+D326unM9b+kc0ELBiyDdYQySAsFqNoJMGsusv0S41sGiBGqTwTO1ODYStn1
HWjRnmSbTet7zKo6Pynqwk4q5XycfylploQP2LdqKqUcr3JTWnlbhZQlJbXhZKFq
S2oIo+5TZtFKkPQAvY+uE/gCpKLPvp32iNkQWfrZYV5BUa6IlWRZNh77ZZXTeoeg
nmldmQQpb2OGizbVm9eRtRSX45HLJ5eEdNYSeT8/+Ine67LNw7W//GpXh1f7AFii
KF0i/XlQeIpVCE6Z+ZKZKYZsJJJg3IIreyfP750B/i1tvNeyPy0pM43bphPY51nB
fPkMMPHs8OsEIlWXEvDxL6wwYHwed1bovQLSUCR3+wcYYVvJkyiNlLSagix3CV/m
rtnR+n43jMCDCrgMmXfmPAGzpEH8dG/pA3iVOcCYRYvUAOIW9fHaNRtfGPwXQ/Pp
tqv7FQubQmIfPo5XXNuYJvx9JLhJkvTyAZfMrPmNICBHFZUxIAGuYZnm7VtkO6YO
4LYesudbjRqmhAapN6vlIcGIsNtecDMiEvcS859Ygql4cmxIP4DLTOnDzpSip0Zv
yeIaq+Mzscqk+SNqzaElLkc68A6bvDspQa/ydy7z/k3J1v3x64bFudeSuA4BXjPS
aBWbjjD55Og0dzriY4PJ8aZX2uHqRBkC5vy/yNkinIf7XvATs4eefO4sudQ+wkWQ
9jB6iZ6jNH63GBHN3Qq17dwjw21et60P5QcrMoQs3QxVIsxysvLMcaYbcQ5JnXxs
Wh3MPrKpjXEpmFhQJNab53c961ASu3uO1tLxVwF9CE7fvJhpai6fm0EoguO/OvFY
DTxApTFAy+k44/+TAAOk0ueyToMY2OoVmxtv5A1MzqnueKuS2eWpvGaY9NBu76yj
AlMm0YkyTGMWrBk0Zy/rr8bWSr2Lp1/I+1ECr06x89TPh+9AztVw16H94g4UfMjX
jKIf5nHI2GOkDfMl/H+h7JN9CqveL5noryNlz1FvVn22gYA9eYKM4gb9/ikuzDnb
oI5LEmRTWMg6ClptCROOBO65r7TsoAxcGjg4HkjOGh0z3czvAhgRVRQX9Y5sQNrs
wOkitZgDLvC3Zx28oW/YlifMCiD/IUibk6oxZD8Xj8uul6lDP2MyoXyoUm3oD1YU
ICCB8dEkhJBKjYI3Nxj5UlsslAsFYRI65WQpQdpFv5ICAXholsosIEIHElKg5RO8
AOXHNftJrxntAFdraD6mAxxbDHdVgWbZ6E3VXtzPf2PSNaqE5tgJo6qL7E07tPpw
G2mCkPwLwerhB+aNZSDMokvsAyddKiiIVSXJ7XE0O7arc/jGlS9gAUQPlohCMu/j
CaS5JSfdjEhvVKTI7upsGhoF76VJGk70x+p5uxljVcKSsSa2vVthqERckSTqU8z6
g5nnvEkQYTHMRV2BFvi1gS6cTDI4oZtKi3beOJlXuuIjm+6LYLO++gChEkS7EAq9
Wq1jpLlYUZRlF/1x6RWZrGU/oagpuQoolqpjFmGq024zEd+DsiklYbrNbtj6qW0y
SKuzCU6OSrZtbAr93kMWTbIIFeynoPaLdV6G15scpwtIIhCGtVsSgJIRu1z0NJSw
6s8Hzm3xhIcoM+BlXm09vV0P1E2Eq1cmJxuaGY9iTuoCMC22TICrHN89YIm8xQ4q
uvfl/cPGbYaYFVWqkd5tVGDGOVxs3RJ3570Zoa3VL062iJHIN6nzEA6IlBoSDhdZ
w7X7KAgqEcT2IkmICJohmoC4cb8vz6QYJhS8n5wi8ihmQcMmtghW4+507FXu+q2B
N3KwYI1AwYCuH2fBxGxiy6VIWKMj5qkE98EaJGIi2KQ01/2lrMyAZEdAndtc6nTo
NIAD1skGMivUmVFeRWVxVuViyvohMpZn/qNf7cIToStdqebnK1pF8eRhi0aVfqH+
CYICUZsZOnWb0x30JiU5wPAgbSC7TKI8neOfFBvvnAUPBSZ+641+IgbHth7xzKPR
i+dDM9+jBstM70wuCnQY61lDVyiKgAub0AGbI/LOWmvUjxkCwzOzplQ9BHWUCIIg
BuwDP5D5fRaJB2v/7Hfg4wTx10OjU3ZPZ4LJlwBxAai9LksUl/d0RfYmN0lqoaZw
cGqUa5kdzqLzo5Fm0Z6loTDl2CqPer95Xn+45iIYKiknG1kL4mvP0JbyNS9GrOgr
W8SGE/n9Xnix09RiNDAERJq7UaNf2Xm+p65KacEw4AjmbLBGEQfWBs+LXSXZRYSU
Bg3143wQsewpTNdOca/2VHWfxEw/P/ZBgScIxj7P/f7N9EM1FqkymwJbRWElcuro
p6A08C7cqFDkSlH8AA1qnMTxEdC2yHLRnq4Uw+zPsA3PIBrqSEJDSMV8T+MZowff
OC63vplrUZ343KpqfYxzmLGEOuKRSE8/Rq4frVm1wAo4OcoOTl570A3VPiS0F5yY
rZ3mWxo8VG1KFder/9ssal7b/Qv4K1DpLNOf5plWykyqT+flz9OwpOLMQsWB9vfx
Hsy7qWaxXn3AGGoMbJfd0u/ZJrTpukwkR7FHRnYE6c6AsCn3axPohz5idRskB0rv
iOf2keATMSFzrD27wkAQtogMGVPjy7rbfUrNAip1EfDaxMOrF/J8k8YK2YDOjZnC
/EhnBYWJW4YRqASqdH/J74LqdapjNvAaznhJTxQxP6U=
`pragma protect end_protected
