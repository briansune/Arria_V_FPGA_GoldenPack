��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t�n��M���/��6����k��,�!(�X4!둮�4Aj�~��<5ݪ8��,��/ĺ���� ;g\�
���.14�`��R����<�p���KdW�K�q���9���0d�:�� �u����'��q�'�]$1��	��Kr�I���2Q]ŗ�L��wYe���1�Gx�g*�F�	���2^�]��.�X�_�)X���Y�9�f�!z�B�q�9�{�8�uĎ�Wё���;9���է���
WTi����/��4��X�[i�~��e��+�	B��Х�<�����A��D���?�G�a����U��~��ׯ��)x�֟��6��m�M��2�|�T��y��&"z��u�hÅ5�xm9M8�p��~~�1-�f�,f� ���cT�WM!��	i�z,Z}��.����]��q��#w�ǡ��`1L#kI���I��5rۦ���G�`j�a�T��3z@}�]s. �?� ���=�L��y��5���T��U����7.�2�����,�88o���%�t�6�-j�q��C��:��F�+&~4C&cP`�E�OY*������j	RAf�A�$�z�3�>`j����Rz����$)�E�$���v�l�`/�]�@�U�xr�eT �̋wJ�Y�������)�d�CP�%D4���|A�b�Ú�I����� �̌�d�4�zb��Q��<�7�EO��{$l�[�KB_h�NK�n��_y*�F��73l��$!�w�>;,k˥��4����.�r�?dtiXT�����{2��Q��Mb�`%HYx�Aj�ٲ���8tg��G�ꕃxR���˵�l�m���q�o��J�GQ��j����E�T����� 6�_B�\1X�̵�L�Ql(��-���9�r���)����`%��t��[$�¬��N���ۑ�nP_��z��ӆ*d�8ڪX���#���@Ē�U�/��e���F��t�0�x����#��D*�؏)�x?�B�{��irA�Ȅ�A�+��y]x��	ё��`�g��j"=�qJ�;HFa�z��ɂU]����1�=��~\p����)�%j�ɒ�Z@k�2�٩���q�.�>ً6cߦ?,���8���H�\����c�ک�須��|�j��b	[p�+��:�:ZO��������N��y2��,��H�����?C�]ߐ��-ef������Q�����:*����/ɝ9���glN�6iN���>7��/����T�>�6��1�n�A=��������e����u;bOw1���P4_T�*�m�%����Lia�hC�-1�t�<�U�r���4m�Vd��2uڊft`�����������K'�G�mwX���k���C�����8�w�tG8r�}��N@XO�/ZӁy��*'P�U�q钪{����ɣ�k�o-b{�tt��"F�u���!4���	�����{@������)�d-�3��c`nb��^�X�8CI���Bv>+�1ny�#q��\h{ �Q8'iO�$t�6�Q�q�$�fX�'�َ��w�_��;��UT�~J�bRR�gUm�T�t thH���9:z�s7t^*��a��ޠ�����d��s�*��)a�0<�W�7�Y^n9+{L�^���o�����ĺ�| ��F5@w�E�������˪���N��a�D:l��<�d(��L?�z�@t�?]A jp-�,������.�����!��<`p���t/�'�dq9��x�|�]'����%�"�x�I�> =Eު1����'����Â��x��6���-G+6��_9�I?��K���A����˚�ڂ���d
����If��̀�_`D�����Ȕ��i���g9Á;�m,�M�P�@�`��N�ۺK=��SP�gƌ��͐���m��n����ˡ��jM�	枨��b�� wj�n�K� �x�եl�3U�X_	I5���)y,K-�B� ��I��m�u+�p�P�\�� 6�����I����Q�oe���x�R�V5�hQ�4!�c�;��{�65�j�c/�wsV�>���b�RԞ�s�@< �^S��pi�.0���0�(����fc��Đ�u�}�H�͝n� �]:ve���m"t$�t���n��g��_��,Q��K7ˣ�~�6O�3Y\�W����;���w����s�<br}:J��V��H��0E��FY'��&��LX���m���*=1'�d�rV�M�8�5>%��>�h��Q�Lj���d�b�OT&�4�!�,f��U6�7j������0�=����g���lsG��H �T������۞�1A�N6J�p�'���YO�TV�b=Kp9 h~��ZZ�	X�$�|@͠�R1{�"�=�����E��؞R{׶��=~���^�5�m��뷜K���s��B�By���^Y�����^g*��d�������p��ͱ�O�ۿ/j�m��4�bO8���nF��_�&$�]���b�$oت�at��킕ƨO�@�T����'�6�N�r�7@Bq�-�I��'�SR+z�/�\��k��q!��K18��&��I΀(�^��4����ߜ�c��H\�=14�͚$�@�/��m9���%��8/9��#���Q!�:�;s�w����n���}8VC�@�F}�o.���I�u�$]����K��W��Q��l�N=��*�v4t��Y;!�����J��G����4�(�������r犏���C)�ҳ�@U��"]�Ge��B���^��NcѦ �ؙ���~��Ԑ��R��e�٥0�T~���4�P>�&q_;
��{�(�bʇ7#l�#i����r�9�u��'I�b�ޡ�;�j)�H���,�p�<����}�懼��2W��"v�[�� ���lL^ce��t�Ũ�hh^�u2{<�m2;�P������oA����)�#VX��l3���/(_��c�^'N�����Z������T�!���qp����`�ź�