// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:28:04 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vvsvv6UCGNRndL6yf7L21DN/sdFnlLbBySPvSr6yLcvTWCcMg0qqNdimc3BkgMKY
LUoiYs0r0cXhOzKmfgXaloWngl0NkL5MU+BbPW8UD6iL0PgsDagENeTWlaA8GPfj
QB53bJ99Rr1jtHohAUxc8faV5nhisoegyUthvPGpv3M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4544)
8lEDEZX3ejCEQHR/weGNZG9xEMtcigY1E9kUBk29o1T8go1FpXkLfmGG3rtfafNP
0GyF+cPdy0OZDAwOg19yNg6mRJ8Zl+01OS74kL9V2a7nKbs8WWG7441u7prWCGr8
3sY9JOVChnQxCQJ/hL5vr3j9QnovZJ7VGOv0aed2Gclk5lop8a18y7KShzFikgYh
5IETxChwN+lDxe+1WtqMoVoH3w3G972r9bqd9vgmG/Ho942qS5qBluvfnDgHHMvS
vUlgHj4brNeDKN5hbmKp2NGeA9a0yv9ESjaNS9wT2qEzgl00fzj0TyXOB7Miy5Y+
Y6bULOIV6czmDRMRWsoObUPa455ngMiErsnqlLPojSog9S+Dvw0hHbrzh69Q/wdn
gHMuhJUe4Shc3VgM1B/OrCZ1Ehli19xWA3kp5Wb1oZ8faicYylGNl+GLZHg4YwPm
6WCxqobv80Y8aFNMorPuYnmeMxwT1P8VT4jVPZMg/Lph9Z3+MQ63GYPreoWygnqn
xiVTbtvtF9Dkm47iwFQMz/wwqGgixH/p4vNh2k+1kbOmHghjbUuHgRAwSFSgHIEP
Br9QqPyluVGA16hZkxLXN3hy+qVDIRdabLXzHZdFyA/r2UG7MmV+LqFQNP0E5T3V
3C1yAngaTpcmfek/z96QiJ0DD2tx7yMB08eHjE7lhYP3ZrHd9hLnXfdBTX6+TuDN
IpqxqKSQXtKFA7Koknk3EDZ3Pi/tMqAfSaiIgN09/rDbLeUUeChocYSXUwlG9Ntn
I4t1YY4bHXsyZ8HmVDAOviWLhFxjW/oIwGzsvH5DwIxuHVUP/KvQ09CqgpPHkCfl
EmwuDVFtEiAXsl0UGl7v9Oz0Sck5Vp+4C7Oab0prlI7j3XMO9mbkvTc7NCs/v3YW
c0+6/OX6YbhLnJltFj3NmTzoXreoFi4J0latKN2LyfTXr/4ZnY+Wbm+WKR78QIMj
enpjiGLl8alu9AesX6aiKToHgJiPLYvGzAaTY5yQ2f73kgo4/IeOKmQu+99n6h6L
bNqAviB0nyo3Q+eTrDUaviQmaimpOdiTzpPRTujpv7uWv4WgqksMRELgk/d2JDq3
oF4iK1JZ2CNXe/TFXXNvWAMW26Ds1mBqBG/RsgocTCeti24s2Thk4EBprfZ3eGr3
E8YCYx96a4bLn1Bki7fQ4YJdgCLH2X8Pv5thwSpxFodsHi2JPmqLMVVtKnDqpRH0
VRAQjcR2DAw3MeuUSEUSP0xbUe0wbONQFuBAK+67XxMdq0HYmH6sroNgGcdyIy9B
PFby3SyuZwEGDwVa1CSWptQuqi6d5kmCcbKZ1v6067xX3473WXiGpUwATyttzTA1
cz5OiSPkCgFK5XKmFjafr4KogkhIgDalGv1cyHVUlDYUAljo8TnQFtRs4ufBYcq3
TSdgLY1Ezqy/0e61SMANpsXVBaonztllLR4zBytESBaPNI/3O8TbpmqdWilVkbAW
eTISyG83uc/Bfv1xHMaqApgBp1CVmp2TpjIJwx+22hcus8BsgyXqmbl1j/mQZqrd
g9Krv5lQ3YZNtoFk6Hu6pBf3/g7eD+HbX+GbnJSVHbb/Ry36/2ouZO4K6umAT9TK
bWMi3jVl5gUiYra7Mg2pecrmkxVoo64mfKUA6CYEEEU8a39fzWMrPTA7xdb5MaYx
y2Tgi1zpY9FTZrJMmaGfKS3zXCLOnhEYnepXnnvVbyKqhWonhpu+UQzQ5EtIA8MG
cQeH/t6ien5uvTZXlXcoZZegWNyJPM1AVv2/2+Wva550Vp6mmd2VAE6ob7xV5V5R
/rq6v8Y3xFOGng7pbCGZTRZFlcilwBa2YtLW5MKZWgr8lfdryM1R0eJ89JMGhO7R
U6+KWSUWLqJWiuHEIkmLjqyGJszb4+W/Vti0o0wLvNESsoe+SbehwC9px8j1AuuY
gCdUyXMnaC4+nXn9c1TVvEPcOSH9XejFBy7DAqpVSegGWMWfLSOFJV5gXGL0qdys
gky+EXedvJq94OidrvryT4cPHWlY4JPTzT/FYv6/zkax00H0TsTnjGHBBZYe8Grn
wI61XT9mU10krVRAY90Hx1mmgAJ3Xe8cXscHI9KsWT2VsNC8tqBPRMPtFO6+8B5D
VS+podtbM3nV7hU3eb3jWGoXVIxb318GjlO7iYP9ZwtQkBRrgpOXaTYaMalj6qCG
ucImnQQd0s/AvSelqsyZoydOQ4/9sWuNlonXIM919hb08CkJewxTaVaZfEvSj7Tb
0+fXFCywo2bDQ4Zr2ZuWSzIM3Mr3nJBZx15dWyujAfMPR7DCjK8/dmtXKYezJH37
pZWSSDOjjhuhQYChLGxBdVYh+P1R2/S1MW69+Jq5SC253YJgrLaOshOzkzYQIIwE
MC7Gdcs/UzJ4aELGUKjYi3jVOc23279f56B+i4SVYpB/yztQXgvwCUzrbV9kxuDQ
DrgLBwajN7QfilFO5D438oNoavPgdE/X1vi5mbHaSAnHOdZKNPhbPX1t3IbL1OfS
wukCBXLsU2eu+cmjLxL5v2VPMTcqBg1ByCkZ/1zhM1mjYDy3FvEZI7w2J5FRE2/t
X/lchW3rQplw8Wlkddhad0ePE/D81rxgg/NamJMVb3wQswCEVivnCfmqgffMi5Q1
7CcNiyEjJgspxjROUKcaYZtJTXdYSjLeEAT/JQEy2Tus0yDCe3XJWKKX82CWGjIJ
fMp0JHXMx0UqAHrx2Oxq0AJ6b9V0nziQtlsYf1v5/6tp64tS+Sc69r10cz+16VAB
57QyBCUwpeg8uN2n9ggCePlSw40aSlFWr6m/TOaOrayhyiqJj2vL5K+zWuhCMlD5
7RgxdvioukgFxRGRjIR6pzC3eRgZPx0qz0cayi6BYzy9WZLRYDORKGP/qTSkrqf5
gx4hG/1QZFP3llgfWjk3+2NMxiUfhKTpFpW0rirpFlVLG8Y6rMjHk8GKXnCiiRGv
eetldq8mrybNe5EfYMNyMF5+o9PapFEWGLPd4OxvRKKAk8QCJ0HdRkb8DJUCKIgY
3xrxGOTEj6dw4+Ger4q4AnMbClKsT1L4ppMSBEpLTNWZ/6yvNGJQzpDisvX6b+am
nJTqFQppxkOJ15LBBc6p6f6F/LCym0HFmyqCceICfo/O9ERx/DPdLvLssjRXqa+k
g1ClPQBTeRq3VLB5wlTJeIHZ4pPN0BzbF3CepXSTL+Sv+UfE6kTs7DXyW+0Cr15A
8Hj0GDQ0Ujxi9ad9HCJZ3dq5oCKobaArMTtZe3NOOVIgB5nD5IwIBFR8eqryPFH/
7ISpZuaNmzGQed3eqIojxCgXL1W9MqCK69Legy6+XTSImlIjq2cVJDCp5ZzE/fim
lbCWsEn61kn7d2jgABpSu0PKcQWW8DHBu3tu1J/Lw1b4rSAhZ5lxmOSuFF/0gbnl
PXHf7va897xK78gIYO0dif8/uLjnUE+etmh3C8CLfdFJHxC+weQyx0bZIMBtoeY+
kiDNftwWVwfcXgJsktgkX6HWC1WSioMpBflB5dNA9Ir77mq3sEOu5o6wOcAbZ2kV
xiHejh4O5fcLA66G0vekVP6oi+jJC7Uw23GP5gTdE9msf+Hl6I3bufwZTVVWO8lG
h5TgqkUT2Xu8RSJKw2u25QV0flvJ5xWuitHjmqbZ6orQEWP0Ca7dRZoU63YEchrf
GLHT5nsifgcD/pC9gRcLhJJa4vuZB+I4fDsUn0yfrx0W8sLmLXj2Qm+ucRLDgNyF
KyzmXDy+swyPtbMEJ13cXOirVQHtdM9YOu1MUOQOY+mzbFyWXRsmIX/NRg8GsyiF
Lfp4RhpLSa7uoQz3UvPCJeXKdfKhLR8ZYVIf0U+FmCJNqjVTlngxiyVvof48N8jq
CelrVrjtA386Fzltnrb6OQc80e1l3W8Qo0yucfVnUWxLO1NrBOQvQSSNFA2FWtZJ
oxZxh6uO8mgO9pspiJ4QDvh6Rd6R84X1OClKDx3fxr65FNdz6mR5ngXJkYq7VBwq
PV6zEanlY0ZmZfiTMJPksCKjre9stG90YFKfY6nlyvsimy+8Ej9i0SRYFh/9XYnD
aAAJ0B/+AvE93jkfzsfUQty141CGkqRB0uVIrji1lkEjaq9SeCuSp4cCyuZfM7VP
cxnDPGxOe8bAqKOXprczzvpRZ6agWhE/tBunivcn64FHzur+EV+iwzL/Z9hHZh+g
O2Qm3q+z4G1NKOG1CoPMJgo/Fm0QoIhrWjvBD7y49ciyQVDiP+idI/ICnPYy1Wjf
+XQGBpTB/Pp7c8EVa/TapatCURWNzFrttkDyLHwLG4fcEx/aTLZRrTCY2+bvgyDL
ddTeRQZ9tv3E6SNjbVp30ZiKlBPeqg7SSYb8iuL4DT7ESbUckMWo+McucRPQLnRG
0qfmn/yMJx2ijwhRgVOQu/nWtiOFOBmokD619xQNHfd62UQzO2B54hihD9mWj1+9
rBWkF/KdnwvCIZRlE497dpdXQ3RczE7Obcsrkr0UI5fYO5zkd7SLdnQM9nbcTeQG
RyAPTB6eFriFF/WkrdISZ2sMpzJ8oZh8ShRS7IIH665UP2qvkBfuDOGUDSliOoCQ
puHsdYtnZNSDFGLERfApTdKLCjPTgbpeAC5d3n8bolksRtP/kw2RHY2emww27tOt
Lq6syb2Js5q3drbistzecsrjaUezWILOUXdX7TEeesfKs+2AWDu0QpRMMsLdTYcR
dtjvTyoe5K7ibf0rPKdQlbcznKND0kEvz+oUmIAEXe6KFOlvi6xNTcCb4zC2DCIk
rAEfFybX7ka8+ryQF56ftCsVaOAqH4MWo8hQC1BGcI5A5U1MmCeNK35n6OVHVWk7
jMDmseVN6Wu1ynApkiNHj3xIWBUz5CIStG9eFJlPblvMT3aqtlsu10A+lGrhlomN
p2xOhFsUozJv2dOF8aLV4FsXJqIvOQ2XnlQmLP7dkKDLbPXtZ14wX0F0yaWepXMc
hnMtIXnI2jI0YMKBO1/SdaTZEB6swNwXyst/SbalAOBqAFu+mSCksQaZH49wKxGz
v53kcBIWoSKb0arPmccVdytOB1CtfQ138BBMHKSJFbe2dzLqGVOUkbgOoGdrkkIC
1zJLBAJMwvqZwvjy3L8Q3IyAXi+mmqIYHjGoqv/hyDnw1xcsLQ7WA7Qw19qhAY7x
rGK73uTWfBCREhAtZUI5fMdaWzv9VfLndvVjtDkI4vE4ZdJCtQgDjf52FVAoPhu8
wdWONndAKaCkFyYDaMw6WmTLK2J/bCIBNg7XDrmjU5QXgnBq6x1Q9yX2I+c/bAxo
ISWD9tx6Bf0/6U50/qVBIBrqt02Me3HWlN0mxBzdYgVrybLFoU1N8hya6IB/lgUk
P/DqW/ncR90Jjju5b2eY5FWZtRXk2ptqkSl2srvLJOresDwmRRVUwZuLqQFlKsVo
IGMAA20vDahk+Wgzqtv7YM6Z2acFha7hODyCQkzxtI7Odv4tRtWaf8B9FPxvRL2f
p61KuYP6kFA+hkExe3PViYr1+h0KGhPoc/zb4fnIx15L2+tukFhTFI+gOJFvAcLG
TM9/4eHsci8rZWwvRgH4ESFmtfPkpR6QRYMYsvvxm1yRvH0aLOwKxwUNxaWEJILC
DT71UQzaL7P+63cdHA6/Yh/cLzIYYZZVXWQe4JbFGzNDgVVdPWUHHHNkYXHKJm6w
6SFQLCHvjMsfw+92+zE9ccJ6rBu5ipTfVLhbydPV7xikQPiN7VDg8nlD8rW+TiHB
AkUI8OqbfMbFmsDuXyLQBxQqIZ+pJikmSRx+GvNVSLrIOjVSaQCigNXHK1ui0wKu
97RXFeQBQRd0C3V+sWvDvlzvAHgkwrNkHLwlYz9UMyuSnBoRxduJrCC1zQp5+WEa
mRnpb7S19xaz/hdl4OrBpO5yngu/Ta9isUsuNmH2hrCi3v4wcw8PTBESecptXvYc
TXVD6KDsgYFwVJF8uIbi/YM2r8kZLeSEoVSBF1DOJuwPO7hYwI6GVjP7tKzCI8mJ
/89mjS9pFMddNjAv/cYkMrbQG5Z6dqT3muHk7eBNCTjRXJOzWvRTCY4fvOBBhBbg
CWCeEDjcxH3lzm1exnU6ZZfwKD/HhaGvS8DF+0tCsJI=
`pragma protect end_protected
