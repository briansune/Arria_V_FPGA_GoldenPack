// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ce5rptDAXnO3wZHgUTAYhG0ADS5c1MKvZQk3iWcvw2BeC7TzPDS41JaZUXv8M6IPfVPT2sCndou1
OOT9MCCa8o+iz9IKWD93tlJZ0fa7eLcidZBA59HrSIuNE9pQxx6PAyvoQ+1p9hVS82bFw22kc6D9
uYG1bMRmkymdvi0kNaNm8rCAnNE+M7mkjKUpDAx2FP7sIawflU1qplOWERjf+t992ckk6gc2nVZQ
26pE/aLZe4eOtD+u+rFa8o7QlY26Oh97MAgBuBM/KQRt5dwJLxNa8ZcYcPsOJUM+hePZaqyEUpK7
NlwWS3SaHU2hcsQx5KjVW5nUncjWwGpwR6RxBQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4464)
5iXH7Pm8CCE693Tf5vYGxJGXulC0npsbcgGdokGD3VoQlJxRySrJQqImaYue4h7NJOpj15u5GT5C
lmllvWaE9lyR8zZPcDXYwg9GPOvXh0QbMjzYoCDxxvwUIKGW14IPD1jUd0XYGy3MX3439A0gHTJX
JcdrYFEt+VM/aULdiooFLSHY84QNjf3c8RFtzk7FcduP7Cx3BpCcECYOKmCLChrNfZ/wRBGdEQ9K
3dQ9FVJvEZM6FPfyl7wLchMVplJeFdXbYFeAIq0PeM7r51UT2b8hictnqGiuUXh1HlXb/W17lUYU
xFs5UtW30BbwNW/97g0Cr+7JKMnRpBfP5d4YilT/5DB0dRSP12Dx8TX9+sXMaGdMUv7FvZtTNF62
Wibf86dOPga+GJasklWw6X3kvuCLYUuUo/k5Q3YOyFSvOA4spy8IV2gKlSAAELLV79sQcxgd+1qK
EsveSn42FKj5Y9VAtO4GwBaTqmgYQFtAdPV58TMWQAWSvmNtSaMZjVNJCyNlbToh7D8L+KrOdtrX
+la3teH9jUZdWl15zTo5bB9745iqFXVi/sVODg4hG4Grn5LV+5Mk0haCHC+yNtENdL6yGGafehV3
c14KGudeLa4Dz5C0LAabsau743yBes3r91iGQj0tpCfjRBI45X/5zMjO3HuFW4wnbmB98g7R+K4w
CnrbGXTlHAa0THSbNCzY2fecoUaidu59LNJEOItIQIi29JkbP4/J695f7w7AsX1v4LmiODeIQ6NO
BZM7MmkrcB48Sg0SNHXRMSHgsh++M++4aSxJTN4lvRN+V6NvKm859Od7pa6DiH/cpW/hS+GqRzZd
6c2ks9yvRqRF3sQ10LW85+bkvuKNGuVVVNIhG+5Pfp5vHDoI1Fa3jn0XHnAGE9ccvBH5Se6GAbRc
XVlf0XJXKUabBy3c2AiGBY8qzhfvFmV/ZfeO/juUTCMISJ5ujbNJH1SMfwG1t2OXeaTpM7ySi613
22dQQ8pfZ6Cs7dXldarU0rRHAlRTY1cRJDBaaNbRDqb6B+gj+77dV4eQ3YoMgKz8nZIjf/j0hCnO
JPN9EbaVVTu9ALnqZ0YsUjo/2znQlHlAkw2vEFVwnPNGpeZPLeogs2jRD8Lij1cQ99OiGjDPHoE+
3s9DXIqyNapz4dkO2/XwQUMrpCYBspdMJ8rb2BID1rKoNjdLQFQs6ljZudtwJpqQ2Xv7LHAEOOHD
9bkwpGOd+AeWXEqhIfrQaGt3UjLibZVY/QoU4U5A4B0/UIW63KN/7ZX1eWgnd2gccyQ0iD/7UaVE
8mOGdT8XrhKLXvDjS5KOZTjOyHd+997+vRjSOptvJaDBqmCbcTEm5bJS4qRkfF8KRQ7O8Xy8ff+f
8BQvEwfG3evoCfMWi3mt9sIDLCKgyb6q29eoXIfGkI0JG403+cTo9pTrq+j+Dv/YoOFiRWcrG5fC
DfCmNPiRZ6nNQwiFaPHVlIbiJDkWcduf/09qvZfxhnlhhAoG9KhyurdioeIJBx34ELfvSQMr2PYU
pH56MNGkOQ13Op1eLjJjnpBiBB1WTrN3g5FOV9C+f3/ytCfnv9CqFZZJEHDWgPCJIey0u5NxX2Nh
5mv6nBoKyJLaEeHyp7QHhYer4VOM91JuiYT+Jk/iS6nOD/2CmAfXj/2EywGFLwxwTKBcqqG+3PD4
5qWALfnXqxKYaiE6iHvDuONrvXGLVBXVjL8JZaZSFqiQBCzv+YokJr1i8C0W243zgzUR8WQEoB7z
iLm30kcD8jKziX/JGXLWgmz1dFp0IuoXjSvXARETDdtf1Fvo0IHJ/QDLeAKIpTrcjkWwg+OqydCQ
hguU1p3VDZQl3kZ0og4QK2N7u8+fdRlrgjV0uSjHatfttvf6DTBimtyJhyWH3xEdPoFCEZeKdut9
To2IaOIT6vHMKxQ4zY1tVSoUzfmYNKgxVjymcsCyWkDY44++jJuaHStrPoC8Zv+2yWQAfjQcAVBG
jy9bJVBGvnwFUtQ6iCbSwLstaQpYyv1KRQyeKW4zqZJY46nbDuaWCY2GDgGWjykZpXTNP2iD/fJU
Sm75ddW4DK+sPyjuI8cDspGbxBJSm31ADJcZDq3qr4x+KuQGzGwl5tE+HP0EAB9o14VAWgHLf7z2
EAL525p5fP9ZsFKI6YDtZf2RKmZV6kDDAQwYgDJixWfF6HIFYoue1Xe1653kmOCL4cbhfjHpN+nx
KymzJKaIMNHJ4F4p7PqkhL3UcyDBOaK6OUUDNRYlPLLi/B+EcwDy2iAkeRq/pXDwtSPe9XCwHP0g
heH2BLZp78ZYpUwQ3pF4xhVckCgUdbFPjvRS0QLtiryOXmD41GkuQhvjYrKFOtNA+HHxyg46/bNP
r04SXVn4JI/LGy7NufU/Tz2ndR4jk4HKxPDRUMa1curx7/pL3aSbrAOkh9HoNo+neKj6Zdd0CWJd
UICINNqDupudTst9ShQXOW4PM8TZwnp0UNKyTCmUw4MrRx8BaQ88vASkI5k61ISaW3XSdsf+xWUg
m6/CyGFIQtn4zo8rPl7svVEOG4+7KB39PBilnZwniiLA5QKTxnXsuHvnlIe+zOWrgPYjgOmqOSaS
xQxa8ApX8mXNassmCN/mluOV1kizyErbLPP2Wgo5/lEks0YbouluXSfgLJwxU9gKEOC0EAp5trGu
qLqs00FE4rxh2XPMBlHmtUe/KefIoBD4KoYH5F2aBPDZeOS6TD5IMQ7TT9NGNblf2rA0KbVvEL6B
WgmTkMDRMQ2Qb8c0vyN04eJCkfZhd+2U+D5Him74aOK0TuInXP9GlH0W+nKlKJ1WF0YqzmwhgFRj
Sdukygh4km5p8z6DoCn9n5aJVkYL5ww1+xx8u/FR0JncPBnAxnJbG+q6aJAIva9lRk3lbXQThXgf
DzJ06a2QzOMGU2NNOvjH7jN5wW+KJvokiY7gV+4X1D0q1z/5dSAyOlnmlNxixsBcAaAPO8qd8Tvg
sUq6A76Lm4hsJ1REUGW7ZOrUM8jgfwjv5v2uTkSWkNkrAgCcSyYG5KRdWS/kP5LmvW5GSNS/GaL3
/bhZsRDBdUo9uWxbEBeNcOaCqefrrMoyFNbt1om7izRKyRJ/+e9xm51uIa84efs+Tsz4MtFzevw7
8PW6lb9e6zYQdgDUKxLDT+0Bm6j+aGGgdmPe7ia7GegNjThMvxgu0ZnrsqrrmbCGfVdaIA3QxxWz
1hYItq+Cxknu0rn3F1QdfZ9/NV3IwF61oG/RpwJTOhwTAwzCX7BT9pgoYfG+fvWk3zONHejF5WtC
bLPgoxpYtac3lWpaFEoe3tSJ/5rLTGf2KHZsyA67A6I724ogrQZWPYEBGMXf17L+1WAAreRUiTTO
AaQmGv/G4woTQMHZVjK0/CFI6+tZmtU3BkmA4mZicm36tGcQt3ZKqj+GcQg24u4N6vjHKWaAQEbc
6it7tf/AzLeeWXgnWO7W9fFtrvZO0Z8QT3PsSvTNqGpO6v2uiFeqfae9qXeV10WJXMelsjfoBYYT
UtDF/vHQ31gkTos2RC38Nor4dVGxICd6r07dqqI3QfclX0flAV5IUgT63w96mO+dBlwGoq4gZlLE
rzR8RPk1BRSeFYXG+CBfrrNI6pWEVueDBDyx+oz2zpsw7XUvABhBoLbCSTCw6niB5YjIOwPtFtwf
/hyWHIkwB6X+sBfWSDi330gjg1hZzpM5AIhSxGO/u4p6hsggQ4A4eJxejV+xlb1y/t33eDxbW1t3
RynXVGJi0BBeFqAoWHBqvoksSyMYjAlgiaq02v4pmWhSe3P/1idL/N7TV2pZ9fdsvvVLR3IwPm1b
ICVynEEqiQxpsVluO6CY+6pVlipvRkSQW+lwLOangpUMgQAdSjlGLUddV2MqRYsq1QkrkYqRb/TR
Vwu+qefJBXIdWbKB96cEj+zMJtwRo2kJFk5iPDY670Xl3+3Yxfk+pCGpufAu4Ta1Ai5j1Tec1Eev
otKMxEY2gXL6mdP1/2Wbs1CsZlb7V1KaFMmvwVdqduK0bPt38CHajdYVOuLu+/PszUKFKxvugDBq
QFlae8IieyqyXvcUHWMk4xc4GTx6hI4e6C15KeAXZavWmP9mMrXSoW8FWfxP8PG//N3xEsRCa3Xh
s7qQdt3hz2gUztUIH5lh9Tcjvgi6oUjdo92td8f8BkiSIWjKM07/7M7/kM3TD1fA6G0x2z8rUD3l
/WiUq2HbRF8P8Av9mzAI8WVGjWzqhMXO3MZ5gTLKSr3awJQzQIZsCB2kxviiclwuL95JhKboc+4A
P/X4syY4M1nNnlOznFy8mlLFh/aVyVkjE0RLf69xiigqJ2rcQJ12yGA+tv58P8cUgnBoh8yD2qh/
c+qMHyBPNZtpVWTf/F3ntL0x2wQsURnbQ61P/SB1+5gHlBfdgK5BZFfSuSHPRJ8QpoGz81tsLrhN
7GwgA5ruTc0Nt8o/D4UBJDathzdP3hyj1eCFlewuJU5xBZDDfsb9De2HkTAcy0KlzEHmNlBAgQdV
8nro8GHUILitTMI4Rp0nBhsoDWycsIMBpVSqnwrDtVx5nZd6DXXAD6B1nArLWjh48p0JstqvbgOz
3WI534Gr6Heump3sEDx/Y1a5R2hYpJ3mkA4MNxdNbm0dOrV12DFaQsKdTss+NOfMDUfYq1KIgS3S
jNLI64qc0nEv+0s77cfORXSOB2YScaN74vfRqOaDti/9dVYMFa2DoVheWPHrbXWKEMRQugmz/L4m
DAhnxv1BB01BrxbqeK0cx3DMEJBkrzteLM+f9htE0wEUvx1GGuagRKRhVik3zaoe+lxdfKiJ7G1k
VuxAD8qoNiACIVw+jTnumKdbXZaUV+ZGYccwCB1XlWM5HNuZhNlSFWJAv7W7BqD2ajLW2ACnQQW1
4xKLlpcHmYtYZJZnFXdCKNcxOg7V+nWzeY2GIxIcpKqN/7hNhAqpwk7WAa5wDgHv3CwOaEs1xZh6
OFsW61svTntDD5dl1E9xOfR162yzoxJ/LdnflW2odzkP89f6Z8TTyNsTBznib7N2n1KWUtvu1SfZ
2HpPd6yPBLWH+Rcf5GHDfMhdU9jRpzoI4aflnENJbisdmAQnkUQU70HnjHzOU/XrJ27QAW6vI3U0
Wvpf1kMHg74bLG/8jl8PXZzW3u/S3amSLj4RILWT04F2njwF6fNholkAKiH1ZJf9euG9TDX3jXos
IYPL5VtUQmlO1/bM6BJvo/5lv7GB2jJ61HUbgoNEW2z1VdTU1HpSpCJ/1lR0NL4Y/Uw8TyBvFOdc
qCWZZgpURRd4usRi9EvI3IZ2kxvdNfjZCXo+uvx6tJcrAW8gbgsEPdyZ4OIUE/iX1TEMChc6DsGA
GxDRezGCI1Vd+kK0ca3mmmrocQOxCXr188m71A4FtVR/UdKavyfNktRzCO4kgTHPsHQaTNHvW78L
46rreoFTVFWyL0MD+8IhAtjdd2sBMUDaPYYCQdKNijzrPcys7G+uTHUuaXOC1aqD0Ka5RwIlWwqn
vYa2JuC/rQ+RfO7lqp8ZNqQttkJRDLb0mAbzu+VNJ7ajvclNhbB6ezftIYcxYcU+rmIeU822N+qz
lYhjBEaH+dcXd8MuD1buH71Uthh19FofUrI25IZdmpq7WyVTgODehwpIXEiacidn32nBUt1enNYF
U+RwleYkLfwP5+mhZow8Zben2ChkrZawAesgptXPQLXG0JdBQt8Zc2IrhK02ANDgHBAcNqNXorb+
mZoUQDH9D2N+WFSaqqneINZI/HfxccWWGYfXFu3Cc6hjidQ4LOANwJpPt36EGieQKLBnzMlost5j
aqA5uPvlkyMdoR3+KimbNU+euPFR/vb7SZiDcTmbRwoDJRx6jZwpRA4zShK6EsmGwzL1fjIm6RCQ
2dKJ7KOS35KQExkOvpn1avM9mQ27YO3VKXE36yWYvd6DXIq5nxh2h99QQzrxDU4qX8Fmt0QcPQoV
Y82Gp/Jo0zykhAKPgMsxyVF+
`pragma protect end_protected
