// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:18 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
plJ42ReiM7Fn42v1UfeBxJ/B2q00I9CFbeDuUG/daROQg98OJ9fLOio4sU8Q4+CV
3nQMd1PSzASz5JDiw+2MaAu/YlBN3pJgRgH07kDO3elpfVRZFsQm1wQCAJB++fyZ
7p/sJOFR5MTladkotqPmu3sx3Akqia7lVPbUJMai5MI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22368)
FsgkSV/5fUnbV39AyEWWaree24dyNmeeDGiDZCSYUS3WEKpOiQaCngpO7nepxEoU
1ArcO2rZR2lHkkQkbcrpcexymHVU6rZXl7732VkKM9Sww8fd01ok5W/vl3Icjj7i
73YHyXvtr/UGFjdHrC/WQ7/tbiVBOX8+5YMiCLkONyvzjoSfU+bBbvTvFPGqHwf9
WJtDopYgT4PEFiAxm72PeyViDqrqQ6WXx0zeB2RhyJ/G2MuuL7bD2VcIogYS5/vs
2VZWeZSFXZA2fbg/x6DwYcFfnYz5cqSAj+2S5zQDf2dQdmxf2De5uZ3uB8kqbDIg
sm3xBZIPg22pc8GAgdpWjYuaFdk8O3ST0ziq1U9xcgY5Lv2dN10PpuFgH56QIQ73
cF2z59eqGR+AwqnIoFTafWDurAMCUvQgaJ2uBL6jIS9qFLpKvRg2OGX19wLci9W9
++yleuzsUp2Tyb6vTJIQrVaAUJoM+1rq4uFEUcVdIyFnvRtknUHvRnMyN7h+RFqS
TNXQU1NZFtsy4igAcjKaBAUuOHW8bN2gE8b0tv0OiYAVmTm381RWVUL/Dq8LZB8Y
ZaV6bOCRciL6Gn9bMBLg4jhbKeKdaYVn/Z+/ukm/xrxfcMGKAe/lXnsU40p7BJV8
VOszzRqZqiORMNTJ3c1F96J61ycLcm9X8AdM+TprK6pPacn2swK2bjQtXUozthmA
0SItJLZXP/+8cRdtzDulJO9HUxxKt6sebPPF6KuxN1tUC5uKV1axHZKhx/JUkruv
nA6DfVvOgpdL9KninY9xdGZZlZX3r6oizcshA7BHnHAN7zBYwnVOam2fluESMkjM
BgDtMnDuwqoosB+2iNst8ODQ0V2f42mDrT8nCINdcW8WJVET03MEkvtK30q8XWWg
rJ8JRrbsgSyidPHGfdjA8OnbR0eLATuidX6LnUb9dQ6Lty2sKXJxOm7/LCu0XVWM
criwEpTKzTMyX4xS4mmIOCwxAMIwzGddcDeHYdwDiJoEZkN1OrNkSZSA/eo/LtM9
H8rjPUsLdmUBIpzNcIFB5OOhtlRTU+HKu1uk4b4GK5+8dsZZAAg/KlBqLXqpjG4f
zBvQdwZwSS4jjR6EzIsvkeU3NeDU5AmALRLGjjDxnkOTmVRHaCe5pVDGUCTOYdE8
8j+UrRlesu83sjt+GwaDqNBPF3MYEC8BbnZXkgNVDGl0i7YrWdU5BtkQLJQF6gNf
ANUfREahdCJTlDdgQezTeqJPj1tc7+3JZKbm5lOW5pgduxNaZiA3Z+0KQ+DulnM3
gDt4Z09sBMFiNRySmQWK/cEpn6XAHOh3I3NH0XIJL4DfnUQPWuyTWcGxAX/Gty42
rbJXXJi/xU1rhGnVwqb1+UoxglrJm1gdtstsuIOLECaZJpU/L4yJffgWPnUgRBRz
ge2jDgu8VHnCV7uX7zTWWqhbbtH/0nP0YLxTeSXgIrnEc5OLvsLuDwxb33OEnyHn
mZ+PfQW+v3TMAdwrfTmuisqzGCoZ5fTdnopseGNsWHEFW2XF2jKrtCvaRtozbPiD
aNp1DPTu0J6FSs+kJYnK5VskX3A0WT8R+ZO2q2epbPk4l8QPAam4Ojx7oJDx303c
XfFJd7reSCGZxezTW9RF7v0jwtOXxgGATyQnAatBvOduvPsP1gYmJ60qThLofXxp
mrJuyH1m2Yo718TqdsP1DDjg3clRn4zCGEprOeIrKye8tpGHCGxqtLOU7tHR9UF/
SphFj00+/eD94Y0rv87PRsQbrMRQvQmmeB5ez5prL+dFRiqUWe5qXNNZh7CMUeMb
0jfq/h2KhKx6X3RO9R/946umAu+NVrzaTbFfN1aD1XOn7GCourBRFh5V2EBO88Np
Pwx0uAxXIOBUrpXcYqXVPpqBDhDInV72aR976B+PQMf79h9ezZWRD8Msjl3pKsSZ
iP4WCWw8cowXVvg2no0PB4L1dAXEqACFNG3qwg4GOJGOPRUoK/nXVWct6x/6UIRb
z9sYLARo2bWPVHHfTXh7O5RjTVd7sK3bkcAvJiOlgIb3XLq1pdEOf4Feygv8wNvL
F4FxOnelyFp//hI3iZcuyG4MUZ8UdcrbRoWigxbQyfUJFvBvFsRmMRIz/e4dtrqW
TRD6rdrC196/etNgw2nwUpg1MCDD9hZyUmyYXtzGiv3IyhL5PLo4trCobk/yz3hF
VSg5grCeqOJ/Uxna9iL3ESpqyXRDLp0AE5KOGJ93ze+f6l9UW5EXoFPKL0+QVhJc
mQAN+3M5YEeyvT0DGGvlVBX+d4yYBH+Gr87XhwyqGwUrOqOw7slGVjIsiSNddcTI
+MHIhYt+C6RmLb55gTg1b9Jm58XNE6oDhXJMh/ZpdVcRIEc2IxhpMLV3KVbirCwQ
mdGxAuWhxrMsz3i6nuzcwAxuICcSX+ZxnJhrkn95sIk7bUTLx70dcOW6fOy5jbdp
JSEFCIveju8U8lpzekgBW0o2SI5T68/n9ozDfPoiyhNFmJN4N+vVkbc3aeQM7yQY
rwb3l31MlU47IepsnBkvz+//IiHb0Ad4XIX7upDSC1uMBwoTIUGoKkXkwWZui3mq
qY2nYm9Gpal5DBhilgJreBQQRGg0PHu4id8P6yPHLgM9rv6LVQP4usNhfhldxLf/
QULnrT/n1Cp2a0kQuiQEQAocxZVzuUEaCEqNliBJwuPe6UNpbfoktxlKmDQpDi5z
9HIA/ytjzlH2gjPEft8JP1SNR9L6Msqh5nBcIXL11MJ/FtxWQ3Mvn3JeyByl/xq7
e4cSobxwLzg74jXbWpzPQcnaC0KVOCp1wVD/jc4tFMgsC07EYogjqwAReG/VODj/
sC9MrA+JOfIUvsYjD7Q9rufh+wW8qsyqRUdLJb+xUqF1kftOZ7OlIMJCI+7Y7VwO
7suxYPXjq9XNstRoel6rC/j/JMm8I/36rySCcv0aNA0mRbms8851guiucPzAZu86
P7Sh20DoG/dVg3zJBUrpwSOsvvAehAVEdfAa/6GopZRXZ9WcEBdF9+0PjM4BsG6E
JPrauW220UCD4WPyxm2CnqlsJT4InVq2Z5H/M+KY57VGvaSFceCCU17wJSkswlep
yKOIoSu624r2iRIa5Zv8oGt2VBNIIhVhuJ9H2N4pKiqxqjMc+FNoWrY9fPtnQPyq
7mCE6tftWJtDDi55HtfN30mPKQxnvxwQHZHXA7FfsOcZcQVMQVprODFq/Y0APGoR
wTgivkJehjy6GtNk6+Z9GCntXFc8RTfaD6o3G+pFXBRtBQ07WcZpi0kvEKfoJYYI
mG1O+I+gUGHLp+In3nT+eKGuRl25TqMNzzen7ZVQiIo2rewxvBWK5v96Ai4xMncL
uLzmcBNCJ8Ypxp4JvEykpB+B9pbNDPeij6CQf2YjKyKhaTm60Zw+PSAw5gcujaME
49ABR1J+7LCiSBFle/j7ioW8JF5nBTSh8+0LyqVlxzIhdXts4Pw36+riwZhrau6b
xhTxO0IvBh5XSorgim7/U/QJmNVznegpRvt7z/oXEIcJ3smQT0Ln2M26vaTLYMKQ
9rEv/2y67Hk4+/qr86mhnQPc7YrbIfgqPtHKwbV0Vt0G+tZ9zp+q/ZniTFZo6ezi
6+7HDa3WojcDdfrJkDr8C306JDSZytqdO5RoLGwlTmKtI/agNUx2+MoaK0CaTbSF
Zy0rzTjR1LCg9Nn7YktXrQznt8OGuZGHtNkARjIIfDvE00o88y+NBkPjw+KsLNQL
XCv3+CB2uc3wO4VwLkr1Jqhw6UVxF+4YBAn5/16LUT+6Xuy5XV/6WEdFPcZzeZNJ
nhdmV1RjIBpTttyh9bwc85px290J+9dF99Ncd+WOuODZbjVtVmVa5fZrCzGN5M7W
vwsE160wUfxaxIFhGOTcRNx+jWNKLu9FGlVfJTcA5rsf2JitJ7YbT3zDT9j/1/9h
EmK/sriV2KwjA8Ih/3kBYVWwWYh8tgWQwyVXPHwZgmKh3/sdjPy+7uQSgK4Gp8Oi
sTh1nA9bnzgsbx6MKV5eXhTysh5xxpeGHZT35D+e0wWKoCTlS/ZGY4GQse3XJ/UI
icW/PYSx8xFpaO5gVjStk2vrwWVvRKOKpMpyJgQ86eyxXi+Zr5KYhY7zKxNTyyRW
58DgrndFZuFe4tSkW21RM5723DijGvurBK0+wUz906EYdo9SQHpPSvE4btiQDhIR
cYqleVqHG27T8ptkWrAJgjoROWJtBr67pxjLkoEUyvDQsZAJ5QuSC52QeKSDF3Ea
W1ZTbdpQKVhaux/T0HgSgMI7A895Sgv/XZOZiLHXlKwm2Gyxv16y3qqQQoG4W8qb
KgSMjr9CtdFXAN/hjNYtUXtHa8/ibJEUbFbHysfxaIGQo5ubXsFzbK3Z7G8T2ogC
wxQ1kk1QGL5sMy55yV/tVB1rmrJJnAZsO2WmnXpQwIFXZVHYyy2Euv0jGz/Ym+9o
9X5IVBy0Jn1P2nlpmn5hcN4uhcTl6w0evhgL9W/cVeIsj2/Xcq/NMKwGukjqFAvT
Bhh/acyyadbIm0bIzWx2McXkKFuS9MtTYi2r8JWZc0oeKK/fOIJzQSMGA+5/vC2n
OT6TuI13iBgeINyevX0ykuRR4zhwht2HME2Z/85B8ySdfJRvJH8DnEd2njj+pqnP
oG4RSlDT4+fLbn0kdK8Lvz6CFvni7ZxYKfGbVAtc5g2Q4tAtSSgsbDlkGR3oh9GY
Tg5uFXcLcu45jd/I4nlCul6B8rzyqSDSBmfmV6Asfj2/kZ9D2ek5Ap9AtjFDrhfx
GpIos7DqaRznuBm5HAI/1nhFE71Al4TiWQsJLtaPL4PaTVIGwh9cRdt5GS+d99jT
8BET4fohGY2WcuTtvtN4SjJeMVut8T8eY6lseghKZ5O6fh70Vv5exCE2Fb7dOIUz
Xv8tXDt99sxAvJCDuQi64sAQlP0LrLkYo6UCPa1SCjyxCkTQeRolO4yLvtzD0BOO
CEIT7Hm04VDZFihr5tr4dD5n44YSopXtgSVYHuJuSls8Pq18MTJpNQf95k7PzVcL
AUpIn1tRYPXSyacqvk1JSYLHJEU98XGruz+k1f120JQEm8IJQFm1/dbnNdx/DQcH
97obd+MaFz2+Onn4eTIpZpTEyq7geskLfHYCxWlOaaKQDqRoISJwUKMYIMQwLvbH
IbDMI3kmXO2JdcvDiot1Co1bkRh9S5XYKd5C6DTjCvXLX1DfqNWz52dpnk7DUAX1
Y+mlkVdtfXHliMpYdUzc1Ak/ifeIyzGIHOVurULjdpAYfM92uCSAT/N8P9Wm1GPl
Vc5AoKpZeD8XUXPG/a+hKOXS+wgsGdlmRVlOiD4Tf/8087oVwFFI3buzqDx+rfmC
PDwJ7Bc/g4CENH6s+F72z3TiCjTOvsFZo374sMwEWlayWUC8JHCQ4W8Zw7kxJFTn
kq/SjjeeHy+93svdRt5Ek4aWJ8J7CCkG/MPbnfMyw7+mVhaaCVJw+9m4c93DfwwJ
t4xUk6l6oWsRDgm39wL6Vk1Eqx2SGd/JiWy35i9nxJUTTUwSGuOpQ5UJsgeGolMS
sDf3B4vtGYDM9fjolTEKDS09fl+I2gm+Rc+CK3KfZyajfYsmb9B/ZQFW2fMjpT+q
ocO4aLv/Bjyb2brNvGxvoqMKNdok/CxFkq30LHjq+/xPcSk7Pf5V9/4MS3P9lsGX
oITTeDdokJ5Cvlj0w3marEaxvrT/IsnhCcMEOmBJgGk1FReYOdrhMYXu8z5bPstx
xabaqFHkVeC3oNDnodgNEg2ud76jVKyUvgPqVriXZUcOeVlnYPbgCXQU1lxg6KMZ
7ErwOJy4H751Jz/ujj3Ql7KaFl48VfwXJcr4sJWiRQaahTW3M/35gKtTKQYcbTm7
YLQEZVUBttksPrARJY1DlHix2E74pb27HOHDTweNC7LtnVm/HqA+gX2FwgZs54vG
pbS6CKXKzx0HhjQOwNtbwQjY5aNfHJ8UhUARpC6vFTbQt9ePEpnf2WgnnZroJ5pN
5VG3WzTDZRlqL8j0RVvOuCgArK0oaMnQQdqKALzgsZsvQ/9WiBcXwi74kCNGWIQW
JfeekiVvFhGU3xsxavasSgORMhC/0uFthw/TBWXZphyOBEGaIQV98NAmD5r1hk4g
oUutRQyJFxdgkWMG/nGtrQ/raoDErxV5LaV5K7UXeUAXWPQNjqyV8sj+1N3y9Uhz
PEZ2+Sgtjb8Ty2uTYgPU/g0sN1x6e0997ai0vCXmijEJQaUoLUrePOqbW52hTSQA
Ic8opKaG9A0mpxYwyPN/yqQUL69PZZhZtxOMMmFCyIGoNOMnyqBEHtzklXnoiZfn
Vo7GyLMVnXLwfQzGYO+ZRCha6yu7BJBIqtzWbs0mRWlGfXGsiJbFIvVWgNz9bTAR
4HehoP4H3stBA1v5/xEE8AAlkESTelRRn72zZQpiz21AbpN/ybvcii4CIziam8f1
/9m3oYz05xnvdHJo7l5NtFCe8Jt3sY0QQ0VyTsZZuR2U3EIO4auyFAa0p9CcC2nG
MLq/JBgW3FVzU6l4O8niMG/AJrajIG7et6+y4rA9G2lfWr+rwkuIW5AngQhOB1uj
LMf3XecgXByRltYi0FulKXaOZHAy76uId3DmK7kArf6NfsX8hznozmlKbvnLZTuB
g9r+2WMiMWPbgJ5EolsV98BDnCVtKIuJ+A13ruu6QPTTwRZQ+B/dOtwwg8WhVyx4
x0EIi64fOy8E5zw0VvymEnfMoMlXrYoCOA0A7bEr1R4gQLT424MxQPemsMGGVmyn
R6EkevJM0Wr0dGLVchXcnQpQyG8vXp65LNv1SjAjiimP3U/6ds9zULh0n5/e5mF5
bGugpMDmW3KQlSsCjaWLl5WCpsrkuXp+fc68pMpSKjsvmJ/l69wEJd4suIaYrVXr
TthAT/QPsR44lBnjsOZlxK4zgbGtmT1lYA6iXyUkaDix6S39yt4HSH6JBt4R0nyx
vUoBt/aBGhYz5nMrHTr/UZYfzH+dEGHDN5XBV+ror4sBGZzCF2xXqAFMfNVLjmua
WvGw8HJsG157m6kSJKydWGMVjd3+0wAYre+r1bQeGR8tGOWpcOwIxEPvMCrpBrMP
Wf3F5yg4PgRNTnqxhquO+VXPnftWD4de+OV1BML789dBelEAozxYJZwEsbCgRVT6
Y7c7qrYF6Di2PUYQ7vH/sMv9ww6DYqkPK0QV0ra7tig9PJOOAAhN9LIgx01NxK9L
QgNH9Ng/i3FHIe4OoVwVuSn34Ihiiw4GmOL+wvNAb3ZCI9ArRvjHPfqAi92AMhRP
3QGVJ5tJyxXLfMudOhg7NL92Y1ainxTYoQotAYwK95z9tDv+Dd/606eU5HgCoUo1
7FOrTZZ/wfkAcLEa52NbzLt2J89yVhl6NzQGi12iCGOMLl1muNYlv9xR0exLqLC6
eqlNG+efj6bg5RvAN0Ya3IAjrP9sIz1WZkHRvmsCiRxTjSAidaWuOvGGErkLD/I1
34XpJBQiswU8XbrYWzaNtKseCHTBQliV1iPuCJ+/jSBR4Vod7BM3guN6ChOGiuY4
6q6abXnm6Y8EsLdasoywgHKdGdTjiSkQXs4nBgj6YdxuiSpurMbNh0UGT4JkBtTY
96RVOLpAiZVNRAcaNp3BsIxs2OH86vmPnyinutyAkboMZGuNCyimLwpAw95Od9kc
AU+p6cWtOHu82YHoIdQJJtK4ePlPL07BOR1jHq63ZQXU7pAbmGM1eDl0hRQ6V4Zw
JPkOMU8JJB9GYHvrTvxfrV4DggeL9yVOQawf2QQO3zN/Bmb+yZ/q2nz7kYojXffW
g3KIMe6jMGCXidQSIULhqtkJ8zaZAWBto7RVP6Aie9L6yvqVqpNvY8KD9V4cM5eO
qsKMofDQhc3MSyx8DJnUXPV8Vb78F/ZY7sFyaPp3bfFZ6cvutmPTcGIFgQmGFCKD
dfQGhL8WQzJali0ydggEW/4VoZHeB6vmk9SkNxE6f6Nxlb0HAhS+jHZFI6ZEmEvo
XXod2YswU7mYdMeDHLpKSPkFWLhqiGkNIgzNfD39sX2GlR19D1uRIoX8J8/UyRuo
g0DPyuzreH/K84Z1UeKRsJDDeV/ViSrB9XRun9Pj4UzWE+VijoOWikqbBSb0XQoj
03BUuatfZx3WM7atbsamF1kb/WAMxhNSoDpoIvbjUxf3Qb7SikAyyYqmAdNcUPyZ
VCwTZzP1LGujhvzpH4UaKeiit1p3Zv/6pnL9OupNIDpvYdHVkp+I8bX5alQyZjS7
yFQPWtZB66dVrZujJ83I+XRxdk0UgclfKxJXgR5niQxgAHYmYvvzTcdU07IZgjUL
hj7NkUJd8xXg7hGgwCznbJMslZPC+x4RtPXZRyohO0ZcA2yNAfW/1pUejua7g7k6
3I0DykRuSQUK8zIj+90GPM8iGpcWL4BruNk0AZqA6M145bjvHIAAGlgj1uOBAlk5
1TVxx/IRoliDgHIq8gQ63f0SjWCB6mMYG3yUPebmuFGcuNQU0Gin4kqf8cerm1/o
Vkp5OruGANRr3vjL0lWSv6eh9YVWnLSUuyDVc2iduTUBx74FcNVhJg6RRN+D8nr9
vPbtD0yLqOtGsHWHrXdE1RVTh5VXsKzb4OAlmHBtU5+UHBU6a7l3R+PnXMxHsIM+
6y4Lx2/v+8ivdMR5Xj6ISpB1+ORwj/PieuqlEwfECj9q4JOPpLUbkARHE1priGKN
9AWX0kWa+JytILDXjgcmm5aJTO8HEXrZPVI8WnfN8MVRy2E86s6RQrmVIXo6A6V6
lN4vEmbSXWk1+KIAslz4HYFmh0d3+MfY+yWA21M0gCBmFFobSN8T9zt27zaQWIUC
cMShLAhm+4J+oAmWM5llNqaglhuevzzmOQe0zWDONvrqdipJ+vOI1qQXEU+mjBoo
H4Fj7hHYuW4Az0AO2RuEW0n/vsRq7+XusqdGw9UcfjbfjNdK4IrYAKRJTxPsJiU/
oAB+ngH/CtM0FCAvx93wSApM8f3ndCThmLCixJ+lIztjUrkl4P/Iy4CL3vuzI7MY
e/0JopGY3+RXBAKam7OaiS0vOSxdOU5rXXOP19eKpSAzYqCXr0Z4OpW/Sk0xHAQ7
6wz4ry+99wFZ+Ta1ZLmm2mZVD1ydA0VHNaMaDbsDq4KEEV8PTpi94ys7YLSa3K0R
jt1cEEDfZrFZyXjUzhUabwrteQcVgeiVTcDWG2Rh5Nv4uImp/F2mnSTONoPHrAM9
JbGMLh6ao/kOKBAmAUroWVyijSO7PUG5bBfhe5dB3/5T1Q8+zAek617ZJHe9aQr7
88EVEthwxifOf7Ge7EAGcvXkOadkxjLM413jbRc3ULL7v/zqN+JtyvtEdiatOnSS
f7vdMfyPme/9/5LxWJXTUen+ljvQivPUlTFTvHgmByLE9XS+0/JfHfYmo2kFDxT3
bmuekfwcN+V/jdVxzYuj/ELAG+KciNYk322e5GTMSWwmlL2dGVyCIO2bqWdjkNiB
paWamoP8Pj/J1azeaITEzYVBhlIb7sFNkvx1OdBVW0YWdU4DYGXwt8CqFkGibW9q
oqP/VPaGx3e0vmqOfIQ6UqD1G5kMgKlPdNeEdq3hzYB9JB9T2AwoAsGEug7d1rDM
13KenioAkw9/0Z3PCVM2o5EgYUWT0esnD9GtR6MTDIsk5Xa4IdIBAniqDmlPt9m2
QYY/GLy1EXPt02oWFsjojvQj4fG7FWN87fL2dmIOPhomZU6DxEjW9wtU2+S43lMj
tHZg/jfwitY+Wup/zOQjrtGmZmAYIDKNNGSe+8EMeCETs6kR7UzrlPdcAcBBaIKF
sFWcKvdZQ9vY05NaTEhyKHgVl/3LMUifRnzIZH7BuKsPTA/QHClwWVhrmP8hOtpr
biMRoiG/o6/IsGpD1FZO5rCO7nfibLZWHOIejOZBt4mI6rE4YggZj/6USM2d0k+r
RLW7D54+kyT9o6bgnSP9SXvIU4MB8EMCt1VvCTkCppVvIUE1e5aWQnsMbT0S5x/3
7h0etKJ6D2RG9t5c9/dRz2x+d89o2eyr8VCIL8XfUQSv4Rvanly4EHQQm3GJBF/L
gQNU/CZ/DzT9vELfndJD/CWf4SRjr6Dinm4ZjgQosWFPlzKwEWGupvManDpJjv7X
3eM4726Z4qctKb8+WDghk0IjOmMakI2JuC1zBJhkud0Re7+oRKUgIsjsooznS52p
FU6/Uf/IOv3duBFZvh26338X+ISGxJZQpMi+XS0WCh7GvK7jFtiz3A9L68TeR4pF
yRA/Dq/L3u1FYmirIl90/dkzNxcPG79L5a0biL4/Cr3VqRujx6GZFNWMGgp1yNLE
9hEfPwV31m7sCR0u0lJIlH/fNTp116+aMUlABptw5V5OewBsxCu6kTYl3+jiYBhA
0YimC7EqEdZyHOlVakSVby+nnxLJjjZHp8g291SIZM+ga/AfE3RQJDb0ue/1BbSs
qciXFnGoc/c9wBLs+3QCm+vZpnfVZCdXr6zHjxODAXriJDonD5t9193Ej4ukAeqj
cCYA0wbdmhApacgVM/0lGztRyN7Vstll38LOlfb7b/Q6ZKjT0FrO3GA7MV9EDEC8
tlUAaejMcsBbQN+3x6Jbvm2QjEzR284a3Dmg6dr7Ac2nOeKgWqb2vJxJCZ+zXAAN
AbKDAr0sroSyySsu2MXMvJasVBGWztQLFmLIgMFMoZ/9EFNP6yHgKzjTqWwnDqL5
HK5LYoycluUn5V+FuU1YnSTf+HmTXQ2fOh+uyspz3FkSGu0oLkhkcj2tPaREE4Br
BUqypH8tJhUX0N/jizBh8nLEi7X5Ed4rnn/bnBllVg4v8Fyh9tOEBvXQUEgzzD0h
nWDyh6K0/iWcwthSi8DndNQD00q28M+Wdj5EZRNkyb3MKqm07OvDGdDfbdxXpjJu
sWEDG6ANZ/u2i+og/N1nqQjucaAFXCE00uaoLA56xL7KFoYnnNX0IE3m+kKijRed
fqp8+Fl0Vvm0x1Fy312+oCW4ZN8MQi2KWDaROjO0uABP+LEbi3HgoW/CxZNzq5js
N3q2wxjiiW5BOY5zmpE28GiMVN98HFvUCKu2mavTBE8Bzt7n7iGcmmpWTFgs1Ho9
08XCYpbo/4CoflS4keqtUpVnp828G6UfWcevfWk/TTgq5ib/z26iEcboWSZslPBD
AAxqJXFaaQoeoQonkO6dqeBJBv2M/xdvV0f6gHD12sucpG8WlkNOYBtTNWWxGhfJ
ud5qJUXWaFATJYmZhXQz6A5hw3kHPoRvBbeCcJO0+fQfSvZPty4Pg0zfHt8lAZ+1
vRaT5eOURCeT9rOVV+SQZ1/bktBew4c46LiSAlXcpEkiNBvOlDA0H7O1Q2AHocxU
BW42+HC01OMTMJfOcYbdkBt3eQgx3x4cva0qcktkC6P/2u0qJXQIJrx2VEinLRUy
qSPQ3T3QnC3L9KL0bM41ym14dqVKVZzvSdAW6Q4D3XtJeUlxHQx+O3IXQEnSCizl
I1PufUkmWC37pkGo5g/MxjW655NG027sEqnwDTjbcpvOuSo1/lueRFVT6YcXeQP1
A3pYwl/Pe+3YHD6Lonw0LYUd9ZXB45ASgZHbHVXvWz3sMQxk2CnU60euOfDKTO5C
kbQnXRiNolKMdxNC+03+L4KYXzpNFMKeb+WPesKlwAK4P0lzmY7YxhoITwoI7I2K
thUDZCgLYPKoySgy8L7Jd758xgWsK1iz2SdtH1LsIFNxKREbQIBBS4eKnQ1SSt8/
NfoaAoTzgizF7Jn9XsQkILSvAsFlWswIKBFQo2bMZT1jME+eUTk1UQELgmfeMQ4A
TJ9YRkbSEMMWg9CPdgeAzNk+IfHSUf+qwyJaJaXzFqMBicpHmfkfzhM1MOvg3tip
C3VucehZdb4UNcWGJgyURMrwm/gOyuhfHLGD8mGg7IKt39dX4zb3NMdh3v4DluOW
2gB3CJkVUI74z7+Liz2rcltLFrZqDMIqNY0ZQUxKQn+LI5kPCUTdRVFh+pFJpvfo
ObrGbJ5T3ShcVwJnQnFI+tUSiWtjHLZTc/a/sF2z7KcDpznMeUySy1T95IzdEGZK
ZmLGjhH4kBfH4y9HI9+8L2Xy+2Chh2P34nvR9AcHx60Mb1eT8LudiOGa01Ms2rmo
/54Pcrx8d6+OsoZj28oPmhqPWGQmcXGnNy/5d9RKdPim6PrOANQKihTaCHgAztZ4
54SWKQ/xO+C3z+DxjpPv2PwFE2USTbfzHToBEgnK7bBwvRmW/OsNSun53akkiLyk
f32LTMWES5RDf4/0fIlQ1knxynVAQmfTxCAAvT3r11DnvZ6KKf2CBwt4qpTEGj/T
TwSLlLEBK9s2QHCYfkoe+/e4hT0u3PxEnSeH9xSG1NTZFfndK+eBmtpFQ0XLWk2v
zEnwwBpWGScAIZAllkhXwVilyEYhz/cckA+DdS4eiazTMkXLrKTuYvReRhb/fiCd
MNF0eIcaEBZelPw4zekEgVi1OmIAAWadvvLBMoI0cU0smann0xz8seKZ/DAiUZmI
QrhlD+gpiNmC7SgoWe1t9m5mg8oG8p6C54ZMjDpJXdyoSEETQhKUyfgaMevTUO5q
hsrZvLKD/+Zj55nh8TPtLTULbYGXR7Ec394JpGeIUDwriPAWHZu5aaKeVqYEaWeD
B7x7LI3opPzb6UMcyWnkwrTSPlE9jgiqtRVeV2m8whWM2ekj/1Z8lwXVGzclwIkf
c2DEAdZAmcvbJeRFu9TTgStgJm9sFT2JpqzR7buxTC+F7T73/fQ2Zivm+4ZDUV1m
Sh3VIbjHG66AewHnivT/zzq17Sh54ErNm6zCzCpsp/2zQ3J1PiY6i+vTWSYSB7w0
VRMVn0Ik0lfE2v3kOnFB7y0h50ForkaM/iqZcw6qxXA9xD1V2m7I1F6H28aoS4GC
Th0otBNrRpNtnQjOUs1+m1niz0NZWr4ORmEJRiYPjqgwSeDW/ff1NwwUsX2+12no
+4yRQHkrg/J+XZbARVqLgL6w7Ox2EicWcUT3zBaVtDX0JEwKs8bO/6pU9y8Oau7F
RLkNKShaFzQ9cjrxwx8M646y0QBASL++g8iFfGoBhR04NBi9RPj+TBHmCrobdy6r
YMBrJXVNBtxcX/vsu+FHNz3CPHIRoWXT7AZqLCmACwdDGwWvZuRAdi/15OnVGkFT
pVK/bXj10BR3KArljSGne1Ih2Ceot+DIYsJbIpsZXL3n9AJnkuXRtcdTzIWswKmG
Ed2W/vTjiV9TloB078FWjVo9c1Nf0kbLfh+YzmoEEu3I+ID+YQtlAdhA8LCGxoTw
3q6sCgUwL/anlgsZU2qhTwnC9w1OYm5tWNJYMhRODtYTxuNmDq81RXw9Q5QV/hrE
QEu0JdAHzMSF+YJ0yHUO/VZhhTLI1npOsaC9GFPqR106ULiiu8NOCpYxeFy1nH3B
HdxmHhChvkfEMQdpPakgNxKS430DQ9RuUCf7um1580/F1ARFMcmzqYL8CpvtuRxV
vGIUccodHToxi9by8ncYDd2JCAnvVaiFcEycVq9jYn2OucXETFRCtZhLQQPwIeY2
J3QW+SsoqjLMAIp7CPfTeYF3PM9BhRaswSl6+kzQs8OR7IKN/2xZAbicOzlrrA65
tbYuv/fsawD0uXTdyZzpH7NvdPoS6EP3t2U9kyyF4uArtGrWgZ2wDAYBl4bU914C
e2PmN2piob7zoSOKH4QopwzVL4ufqK2n+/U5Gvlz5CFg2Yrkopk84sAbCY+MjN94
gK6UJYhDYVNG29YJ6Lxk345YkaWg6CpH3V5rY2yPdYi+zRjQ0QBuitLooWrSeJc7
Pnf5ZmjUdVpKZWbvMtSkv8Ty4ZbrCKwQStHH+mx+vLOv8jKrc1FeKR2qUdZ3fuSx
pPF4eDjDWgeM6sjAriTXjovj6aYAzn4U2f/vPAHLnlFPOMKt7JNu6Xm6z7ne+v4A
FretiitQuqPNHuMvIteFYrRR4yLtHHwPoF4f4bf1746fP2O0wt8aP7MFzIU4jtdx
T9OKO+FnTMF7lG3s9/VhhkDdeX5o9pNF4iVNWKtQOjkiRhzQVwUHgi/+awcxVhSv
JwOvVrSkuucOwQbiAGqs8o+se6kUuFJzFTruqXdUifxHQb0Ki5xuTt82auIPJjOK
5/KMK0+sznGFzYcJxJNyjZJoB1BnPLEKQCu/VjOpTnd64JfBqGzcfuoTneeW6A12
F3Q8F62mF9pRG5D74FZbeYlAkiNLS70/syQqakG3WI0pKAz7gBszkL9Z2O0eOq/W
9Q9QnsJyOGSGMkgLYHmZWssisRGqAGpevuPZjj9wjKQfSsdGj620l+kvnXUfmpBv
utuG6z/xRYyJEQr+5vTkeHNXXETNl5+ZhVipnOJJ8m2PSkb+oyvuOrT80XBl7c0h
vMcCrlmVL44/S4Auc9qE9/7jjh7ybjVmllys0COl3brasq6wkcVQdTT2kufipCzj
YkMdCUqM+v8WxaZEvdQg3JIme3JkUO54Bmzlu6NTj7cWhYOU0Huk0s3djaAvt/fe
GAbAW9zyjoXGppA9+rJDRoJqCI82DzKebip8LrJI6PNudv00O1Qp6m6s+Ex/hWOf
summAK+Mnlie0H7n2NrS+8aBKm8ErpIM2eARK4/qiXatErh2Z6eDHpX8fglWbmLr
RRpjQVZiPmeyAtN+b01UQjkVpyzYN7eoAADksSRNyqi7LCnGDB2mnVYw9b7ls+ub
JX4X3l968fbUCYbH9HwM92Or7SdhGJDXYT/aC5CyYnWbPV5veNdJYSF3wsSa4S2m
uTqnHrKZfo1P45sNMIxboMT/FOJYBprunxwjlgZrw0hnBvUf8eF7xZP8W4K/TyjW
QFh1uEfBRfQwtaMOzjL5Jy27Qy/9HgsvZsDpWQb9KOwLRrHUY1XQgEvMwY7U+3hn
pA8MJCzkgtAEXWL/6nRimS/O0mQcIVPbVICBCOjlqc3OXQHMwFCUVID/hU0Vs5Sd
xAVUC+NBMRCfHKrvN+HagVtK7ihnXT6bFTYkWEbbL70sDELNBx/4n9XkTDXpsH8e
VmJJS7HKSyRa4RIa+sQnNQb77o5jCeq7d13NJAGm1Zuo1tzWXAMsneaTCzSWvgkh
cq3YalVSQC201ge4bplkjqKRBlw/+31xISYpJkG1PnVXzlhjyZvf+R/LqJZRt16r
aDwiudkQ0fJ8x8Iykf8J8kPW5zwGcqlLU9sPtYor4JSbT0Q133m+scMRNkTIBMMz
5MphMNpzBw5ViOCcHS4Q4Twh95w+C2VTxK7tXjwJ/W03SfKOib4KFu4jHKBUJLpI
FeCc8r/nqBGkz9199AhKZtOv43jbHyZNMNl81hVOon5Q+HMkU0W8xqj/jNRjXwGL
qT2Wij/1n7O+v9fIgmTt0vJ2BqR4QmMjN2akZbMSqUo3AoYtXEAtjNozs4VOY0aJ
hrYRXw2J9Fpi4u2Lbaj1iwEO3GtKk+t2ZzJUgX4aNdNeHh+WQoLiJtGzDI/hDHwQ
VMvSwuevZRVGEMrIaFE29VcWzVCVqqd7FJhuzbSe1TGiGMY2eW5wdEKggLJ1PQiy
XzUT//hTAfrayFVxYpKdAjLdKJ55qLJ4DlQlxpUR5kAGL5DGgfF8ROCKoVKVWwzM
mWJelAzv5lE16U5+lLwvtWHE87SkJUiOAWVdhy7AXZLToXI5Zp4LGn1TeYdnljtQ
o5gSG8oXefo+0kf2LeveEOzu6OW2a3bnOZeCmqaxP0YhwsCtsi1nT+/UqvybYGLb
wrVcNHJhmqb1QuE1z6efhqcw0i4sQM06us9m/HEnQD/Wp8k4s7rXN8e7w2pk02OY
FKBfkP1sztipxfgamMslxsnALzpsb42G2nOsTIC8sOOaSZSmHn/70LOJ7in67/Ri
9TlQnfrOwXkdg7D0SUhZx3huQUEfL7U9ni9ia3qB/gNa40w7F0dJJvBL+0xjMyem
QHhhtlaswKhDHUFpsZR3qbIEMyIwkVPARI3LATBSdYcVyZB2mk4AoC481ag0JzsP
hN+IlB6/lOGqeg4uO9DCCP0EXkTXDcochEGTjCS17KzBYjC+sJVstTgFg3XwA9+b
I+dx7lUJ7XcZqAyE6PHTWhHO7z6coo858JNRTNlXkhJCw1/XZAOG7VuJT9pnNl9X
72tn3P2iubv+t78FKytOqb/kMYeAWdiqmbxL37Il4RXvQ+nquTxESCwRV0tojTxf
TotG/Dyf3UXOrKY+MvmO6/wOXoKIE2hizK6jJo7ut8VJjE6kRHBCeHa+mTTHGaj1
Meo+x34Pud5sp8R8isnrHJWlECXcPdZhXvRQQtIqBuvdSTrTmjw9Rtj4hDwK7sis
QyntexpFiE57IpisG2eL4lEix/ppYq/z/6IQls7Pp4kYDEk0Vp2nlh2H40m8ekx5
XmLT4crxGnlRYuDqWYfDBT2wTJy96oXUBCSVFqZdayZ9mVZUqOhIhSFVhCx42jFe
6lQVq+Z6Bn+4bIhNjOYbfdWWmP7CNL9C5W7Ggk+n4V1zKXZiL0jgOWBgHXaf70il
E76CAP1v5DmKRZTfvpbSDtNBKhnq7jkkbXW6KxC9HPNIYKGhrBUawb9UU/KdeFxu
cjF0AQ/SsrNXbTFHM/GgGM1QjNtJlNogz3AqjcNMVHhrv2DxgNWQWCu0nfS43kqD
ja126+lPfoJqdweem5z2NOBYj8VNAdN+I1H809W971S0ajbisR2YiIktGSuVXn8T
bK0CBaFZv/eTlxcHD5DmpJFJTt4zsf1fmmHXIMxdB/megQLTVaCqv7pDas+51r+B
hwhModD5Vpjy4j55FhGsYgI5+47zeFTN01duvrnlGkpY6FKVmU9PqThwLfQFWiWe
tFnVa+rc5PvigEaW49+oGufrJRwiH8N1faoemup8G/1BkEm9OOWnasYcj3Vx7fF+
5jV/y+FgtoiFkCViQ0ehM6eCyVcQ/EBImX6UT/SU67mCHIbXTLJfXNBcuJn/A1mC
gsvYz7Qni4RBm1nbpj5mZf/GefQi5pF8CN0UPnQaJoBc4uKVrgdBaZfpSbKRG6Ui
RFYd6IC+0I2O/XflUN7/fDDG8zMbKGX+P2qKKCv6Iv8rWJuQ4ob33075EVNknNOE
n+fZuQyUdy82WzKuKI+/Piy5AmWZohSLcy+Y0sLswi3/KSiDHGa6xYnokp92eHXO
uKxNCHwsdQkvcxPZdL2ocHjd1NyRgbLpXffFNzl1k2dRy3RdVkqx5rWyjEW3Waks
zRF9JY+Tpc9WEUivB2n82get92ujrDEdzeqHA7Fuv2o3cfnwFS7gY7yzEX/q3LFm
yHELnyWRc8FYmzLuwlwAWY7p3t1Ao6U+4JQoFWHnR9wQKT+KJ7j4eCxaOMvqpr6v
BiR1O8JEpH/gUIjfRommL7ZJLOXe8joaQmspZueQcJxIJzmRyr/t6O5elH4Guk0S
mkwD0tx+9I1q82l7ayr5vjKA5ZClS9xpBjk1VTbsebAM+RHaXQhpMXEGN3mR4/Qm
LO29/k7dMW+vAcDjcK+MF8L8Auk7+7vlv3dAQUrJffAnbNNJMMKvyi8vAjeZ6j67
r6GDI9rs2BCfWIKuDVRFfBCkocIFn0RwXr4/+tbir6xdAT9uouj+o1dm4iOzpQpl
YPxW2i715FEkO2EzgIfdPyfeUPlUfuh+bZOKjkeThGioqal7c2vmIZSFS+BfDFsX
3VHi0MP71NOHprhVxz4h461gmwKEhqMHyN17wWLqel657VEgH53/G+zKfhm9BiuH
+EGJL5AhqQySKCWXNOn/xgcFrvWEVRRE+rZEWlVSmWU6OGD/7y1wjTp+vRrmD7im
fHu0ymUSdiymbDUUd/P60X5XlymaaPqWL3KxH2f2wGddTNphWOnHfArGlCmyusCP
JNFMImZbzagDraKna/ARN3wKQRNeEfPfA4eLbC7VNA8ODV57BC+dhQh22FKuaXNN
22GciIwsmp2Qi3sCF8uARnzEsv11K3tEJhaYVsbFO5AMcii8HNqfCmx0502UKwEJ
l3pwGBFGGSLQR27u9kwPE0TiqehC9FC3GBXJLqyqwD3diHf3m1NtHfGSYLRkLq+C
C5gjSRPdDDq3d/vEhh6GFo4Biz/3V7TF5IH11y2F7ZFVTUgJlFuK1Kwbr34R3QOw
wgjXEXdZ38eTdPVM7LHelffqYsp4jm9usMwy4E+6XskFzyQtB14cR68IIqsjXYx4
Nly96BG93GlYNa4n+2nyAqAumN+cM1tfvGh0gKPMx6W81mgpPL1qYYGuzUzBUXfL
jTQx4CDuEjUYIA0itKeArbvUSWiW6eXMiFuiYV5GsBcmD9+TsM4mzBYXR3K+gZpZ
NNL7nbrSxfx0/u2MgdktnzMwHiVJ6CE1EvXVyU3EEPOeqwDy2CVlJz3TzC8ij85V
6yxsUqKyX35Y1KaQTqHXizRaa0EODOXbhVRlCDD3EesCJQ1ZuGdpgqQ6GJdKQ88f
eASFyBKA7HGCFdvDkvQzPXo0vrE/a6wWnP3EadaOgQBQHYeyI7OnXnIHpCp3J0q6
Ssv/bIwWNjiLfn2JuRrxi5pgmHLKxB9gZBUnr++NqE9ykMqHzefLYNzljjQU23EK
hMxyDnWaFFeFsTKbn0UkpjTwev5LKPMH0Cuvwu1XEIxQ6X65h1nl38/5XF+smfyN
ZtCCbEh4pd9RmRlMgKisNkyCXLCVQH0nh9pfxaEKy8cYKZe+uk78ELV02UElV969
WwZsqrK9mU0GBn2zVNRSLPaPRRWcXtmjuLVC1y+awxZ2hV3/NEwKkan3Y/OqZqFq
qFCFdch4kZjNLIPOc7MBG1QGuyi+/Ngq15ob2SlShqYCjiu3TIE1dEdZOmZXqATC
IvEsCeM8I1KHTYgVwvQPVatXoyH77Rjh93L1/7ztvQa+wZZgnMVVS7ctfuaCsmli
nWR4yYv4dOm19U9HYZXydnR8MxKljtE2fFEP60G6rITGasKBL7IZ+bqfQTYmqTWg
n/hiG3NqNg6GU/l+KMsFoLxBrcT9QjykGGeiJSQ/hzDUBH0QJ0EcOXJtBY1/UUnq
nFTzEMS681MIhsar9W/o+ThcrW7h5YJbw8UaaGQmIqSzFtOyP3WA+5EBxbz0E6KE
YfT9dmYCajjTXIOMcvwI3ftwWIEFqUBxMW0hTrovRqWnAjJwfLtLuA0yO6JYTji8
AbYgZRQ/2J7sFyPOEolrcBt4K+sLwaQTaZyll++KoxwdiujI+ABAsMipk6RnVfFb
aRrANXkyAssiEtLRmlN1FGrOaB81XUCQW7jguX1sHBWvq5DvYjFdr2VXGcCpKlI7
9qfYgX7z8t8TjRZVEFwelRjH12EoCxatsh+cC8UbrCFUNy0cZyaOm69WVlmv38F9
ZmJiP7nihD8Sya4BCQR2ZoQngoDmgPRz/1H8viyS1GlO56WWbDdi+LU9KbS7eM8P
2+S1IxNqHy7U8WUEcscQnfcVFKBjDxSgMkKS7MOjJUkNOL9o0OuMfkiyZf+QTVQ3
9dTnM1dHXNxmJ20Ez5PUaVnIgXL15klGbfKRulMlosAiYDuwCeQLVhDB2GADunn0
yKuM97wRooJIUtxlfwq6rKEAX79YtGZzG6e2yrTLpJpRbbLBvOBwwpJOcuWywEDD
g7vPncin92xKDr7vhCJE20Q1jBd8tlMfSWJ64rWYU44G85YiigGcQx3VpeWR4yKY
9q08DaIEA3VFznfvMEfM9qlKM6B+b7pcxt5ZyH6iArJdIClhYVGdGiVlFfFDB6YY
dDTKcTeNjErxdY2sh5ortczFTsLYIrHbdXdcpHptbXnKgAH9mPKtPq6YRzPxqaVw
mSqSPmFlXbiJi+MUStSOPBoTQZ/qQI3Bc1LLwGTX+Cqmlcaf/nnrrKWGReYDNmiz
F5p0CzA5ldpLQsjWapx9NQeuJ3GuPegvULH8StBFRRyxPjyY9nbR0v+/gMunc+kc
1HXPYEz9gAiubmhTpcGQHFE+P1KxIoI/frUbEU7tSJiXX8U/zNJISxKBT4Z/BCmQ
MwdKX9BA6Vow5az1jTn4dS9yD/vTpBbVFEmkGcnZkpxMDdHz/SIKUs3A08pwI8VJ
Ey9AMi5Cyyw9Run3H9zxU8SV1zgOvFiuICe00KzIIpS3UPsQd82JalFWkwEtggfE
ApukaS5JtxtCl6ydBhuwCfMULuun1xF/vIE60LrK7rkoMou4VeAbJNazS7I7PtGJ
PFiHJsH9O1Vg7+JLRnY2VDvyfVcAiZc/X2rrn9qow7s8qdZfiqqEPOg85WF6HTIX
iGd+8lOAjnuCCj02Zyg6jAu81QllUg6t89EivJ2csZ6S6wvSW7Q/2d/6MfS59+cu
xZHVr0vJHMIPCz9zPgPkjjEGwVbKl1kbCmgvT59BMdNxU8Jjo491PNXNOGhJwuaQ
FuAkQdSfmydus4Hv+RIu3E05QAfcrj+iHDzyne53Q2x81Rl2h7QtzaCUhiAPWz7R
HVf2C4tSLXucSlMRvuJ67pQplADtW0lDgl66XDUGvzv96U+1Jcd4nB3o/J916I1r
RG9S/PSYGu5tr6JO6S2GE22GnQ3y9hChXyOcFhB4mWppjoA/Xetc86sVKfimKYnV
J+f6Rver/waVEPq91qcYZPKnJFPf6QNRH9dPkwoiXNZzjuZipW5xGAclJn0+R7/1
lNpL0zGeTxMWx+J6L1uOsoA6Z160wE7Tm3P26hnWpfN6RuZC6p1bi7xnH28CnfMS
0lrfXBDOQVmIXHdOLGEV99NLeflY61SZnHX73TjIUB4Uh0vmJcD4JL7mpNUsVMQa
cegMIX5HM8y9i0uxesoEon/UXUJ7lkPEx+6BMcRIJn+5AUqK4kzoPEvzhqFI2fl9
HToplflcTgVyTiWJWlcSwVH+cQaAlozGldOsNQMfVH3ncOt7rnRC9a79Aj0UOU36
unb4keQhXFGvA3INU4PRQUW2aF1FjrHHAcSrgO6KjDK9+Mrv9TkkJF8PuSJ0kXH7
PNnJIPZ8bo1WtxxYT4r6/d6zTTMG9w0Ss8tm0zyoO0gWihshFtX4/Igx5eSzmvJi
2lckZpDeytimL7iyNDLPIXOB7Dbxy/hn4CdQHUQ6YClbPSwTpJ2bNBy/+B5ssO1k
vn9x4PGattEwO6VziZwmvTNoYpfuy8mg5W49RFXyDiVlNr+h7onz5goK+srpi3u0
mV2LCAOoVWG4BTrm3tsc+i/jD6QGirNamQtGuynTJA79WkSEHNyZ50zaudI944/C
Yy9UQK3pobFE5eu9IT176VZqnerXKU0FolxB9KwGqWXjFZyeMOOd6K8lbUs/OEps
ChUMzdTp5kCxGgrU/jXK3uxx4WnyaLO82q/+KyjdXB0PwPipHR628n34FIm5Cl2U
yanH0AsATZio3WC9p8KJy3rp6ib/pQCv/ydq5Smzipct9Meg6pU/u1LVN/MMvqiv
yssV2uZubuHczr1it+E/OdxgXh1LXOL1k4xuprkk1TtcoNz8m/RwksmgbtUJ0Qdo
DlpeZYgSDPYfWHhiWpLyUSLB1lYdrXJsedOk8aG+/IgX3GfxdXCpoFz4VtPN9f9R
NIYwN9n8blYzESoNqjYQbzHTiy2OaDJm09q1m419MDYsegW8QlR0RddCMCBehmTr
qPjVOtCLrd2txnpZxA00iz+PA4Xl9a7t7Tdq05aBhqSTqQRGPpdTmwqZrux2aw1a
EkaCVb8IputGoK8F+QZPxXy4ifeJor81nfr02pnhtmpciPWuOahJB1+15sOT/qby
+2MU995EF/FymmQtF5/+pmHKxvD1JloO8P9IaE64trcD66A8ISvaOM0/Oi5BUy6Y
YBuV112l0I6pU/0Wh+PfUmzf8T0oJCks52a/GupYSGi0EwjgN5qDNp+ScpARLv71
7AMNNd8tPgpWcOHmLB9fZDdovDV3A0lnXgAQTEstFgKZezLFy1pPr9ymR5lu3/c/
4HQS2B7q3EBaxsfYCiaCWWWW7rvtu88ir0UI4w73JbHljXsbuP1p1Vghaksc9heZ
C3fI8mpO5ZSk06tiDGqjtDRLP7RazLBwdXygiSINHQeshCMjWd/mvk5RPFSjomDT
r5QxhQs9dpFRTkKEt5lb3Pjf8rUH02vp3TJ4txADzHRl7Oc2+QsrpFHx2Ttd/VYA
/AW1YU+pY8MMBQWfJEgupcLDLm+7eLHRNIfrBPqeZcOccIEx0w4ybb402P8wZi0n
SBMqU9c6sNHxEHeKC19HDy0vV3OFTYRD+kyeqZ3aoLpiKwevfDSILPkYwlcdmkZZ
1752plT+dRXwjVYs2UnrdjSNHcTHaLiDlpB/OeGOWnC4GGMNqqsMcjicIMJqMKQW
yUxIvlXeBFLMPufKzIQnbXSzgLIsSmaOuzb+aJQV3BKujaAI6PSVzTA6/cpap3cd
G2+ykzT0oeiGMqDDrXDNlRx3uEAMZ5WtB++qcP5SE9K/08DdEm2hgKgw5kTwUh/c
WI6l0JXisEJxMHHt2E8HeslrtJZR3V0Ohq5HMrNUwjrf+uILJFD2wUm3ACCoOoax
kYguJEdLXXWyoYtE/qEIA5tSht61+Nap65nifXGD51sYGWllq1J/+lUwR3xG5T5y
20WadVACoBEMtyf9z7MCI7iFFSRQni56hIa+IV7TrYHD4Keu+eNi1koDywtEJ/6O
jnRW3wqMDlcIG0Uje7dcz/PSejjk2mavl1o1LrN+pdqsO54vxUk0vws9k635n+QA
V7aEXcQvkSd7R8CqMxbbged78IGHUGWOIAO2x61TgdW9vBQwjnPN0q7FDWblWsqX
4xcB9J0G+hvPg3Dt3Kc3XyXqloC8812KJdM1m5RMWin64JIN9dwM67tAP/sGr1k7
GZ5u3jtb3FZGLj9bsIyPqOqnJZk/QMQovWTGJtigsez0fRcxOczmOKY8AVRiaEJO
lFq+gNRiI5ZVM7qujXt34vUA9fwDerXZx2It7B9g8H9FIZmP6rNG+PWxCfE8Rk5M
uhUpvEBnfantbketzB75UdrojKIe7GGl1hPCzNmcrJBFSVVqxtofoJz/emPWj/QP
Fn21weyN3RpU3tNfOh7z7Gxd4P6rzJhhz5NsByQAwDxFo44pzL9nORmUrCH3ZmNj
faE9XyY/IqLaFzSSe5KRSnIjsws4xEnOOlxXjhSOmOTz5pBm5K+vDJEEOO8o/nDc
kZVu0we65D7kcB0p8zZQRtEQOkIrCbrR/okaSRAgzSfCYRbAZtPgPQEF798+/in4
GoF0x43tr79H5+uLIF6LTfa2uTP70RlXU6fwglCMnV6j/kOskR191GOpVpabvj2+
WQzOOhg11oUIFRxLI1esff5uNU/KqYrpkhudGrFj0dsf/G02De2ugz8uH4Lqyxz5
VNbAHGa5Prn+P2foYEEiBP0xanbEruG8NR+eqrsXQ611nYDNecP/t0BVrMh7xceE
5fHxK7HT2TQsn62O8SqDFERSXx/VENvEmkWKWSBRZx29jWsMJHodDcm1wreYpFvL
0N0NP++Rv615oxzqMSUB3VKnzNzWaPBE8GmpV+MJE9pjgUqN+TQCpX7cVfb5f4Vp
Dg+xlSFGvUF9+RVhH7vgI7I7ngQ2nVNIJX8+07ZLs0T61Y4bQ19C8eD6XyGUoKcY
7CvshG2O9OtEZnm9TlUPyY4LvapBgNwh+u53oup0gMqq6p8wltvUiEDFyAwhT3vz
tUTydHmRcvrWk4BE4vGDbJ1wkxYfXiEm+M248Q3BDy51P1iH0y5UVA49k9ayOExn
o6siH7Y5yfXvoN1PjY45juRZqFAj67xRNLudD2gNGfrPRqRFowVBU1mJYsyUo5l2
XZNV0EHqC/7d2vspvlLsNdjBRG8lBG/J9tCBpgVYXWOFniTdju1G66VgBqk0b2ww
RrCUT8MjekxhnPtmJ7apS7sNjgmco1AiaQ4NPUbI/mK8gG/iseLb9b88fNgyWfqA
pMzpk1bmR2k3SW+fIg5cY8ZGjTeJXjiq/U35vW7z+PsG3rPUzG6jerl0ksxiZ88Z
qFAGe3TJDcPxzP9MkL9iu0KoyxfP5Ub7EWscvoIx06GzSg3qyIGOz3xlZadDprGU
BywVarcE8FO3URPC8ejfpv/euLYvT0M++nRbSRucsMz8E2+2Ddxa9pZ1cQdEVApf
jYVgLC9sLO5hTQ2WuNS+4Gwp2Yq9QLDgFGBYZ/yN+VKdQOCXYppm6ZOGhrxUBogG
Uw3wxQ1sNWTC91ap7PO4evrpJTx8DtNvFlNhhY8pZTFFamI4tPh1Jc8oUoTM0Pmi
MPVn151Ksxm+6dN6zwCUkj+nBJGJ8EnEgxm5AoiePpna6YbVsFxcBqePJj+9YrtS
4SxVbYTRxBHdD9YysANqDbYevFCoNxSSfrJHecW6oLiCVsBgzoSC7fR+n7jjPZPM
CYRQVDvSnJ+uK4jMhMdkH5sbOUheXlAJf3R4zXSa9NcGDlRjvmUhtrUftsKe4KI5
5JZSaXJXhYa/Kf4Hk9lV6GehDg2ztXMTEKDJgNlD+h22x3jkLWWLrFt3wby2t+k2
7n7jur66yswIgoe60DqxLoSrLPaFZvHMKv8x4X7ABic3t8TZseYh6FbL02Euzseq
BahE2LsgE/Pa4OEaBRAdX7vRZBzAIjIAgi9q4FM9jomR7lVFLb9aDJdINRC/1HMq
y/AWeFjZpXTpl0IY4P/ULvsBsEtPLbWyM60wUPS91n8OcMCoEVteAHOzVCwoD+9+
yQixdwvnkUKPcPMnNxszDfQodqd8MzRMobU4OiRJyeiqCdgV4xZzNv8Z0DhXP/27
8e3PL5ZmRvYgV8iVMwUYSGkkGog2NvSPqRdRSE6k1STYCzbxnN0vx5BV0JMXtRUf
GeYW914qcow6Y/6JK26IkkKb78cDyQ1MHanAnQ8+qwGqDAP+n8Mv3xCFW24L6k7U
I4quERvYgw1mBzVpIYI47etvKfN9/Y+otJ5u+ctUrbEBBIbgO6BkZgzOLorNJKQP
LCCmVtVxz44frcdWJisJ5EdvbtB+28NqjQoviT0924E7LuXNqracgbx+brQbdLJT
NG+9wC16gAtp+lcPx62Mz/DAJJ7q6nGco4U+WyB/Wao9CRC/VHCUWJarlb+G3W0d
h6g6HvdYQSJKuP0lohch+iGVvCS56dqaMoZLfhHvABWtBoAvbuk27ZGak+zLjrFd
TTt+FyST/ZL+d15QranCr2iTRZUPNLWjT8EdmfLkQsSBTJmrrIUTcalZkrLo4DTp
yZeaENbwGkLCTrErDl5BCqFSvfxs9NSury8kEWs3LzpAX0HBEULksYJKYHz2kuO4
gubETag/3IVw0wIhcOnb39cuDu07ASdTcVSgsT22bkqtRmbStJCLTLjxU/0F72/F
UT8G8S5MhXJ+Xq4cq4Y0pEpryU572tvVg7pbsIIwUqCBXqBCT28xuuzpok4OtO6r
RljEk/b5EAbpxU7qjPBfTQEAE5pJk+C+WDlU4uzYUrnlvyQHQPUlKzZdOBc0bf+N
aUuR4C9cIkzJTczV6DmiIs0yhi5QKQPh2J4ebCWPPEpZZj7SS8ETs4MG05URMNaV
ClqYAwQ6jtL4dasx3HW0MIDe/KMGOxbBg0Hp988rJ0/fwUASpLhcbQyiP2x0n/Pw
ytXYX23O4TN790Xp4xP2GxS+U5sUAjAoAm/etkAYTN8+N7WKQKgV/IQGvCVgwsuY
lfl5rojMOWjdHwRfQ9LQlhqm1f+QzsTVeOiOydNL/7CKEhXsl3cpcsZ5j1tAVefc
eoYG8kUrDx3DOubUAFNdDohq490VZRuW5bN97QVJH/VS3MpMKQi5hpyaSISxsABB
3hks9W0eV4DasR66CDQhLPSYy9C77n924yOAiScSm19Wl+h8g82AtZQAgY8NO1xz
q8zWSFmMVt+he4gpKTmFAdnXmKH6V6rFqrwVVXKAHdKMgDPV2et/HiqGOMoVf9TT
L7rKvnn6GEtKNUBQ0RJGFAaAAIpCuGbibvCvZecz+ptWYuhWY2mmewfBzIuvLVuG
YeldQ/iJzf3XoSSYYzfBcaBYtOI0nHPOmW8OXxoBjFELh/k9EYwWns0owSdQAIX0
rwN3+Dapvse+zjqH8DX41NN0pa/2Y9JhvEV9dLhrBaBHghfrQ0WrJ9CEwcTy9ran
Wp7freYr7RsUNeFwJVaODW7lnuCzeOSBAuN3Tycej1qCnaJuX8HcrD5dBc6tGc/p
ssJiOekTm2V+izbrrgMlRvG5wvvePLZf2igFYdmrtJSTtIEZivnUWBlKzwA+OGwO
hrsPoo6aeUvRHLwb0gNqGdjOKmv3mJj3tOD0WRf6sntYCoerRVSFJPfxCiKCdx51
V+RGofh5CA1wAAJsd3T5JjUkGiWWZFGCghhMZOvMFGUWsExXbQdKod21jI7VfOJU
byraERCyNA8GxTo3QeSXyiJIqLE2CgQ+UWzWU56rOV581a5QEjgn4buuSa0U6whm
NxkbpipjKqMmo82A4AVOIIKJea+01pfka/g7ZAAdER0Tpa6FpNlil3z8OzDEkbmf
acr4bHu3pDb3vpEZP9b2jdyAiSyblg2Rtbvls79/+YlQzTc/OLWwEO8q9JWj77Nj
rnwvezXXhuzDhpaTy7auDeC4NPD8raEnzCxPe2llYkn/WxAeKnKqCdZOZePi7dL+
I/JLSLSxR/DrNk9WjJXxAF0J/wjOlinZThhPGlHtJWZeslcNCMF+Bau5sC+mC+nl
s+3pYyyNJqFAQJ3wCGU3HZ4cu4KC2THRpdPThPzYHNJ6dXO1PMlY3DAKM0m+pePf
cb7kiAvgZkiksGSxLQ9MH8dEILI9S27BkWAxmvLh8kdBY8/feJZwasOhxoCUTDWA
fCs3MvlI6TpDOxvRkCK9iSz+5EwXnVjIDN7012+xXhuMm8B/HXKvV2Osqg2nN7k3
lSjBhgm03Gj+gVPHFzTJ0wRZn3o+o0+8/xFXXJ9GjX4504hORF7sIE1HdvJj9Y7J
0ETE6lm6FFlNR6EgE5yHItC6dhaMCqeK8dwACCi6Y+CTljW79Z2J1oVoMkvOcaI7
iyruinP5mqYxTH1WrFnhF+C1DB0ETFW17OojS1Mno2ddFGMjwRWmErz+3ylNYUQM
RuPZzJR2R8o14BWnBKWUKIwumeea1KyL3/bJmixPFnZQFj9pq3hzlsA3YBSrytOf
i46f0FO/H+4EgfmgIs1KhoKG92B/Ld5q8NTUVuo0bdGajBQG9cQpXBP/qWrOa818
E3c3wUPw4/goxdNF6wMbLxgcyUXE94TrQXR3rGir3tNTYJEv80uAhZyASssDXwf/
2Eqz9ilq3Vt3jat1qtCpaNqb/aLtdd49yh08yto7vG8yc8TbToMwjVityXt2d3nz
ynNJm6osUjc7wsJKw79FCQnpkm1T3oa70CObhfNCRYn/evp1W/xOtaQKxbYm/80J
AOfPT5skdzyKDr2HO36k5Ovbj/jZ3omMTXm6vh5HjXrDgN+FnxzkrLMbOQGmxMQC
jikyVa5fpFEcS852MQRr4/BbHB0W25U1SpWyapx9XzDYad+Iy5w0SsUMV/y94QtG
/v69fNvuKdL6YEeJD4inKGBY9HrE82bNXAJnds+7xssZS7B4zLWCNF2dSRNQuvOh
k/9RUwv2dssSBaWOSspIrsl1PnlhKemAU6SPX/dBBv9jtJDxl0RIitol/9PUkkIs
TcmnmikrfZeewp/aaxunFVvRXJA0OIB7SrYQE9uY7mvFR9nZcP5RiNNMTN8jZVFO
aIDE6NdGwL+NxX34DbKW/TVCyPaa+fWOQ6fEryKs+JPzQ528/Uxp4ULKECJFHIOs
2laItgJYqEzqU5xIlsOdmqq5DRVwzs1xZhhMs394a/wZ+llxFUS7wIXOr8H62WR9
YiuYXgzSGfiEnflQzsnMrrSae7BoVnJyAJGdKmK8irjSzYIyadxvPLSXRySkrH/W
43psG7VBA2V5DBMhBtNrSGb9KTh7Ky/bdO+TKbKweENkFTKB1xRMUNscC0tG8fBR
hXTkHk0w4ucSp6LNu9+NuqBEB/UTH7qq7zqC0ppIImhnWQgmbVB9db8FU5fH2LT3
5geV3tjShL0ILZdeFAaWqnkZtnjAP9QQRTJoFJFOQslrdZVWw2rEayDY5elLawta
0iYQriGgGqBLXz3mSbqEHAz0QzMVi8wLI5fgvQPYqc2GOCDZ0rtBg1Z0yvk8p+U1
dM5SLKpZg8w0D1ANfN9CTiPQBlGVRI6kKaFsoi/Kvk0Um88TBF6EeYkkPNXTVsVw
zHntHB4/MGl/fsHxcHmIV1/guIR7xKpFCRryvd/bqSVXSj3TZjWsxgthGK/3/yN8
Cub/8vLNhNOd8QhQX8ZuzPiK48hRVTxKBPLezwgmB/czKi1qaGAHqYiYUkrT4I5J
s8P9io57qM8M8gWM7vI21iJCRMSL/XcF8GQAXq4y/Nv92xH0BjCmr14RGMhTwbQe
+vUdfYvtrA68oSirs4K7MELDbmPVS3KJQ/02A8clD8XUSIsQbA1GHjoy4bThrkqB
K2p/sUxjZ+DP5tyN2DJ+OFrTAU+auTVW/TY/KdZqK+Iiq4TiyirqfZo3dUbr6NO4
wvin0gLJ4X+aR6VPtjbhUePbQowr9MRAjdJ8DNxtO+JGmqniBHRVsW89nW6mGjFb
iXJSiGBZjjAUQ792K8rqHItbU+H1nxijHel91OQm+LIFFXqtLNZluarfkmpNrfL8
PWUfwBNk9PKUTZE79sFdKyEh+8cQuLUsEBX2Ox877husjvi4JGeegEhF5fqxD2AC
yW2DE/rotn8VtuZe+6iWM7uRumWLqlP6B/RdUrWrjlvwVYykJsLK2S3wKEbetHKQ
CD46+WfJehh/TGU61SbTwavYlIzQEzCYvwWzUacpIbI+ZHXPWBXMGUX2/ouPIS9/
6o7ZZHocX1LuL/khAA358X7SvR30Pdm5/L/h8KKLpwF7sq4d5WvkQmENyD3K5d35
0+l2M5Oo5WGGScuQGAHjhcns30buOnuNPptA+tG3aiS6fls1znPhv76LbG4/jrC8
J9JtX1CKonAtbklzH10Wbq1K/dc8Xd1rAAxw+y9FYtZRj1gQTofQpKOWRilN+Q5I
aOCbu4q3Dud/fs6GN/V9UjX9xQ2e5hX0vU4jeZH7s66Rkvoh9/a/I0tu53xjWFwb
Oh0sTMk2rveV4KlsNhLxIOQWJXnPef6GkSVBSS/iqU9nh2Je3MHA+28VyTbgpO7M
O8fGCf46/D0eD3ppVkRLnfH4/nevmdHI0HHYuUtcv/l2mpOEVpYxqIorh5untmrq
vOFROK3oWepLWWvqaumGgdzNg5eqZ1NrqMUkfMh/thgIh8mPqeE+x0DJ4k6pZkZi
ioE2hHbNejoXsyd03wtXXRPiE+IelTAPN/XxtaxLnLuNM6ZdfY2/lrPsNbLdaY1B
Os014mxs+X4D9UhIb4PGvlMRytSxpOTIWuGJ4Ietm1rZnRgRFSeGH8rYxwExelVz
XFci+e94OJTJ9ohmblqZYC94vrOBcMTOAQJDdT197MGa+y+QKvvm4v+iR+dETPRa
INRPaMb4tLsfl3fgEhmHx9Vul2PoWNCvJ63igfmf26FKjjDMtpvJGt52SwCiSdT4
jY9vU13JkU7xXq8AMecBbhfhZSfN8A0PRkV7NKqGvhnfEXiFCxFSs+r4s6LtWuDP
4Eh93O/CbuXLha80+fhHkcy7dUFXlxW/0ic0nZKosc9u2far28p/4ngXAQgwZl9u
IQzP9MgEZU6FdKNzcFojW/4mBiFuBAII/CcN6Op3lpY+rJ1iMgg6uBsl8QKKPe6I
zSt4yxoYYSYooimHam/I+v5DH+/cnG/qpp+M2cpksNVXYpsn8pe1yggobVThmzmV
E/6fct9iXlXi5Qlbd8S4WE4MVqJdW9TljJhNhjuc+U/aOi1kfg0rabLi5oElv60w
bWTS2b533lPK9ZFVq+8yayykO2GUAFt/Sn2gDYoVZwPsnfm8rgflK54kJ+rGVhKr
gi+7nZQ0YH/ZttBDkJcusyAHQ0b9+BITbcnqWttY67EaD48Wfe2gYIUVW72CugbS
`pragma protect end_protected
