// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
DyNxSjVFSZU3JOb0CJYp5ATGSCeHOvBimTDymxmOd9Ii8pwu4dQwp5bbHELhlE/m4quwY9doLSN4
yfGJyKksiU4goNQvfu3VeT1SXcoWJYm17n9VNbfU0J++sGOERE7eMfdf4A08hsu4guFX36d9uqMV
ClewbjJKrx4E3KGE5K8V3Zff3HTw5WqAOTXXcmT6whIOTpULv2ouecN9pbLZZ8Q3q27/77hLs3wY
7nssKbDCGQ09tQF6IrvvcyraS0CsElfOJGtRB95iP/luqIHt+WY+NLifk+MNDB3LbgEgn/OfSuWw
cr8/lC2tNqCELdCRyUBBe0jTc4jMiZMTxuq2NA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4944)
8p4nEUePG/4s0f9AlAZJYsS4Qfaq3UrIs3SQwUBb7vCtaNf25oZW62yK8Uo7cfzHYpDAtO1rWu0U
v+QWdbtQSMNUkHOFCd0uccVdQYzQo5j2ktOcDZn5TPlWopPr1SsjvqtAgbVH+KLufWB051j6byrs
ELqfMR9pHYYhi59fzftOzJO4D4dwqpge5v4H01CcJOQu9jmFqsB0Gh2YesC7w0pmtrmsZrORgryc
xANuozjIsrAIfmUc3bNjrNDyvbv1oSX1/5sbTdxOCLmMvRWP39LmQ5ikVIZ2D59ubLe6MEeaLc57
Qlujbp0pHntdHGGHYtoJzUygq3BfMY9VvfZX8Y3V03cLx+HKjmpRaQimmm1TmfXH1pbAGP7SbXSy
YTITAlpRKVl8yOoxA5RqJFbQNyHW3I2AzE4uvVGh3Uha/u0SS+oWns+6ZjqPIP9yfDVKl0N8+loc
NqLhwHI69c6fVgxBEVG/CpzcCJZBoD6uX1+iTdJ7yFQ0X/qE6G3I0Tb6WFeZDUIF/3FTMA6Mvmvo
5njF9QxPjqcIoXKMSvH4YvYKiBNzaS9mWLZBYx/5GhfCpWH9kE495cGobxEF7rhsfs5z6qbrwKjl
wh5vEkuLahzE6Nm6vBlYjpjbvWKOJW1g1jMnu+UuRX2aFGDnlHaG50PIbg5+MMhJfTn/z0Eu9sl9
LEWMPxxslCtqn6KSc7jKC2qYWQyLv+T45PD365SIDT9iIG1qLii9t1K4xRBadI4U4qXPY2fPPwvT
gveB0CGvkRHrwgT/nnTUwR5vwZpvKqzcvzVkm1aySQ0bOTP8+p2/wi68rF6zdMZ2wP5/IBwerJuu
cGUS9aJ6wEAzKoWXY4j6lLKisnbpfbXax3XbBmaL1KosD2978DLzabyR6QAP+6szgAImuZgTXQF4
eaIHC06V7k/Wpa4+/s6rebM+UPk3NxzgoBs5HfysBNJnJHo5XBidfG8o54KbgzohtQuuEKH+6VUP
bLB5UT3580TCpaeClyGMqXLuU1zI97DSE97slgMDZ4Sbq79IKd0purDe/Nz50oOU4CM0qsTRni/s
Q4xeAeMlO0MICyyiR5GLWIR8xqFXTWAxAlr2QyIKtpojJoiyYAC0gAqIj0Em7IZrZUgktxMd0/hF
EVfMBPunt08L0BbAOFgYdqWEHSqv84oU0qWk4QGOFI+/+imsvr3RZe8+tVL05S8nImFc01yXoRUs
jdyYhNtJHwnI4eaz0nWX1UAjcTI9ITBPHlCt9GR3AQ59PIsPCo+dCvExZawJYu5Ilk8Ox/S91k0S
8Rd/zb8EQnXLMnt9bFLfskLcjBCYgzWP+604soY9HKCMUeDDiV6d+piJfFeGU1E1NhKWfJE3SkWR
nTG0EKjADXCP4XK2EJseZD1DF7h8y/+jTr199ZiMgr5ikqmkO9xqM06InlttIqk+A2uWAyjwTrsr
wxYoUXNC11E9G2BXFFPX2Q7RTEy7ZolG/XQR/6XkD656nXmL4WiBl+153tnds5k44RMDLKwblo2C
wiiwEnYdurJjMm9ZbEd54ODuzZN57hcmQKVmu2Xs3xqkHBu5xDHzp0Z3fJmKXK56blskAQ8NuKtZ
BZ863tDHVFdfo3bdNM0Cn07iv/tryqr281N1Lx6JQ/LerlpQ6DFv4lboqhj8HgfQRzj5ae89ZzpV
22lvaf/SWNwkBGYtyII1iwtyzAYjl4uB8iVJ6ZkhogHKpvvWWV6JSAnmLf+JiMe+elZiFYJ0EGpX
dx9UvBcsoz5xp0uM8BAwhMh9BEF4qWtO7BMwh4qkJGtTiO36BRWokYP8WiP8AckwFUe7B/JXQFcc
Ymmp/ebvWWyj8IfXXJfc/aWfS05rr/OY5ox7KoKsmYuBVEjbkIK2Qssw85tY3kww4cQ5Yf5TXCvp
SiI6V6DUeap5elBVXFPVTkYjvHKyMkoN5n7h0OcgS2AA8z5tWyG1ZHp1FQ0q1Vg3b8/uZiISJG1D
13zrXVMhScRzJISF/xsVhlC+Zb6zmwzr0wQgcXdhIWvaEj9nNVJkVLnwf8m/78qC8tG7dk9wCj6+
hlKE6QOk0p5TQp/ZZFwbUOzz0pQ5hFOlw+kFHx/KBop/314dgyPmonHcFJyhMmRRHj3BCfWnaH7S
0bnla+tGqpA8P/9hF8EG0va2Kcqq1aiB8xRl1vroENdvOD+XnqGqQKiU3AsnQuAzq5PVry+aZWTc
hydIhAKq6/0nvVVERKXZquWhDhN0V4Wp422zcS68AD5TDfmJCiomD8eNrEx+137bTY10ayjjtqlW
3Gi3gWcdd3I7bxVh2LRbsuJttp7+VhoLJGewRkYOjF/pZbES/w8nE7hkL2tubPzL9o4V5/cHrJAK
HooPimUOmPR7QUZFCbbyLGr0InYYe9odOEKPDnYbSa9WguYnUmaE+iw/7ch2YMJbWHgC4Bs6Dyz/
iZcs8P3X5z0EXdBKqaD4hsO5+ZoLYVJu6ys5mHGQzig9F8d89sHTMfJlgC5q3Cl+ZcX8KNbs44mO
99bfDqFH5jENBAyzsdJcYEUqQUkijZA7avmFTaDRexXyNM4oC4dqrjy9RraFGJJxTdSjyQS3NhWj
P0aO6kHEg2bQRlQALZX5TjNauaYKdEo2PHxAnePosc6EQVfb8e0OZrxqTXRRodc9JCPMqhr0aY7T
GMwrdwwhihbn3uEk2QIANiJhegtyxPC4hgf0hrQjLeWz6hf2xzBVzJK43ZKi/Yiggrb4ndKv1JdX
sm8vF8pSNaNLV5E9Y1z28O4Lb3Wa9l+tvAF/GSRibL1RmSXx6Pu6OriJ1hlN9NU0BzOG4of6zYhX
0YnX23c+TCDa5nwqscdzgI53poaMtu37o1mGVf5C+LI/x3JVWYp7qtIF0PqOAg3XchwMm1neZDho
rjoXkWcPiHfRHMX+HE7dA8DTDPirZd8xC1oBcU2NNJRaPNLRm2SpCnQizKeELhdNYlNMnoTSCjVD
kpBOwhHlxKUhKdpd944+o1CZGvkaaM49xxTuDKPzgalK3usXPHY5ZJXGJ4oVA1PEbC9XddUYAEqt
6osicOpisthkKGG3gmfqnozxANzDbZ45rjjjCj6I0eyHFEhaNysmzLdeSES5jNPhgIe+74AXMpf9
SIkCwpA/N3wN55nIkGqroTz6Y6dMtKx2PbF2uapRhGD9eMh9yLgzQRwPkp/zzwztVEI/cwJvQpId
xKC/OJaE8ELXoJjiD7YWyZaE837ftri7K/4TVH75AenEuWzn1xyDDBnSRUcgPafoapjz8XW9k1jN
bBN4mjHi4XPsrX4TUcdayHVanQwJYBWl5EWth6LON79/livTTUAXnjHhc6W2dFcUuSCaxMped8SB
gIENtOK2asPzGxDLeGzhpcrPpR1R8ZQNF0oduFMeaQv0ncF9EqK2n+UxH0RPhXLRUmK4EAGXI/85
LCGTUNY0gCPZ7lKRXDeIfdCYBZzErBdj1ZeIQLrmnWBwnDd5QdWJqETfJBIxB8QCp97OhUxs1GDx
6AR0zvBqajF59iO/HoCs9ojtcuLipvQkRAL/GHsAM3f6rHZGnub+Oa/d0FTOtoUCbVjqFEVvyyRf
bSdm02ixDwkeQLNca5+6kyP09aA6J4rUsfpSjLP7n4hUnakY5jA3/uRPa3z/N0sc7JmC9xHfuq4M
RFSUG/KkC/pPPhiCBMk+jACckWl5J+obg3mgHgHkdBvdoRjlo4gP+tgf8r5AVSo56u1w12GUfAyL
mC5pOteSLkiAv86Gmagt7OoE8sYNkZPLRMQg1qMTBKRip7ssbZJPGZy/vbOM66elSRWLR/l6vA7W
sJidGEQlMp+dLoCraaqgb2JoW13MdpLMKaPpCrDl0d0ebUDsesGAMQcUskRPFTZ1Mc2E6TIbW8YB
MvDjBKBgHyh1f3EvTPG5t1jziXpf5Gl5fXF2pBaIHsZFCktfaafQByEGp6tRds1dB3pLnzP7XCay
29/49Wxq/tyC2qu7KXN7d8rULHfW2dkcAdJO06QlAn95XJt+mpuolIPxQic5cQ0fqaTWofdZW8Gv
IXwpIAWAIiczNvkP4sdhY5IvgUt55kKHrkZb+atMYySW3DrDPVFbgVi2PRd9rWJslHbHjg3QhxfH
2TjQpyyb+KUH8OCfWEK+/qjJArWQrKSECZDlNpkByPbzz3g03X/JpMra2C9wXK0iTpfvPqg176RH
FPL9XTsEPHkNpcfaaDsC/KOuxFyB8/UOsl55wAY6HMhzULjKy3RvP8cI3puyioU6MxMB+VMNIyqr
D5lpKUqX7k+i6wkNV9nWwwH6YUzgiPt6YLLhh5XGoyl8Yo3gNosA8AxnAnHDHLi3RMpgwVQWDBHF
7f016kTaqy59YQIs5zd59No2dAhmHUPcar1gTugU1jufNW/gwCcg7OKgj42l1QC7QEIZy+pEniYT
Ln1eFwNlb5yxvAo8Z0cS+983RGGIG3I8Mx/Zv9WvrBhuLRjBDSdaz0X9EUmWileaRzA1m253+/w2
UTHRqxVGEp8IPTeHgb0wDZm/nl+DdRoiDLSOx8vP9YF5CPrOKwz+l1z86SulSJz4Xcy3vSL7W49L
XwMsQtk4QvZWfaWhyuI7Pd1vbSZ1FgnCEC4/mC8zgtXKE9unMHPSRQ9Vq5CqefvJBDPHp6wKrgkV
zgI7We7l71WeKUwlCRTAAo9zQkwBUYCTEL+f1i/kKATaOXpim3upztR6+2nStG0L7t2h9wHAtotJ
uhrzcv8xz+g9ZPklja9qmVtgqSonsA5127b5lKYH5+jye5n1n4jdts8yEN646/mcKUqz3JRokN+Z
JOn5tmVq9aRpUeZjHppr9zQEAySRWNiO4kPzz9ZMlwRgfBvpL4wrckRZUTuJP7C+fq+/9qq5TaGk
yRxjjvRMgN6r3tItEx5BCqpDl9gJZuHHHFhFIF9TI/tADdUhB0BE7nN6tm3GayuSjnweFxNJklwF
oZZFg/nNOZTKqWTbKONGTmplsNAoR8C8mlSJ5dY+XoWIUH3ntAI0Y1fZODSvEfXFHn5wLZ38Lb6O
frcpbXSS+z+pZXCjJXSkbfosLUKcvFrpiv705tmutEUWhz3KXZ9H6UPBI3WgeHU7s4bamUhQkAdi
8eFM+T0oUgUa1p+xukXwQmyUt9KTMWgXFMcBVxUw2VXz7MhynJMYUCRDsafRBDuHYGzXVphg1FlY
7z2cVPbXg8fggsZ77CbWO4L/MBiwZKvnpxVzR1tvPS1PS0ZNunrfnRrDrkXpH2NPYJjCmHMxEDHe
y/ILwCPyNbEqoA95TfjI7Q/GSng6HrW2wD9nXvWx3udQPUnjk0K50yq75R+Y9QZ9vRWiQ70jL7D2
Ik558a9bnBHC8nhN9RwaQIph+dsd0mOp/ybqBgo7goRhu+BrX7H0/SpdrGzwalEZK7Dgf3BM1vQQ
BsKE7b5DQ1IsrrOIiUVlSFvpq/1jbfwYojAtzCF2yZBly5HF+W7YHB6r+gE8ezZVnVOOX7EWkDFc
l3QbjFIbP4EigD4wAJGYuyrUovVuPHETj41KH06rbGVhpxo7sxqM0nKTkUsVV2ULFzUjVl86tXfp
O2OL62tLPQqs2yncVWDlm3QH1iRyxmWVgT2XrlKCLKjKit9gHzCwW/G9SDubYV310Fx9WSzjndIc
HUsnC41XD6zmiN/85nVNTVI00cvAPncyla4j+ji44irtfrA9/bMkiXlCwtM3JBbC8HBdds/VmHKx
u+u9kGOuQQMrM8cJ/1Hh0Gnx8IuQlNttvKmKlPBSHUsisQrZRgx+vhhuyfLdIla2GGXOgus+rf9q
ipREmibjV/OfGaWGtOHfWqg2rWMkGqB5edBCqxadACYCeUwALXZRTI3fO/jXeZBbkCYAhaj4Rxlj
buG4pN1z9Dm++CvXyWAe0blNmIs5xXL2HuvxXV/EMrKuFh6nxrFM7ByvqDXJIb47GbwB0MBRYCWr
D+f5MAOifPTuW++wZ89mGnhSy48Aa64txv6591xtLsYWNFCSByQbxznORYHuyINUKfb9MqU1VKEb
qdMiyjOEfcyDXT58Hwl7m6rgt+UgC8CBuC/6RtCyOjyDZMcomJRteGJ58WzGgDec4BGDmDTBvE/T
ZfkPegQNpnAZXjMtkBL/ZCPEJZSshQT5EGkvEYbt+ZgWKJnZdOdYn9BQjZ45n6ndXnB8aXxA7dtt
U3CNMkX9KeLxpOVsMe83HCxCr+tPZqgMOcd53SVAOziADyUBOCa4861dLK/GU6l5K33L7UhY+ODh
ZiToZ6DRGfqk9zT6USDfSOC8zsnu/Gc1yBjalrUAmGFlRWFCPZkLt0gh06stckchH8EpPIFxLw5R
RKsfnyV1u9mg4ggp84sgCFDxdMZQn28/lsQ0GAy6iV0D7dbH59h/1zGiMDpfwmMTat8MyAc4HMys
5uiiARKmwQ/Y6ZxLvAkPQS+dXgFTXB+H89ra+S8w4p0ly/+Kpkl20lL5+aLVpzx5BapGiHKK0+K6
Y5g12HFOzjJah+QthXki3yif57Gvu182mM1+6Brq6srCNF6KzFQF6F5+yiXVI73nAjiXBP10Z+Ay
vpboD9Y8VkXGQ1bzKQL/blPGJPeU7DRZZMwloxaotIKN5H0SXP0l/Kmk
`pragma protect end_protected
