// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:20 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J5hGRx30CqAhY5kIPavi1ZpusEIDJmJpy8cSaRZq4IS2eqO/EPvi7OXPV4cVwY9P
IGoLJoRZgJJ+KgpsnOdL9gtxNrRS2TLyJqyT/+pzU1tlzBi51XL6ZHzJaZMby2T8
B6cdH4PlybEyoPcqbBfktgahxaBkVNr986QaFk/tFW4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
OIwKx6Di0lYsK7ChUDAsaGry45TQsi/YTZLsGdW7hFVfksy0ZecSjAY44Obz0KDJ
McDh81sbUp2fmYnI1kTh+4dVLbowaqHmZcHtS24cI+sheUIbbBAbBaCxFTgz6Xt4
53n47LtMpDxuM0XuZI7XdeG2eFqM1/gt5IlUhhHX4cQRwPjubm5uC8UfFvsmwr4d
PgLNZBXoQf5pIpbaRvx4bFF1qboqKlBDDm4o7WAJb44rmC4CsvstFXUKvtApt2Qh
Hq01FttQKG/CD4WxJVbw6Rx3fUtlSrQ4L9KXtwkNyGdNHMUW7YapU3uvoZg4/GKY
VE8DqHvHnBHfrSQUBAtwUial2Xo3Aqs24TkdR9D08Lf2y/iF1uYUuRBEIxdqEmkt
xwORdS7fTZhMQjA845kYpuYemfG8PFgI8U2TZlsBCpdK9igqTyLLbubYf0NcOzT6
MGbuGW4v5a6raseqfPuk0JPCnvPDSRR14YAVXs7Kz2PvK3L47T8oVk1UNLuKwd2Y
BUlbPyVRFdzKHaDdwZTFv8ny1EJtRiG3avpy2J2gZVnHTtQJDXvvbw15ywn8EaRI
25Jgvtj8yLXF3vhXctCnj8HGWN0jrsb3DsG9bui5pHsWRJh3eLp/FSCBx8XD33eZ
gKay7bw6GPdHWPoxXNjoDzWP6gGgBCqVMxafnpOatydQAMbN3T/yvIeNkz+gk9lq
EQCGL0RnaWjQ5xa6OTMIx54jzwerORbPrJSsppo9TVuiMlnV8sSJqd6XQfN0DNI4
YOv6z5GeZrXvtx9ybrKHEV1Jw5eKQAkNC/xAUdwgQxqlKRtoJzkrnu6utTV2imhJ
1Jo4Dfjf9lsgXhdMQkbiWV6MmNhKVt5OiCG+IoizFdZCkV8OhSvf0GvT8vkE8M9z
0uKTN0z+GqP8Yj4J6zEbOAY3A1f3SpVox159zpAdxLVyJsFub7tXoOO+oPuPO2S9
mKBQWAMUM9optTFuw/ZIIwL3VtX+HOIazDcBoTmktIa+tY8Fu1pS/Cvuu5NMH4t9
6O3ul71q9D1JPYcfFIBtG/IEeFB81t8nVIwP/dgOr/cEDaXSQyVt4MxKJTvw2jqS
xFOayPe+FnjdyllnxhfJOkVw+apg82jnOknQpXyOS37+9na0AmYSHQ43uFK6Mosi
8FDTVY7p8qO+Ti68IwLBGAdcEn4eVwvJBVgcAkapGHfkFQId/rwj+mxwwIqgu3fr
iH8y/cROag+6XBjYuWUSqfrulofYNJ0ruC+QigvcrENts46rXnuy6JPv8klYi5Jt
fT92ceRfGM2G1u1S1cmGSazhBcmYRAqp6Xawr6vCR2llYqvBh4eq2NTuC6f1AZlV
OC8FXZQfgKMimFwiyTmn1bMmb5ZvTwQpDie9r/I1d7EdPqshYAok07dPAAWuu+S8
DcM0NzcHBQGL/iWblWWrjQ9SEFFuW5SSEF8tmPRoG7j8MG/gGt8EHy+LcOlBy6mT
SwkghL1KBtbLYHW/EksBaoJcwpYuGfGOye0cMR9FP+VCYY8m56bR0noKSnHAoJsZ
xKPUFdJVGNUNIuLP3tk4E/EpCgPsWbCcGgNOsaImM/8CcbsfmKnlwN7meg3h2zgx
5gPIcB3rrIYFEXQauEgAyVgYrOyvkOyLSF1l2/aZ0lWu3uoOLM7aqKBf1TdLQdvJ
CHpXyCgW/FQc+XMxhaedImeC7L/wuLWLtj0lsbjUlSOvryB+s6bDL9lCSHVXfm20
thK18d8fdPtPNdAE+g8q/4RTsaSZQ4vBeL9qymwBE7vXb3HjmtJQzIRq0oL1b6Xr
C3jqTj2WCmQqoQ4JsEa99D5Ku2jXZRFUCTAFwDHrhW6ZTsSwGQ3S+K77/spDOtVJ
Xph3dff3baWVYq0Tz4ZesS7IQBUcKr+hte2NOrAsPJFfGNlf/Cf0KP2cn4JTZu6+
B+NCvqOGwPoqj4PY+4rGh7QAAGE4D3kYu3Aft6287x16veFXyFHB+H8blSti9znf
tcxWUH3yuq8GXFa9OB/Tpy4LNVF5bb0lRFjyVuP15z+pT1op+cm/pZI94qT2t3uQ
TIWlgmAHEnvAreFr8wMo9ERwJ6V+BTJXO0pruZcgTknWvkXE4uuIDLCatYFpkwMS
TvU7gmU4Sviyo7MuhOgL9aSSwkZa0/gSJmcPa8XxdeEdGm+lGExTy4a2WMuwp/D3
emuQWLKyy2BisP+JbJXPK98xseNbR47Uvc4xh+rnrIKFnwFyQlfbkshp9HsTvqgS
SoyMhKP1KT2cKJ2iJD78J0aptsJdOV4r6kSowI99ks2q690+2740pSTjz42GHji1
fc10ocMMbssS/DflgYQ24zpjKUjxhdUZi87rOBkBZQ+iwxaXjYKaRMvRfS6e8CP7
DFug+CV1Y+sZIxGao6vwyoqTd/L2oxI5JNfLW45mN+W9yTwdgKmVKm3ERCbrAe/F
FEbRDmaBrA12sukU6vRdpkmAKDsCFwNqf1jMa7P2AEzbQfaQM2UJf5EgD6vE7lHK
rWCQdfbeT3kYD+SWhBUqUUMVN8OW/4rUL7kojDfRaxyMgEYRrFNTxnaQmZ1fLzJc
opErz0+9qifcDApijTnuguCpGJagpmo+wySsrS9nHRIBYQODaWp7fvDAr1PU7HtQ
CZSiZkHitfTJERWNJGUrwEaW8XoJ5rDJHp4He6oJrJszvsVVXbFKzBfA2FY6hTOe
AvSZzVLOp6NaJ7W7x1v3moyzOOG/UbIGBQZJ7UmmsREmPLYGyjnZ0FGtP1s6x3Sd
eFlFpEq+ljw5RCV/Jm1WyaD9ozlE7OnhH/tTGYt1ShxNm4woFqjkIs3sezxrfvbw
Q+g8piTWeoRpIdrQsLU22Jy4UGHegODB2NUuFW4YQCkDFG3BvBUG+YPEGaQPOTIj
LmOYdnnY+9X78RsZCRmwAOnpSUbM506/AKLkalGL66intYyN2LQyduofZfBjKOt0
ppX8AwhPmbrJzXEXVp08yFckYn+f9/i8xEqV8iOMZjuvBkezd6D+HWqJTfROGpOB
g1AhibeqFbxVNZbhvOu4MEjdPsQnHxBiPMFAYQR0bRyMZD2dhojcO84OC12ZO9dS
UrdfkKQQTQxRn+vgdGlMuuo3PhZAj/lW5r0iADVd5Wj44+udPJDCULbKj0sFibww
RjrELCQqYejMGKbJlk6ZgCBrpS0JTWFkz5CpCkuFyccNpXV6lck5CvDKFvUlaJ3c
I8unhMIFAGT1FkfvOLu3E0oJ9kBqiNXzOcZ/DyP/ben4u1rCV24p0gdzdZ1bDUC/
Xo5RzMMI+Fo+opskIZAyoAEFDqwlt8ABD/9R8tlGvp2NrI2yT1tmvyf8miCClGNP
XBtQOtWhgOYuyntUjBtlYxyTKm8FBlmKQ4WAyYzFBXhzg1KxsICTnFwGWXE+P80u
B4fsSQ9VtN6KduEfibz1tWH0Pejnjh4Oq8E9kOA2YVy7aZGRbSQWY/4UdjI2vPMk
ypm7xmpWhUxuSN4llICwMQ1N2w5HaScePxqtKcVRUICJqESfysn6lO3s1KQgMZCc
rfNwXzznKggzvp8F6SRwWDNqGcj4VJNlHY2tLC1zhofsCe5oly0se3czQpLEaJx5
QAH6+bHOO+TeZHEVW1sD5CQO4Bs2X0+PaihNcEfnBWMgKsCjFUYC0TbHOPzOWrJq
0HdXoWdBeVlsbElqxflysxrG3I2VzjGVWOjXOxAEe7oSPVIO74ghbNulOK5KRMjJ
Qo5zASyAGZVjUKEHO2f+FqDSzt+MqTXwnK1zO61TvJjcfyejkCPEDnotyx+MFOFH
gIfLOBf9ua+Eog1CbbGkOwwyAE1Gr9lYfllEPRbsRd/BviH50h5/WoyfBAqbzr2x
Ywf3YiTkp/HwT2+EBR4govUcqQ8kzfHu5cD1tGXveti99W53+CNDo77/Tn/ierbN
wMeH8GrDzHQTe7fdtvc+Y/wbU1n+gwI1QmZi4nvLcs2nrhEinBt0gTMil8Otb7Ft
lZ3BvCTyhK/C7Qfe53zrNo/RH5T/TQwTya3Vz5D2YMZfOfCbli0f3aMQ1LbF44cc
m1dV5tCYDnDIE1ofYYA41Y5Ad0txX/6beoFAUSp+stNHXawOoeFq5RIKcknHbEU6
vOES1H183JTll0JkCZ/+mcQjiiev1qWHhgIr5fOaoqIBN+U2xfd3t1Xa+XAhOxvu
a5MfeCBJVqO1qm6M25wGvZLnW8RxrylM+8SqUh+ZUHfQ85ZjviO4JM92rXWBVGpV
VSJoo/I4aETuTd1RDhO9+wLqiS7OFEjOuAglXg2YOYAIZnmiM70KWzPxFwhc/y/1
cHtkJwqtjIL1Oy/6A//H791GILTrG/URI7+Tofttaif9LxT6RY9CS96WeCcv7sgp
woh/wKpwIk/Z7TYbQa2PwcaiaBsTu0mr1Nh/qDKA13+HAEIDtvZ6kbq7dHHS9nxE
9xp/Jn7LY4mvBXki5z8zXT3Ub+fOvgkSySiuN1P7bXZHG5+q3zr9vIsCqFukfH7T
ufu4Bv6OaknopYg2BMJM2/OnItnYvaAMO2R1PRh3DK3q9E1wD+f58hoTsZ0yASM2
HEMnpBGOBnBeUi7bc8o7Sha87RDzOj2N+T/9hhSFGVzOwNNGgFifRjfsKKhqjllv
bBb4pN9Lb1jbpwDsQSNiteq4wKtXbTQp7BnoyB1YsIkVs+dGP40lS68Jm2cI/Vpl
yieXgliXzwAvsD/pt7+ClmNy/Cz+7JnhUQIwq9dcr1DwKx/fYiudVjL5/iP7nLUB
vH8Nb7kj7+rgd6GWpQhYVyWvCQv5qrSYj7J1x+At2VWrlHFUMSWlhpKGjk+wMkBw
2zsLYxbDbSb7LQRPdvsZp0HIbVS+uhdoJrxcBeLrsQR2zJogw0Otyh3HOQIPQzc1
w1I2/Lka18VjbksdzScDe8ah/O2TI//h8/4yUVZdDTIcyK93JnlC711Cxvyu1GN9
xvTtWFtVKYrWNnhnuC+65mLazoePKkmEslcYft6icMwWUqwItMuZHl68Qy2uQp0E
NYXXXfQLXAf9+I1H2/jMFWVuzoAnrJccxc0t1GOMaJbQBpQglvwgOatPsiX+1Ez8
d94Idg2HWnA/z8RIO2XyL4BGLTpgtltGU2U1vkI1FU+QGvnewIK669zGZWoOdHAb
FYy8HSlrUKetcddZOuTkKYz0mTAtPRPpPRqWtY6ttl6JJ3gPa75Mt1f9qnBSW+Sv
vrhAhpbdfJEPjhe10adYVOoLldMbu2+W8WnNLHhJiDn8lebziW6UHHMm2aPtwPVq
QxCspqzh/rArHwGQZxo00AalFiZgYkrGeYDEn1dU3Xt7ZEFZbuvAauy5mwnlYACW
+6XUIUeZ5QzjeChNezjHxRDIqeuBt2vVRXGN6b9kKvROOHH9z/CxAWz5DyTj+ws2
UjyB5/fvclLoTjHgZ31wLxmMmbdyVDrPmEXnmCrgHNuD2ISiitKIhJhmohgnnpqK
hD4b2dfnnzbZseCzjm4Y/Yxp03zwcte2nk8XUuF1w4Y+E3VafKZddgyoeCkAR20B
wE1+jfow3VksZcbpKWv0NWlIM2cwoDnhSwjKDJ27t1DNcE7zELrqNmklMWznT7OQ
p9ZdtlElc+uYJSUSGs9xPOXYOu6wC5qBy/D6v6k4UFZFvUcmoekbSE29HC1pROUH
HcjQqz7kAG4mH516MYFjtUxMEBftKH59n+WMfVQt3rCpLtI/vV3sSTnMAsglQeT4
Yr6GTkCRI0Z3Lb/J7bVr/GDJHuCcYNNFXLpElrLAME3Dvq3hdCgtsvaPSixYt/e/
555bwmekspzcj/8hb6cQYIJuaUTEGYz48yOM7KiMQR5oIb2OvdfXxUapjGL3QNq1
rh3QWljvoCKIhYaXCznMQfm1MWzUQ+pZTrQRNhaZS9YWfghpTZI1gZtt99MSEowb
/KnM/cGKF5kDjClNpRxXmhh/t9hZnHWdA9MtR1sONglqUKvdrlSiNgKsoekbjsM1
MsXOtlSURaXHVh5gGRuAtvV7RN1z9YqTiJQJrxD+0h9Hv4Wa77zUnNtgRGRjguxV
7u+SfntQCMm9zU3RHv7qTULyVhiH10YbcIvvRB0GBfMS6+RvoNo2M+wXM1Bekc2n
LTMmsSjk/LQeQQv2XCrdvQaGcXD8ScMXPfVTLDxWy1VhHqClDQdVTDQtEB9WxltE
vRFEB88I2/YHhMtrdbqHQ/D6YWYR119hKXtW6DR0a0/F5kwSHVG3zVz+18CgvFtJ
1fBxxbSHF9R08UYUPio+lsmykmkGLFf+jvcWF+3oIa9DSikRqPZVOMO2jJ0mYL99
kxBQi1nVWfrIf/uHirJvJrJZ8ZfgmE6e8O79LWSaoeLYXSAcrLlK4TBeUvJhoe54
U0SFvEnUOxHFKQAhjv1efQJO/WCYVMDNPBwVIeu8nCv4mlW7PdtoC1OgJCJR1Eha
H3+Ms/KDt77Ocits/ljv/gAinD9suJNshR+qLm61u/U5ovMI09avnP2sUUymtfyl
+YnN2LNrzoEPBQu2GLnACaXIgvNXsOYwfggoJWlJh30jGcHWWN/adod5TvOz9q74
hhRunO+jKKKkNgkqGbxmL5ueVnMBoi4xRL0fp8HQ6Dz5vTJBkjZiy/fMyvCYcQGh
YaNZV2JnBqRZ/OrrpW973Bbalv5xTuJanBuVKMXfWGm01k2A1lw0xZvxUsD3rYl9
+fNM8h7Y/YqFG5xGWo16ZLP30tnEDbTDVWho5ZdQWHDXDVVpHimDNdkxXXCk7NhK
vZMhESFd61VSfRTg53+70DoUJNtDOl5MybVEtNGh7I4p4jqENbuELeiXXZwc/lTc
VJUZ3LTiplqKKroypdOdvzwDFqidoUbdcvMYWQ6kmWWJ9qp+aBYbfAm19aPFXwFF
WOEB9hJyViPubw1UamfxB9Ytz8NmVj6eiquqIMfPswq6DhATkKaNUCxP1xt7goCv
zENrZEaC+JZjvFje2k6QSzgjheJ3pJYRdqS/ns8KxbD3RBtk66z8hb4bspZP1u9x
b+lXBgs/8c+L6vMPeinevjFWXubJLHLV0RGjdD00MMijWQdx+aCMnCWlUw6CHfFT
krRFcYl4uTQE1zimfQ9sPQtUZwKb3G9DWQbOXiLWmVfjD0ILgEv6qqxLnystDPkV
hmcCFTSEgI+vvCbDDY8j5y42FvKQmOGCVpL9DC5HOxR0eowvFF63jTA51zVEwvv3
DgHdU1Fjy3jzZu4BUZeodVQuVzXpPlAf7IlgYIte6VXUP6cG2+9ow3eOH9KFC8Da
7hi55ch5ESo5/IRn+jEUyMU3B/WlQXMDoLVcRirBYbocet0WD6Y1aiygSugiTIma
H8p4yK8te9PvtBfJ1j/xyXm2Mr2/lsBRaHxJbDDfpskTe1mc/gAmrPovwS587adA
S8OIlP7dM66ml7zRytYFhZ+iIZ3cj59I7dA/dejg1tAbtJcGYAJYkUsPS2L0q9Gg
80Pht2E2Ys5Wsy7vwdbuIXWBSN1syaGhQRAM5BE0xthMYfvm6ZlXWkGlBGLZeWqM
jAgUGLYI1ARJC3T7V8hLkL9B1xGaVYnX+FBkOaM2NldiTAtzK/bDi9GTq33RyIz8
i3/vJzjje/KE2sP6RBSWVdv7FCAY8SOOuwzZvrQbFz5iCdOcSGUA9b2stfpYoF78
66VdkL9mzFKzOsHu9ofS2gDT0HNJ4BNZz0lDl1K5Yq+3Law+9wGyx2R0x0L15eTf
kq9n1btmPWYEkMmfIlQ5PnyFqHyL8WWBZqSoQXQfy/i2+MdPkX87wJrW+O1Swz9h
fV2T+n4/m0Ru431LOtn6sIJFRlIXf0rC0qSsrdBJhdVy1i7w8pR4RUdjrpElRMCU
/4S66RbVodiD3D/Qy5aQYEPU/M7s8pJbNTSNXSTraWbrvwYC4q9FudgK3DSgzE0A
1xlVyshJivW1JOWqfj5NnP3Pe0rqlVt5VQUADtaomUGyqVEgdNFRicgDRMzTwSwP
ZhEqV8lYh9dGnIlBXs+SLRgLtHOxMv1IagPwkd9PWfLQ1yyIlNHyOEmf2OSGWYw/
wo+tzudQOxyMGsF5LeSogHjTrHDmao4VxeUbpsH9Gd89eqv4TQJh7CYjQoTo7YC/
QfxMMkhIMsB4Y5+PXSsfCzqoJRmTS6L0PDToMxv2Icz0k+1qKEuuLLqc9knnSW5S
MMiLMZpZb4TZ6/kZP/lqxkDIVbUVC5BCFDjNtZqmmu97VIrzKJd9zXDLx6lMAzvR
1ousuh3i3jDIW86KwsuFdkembHCu3aXSi+2vLfUsg+zt+k5iKWaficeJyT5KG3Zu
YtMqpORJz7Ikt5PSiLtRlUQcQx6xskKBqyRk7Ofhu5lp14sJs2LmcWoYEO8eKERs
YeDf4mTOBDzrDetjJt0oG6FZsoSP+yMQhodcKkQSWGgai10qDgXcASeKw9O1mxo2
MPuyZY41NtnJSvhfZ7gt6roz7BhJpOK4W0yGCOikoDCJGaXSfAQ8Y42H5byIPh1q
1Gaa9tpiKNHHlxMhXOGh1IEIWHdbLpoaDMWuZ6szyOo/fTFg3lgqamItNbUTTVmg
RDnwP48JMM6ROuYCOF/SgRH1sj6RRLSVMI+IcQ/5QOp7RjbB3COebyq8blWyiUqE
8nHz5uwPArLAI6OAS7ujGyw3osjyUalMg6zpClLTlo9PXXXl8XhbyoaAScrWI53d
L0eTbmUX6MQGVcA7oGnv84hixs8/RSNv2JEoIJ6heHJ/b0Tcd/VVlhjfdULG1C+0
WxdgV14WPtroX5vF1PXd9Hg8lVexf8robZ0SPs3EBLJPTkMeAcv3BRALJMdfL213
O76LRkKlQ27Zs7QBXSk1+MS280US3Eri+DUseHZfe7+scKVIU4FJ9Bmrj1VTjonv
HfAkcp+7+CY2v6BMCIP0/4HFjkGZ4J7gMWWSqO5IkyJ1Sdt7SyL5ZfFB0QBvaQjs
aUA4F4Bd4DWbLsetCWgtFccp5lui1Gr3Eb/eyGIW4qQt8mjzz8b/rUkThqKOu6lB
4anmuxjrxvgYpSCE6h+asDvyS68Z+NFs3zBJW8L0BqL1LVBsivJ05dkY2cc1dmZ9
fGZ6gVHzISdnV5zR7u1VpAlOIEBRFEfQ/zxFGO+RflcgvVw6p+uuNr8arvCUIJQZ
fNARN3PpRBirBNl0zxNFSMV7bcuylH4j1R8R76SVuyYAVsa9+QF3ixTFOlkcpyBa
x5DbN2TmDzaKKFTdC9900XHlPx5TafAsCJ2gi7nfqDchoW2EVkf1hA/ZXVAcJs+H
0cmjmP+q541K5TB7/GffX+YyOXFMEPAPzg90fEZWbadQTWKnZDpnQPWTgsUScEzZ
WdlrhDkgB4BH5jxjUGVhhypeOPtaFSAboOMeD7UNBWKEef6Q4KBn07sJeH3gaSaf
YKdko4lcI0XZMNHoQgUwbJevDT/WqZL2c3gzgYN4z+pjpCpKQJb1xzHGD8Dj2yTD
0qaPg/a+0Eqj5oXI7ohZoVzGcJmCgNXC5iqLvuOcA9sEYnIPPbJcMDql8FwhP2Sg
/ZIlsuCNqHKrHTwTYDhOKK8ZPMeOl1Qo6+WevgIVl/2/hbrCbp4MmoPG4kJOEWjQ
Lht6pRIG2lWaWlAI1/w+fDg1IxzV1Zh2NQnSW30A2slYVNOUYcwrnY+XdDKHKMcO
OOmI4/cPifxIn7Fw6JeySYGHhXOlNqEzTYg95rlxHlnKpe+34LqZ0bTvx225QINY
xEEYbFdoGPh3bo4oIo6TJTIEfdD89D/+vL0uR44HeMWsP/P9dFWTtpRY07q9jwqJ
fuyBRFBNH6/70dYiui9NaphrkiXQksdqoBUk4GOypn4hemagY1rSP+veoVaci1fH
wjRChk/wi83FxiG4zM7t/0qVv/sbIioVMzZkzG4dMr8NTu/kQRTUQZ7L+zy9c5o2
SIENpqlT1JcuFKwwo7mm9MNwhSzArh2+/UyP42FTA8a/0h+EZSYMzrGs6COJwEx5
vAJTQnJyXutHoorOQut8gM4TZRIQ4xoYJ9ANU3W5OXG5A5z4jqJMZgggHu8nZoW6
4XOJdo8GQTcFghgqqbeoor3MrQ8Dn5pdl7sOePZwRgBnDLoLYELOD7mxE8dEEmed
PYh0+YukhMp9tcw4WO8CJf+frDqE2Nu3T5H9PpRs+8gByNzyvxdqqxupi4a4avyV
PvXKTr1ZWSKT+BYdSiozz0aaUAf+KJpCoEXPQ1QML21Ai0NURVWnXO6VqV1/06cG
oXt/u+jCChx2U2unFkZW1JP2kqXISBrDWI9bKzciubi1QfQmbOCcGz5Ax18SL79C
i02/zKS5agr49VviuYfnvav19cJNgA57D8ypvC/VjwXIurkpsJ2vo4pv8Ue58rzk
0h1a2ewFbpN4xud+w76AFZPcS4Uv2xWwV2TnE//PjChvgH9G3O5GzSo6q5vmwdxl
JQuOdnzWS02NpwTii5mUb5yTLXsRRn+XCs2WepnPt+V5wnfgqo0FgW73iT9jnAaq
9s6xtEyc5fULkDwwJbp6xBDq0gteBNyvlpIF+7UY8sqqT+IGsl9OK/yYPe2c2TMA
/n7/xO8HjGZOKOXujm664ztHOicWmdyxBMPnY0XPtbZwV65xcdKRaFj/BBKCyiY6
5M2HaYiYVDxHtcA+PmBrCuCdftARPnhO2qIcIoVCX/62i+4SXjfzBDtEnq9AK5LK
PB26PyYHgEs7NI2TQd1OlmPOxns1NPfScDG8mfwXu+vuS5hQc5Inv1XbaOWkWiTo
5AhuvPnMDgBlvQIatEttSKcJB6xx9uo6VwOcIbxbSMHWM3VVxk4xSpbXqXjprSvY
OYqc+PMggxIc3TkVHY6vSDyX4h85JOhVOOYrp5+nrXFGYwquC2tHIQSoYnfNp11/
vvNzQEUyDxVCDsbZrJ23OeYczhN8kPNPpfAtDz6uXQeZguvyHK33W3VLKXdS3pW/
YenN/5vbWKGGVjpIrx1Xs3/1ZeDt+OqRG46hBSXcRpanlWJOUY5fsjfWXBRVbhif
vQImDZlDZXWr1Duy1OEm3DKuYRZzB592sZTUNFTeBLRWhRRotRI99aeHd+Ysk7YK
QUKT9YcAHyhxQFFgxpT4YXxCvTFF10vxN6Yyj//J7cp8VEO8oOXPv/GNpwG537vc
7nofvRXfOTUu/wXrIyZnne+8xP/UcTSu1w1d0zfsKjc9OLGCDTeISo/Wq0cCDuIc
6TnCklUVOKyd2sOiZFxZhkJfgOy8YwP5jqSqH9wes9mcBmqlPjidJINYgHummKv4
wWwnkwNKgKlGySFO+bpFgfD4IuhurLG3FoGyJLuLPgMnqNNWbKi7+6OKQSgpspMi
arbFwuYgkvyKRq4nvOzYxmuUDJYELh24/v7UVAPgBRlBiPixnVHda7iAsH3U8LbK
8GdzJ+aFiK8EeeiBdyS7jnzHjRv2iSXKYAfEewuWRFEacb097QxPdwGrR+SHAc1h
+bmr0xPh79pM07Zrec8EfqSaQSrYzhI9innD98NynRauqSZenOziXqO7/h6U59oI
0Z+TKkV0mIg2/hTbnY5y3/hZbRWA8jVFi1Aty852l5YevlfJEL24iOP5nlcMUsbW
1L37O+Rl3P8WpIBaOsI36BXxPtFP9i+GK3KFndEGk+yEr2NK8AlErIY7FxTMqLj2
3+gYbSSnRVgpmd0yG0FU5HLEb29otNuvKRG405Bp9F1JGHHOWvhO7YtUUQIOZ1dE
0Drk+azTmQpszyYc/0b9c3KCXLo55seiphBHSsSLf/b+U8c6nVZ6Osd3Qm4LsHZI
pxjCf59vQFJgXT39w9XqraMvKn3O99QC/WjSI8a40piA05vbGQRMlZ3OiFbfCBsE
34agqcr5EHLem1OcXa5w/kavA4uA7sq8UNpqaLs+eFaiy+b26ZxAXUET5KxYP/l1
8LzATq8jFCdi6P/LrAPLhVAeg9b1cI8qg4tKGlCDWjKZHKg8j3/Qxe75wCR3Fopt
lsq7UxrLYZGStyMXRunOfbMEVQwWvqjvRNLKmK1N/561yfbHg2d1w/tPok1qAjM4
RfIa4sUpNPrc5p8ntA0SezsgvCeB16vATuvYIOVzsVPeB4QmmzZfk7VYcVy6zg8p
+WMiCNcDtkzVm4yBZS9npn+m6ln5smT4kymgp3pP6UKydNeHGgIqi0gAEHxt2/Od
dgf8EnESVYgh5WyCu13CZqErj19GtV/cZQuwI4CVwaaJgNaOqRoV0lPSMl0G1uRJ
rNhoyifdJ9c8WkbLfCnHT24EqIOCFklNsDIhpBFuv/4RxO1XBd5QK75cXXPiDFNq
KLRDUxhns3SHc/ntGMzYervzDuyQuFxtcz6Rd6mcBXvb22IS6BCAti3EhPwHK3IS
841UEox2xK8bTAUcDYSLtdt9OXZXbxU1K9A4/z7vRrqiT8hdm35nWqubD+k+njxo
FOqFh7OteP5frEUfLj9pTNr9z7N9uYpwk6qdM52XPms976/2Y4BvEUmTaAHy1OU+
i5uEMgBcIdCxuASQTCqeuMjwGgNezChgqObVBJ0iZbW6oVrEyv4z2LzfuBwb5L2H
q8hIgdoazD+qZfU19fTZDvAX1/rNI8H79/sGw6TL8VJG0/i6Q3coEouG+ibHd3Me
yOupDpHRSL7Q4FbapKjDf7LktJ/wBaeIP1vRlfKjClxMuww1yTkhTX2gp07rrLSN
Uiwd+Hvh7jTVuefufs/KQGZLLryG4OuTtu+ngvDVL3BRThzVDyH4syP7Ag8jQ+Zy
MZ7hXEDACXTaAYzgx0kzAdk4yWV0bmHeB/q655LwrT8kK35XDaprzynJYjyNZ2Zg
Gl0SvKzVhKNkzLUgPMi5Z10yAoF8fFmLV8+qaZCRRB6e1sjIPEuAO8WqRq+hjygj
OZ6aJ1wEIX40QSWlP/9BWLxaTOTYN9br6q3IjdDdYTV4qVXb26lJBEqcosu49fsb
kiOCd/rvEbDVJScqHnxxWz9075Hld8YfQB+Vox4Ua3Kr5KQ0P281S6tHy6CL8mDF
ibl14oUf9txZ/om8gR+G84AwIqtXIp5wkdKeDggOLxEH1A0j0Xuy+BAoBM/g10b1
pd+Jafd0Q0PomZLmVxZhjI42kYJ3sDVW6M5q/droYZpEmNB7RWurOT/0gQlyjwUc
8qMhygvUjGIF1Fbs023ja820139eNbPqIX60pQYnf8O1xpAKTdBz2/z3uJH0UGP7
pq94dZxebRtFwO9Xe2RWGYuc2ZVTAQUp1myQrvGnx6aZJwJI6pgdNkZz0wE8Awry
Pqy7WAyWv8upsmXOsqkTU9fcBESG0eNeS9uJcuLQTTUOXVLv4veHn1QPPYLZ8Ohz
pLho7jhsACykRT33ng9bFE+3Wkbqiey3TLCjiaZmkDLgxZyA5F4rH/5b/68LeJIz
rW7BnzJcLwttt+jrFRB7K3GSN/rBCCzN/vh4DnEPxwXPKMqk1WxMvJugAuYqMHau
y9Orn3X/UWm6AU2GxfzFDwZTFOWpiyk5dh9yE6oxR64AShGsZAzGU/yY6R7FTaKx
wp0DaBv6MTb+anlUHQ8sDGUoR9MZ5FXMRJymhpfTKlTGH27R5TYE9iSC/wd92rLa
ln8e4HEy79YwVC2ghKRjtKvUc4rpmEsmIarEn39zeReVmSfYdg4qoWgAJA9ODLDw
8WcoG3pvIS5oY4Qvmn695C/wps6KmHt0fEdFyHV4WHcbVBbtKfPcargNOkIOAC4J
baDNvwhS2NQ7jbsx/WtX2nZz2wWwqfrudd0GhJgu3y41b6efWpcLT17mNzeqOA3n
SoAjbUt6I8t/uWC78C7CFv+WW2jGteIIasLFzXani/YNDdYlHGhwnTVCBzhlQq4A
eBQeiACA8FUqaD1Iy5mukx2kt+1IcmxWNQLc1RU/SZ0qbkLdsHNRKzuAICY8iChK
DmwkPedEthSMZk2gJa3VltnDwXChOJKLjKBrNGcQtxIQV3gnAl3FsFzuW5A9PoGa
rocigKpOC2YKtxQM7geASTwMy6MqyxU6xDfGQfwQ+BX/4YH6mtHNnL26fU/i+NiK
8dq9/B2j2HrhFvNsjgP3z2IxwvKgfEiub1dc6EDgeW+JeHLVOCkrI4+INryPwO+T
O/g8uqOGnKoll/lEiPUx4+X4/gb8mcqPkTEcXdBNkbex86ECC6jkcpwmqFEyMMGY
w4tFvmA9DxloMDvR0Hnb5Kk6LVtoyoILVGH0Ti3HluWQAOPfM8IhL3m3NCQckozD
/OQ00TA+TRluDwA6Z6evZHj0i9zJZhe/ME5Zd2G2FowhCXzFAEgE8StILW9vIzZW
0M+ROhv+MxtaS5VU+7EzR2JgHTfRdtpxlbbcR/r7OXRHTCy53s4VQG03lfVo2CjD
71CyWjWgM1R91niHTknK9hYTDcjCna0Wqv3ochLUslYDYxF4vO3kdfmdx4yfcNI+
cIGHA1bIaBXB7soCA99elOjAPI6vA2Wg3DJL+YCUv54yyGg6UOgTG5yFOS5R56k3
CZO/N3jGhKREM6aAsv2//duwE6u17Adl0dttQY9PFGzoJCmCHKP0UU4v6DOH3hJb
zr1fQgpfp0nl2ejYAqjbPBMghE1AGl9N9/b0ffXWRuYCdE85l18boTvVhrdYKg2e
nOE2P2+qAb2GYWgqns9XzWqoKHWymR9afcgh0OKuLT6dvaqJ17G49sNT8V8YSDVc
MAvqRjSPuVaAChcKbOkFhyziX60+eFwIAdk2IWuyKzlvRUDgURR4rRf3YwJB6TAm
G3hRBOTb0EJLSpxb8/d39ra3sK7h+rkyQnII/Zzx0LycKqD+5kTOat+09/WpwsYZ
CGcvBunWj5N3Ott0HEIx9NqeNSZpj/jOmo4jhBKUV1Y915RxG+ZKO9NqBldytimE
WzzelrLnkrMfHr+S6V6XB5aX3LvmS3P6jSpfKFc+jXxr9E4SF1+4K/55jEJE2Le9
Jf+DqsKom6ODrLxHSbKuyplhyid9l/JuzfA7qkCNBztrMjeyfGHuzLS543MfMnhZ
E7hYuWOI2sd/bulDN11Tpl/GUYtxWYwBdz2TvNAJnx0gPifEf/KZg81bMPiQqq8H
lZmHJZ8MCxXhVTG9MFrxD90mG7CNupJn/JjlxjEWKN25bRT8MdBdeK7rW9OOse06
FpgBo3ocW0ZYwe2wmcubnH57snaJHXnANCWCAqpKlilTR3NZXelKUDicnXXf8lpG
nUtLH1K3/uMmHtSLjODi2scp1f35DKSDzrqiVFS5+MwMv5Sphmcf3IuCtS0GDcGs
KZOeXlV7uxRWHs+Cjm6q2w/tGSlUVfaigFWlVrT92NaJW/imq9hcjLvrF1zOVzZN
cmB3yQOlkDkz9j1Cnwwqbh87SPr2LYkDFYeCvf8Vfsm2DhVsEz1F2eGMZmgWqCLI
ZRiO2NzfTvkPjA4PQIIzvA+jbzVEL0J60VdbSm8L+nh3Mcq4oEQzMfYBjbJSfHoK
fHjiPY1vRQrYn9ccNmFKknBu6eTmu/i3eiOoUzkj4dLsBrLG4KQ8sX95+mWqvISz
+7VZuHqI2H05iSMkSwEaiX2xKVzHbMMkLCHedK3oevtZLf0gea6OHnFwIAoBnpze
HnMQofMw8GpV7znpo3kqD14cMpRwe/pRIkdAzI74FFN7rDdfC80S3LWi+yc8cb6G
1dc+tAFksAjfqxeaSjmhlky7MMaZashyR8hBOj9G2jHMfOxyEAjDrUumkMZXacJx
4l4HE7W59CFqys45hdzJTbJ+6C6ZkT0NKpznzsZ8vN6PfntCzHUZ8RWm/Idjkv82
XsOlXEKZTaAr0tQopGlCknZYLjUk0w/95k812rbXaF3KSLcpYDNLxaUnBc9wRKms
WQB+1NfphpwDT3rc6QYRJHWyPLifCHTEwmGEkhwTvtYX1E+3cQY6/PuBTEBvaI3J
1plJIc8X1cJUISrQz8r1tz7ThnGnqBgCwgByQz/F/tlprTlEpP/BOQ+eiVzzw6vm
IesGjIwgZ2Ej4kVlxxLv6drZE7xG2CiDc7sALpJdb3avgofEG/0NyM03elEnqk63
Dpuf0btJtR14vjAo9Vg7NlDRrDfm6Pv4WWqR9nPSXymYkm4bu2CFu+q6LjNQpgoG
5+XzWAQzMBf6xYn9jGLSDzjlP6+x1bAaDdHIiAKmqL01Neo+2DW3S3utekzbXIIF
bdWC6Yf0OnkUwrveEjM6We1OGKlVCse+dMVOQeY8Bn5SSz59aOn4cc5EWPhvhAVi
Spl+2k/VpF3bE7vSmeMVM9yDy7tU7ZKafTzajfppGcpXhrXLHSjFhwlyw1pOTiy3
mQWPtG7W4fX1W/3+nfDpC+ZU3UAwQV9VGUDmxvtmCyuY2vcoRsRBBkUW6mKh/epV
suiUloy9HWExH2Y+kUIOd55ADDiuMN2RhzOTEDM6LX5nO8mpdky7d8l8UGdZZoMX
GPeEUobIlEf9ZS9ps4DAFsAf0YBwXSjIey1wcC1JCHWbG+NKMQNeKtxathuNj1B6
OiPps5C3v+sZBp9PUBTM8S68rOrWij4XylrHsqMllC8nnK0dqprV7qvnpQX2Exxu
wgV7bzeE5MN3Pv6m7c/q1g0DnVnS2IIWZlKJjqvdtuBnNb3XviObSJvtRO7hWjeC
JoL3PKesQHHD/syNGiTroHJlIbzx9FOwtdAOT1kyKEGmyCcaM3zOXUUK7UFNNPM2
t8P+TDo2Qk6xHc9jIeqrOJFhY9iYS5tk04cCOfq9peGSAaPGoxEZG5iC8kknKV4i
qPKj2j88+zrw+/NIOqxkxwybG+am7sXq0L4CdLv4KUr/XxCvMCVK3VXWjV95PU3y
8EV/QHTwEuqY1ufZnpSNP2tdtSOGVXu2z63/Kiel2iWIvmCnZTkyzf/cKHAgM69q
cQg2QT7QPQfzfVvM+K/CtJuUhXmnd3AbR5OnKjFFZK2ds1Q59DRAtGIaTUN2CqwX
QGO8+UyBLOw5tIhp1gS8PbR16tBzL8jdgXpIkO75ttUJqexfz7QdVvDbKyD5wyFl
7rzOwrRBXZ/fbw3CmEH+X9GQwGgl1BTob8fXHk7qS9j/OkQaoCFykobfRBCv5bHG
Yko4l6oODiTpyw1TbJhJVHZAiLgeipp9Ap4AMPBbFwny9PbW7oRBsc87XAcWAwRA
u3cGsUsePtGqfqi5O3G05P9eSrwMyErtbZ88WHA0TSkCdrzpMmG6nfMdDpHnjsFp
UyuHh6MxgY0d3VGtVsUxEqqlW+xxWkw6Gsn2lH/5TGrmaqXSQjTu8R6HttkEE1fA
0o4L3zkaq9qM7t65yaDJSIeJIoXF3o4Fo9VTGO8BwyBOkdWVlg8r6A1b8IN/wAks
KAg68DL4AGzmOubbFDjbHpt+Po0UQkNWdHIXsGfo9mRDoL6CXAUhlL97Dk1Uk/R2
IZ5z5ToRVf4x7XwINx1W+wWSw13FZl4OOSudFdIiVdfMqfH/p6SHTj3ickogfWvJ
XFm2p0mtPmm9SS+6wbt/ekC5mKpzbsx3BXTBrl7Q0abUpxMNK5i3gJJKIAqbBQMA
s4gh+8vxG0upw6F8/nKHfzTVWXYY1sKamWoFKNX+QSJfrjVzBPnLhsR7qeJEMbua
s98oP0RJ+86pu1B9EHpMry9u2T5mMFWETYqIqsDJa6MaR4zBgoztxBsZmKaLOChZ
7VtNZSj+qK1j8rqOA7IzZdcyDP223l8FY0Z5OLIHGzS0yR6sNpp3zCNWztzllWZD
fRVVf4ozUtXtgxQbRYEL2cktxneJdWvTUWSBMxIk8OsrHYIgKx4X4FhjakTSkIBn
XJxI7mP8ykBFMJRI03D/xZ4D73bwwf1yV3fY1Gq1L1dMp8ZvcsAg8hAlsT7X9vQb
HphTfA/ESLnzwrccMoaNUiYgARKG4flBD4heKRP1C5JlHqYs0qFe7Oisw2/NgfKO
+Z7Po8sGq/UJhVP/NxXchkAWfWjlL5kOqTvWBzLzMU4Fb9vkczh0ZWnamCxCSpFz
/tkqnkLOeG4wZO/wFLB7e8Fs08lVEiOnc70GssfT5pMJFzUc9FBw8gUy8AUXgNW8
Ip5QpJ8nmtUI85P+kx19iBr4RzfsqN2Nz63pMrDGhAwxyqC0eHNCnUsHM1IMwzGn
crInIZamarHtm+O9feAILENobyI5Mczw9xR9lZDevBiRTkuAIhup76ri/ppBFyvM
+4BXw6vl+rMOQYj0zBocSNSchy9+4z3eRe2UIwRHvSXNdERxj3TJ3AYjqub14SWz
BAILR9qULHTN7jLi+sROrfoeX4u0eroNQB+ZVKvauPMSA46sCkQK+Xrq9q81KAyQ
iHdwxbIpgrb5rl/p9rGZZl8ELN3GMz5TF0OR+vQ6p8t7jzJw3Mgz0hlkJjLXpH97
qu59s6On+/3bghoqWuBhvQJcm4M/IyxTPJO31FbVGKP+9SvYNg+N8QdQAs40WLN7
Ndp/azWBUjNxpnGUEp4bxH40WMCEv+wFEp0UAGo8PqT+F2j4ysFRL2S6YSc/Jv+U
HOyeGKdubqmATur9MupBvb/s4iJAvyeL0bd8UIkTHjKGu0sdCqGmwcdu6+f9d/FK
2MGpV4tTn8bFDJE0BBFCEdk6COdIKVUSfgpUO5Hcj/P2l+FPzjCFhuKPMVAST/HB
6AIs4O29K4ol2Y4Dn0wepjQKA6G5OUD9ojZWOqTZWF9HDDN9fY4rqk/NrrCbB0eJ
2ovoaCf1Lrn+n+2mGQuO6KeIAOp3HSldmEsVZkk8nKjN66iJtiJZNoEfrWyvrPn8
Lb/rgYRSrsHzyXlWnZmIHUa+1GfjGtrsjjbl2ayI75PiCjhtiBc0AQDR3/wYg7fW
SLRjLi+XmxkezAMzUcdRLE04eHtdoUeKrXTJsTCuRlR1dR/00zmvkHMn51r/HQym
k0mcPFhMiFmsKV1vKzhzMp5mvfAZc/RnD6lhfyf22PBGlzS9OLFJ8Nly3IdpUhKg
XGl0512pNW66cN6WubeumpEY10AfaVaKe0WoDAAGADPoeozUl7KLbJSoXNebK3c1
5eR8dydHBZmgj9FQaoezfP8nGP/jwwz6RW018InZ6WMsUPOLDaR0EMJTD1bbs5In
1NqGk8Xmu0tSni/DzoFwcybP0gDcwett379azlUPTDOShsfjZ8uaVWj8+LJpWzCJ
saQM1UscOxro4kL+EIz1dhdPuom44ewO5xic9N0lWCUzExHPgf3bFeC28+O/SNvn
lBpWGLV114FDkjO0FYyERZmdnn22dMvDC6icTQnDdDB7PLBcWYx6i4gsMkyI2rLi
UXxplVoi/to+qwgHdBptNsc/HrKxkLaTUEKGQ6+cX79fGz8wmg+ScaV5t6AIBToH
zFzPhskeNtXU84RgVTYf0WOaDjqQb4KTE1YZJbBlw3JlBo1+wth5Sdve2YiF0Q8l
nly52llYcPGPTuQ9Wsh8ECsOrZ8w2WYKjr/OyIcJpREHlMD6Pe6kLeApflbEoZ08
JEVfAbiakHkLDhu+nmt8ZPNyx2t1xHSkkK8c7Z4PfxsvibEwF3nrAM+OnFSjaIay
Y+6dl3/7m1+oYaU+Uunc6SV8kKW+IYD2/woxA8C6S4fRAq6T0eX8TIGbiR1UyNCC
2Urk9TMq1o6gTn+X5AfxXAVqaqgpsduslNVgC5Z2v0y8awgRzNGPfKR2WS0nmWUX
zFTO7NGji4+6wNK/pJv537IJmj78QBgKtoOZJVykfra6cC1VrxmNTVmzOmFgweyP
4rWUNkROVj7NXafkIFjfU9gtRc7XNxprU9nJgj+6F4NXwQ6uQi3sfnzjfYNRcb+M
j2OaYaEwzHe3Ev1tsk6JRkHLGc9fatWkFwyKkd3rxnnJe0B97ThJSERGgdnRAE28
lFx6I6UKN00BN6JyayEcoMRULlbp7K+P/lg5MGM9USwl2EM8ajpjLy7g5E8yF+x1
rGlGQccQCp9iS+SsUTmSSaGqqYfGTtvGO4JJ+CxREEa4KcrWbAgyNR0AzneLh9ZR
FIYZgG6sTQIzmPV1dWgwE9/ZNxz/EdT+M5kZIbrK9OzpcBmdc2+ycHSnYbJRVZtv
MYOnyPdQpexQ5P2HmXJkfpNF+P2AkU1yTggpqXXXK5Qt+QYZBtWAZoObRePI/px2
oSbL/CV/WON+Xhgc+GcD3YjbnbQf2a9ARjuuRODzKuxL9oNERDudVlbFHYICdWmP
kdu3+VTvIJfLrhSLZR9O4YATyS9O1Rpag8maKTX+kiSURKSnze7m42b7tu1Q0dag
Jfg7ajeWQ44uFS66jYUVBctm3OuH4SPsEB6BKjdfHf4wSYug5yUsrtQjVu06plKD
rBvyb3zHCyhw8BbVWEck3R42HN4yGpkUyzcmjtcwniO6MBxl+2JdN6PTFz3NVXjC
/PHemWQzPRwwS8NGwx6YsJj7dxSFy0xvfGEQEFLK+sCWm5U93dzb6XcTnRA+7P89
2GBTImap4rLXbcLTnwM44xThs9KBn/UBKosSvhRdafkSUg/elsn4Evvqk1Nm3hy4
bnOmlv4MbOFOV6lVPyKg7lnCY4Zii0tck05Y7fLKFtaXMSMDy9vPp+VqSZoEYvOC
GtYa/B9xrZbvw6qdljxsHr7JXDOnO20acxLyeiwJZb5yZzg4EKUZENDn/G/TnTYs
MiUnl576PoEyvl166Ua7SaLXEjjtqIXQIPlBJz3ccB7pBVHiXYI9UHZVVZblvULv
ywFe0CemQiq6MYYgz8svkMliXriOZy2YRKFECLPmORh/GVgIxchfs1REGtfuIuI9
eV/Om7mtG+RuqsY5VAtYLQCPvGm8YkpafFZnHsV7qWlYu7pHAyVSp0z0/HZHq1ks
rHSK2sQ4GaIAA3bD3yqwgm08Nbv2qNnldFmEz2WCZ7lCadnIu9qrVfQmyM+MN3IS
ETysLnwmNKINB8p3riFiYg92f/aWix+2+Oo9mwPkgrgQX+bk9MbTKWyR5jmllYls
DpovVO02H06LWfkysBOYUHEr5EqK3kZOKRcdmUf9788Yg4abG0CIFKXss8M6iiIF
5/FDRksxIdnkg8DwCEIq4boZAqpwKMPIGbUOD7zBWMWRWB+96SiVBVVkisHwDgKc
HbvbIFL0u6DfKAnRu/BY22X1ZnlKbVHn1eovHXROmxpNroCkhQhXDSVn6kc1j1qq
UMYCf7egsjXgVkSJlJOf/nmxEGhW4+iBAFI6gJTF4ImYQkxLLepcq3BPQheJuz0A
9E/yeHM/pRNVswUobRlyE/mwaxhVGRlcqmJ1RBZnD6jNBsrtQM9xX64GClxpXLwJ
0lvWAzfTUjtdamxOpHzulT1BsDu66Ya02nXTzJThfFGkOFvWzpMmErvMKWPAIRFg
ZCyjc1jJSWIU+exEAidbCFtxlWvIxzgjLIpmjFOG5NjUndEeXO+uAC6gKebYaiOK
AEE3l7fNx1X4Lu3fmJRQ953fcc87pdsTq4UF4q0UnQhOtzQELiYQDSQ/tJbnpV+2
Z4+axXXBtNXup9Ieu7+tmQGAuKmRLBPQqYoUW+uEoKN7+UTu96qAfpOscrJcEnxt
qNH/rohqnfrTP/OtqqfdpQ3bDUpX0/OsDcDQAihFfzn4yadukYqBKqbeTdqkN1n5
gL2L6rkeiJeALI5aeQ8I8SiOqz9//BMylqrjTqi24D1knpoLAlBKkKUhPFzcTro1
/EYY+n06cuLA2pbOVON1VzGXcicXQmwj7ao5SmeqKYyFx7qf5BB9MVufytftFT+t
rmO35lt+ABB0Z1BnvW7DzK1TqpljEnfoE8TOQE7ZWpNzSsQ7rwkUaqUfXQBCrHsw
cJbsl1ejLzM/mIxe4TtnI8n8XXXMnQQOg80MG0/v0Z07a7jtCyB5zfNekmOf9IrP
PD2RiSARixfDs4FOUK/4/w76e4kaUzjQMpNfudEQg8R3lIep5zE6JzrhfdFQQFyI
ubs1HQEzQ9vvVBsogk3ObIIPbclQ7FnQZSXTNd0yuTytTpPoDXnjErfNbOl7uYU/
atxChr51gL3uK/+GFSmljrXYf9M5Rvk28B7HcVuK9ngrhXc1bH2dOdwDAQdQVxVd
PH9HD6QV6xZOzn66QIPfH20YimrDKKbBf4EGKqC3PZpI0gCVhvMqgJQXzmOPNVfE
KwOw9AbCetnvQzUHucIw0TUaE9keP0iEreGek/KVEl++jNjz9MCFiEtbChqe1aDb
7bbiALLK6x3Ur8m4jgGIpMjVjTGDm0sNmWi8t0fEq6WDNFY49TtoeitNsjBQzrzp
Sorz8/iuCZdcwi4jchbiq8VI+1xPJcjEDaL2RXPt0l3p8xB2wdy+X6nQBAWfhkFs
viYbV0QpEcxXwZcenWyMnh8sAfqoMnhnLoskKwCkEgNHBSEcbcl7i2t0srnliwmZ
xuqgKpe4/lvxDX77gGQub8FZ2rnmDdGxqrLViBL60mcSC2BZCr6EyljZ5zkS+6Hp
2i2PUzZ7Uk8V9dKA4cWfbFeaGcllOIbrS+mAalkJKA+CzQMw8Wcrze/BseZLho+Q
6ES58+Y1V1FA6PSArAF9Z2u5ubqfN5H8CrV35cSeXBrltYbousiYUFNsDW6sJm+l
WbmmKI9xv1s1LL5t/98JaLsIyXD2Djv2Rzkcm+5rLrBbalTY9e5OKt+rNM0DrurY
pwnkdTlYM6qXI175S5A+ovmyPe0KYFMQEzjIQJ3G4vhUuK1mkbERNCp56M8IJxT8
Y5KHfEFS+vleMiSGOkJnS/Yq0fcu5nwtrlUWAc1D/4A0B7xclLTSEurN3YfUlXEx
CEtHkTA6UG8KJUBkJI3ffDFeWOP/n5D8FKApVun8zfijE6ckR9WJFu2FMvkKHnBX
g8s8vyits0Y2Sowk27Eemu/oOOgusprB3qDYWq+WCdL7BP2m4LU2r+8qyEXc+0S2
Kai+K9qozuxdYH6hY+IhtlT19P4pC9KGmw3cuFfS9GtZag554pD/m1KtoDVbqQeP
ruBnaeJ7K/qiKc/nTGOuLe9fbbFPfeSzqvFdy386zT/5CO6xvTs/Wb6FBHSx8+p6
yfgAsq1ZuD7d5kWR8zdlV9amxhR8bexh1Xi8SgROgJQ4rp52h3wcp+Mlj4fCtSqx
XZ0ekGbKh0fXaUjdJ8mLxlKmh+Si/3cVaVBGel5qU5LRG968R2BOUimoQ1vlb4RC
4hyTydxyiFRNw32w66Z+nq4L3Jw+u2Bfn3gXXGsQ1kJyHhJ3tjK1kqSLEptZnZrV
18nv3AEwuy0AWOEcMuEOHuwezcsXl3+Sk4MTQgzw7QLbiXIuBzZvWEDHhnfTZ21m
DG1/kdvjxFYvNvRKSVxw7qQnW+p8h+uIScGZ6dkAfFZ2Lk1gVhM+xgGIoNXJm3VR
8wcnCVGzuOb0rt7bsZa1fsTsxlTgBqHLjGItmlktLOUhShCe2qqZzQJgWhlnYSWF
QXwFyX4SdUmuJ/uLzZupP6Gjiz2kQTzeOiFKku82eWsRA7aECMtbeR1w6iTJlMF5
3/GraNCXkk8FOu1lpzbNLMLCYrwoDNu245A5SHbVsXyFa2L+ipMgHe4zoie5/VeG
sxk/yfYaYt4vT7zWDnMomj6FH9OCmHo6d+b701BrDMSGVLj30cRmfYKkDIHd0hFB
tTQi/4c16KR45fAaAX07iTir14ImducchJZT/H+sCsLdGedWNCj/mGPu/lG1j5wH
z/j27RhfUAuucQk8PrMzTsYX22zSyUTzF8nmRtxmaBiwK2LE0PU7o8GDN5sBSQHU
N9HqStY2EKEqQX/mcRvzROgdATJxhAyHc9O9ZFH/k4FaUgDtdk+yNIftKGLnuW+O
1c40zY6oAwYFjwXEtecvqgEwucMfzsj4YW0gy2brjJ+5eCO0SUVVqldHQHJdJUd1
6rjy1+3UMgmDr8zY7/nR5Uy3LVOTAnr+KDOfKgJwxVhyHe9YVVTDLkpf7bHlPnUQ
eemCSFpJjix2j07o0DS/K54E5HEpmyRKMvaCYwdHpFbDuKTjU7aTb/2tMyBPwTW8
bFpIG8oJET3aARTVaDoEB6BsJFiiEPpBkz7yXxQd76R65+TFAVgW+jC7oryuwUej
2R6s8FfwjG3EQwOGx8P3f126agNsPClSg2v/Rc/u9HNRn44DwRLQ1wFFHqDxFt/S
J+WMIui/2cUsxfC70ceqf3eoZobi4jVOb89vTGp1E538qhwhi9rkeOJFq6DokRBr
nvo3rs8clS4rQJ+L8jzPSdJ+EbC96XdDdZUez8waMIUV2oU9QIplcMI9+Qp3ueVX
5j9lhFAV/vTGmPSyJAp9jxpuus5BQy3Qjkr14jQsDiQAml9t4ZtlqEB3yHTi6Hzs
vCifaoDIG7k1LDDypq25o5u190R7vQ0jOiIbKlsCAJUjXaM4uA8FzHfhIC1M4OaN
1mW1tohU9zJDgK20xqZtSZhXn6dWEIxvMPbUC2yayTgyrEM27+nKqJbt5RUzzaqs
7FWgjTcIiAr1Y2jzSZ3jyeumyjLwbXjz/PhUBX9qHkdW1lPy7RXRzMm2g2bI7gUS
nJ4BYgrjJVieD0M+gIcejjNZIu9b2948/j+WDhhPhH2JqmTDG2suZBlVsQybrfv/
UgBtvLBA+37Zjb4egO08hEY+gaiibKIseWfMqJMn8Ksk3QRSjg0a8+guCPZ5CHtd
SGFfjj/KglhSHhvgVLCio1LYSbzZI2N2IgKIotaq6ceBnTMSJydwfDztPe8gHsNB
PtC6mxb+eQui+OdGEa88mXoZgZnY85SyKYHgRk/BP+im7xFrUsRDfXhi+0WR8M1u
Z1mULmaF7ZL6EEv6A3vBTK/NpvA/DhJdQPKPiCHPXVL+pbUHmnewQJEKjktkuvtr
M2d+LdJnRqsZLgvvDTMMoE7rkwYfTOb7YThvnVwL/VwYru1a+kY/OjC9ZB6bnxL9
QAloWBr5PRdFdzFZdX1nlZISOR8wn/SiOxV3r15IHjBgHGqJLJ05Kwz07Duttvpu
UaRsGw5XzbPsx8bIcAVK0bgmjs5vsGrh0cqNNAJmldo9t9fsvlf93fKjGi0j4jpY
ehSxj++J+R+tP3/pyr6ue1yo8xgi3S4gsakIwBYUcdWOgq+Es9AjgyqpRj11OhRH
hFfWKe1Xj3NZ4AGkcMgjsoZFAjDDtX14lAJXoQnppuulb6DoqULmpvxDdNQII2GF
eRPX/kKUhnfW3x4r3dQSHRo5GruljK+MiE/2hLwKP+cDTftbWC8RJQI3NrYLN2cW
hQngWC24IPBUel8gNoRJjhA6tjZN6jPUKI+AgZ6uILz7hq9WCVBvp3l5unNZEAW2
lpWRI+19tx+zT/+mPZrggAqGYnTX0nQ1Bxe12oqYiZtNYKgeYSNn3uvm+A5xzkM1
DWFknMBb0sa8VkcyhYcSf+wm/YG4SvwSxMkSXY6NnbSL5pSYzQxOFdPk3+uleou4
wITzfm0H+P7JEoYhImgMXIF/wZIlE1z8AbIi09tkUtBh44AxabnnHnSrdr6WXm0S
qGINtaEHUhHWbA8w1bPMnwGP2tTXVNBK7CI6q5RsC7AurgT6mlCRFRawbzKnvWtg
i1QIs2zcRZ4Era+xKUiO0GqeEN3PnfSKT2c3beQIMJlYDOTJo1oNTMUpjiPgpHV1
9QoE4e6j2ZESfD0oWg+adk4Feof8kUB0+kT/Y+XzsaVndyXklDCeJRr5zo5w/7oe
YrPYgMuY0qaRHInAmc5JFeRjUNu7gEBl80Ar7XbzJaASxbRcoEaSnTHhRnephs0G
dBQMslhXGbtp6/Ah4TCUY6uv0bTA0xCIHr2rYsMz2s825Qm/lreGYMgajuTy2lFn
swDFuq7bJJPuMbPh2D5tQHXwuw6SKWyQitLeq4OTQo6E069sYRhUQbQxkDn/glJj
0pQRXUTTK4p7Uh4NU+FJrHWAqcErgASwGcFXn3gV/yr89c6keuakBwqHYZ/p7tsg
ULX0V/YmMYQ0Ra8XTmbbOTtXY8HTKalZ8tj84+GH5zLJ+NTB5yCLVBG8KeC1CccP
i2QDXlQ+GK7jl+4Lf2Rnauh+e1cZCZjmSprf48nwtKCZuuWYJvW8PaQ0UmOapsQF
uoeLXtnMGmtH+sqigsI5SATFBgveeOKih3dr44z6CsPqER7yyqWGavgveEEMJII4
O61lBwrSUoN21gxhdn7d/L/ianbtWJ/C1L/qTMrahFF+TRUYoPbtjdDT3Ao5TVqT
XHcYPmAsSVIN8YRQXNle8QllyHbH/ccH1Y5oTpjvB6rHTIEHqA1IeamILcjUx9d0
nEqqqpuhwppgQWPozLAzR5WMQM4H61pGrWQQxXDfbe7J7SBojNKJok4DhQajnrGz
PtJjqFO5iWaokCaZsHfHRvclYskFf8clUmp90paVplZdPSImXLxZNdCDuHj08WM3
AG1m4XThlkMMbzbt/Sva2/SrpQkcsvltEoEetpTb3oSyVifoCz1OzC/RStChUoiM
uwLn73nKqrIzSLoluoKayiVfE13wUe1BcZbK8tsE6+IsVCdlacHt22b8S5Vm77uG
yrw/nO/KGjSSC3XGJ5gG9ohpseJ15PLIpSHOLqjoXYlO9tKdyI5MoA6nvvyRGZij
aPgBgS7ksdsbTGdYKUEpXcAtIec2J7pWlAXXVrHgez+FwQO+9ncOAWOkCseVW5fk
eKWhudfCqafvHaki/ciKdzjX9qRfFlBgo3xMdAbJB+eLK9YE3S9QcDLXNAVE/TYM
bYe3RozirD0/8FPDX1+32tN8qDNTv/YIZVHaQ5RXDR1my2BhUgumJbB7bplw9tYz
nKrTzADvVoJZxLasS+aeaVyfjMBxz8o+S1xKVf88heWWHeOp1dzWRjnpYDzPEOlJ
Atw5FKp22ZAJuXJB0OtMzlcfN5Zfx4Gs5+exJ+0sp3LicH24H18Ac4cZfSr7qExl
fB4NJ8Io4YPEG6qgpN5YLmiPhjFiRcdNklrw4pwsg0nY6U8NPcvGbuFGH2eT8w8T
WeU2H4T07jON6ksVHvbbKtprtWs8Iicxg4IwYe0aM9NvhYkDQ3Fne3QUQ7m6AKh4
sZmFJ5bzymffllIf/JyNDg4fWRXX7qycCTkpkOVFexVlcKyi6h8iZdXPyNOT0sy4
6nEFHfkEV0graxZonNvjVqxOSe2drFmi8Mq5S0vkx2DsrRQyFePLF9SdBZqnKEuE
rXeKHZc0haWsIhXKM7iahtn1mJSFFP22bMbpumR5Lf8zbN5Geu/TjHtXCnx+Tv2A
D32YpKAoFGQwFpbZOm/lkqxYlfDphI5Evz3niyuPuAwD8fBDNzZz1gaJkmZepPd7
Q1x80NtZHXeHXUEH4ekAG8fziCgMinp2OgUHjASIJglV3F/iXHPcW7WpVOxJxngG
VhxJj9+nDKMGtSVWG6elGwsEj1P74ueDbKdlcS9Jzyb42U8uC8nMKxH1K6tmE91b
1bFUyu06SsRSm8x+QUfY/bf3I7Zjr0y/1SdOvhLGtRgjcWoZfqF8r21BqqGdhjHu
UBcBVOaixcIXuqf7iZCfzWyZ06eeW/W46Q6Q98SYDXZ4T8fejdh7tMSCl3N6vkDS
qSJC71PsHBHBLsamDGHnJFql+pl21T4FZsEJqrwS7BGoWvdeAt1lzd2NOwwVCfp4
iAdQ6j7LIttiR2WKAyebt4llQK+Rj1JoDMwC/PEIDzEK+EDMWzKwDpnN04tjZb0s
OqfopilVQb6o8FG3OmFKQP9ONtqRHRNhiGqAZzAdN+Pn/3a7fouJJReoRWypKNoK
Yidwljibvz+rtFgWr+Gzj1knEwhcfW5bA4B6OEbeSfLyMGDbQhj2pak+fL2wDpSB
mLsmNePlxwVErqhfB4GlWUWhLL+lxBrexXY/96HkfIRVBKND3dnvaWAq4cTZ18XQ
RlU1FRNAK41hzSVZBweakPFHKiIsR7X9imds3dFQNKtt4hOWBtCvvvkVNyo5Ljf0
QuoiP+M6kZKGIYgI+oauqEO1y0vj35mXUTMyx0qbAuUIp3ASoQVmmmmEguI+5zCO
UDqcwles6p94owAQsZljGYQROcmllbCtmsc9Sv0gjTtiSRtjeuJLpx8CjPUjnqvZ
RuruIhOR6/Fs62GePWjZEoZMQmpDjhn9vE9GAF5oRYhFMKuMhKz1NXB2uGI6ZT3c
gs/pgS1rr3+zyGLLxLobH5q9PAvU9qLeu658sYZgOww6juxkMiAxkXxnWCeowifB
mcb2lGpaa7WuZDJgdIqt1TacsHL3Togjo7ryVJIlOhUM2x2DqoSFljAYOx0rlhDp
MdjktiGAUBFiDPW62dbChKukwVcMWEXnLifltBn+/C6C6bxkDTXTYU9YFhCzG4iE
GvzKS+iBR7VIQBRLp0Qc3PfTTAA1hE+9cZGChI66tAcTQW09Vf8+kRAR2uEuYudA
t8moF3n+U0mgmbyUoviCof4quogIkZK7hfsPYCHWlFwYiK5Zbl+K+UnoxpvQt2JN
IUQDL6UDnWLLE1AtcrcO8CgjeVjHyrHpwsxYdAbUM4dsh+1UpsmuT3yv83g9qp8Q
3i0eYyao97nCUIEej5/DF5KRQWVlM/bMiPLgtfKTUNX6KsW6QifnVXgJMFZ2p+fc
Oxh//9YhzlSFzPLJ7I6yIPbwuQ4FGKc8zQ4Igyq6brZ6BX56mGbeOwvUyL0y0R0a
bpmrLdqkRwxC/3BJYbBqwDSq+2rp14ns5WRHcx0RXsZTpNELyKCUS1iQBxOC2EgB
n+rrDyaTNJYPKxseci/Vug9zptm7EYOvVhpDHYHxc5/24xXNl33GSDGaH+uy5Oob
lNpvJ1mIeCelPApYdUejgyvs71uUnYw/8IlHQ78WnCLPK8KyOYyhGKOq+qYWWr4A
UiRhLkgX6z0NgI4Z03OIb3ghQlyWWaCVuGTe5UbDpPzzSJ2G1yW+URVRBEhv2Epk
Qd8XAXn7/3Il6bTcGHHz3tzpkCxFf7Cf9lbPDyM0cQbqKRtKPpoGlO7ZkefEeFYT
PYiAkJrtKrqgn+Ycoj1SD23cypkak3zilwYAcgOjbkt7gKWmGhu0Q2xcxpWtSe86
OYG6CzP1nUq1SV5/Q/oOIaksoFb9Roq7RiAWnQN6VBtK3sB4lSqCIb9GlGNEMVT6
Efm8lQ9Wew+WJf5i5+odrIUeA1FwOA0gwZK0sxDHM4GEtbqNkPf5k+ns3S1yhCP8
LpVbTnz7khGksALaq+uOJOM8yDCsDyAVAQRYUQJIEQ2TWYl/y0qPkmq+blmzHMJO
kgX41si0gvf8RqaP/g81pXgyiYk/maYbBaSg+JkEx4LsoggPdeU4nFOrO6h6gVjt
TLlXyg50AnTUuhDVjnaYm/I7l7d8AUO6vPcsl1YrJR01xSctm6J1v72woRIBJqbb
wlukA43BmUcCZwPbcUg53lBjdiKZ6I6zXI7HFrqrXtsY3ca6scDlUPkon7i1ZPz5
Ion8VBdxX7DIu5G/K+MyBEEz5NAsrXppIc+bBW9OotpMOWVyANp+TAktWlySmTWQ
wgf1XQYCIHMrebEfjzcIQMCQN22h/HPidSqWoXSZC/rqNrukuMtV3RXNgFCQn4dP
+sXRT1vXvzWHmt+hb4QEXndJrud+znyuF99KqZdo79NiRWquJolqGG+1w6G4cxCK
Lrx3U1t0EbFuBHQqWO1lOixjgRcR7SJhrV3S1BfidWS+76sIlqRtCdRcnXiiy/rx
`pragma protect end_protected
