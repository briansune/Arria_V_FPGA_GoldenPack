// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:19 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Exp0lJLWpQ5+jY957ULEKMbD1Bm2pJ1p3KbEDzzR3Ejtyhu/vQwgrCUs9vVIJIqZ
0gTFvPIau64D1bhWONVqjBjjYawy+Jg/QJ6K/l9SZ5FLt5ETE+c3OfQ/AwB2esG0
SfiYZrBIwk8KwLLhbJod4n+XN41axvDbYuQLEUn66co=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
9NU0gmRm3rYAeq3jlT3BERZ4wsyZXL6UOs/kdCIZwSU05gSIFmn5jP/n7UvPRG14
bD26dDQ84nf+oaz2/886Zr3ws8UTv/X6LZl2lnxLUHzFbD9y3+1w0sJGek0hM2Fo
I1V1L+fPV9YvYhB4obyYN07PsyLp7LMXNzWJP9o8SyMBNYLu/ZGYXe/o4zaC/I5S
6r/4szyLa/69f2UEnROAYYTXeq9Mo2qOsf/dZ0KBaKVgRwe4ihd/fjny745w9GhU
lmRPSTqAqTc2BRx33f5sbuQ5UBbpRAHX85c5TGsvVNr7HQGP5XkTalhQT8KaksQX
SBnpclUAPOiMdMdtl+DcWclR+41Mju5toYdxwA6jH9NGOVshHRhPiYf+FkzcSdm8
nKxd2Yy5k8W+O6tCPyf02bo40FUdhlobaxx+awXpvdzwRq7Bf9OXOCUctlBBLPX1
athOijxW1/JOFWgLf9S/iULkaRM3Qz9XbldQ3fJb93ydVxKmq0sLI4w8dV3Vpvz8
7SsnB8MJOG31ILR7LvF0UMajh4yve/BZUqY8J9A+0uGvWj5AfMFwFziFSJNSRB+B
/ihAETzrA6P7w2nlYXhdS5GcIvbeyCtu8szBnKThxqqQo4MifJVjsisJOzsNKMX1
5EEvSvrfdPNa6PxcIJ1B+rJHRZ/2DFVmU7mcmBE5FbnL9+lCEi1reHK6vJjhT6P3
PeBgtsSV71phdN2Nmpdb6R1ZZvo1duoSraBdMLN13uEaSPY7FaInM2d0bYaIzjwa
91hXeHrh/4tfXo16UDs6qDVoRfdw4p01FmXF0O34IOaBSQa7QrEh3a42eoRFxIEO
AXkqhPNy6IQoEtR9eR5UBvd5oJrpFXZ6nov8lFtFc+RSvIKXwjk3rjVPY1fU9pi4
GIGfFdZMhZ3sfsnolIDjsrndKjJzsEVbKjqvrOJ+QZm/lGzShRJr+4Pq5yqogpHb
v7XF3nRcmmbsJrnpB63QFdINsS6HPUZrUZ9D7Bj8PMjnUz6dVXeSRjrb67nN5Oi3
YWKd1cefdIezrNowKqHiYBGOfiXdAOivNQ+PBuYEc2I1uUKJHKmI6BYtB1HaKNE6
ofOeoWFEmiNHhNsLLpwFlZy9CzqhK5eOgXMAdSn+eoNViRX11t0nSH+BRprpyHfT
XN7E5gjR934MkAyxOibaeGs+LecMscQ3d5/5N86NNrgiwKWOBqUeJCORU8k3Jz2w
j2Lnn/SY7thfCn6hCMuplzkvky0XE+4e5BctiMBDudLtz7wH7LIMfQeiGXN+mNo8
qOqNkjD9v8Hx63vT+DMrv3rnDrtc3Yq5rJhzuv7VybyiOKxJx/VrTh2v5aaWQdSQ
mlJsv4mXWjZI+hVl1tBf/UAdRFHj7BGjN95+gAMC9qvLLsBXNmS+C8c1pp3yLWU2
D0TI05ycnaae0mezes9nhedEkn2se69/Q3WsaVSAyXnpjTJgf+KCAPmM+EhVY3c/
FScP9VzkT1BUtRzcGNxAMRgHnsecHoW/h9n3G2r1c22sIg7iQLBA+MpbeU9he/Ox
wOcGBWGd/kn0JcH7djDbQ8i8YfSMsYyT2PSdeanGRqnSZfdPyMp/JT9xiNyfjmcI
ZwfqT1dJnjhigxOO2So1fm6DfD9GB6RLw5Fs3JwcuK/GpXCvOj1pkcsFUcJPBJBK
g7epdd6YyqgPcEiJeg/KryLIA5rkASA56XrWuBblNG6beKvl4HY1pYKglAehyzP7
NGXYhwOhEzi5UqHL5o5KX1x8umu8pD+wrQDJ99+fteSTSgA1Spz+Mt1zzV9Dz7sa
ljAIFvbKY1+SDUic0suU4FiYPFIAiuj3BFO80aAVb6xjKj6w/iPBOaqhY9e6g2ME
rLcIjHKq+3eVURhwJp4pOMwMOyCq9bQxSwXmRWoQnnJqYSBp069TuFjJ0LW7uvvg
rlDImQMyM5yyihDjnRQuVlHwT2NRJU3MSEZ20wvS9S/4/D5rgq2XFkSRyhXFwcHq
WEEJe1b2LOXudSHHDo+5BySZrh5u908ycD3dwVTAVoWiTchDNS+asnvCPaLoCFxG
zEc5ZNtNYS/6ZnFs5dXeXEXRseIPp/dAeMPu8ljB9C7zoV8m+gQsx0KfpbxGgonr
HxFs+YuUqRrzhmnZqzONckXZHR/4r5jKkdsC7yb46MQy5sCXDCw/UDxi8Svp5Xii
UQycp2vEeTQUkWJ0GkKU7I/e3sBWSCPsnDtP5qHdSsRFganp2debVZfpebucteqw
gTtjQnnRuFe0CKehG/jeFj1T4ltziZwOYp9XzpfIByvz4pIX1L5zHb2VaSVVVvXl
SpsLpaSWpnfRhPuNb6Js3fdS5NzdXDcwYDAsSRGa7uveRygnLHUEncMefdPzIkQI
bmvSIcRTErM56xJ0whq3SvCRsXtgfV9pSabkwiQ9fGWhViz0YiCEdqI9VmNw1L24
Ip30nQgBghyM6YQDNcima2S+X6I3m2DdOnF8srqDnGrMrhV3nCZvU4lm+U85mnu6
SxkXceYHlidW0kHXJ896HY313PoWNePci2hXW7Yv2wSiK6UqwFG+zz6GZ3FcVJoc
M335Znzl9Jl618KCBeWiDLdeuKTUvMjjoOQ0OHevCftEEVw5hV1kyVpZ1oD9L1Im
GG4AXWksib5wISDAEY8xJBIAuLPmKGHsQmf1U+tBnpaTqkD9vuRerg2nT/xUYtMt
mO8HRIkx8VQsf6iF16PJAHq/QNrWRT3Toa5c1ESeILBp5SvCMXyBBMr8BiBFau3n
q15atiY7Dg6g3sBJdOLZFyI9UTKf5RjTv6Unomhf5fKiN5aBkZiH9VlPiwMaQZRq
LdGbXdwNZEvecsN1FiCYPlbgytvVhNXH7myrUEzf/KS9/RXn25V9BPx0XbtClv1r
byEHst39Q1ZFRPkyEU97a+uNdVQ9cZxwoONM1Ztk2EUJywpll0ckQXKbqNm/f0wY
rbiLVTiN9GWyOzmMKUrAsTPfrh1Yno7xhMkwQcA8JaodSW022+PfCRrlRBrcsVTZ
hkCmXeZDEVpcVV4iFVbFwgegXA4zOAUG+N8I0GNNFVtv/ogaayD9W/8/vB9a1bTT
2767iUkf4AsOP3p/JhZldC/CRTCeYS9q/PfPSfwWFXoOD8RhUBMI8q0W6SGnPBvh
dgyVj5uGEapAVpteV1tBfuhIw331TbaHMFC/uBlUVwivRbGhMOvH/3NjwmjTsGFa
35YwiC4Jqur4jw///E7U+mGHVstURAXU3stAzdKm6V1T3EfC8jrpVKdDlK6R7Pvp
Cx1t2W9rQaa0p3PR16HAVBB1IlJDiFwoM8xxZc0QFbGNlHdF3u4LZNo1dY6zwuej
qDmKG8LtZVYp82haGFiP4Iljd1e+9eeVR9CYaMrQGmovwZwu3s5kSPYrL2quZhoF
I1t2hN15879cQ8QoduU4/2nyy6ukyejOHmz9XzzzHh/czK3+Pi2v1/jdsNVNzyWJ
y08NsFzfPBfOAR8RP89eTTkGKSd44zOVzLtqWDS6vXlISpQh0pvjKnlr7XkkLNJ4
B4/w8o5OstzRREzX+b0FRPVz3D/ZPuVlQce9ktnEQmLpjgwVEWzAxSpVF08LygUm
2qNyvaPqbA1ZWq64U6drweL2UGGhMJH6zk2qRCW8Mn43R/L07Owvk45gAGBRhq4z
h2fP9R194jJjqrACYotVFAkRtRhJaGE0Flif3ElwZNaz4z3jJ45+6QSwLrBgscfi
mdvzizdKwbSChJq/hCYGGnoQE/cn6hCD2i2amYYVkcGQJcIsqWB4S5X5nYm1g7Dk
PGZI0Iq5MhNnDERrcaAPhCbTDA4g1hu9QRRUWdnbNRNH60UbqKJUWj+5kjD3Kc1x
YVTvkKPXwBXXV7OtjN21mgfRAVzSIMenj5H5VyOKIhWPX8ahxsVKd07tpKxHbzZm
mtc3FEUnM86CzgFewGOnxuFw6IxaN89A0RjE3eGtatkn8lk5nVclAQioh06yzJL5
QYTp0NSnVejcUrA2q2clI7CnuiJf1hmfV6rbi3pOmuK+xstmhZnijOYJPSkleLmp
HdGKHfn8LP2E1vX/BxrDYmJlxc4kElbO5AxgoADjcu3iJBJWULIyObJaez4BLgrt
xGxS22g0y5bU9cL0TxP3XUWRzo3OUSQVUYi7AT37L60xEg08aVLg0AGxXWJ7EMzB
ww9A1LB/TwmgT9KZj3+OfEzYwL5wOVThBx9rlnrbZgTp371MSK6uJb79181JfOBq
a1ouTC7iVAAn6Mrs2n9M6I+n6Ak4Q7qKSm5rz9uFx32UlHx6Ddh8rrQh6G3iKa7F
lXKjRi+PVlzBgN7/iH9OdZvw8S0K7S5uaaIrlrMuGUuTSQAu4GIF9aiTOY+di4fa
TWlZVnRRkfS51k1o/C8fc9aPj+Sz6akNMY3J5EF+xnkaKN6dFTto7McuY3WCLk1a
xuh1m4VxDmPpAXIn2DN3xKuTUlqEU2n3Vpjlb3+HGMeXERQmoLU5EwAlo+7/p5Qa
5A0xN5FSWBhkbOiQWRqWs4EJGe9PT2HJIog/7/gV2S/VPKDRTjasDPjmOGf1TFgo
UtE7rQ9KoVlNjgfeGITRAoB4p124AeCZP+dGIvBr+zs/XaRd9FLYknBbXnfNSwQH
rgYlE8lI8/gaLLm0j/d1uxC99aO3NlyTI9uzZ/Tp/FV9hHq276TJlQpCPl3NqSYo
uTu1p2B1/7RI6AGl4HzHr6QLc+7DwjugtVM9PxcN2CDd7/LfPEuEser9uyI5E7/v
xnp/HAk7MvemlAqFcIv+axApM3NLm0j08Cq3LCoL+XBCzf8oiyhSZYyCCnDKKh24
HqOa1GOnu/8uKjj58DTmZKB2NPUfgyZ4WSGiTSOG6fH/1vIffyrrXgMyZrSTE6qS
PtBUxu84v4imKYIPBdSntDc2CvO9VuqqYJ9LsCZFrrPd2t5Qle2xE8mojPJ06V3r
GRORdX3MUwldCRPN77QCfTYS4/ZAYQSnfcwkY5v4rH056+qwnGXr/5bwyuTPJKMU
sZkKbZHxzt86HpawNPLwRQl5PZ3Lfij89E47q+kq0KO+3pWguTx0i20iHGC1NM6S
dXgl9npKiXOdnHsdnICz8LyJUpdbo1aRuUwtuirBp7IPpqqciKuDhPPGbdL7IUO0
26NpnhCMKj78o7lkkLiqFsEv0zlZDjmJUOPToJpU0Tl2CXAup9D0F19VhEL/TinF
pKvh4Afm+Zt+hzLxBalFDM/c2SDMyUSSkkBxj5mgirVAwcHrMMaC0LXhd+u81e8K
I8jN7MHFqoyfZQvMZnhJgg504ifKrQNM6RIRkTdDaPiPFcQ2jHJr7KbqFN6ep3uS
LRqcA/IVPA6+BV+rXKfq1iWjsFdMiySR3IG2hmNnprHfzFZ31XXt6MNujpdLMtgX
MGsH8B7mAbASM6y4kl8wEW0eYGdSXNWbqIhRp/9QMUyA9Q7L3BPgBK1tbPA0mzhL
IEWFlxTXaRXRQLYLOMOOhH6Phb2bi4OC4a8nVS74uR5ErDcQW8t279WVTg4QFCtO
9o/PXeiLCUbrvuz9CwGSDjut9durZN9026qva2/EsK2zQFc7FuugZ7XCCGKPrl+m
60/QN/wW/1SHrA/YzGdrc3TDbcMzKSRw0TQ7alxykuiXRkVTmeHU5iT7qkbREZCm
cFgroPKmXllCMXvb867BxXhQ4f2LP2019pjQOKtXw8cQz+i6hkHtLBlXPCCrQHfB
IvzjUbEy/VQ9qV1UhMwMBnFHXfLGbQzZS1nOIhncj79IVOGDt/KBsPqkBoQWvoJc
d1m09MmaP1FdI+3LMpAyi1/Wz5+gpl5cwV29Rna0hbOZ4l24duFkfa9ugipPDQsW
x4bCIZbTbj8N7N0scD7iY7iWQcdTsxnmlhLd0j35x7mGHw7AaTvA4evqw+AEYbhr
Dofyz0V6UKysi4y+s9hQl2EXat4SMyA+s57eh4M/96HtNV0Ubl2JZ1TzZJVL26i1
QEYj0KGAtf0dMXyOKJJ4P+zeSrU6aSzGR4dmo6E/c2qhaxYwTQDI1m8KD+qTO4I3
rd1vokdDNSmULjCVNt+fq+fsfFGDhcneq5UUPWUp7Dr+l/Ul9xiBRdEGH1i/z2L7
y/z1A31EnFyBzSYMdvoJYPPIFMD34dOXxxTPLgPIYzPm0lu8nHJIbW/WJAgh/E19
F1uaI9WJRcLrRrqp2pWzC4A8i5I+1De2jtmw3ypn6JpyIGB+uFp8BFfB5WztDgK+
ygnk9xtB27ZL4XhxFfazoTpB5IVbtSWS3/HjoYk7gWAYwJux06RW4YrrPbg6xAJ+
B/rFQVgRwgs7/0J47YxSdvFMBbiX4W8AccudtQP1t8mvpWaNNoYn1mt0TnSFXcri
6AlKClOo0IPOHdbBOrqQ8XT5Ey/PsieGUL/kawR0BrK9I5lMAgRz0Q0iRgD4aEHB
N6e8ek49S58Kh3muynkxBLRPk3+gD9EG8eHV5ZdCDytJRnaLvE2G4B3MrI2RsYTK
YxYBVgeo1lrR07CEzJkmLVoYu2gDGARxhlkWsdVhnvwT2hJ0UBN49WyzfrstaAG/
D/+SHwN5sEoHJVAc+UEvOkq0draS6lIgS1Ve3ES+SS/LeXFWbVNtwXCIKDMoard9
09cqTtlRDpnscYLuhHXJeDvBfdlsOSod/Zqh15jlZ8nuMMyfm+5K7efTqqOrSai7
lHKNHCs6ukNFtjWPiyTpyqIrAg8VBv3dxmxyDIMgW9bZhSg+P9PTJZqM46o/P/Bl
P20SekhGE0kMLMzUtuLOsyNh4o43wbLfN0Rawvyf/i4ih1Mes9sZ1q5NVwOzeWAv
qlXII72OHHY3QktroyrUA19+EQdp8j/cQUMoyc0mD0LDV/FGRMHKzDdvyrFex2/L
4UWRAM3UhyOTpk0NEGqksZsKIumb9wi8Hli8GaJXD8GELnDrDUq0B5QE11r0kllM
b5OcPRvdsX1j9ZVGucTylb3GLwqBHMaMNKKsrwIGMAaNSJdsD1hg59w1tZIRj/4X
HdYLR8v/MW971k9EiNDPw0fjHTn5vzALpAxu5i9+MSymzwRSXFcyHq+o4tBxR+IB
9H8xcPBHjq7EHpy4JBWDOSIa45BmGdbv8tSDXy+eqpZSHgAJzGfma7UFEf2V1CbQ
mntgPvGAWERMIfZaFRY9GYaxWeoZy4LuHUeQFtWD9QSU1LLgsbpF5BSDZIGxiMby
BLV+f8ZDN68qo0MzYz9x+VH5e9JDeSyHWF5pAHcdMv2iYj21DUQOn8HGWwkAO3Rp
NkA0K2++lYPeiiS4goHDz0RRtF6ptNTPVHuOUjsb3vacqOD34M7VBbYJD+eqZuYq
uEUOH5mtWJ7mBxpX1aWBSMfsh9DBFDNDM64zz8qAYP4s6k9DScTktRgPagKn+eLq
ehYre7pPmEMxkhB9XbpKy2YPExMDMAPYjaV+650wPZ3lhQPGO73/wDnYSB+Cv7b9
OkFgfJ8UJuKlnhjdm9qIt50k0zyuz21s72/2n56SjyoMvUCSTKogvdSUHUogQ2jm
1G+57DBW3HuQSGzIK32iAk1yWGkwyzVrtO4vM8Fw3QWIUfcXRG6ooYhVsxW4IVbW
5xfLWYQZ90SC01PpR/HH/gQ5vpvUoAW7KObz3xF5ecp541tAeBIAKzrAUSCc78ZR
rgfZ836i7OhGh4FCzRWnUw==
`pragma protect end_protected
