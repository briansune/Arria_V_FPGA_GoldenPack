// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:27 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WpGW6kBHK374hFzXij78UmVz9NHM7tN7LSjAeRof68WIwBtSPY8YqSg3zPuj32qe
rf34E/fD3IipYuIKcz9CS+Tqz2bmmDkOkgZ5LQxgweSAZY5R3CiNC34ShZA/dX5R
CNkvVM4f6UrFxGVJC67iit4APMp5eXdyDkS2LkE2b+g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
rO02+PqBci5PMMG6Uq7U5bz8KaGuRy7ERYwCuj+uRU925YVu8vCkZ6/yxF8tN1pz
ErMdcBAwIUeByhabNAQf6NqzwG3vsW5SOb7Rdac/lT2vC2dic1XxTTxhgUSADVFB
35YQenI2Lo05wuYwX1hZaOGjlU3Lzs+h/3hX74JSuoPMxch4cx3hZn6vfAktdQS0
mHEGpyr2ePSCdz0o8YszSKYWIred6efGpjip7SLktGd1xdbfNe5TZB95lSnFY5ZF
cC6ggeqw5ouxysgu4SzVhW7HMLtQ+i8uG38+G+1V6R2w2mxa/uUcohpEDopYJj6M
21mDpguyNX20QEp8YDAXzEktw7fk+HdBX7jVvmHstYY/vw/6zzPZewznjedAbp1m
hH11USs55TEFP+1iqzJv3VyZYF+ObfU0uFNaDIPCD1WZpj9D9q8mGdfamrKoFKbf
L9tp5+624RwZ3nULWeETsjUPVKdZcVF/Pjl/a6SraBzPdZMfWMqWfB3LmsPRnY2o
X1HHhuXb9QSbXPncjPD77uJ0dgzw4t3zhHbk8vQ4LbSPPFCWKKkNj9qe2Crs8rJ6
S/VGEiU4DKgQKgfbsHAa4ETTU/F7JXCjii3RP4WOE1eP/DaUXwf3qkXNSBSmZfCX
qTE3yP0V8si/OZIexizsTG2FxDb3BYF/zKsRA3f6RCD7uG0gsfX2tFEccwrmzZd8
VIKClLNIHqTtXIB11nnBx9TFep1TIufPcBKNJ6JSVv+wk07lDtutvDkFxSphdcw5
7XMKc95UphBdWD54TZLsYR59/hcAfYIE07dyuM/q75tSWF13pTVhJQhSmi7JRpgY
QdDIrOW9G4sAZ9bMRH1FVSd7BMJlHO4ufUWkbVOwd9Oeb4fWMAs/Z5T79tvUAu/+
eZ7C0MJbHzKyuM39bJN0MGJY5cm5atU4IxLyiroFdQhMGMXsLWHJLgY/Ex4bsS4/
nNoWlY8Q7BIoeQejj0v6AwtGlVB2Z3L43bvxjT78/vtYWhZZnzGo2wP+hWWc4pD2
PxpnP+lF93qdReRMrHgrVWEF93ngsWjDFioDKVER8+/nfxq8QMeBi3egm7g4y3eV
B6RvCdjnnGxyCHPhGZ7oRKJuWItzxB88pqPfafD1jopAF1TrrhTozyiROjZYeeQr
KJWkR2Rgh7NH7DWN4vON3pLLAr1iCTCVW4yOf81ZPpADA0a7qNT7afxiIDLe93oZ
n6juu/Baa+UoTQ1j8Kw9LYQ5gYC3RnDSC+XQ6W8s7HFQjGliGF00jSNGjzSTX3Jb
ntdAlJlwvo/c9PCZjAyhIoKXf+V14TpqAx9x4GgiJJJ/lPe/onSCchH5/HLAvIwe
8ZawPc7vA0Dg+ZeGdKB3CH3a9XZOulkV1QeaFIwhFDXcySdtOUMVfB9pC5uo0fDx
hpr7SLm7WjrPH8xbYR9/Ua96GrhSOT02jNQ+1AY6hDMZfcWjMZdwihAt48y0ud/3
GlY7s7XrZqi07UHl2grENptW+NSMuM/YK+YrQYa0CWlJJvjWFI3yutrTBn4YRRg7
1S0ELFKxpF6SU5fabgW9jWQwSHKWAUJr3kercMx36gRYV7zqN/1lc3Th5qQ+EfYa
t9NbAyXDzygu5oFBD6uePh1Bvjf4PohpTMHAfkxis3YiNvvGxesKqHgFEBG9AScQ
j4XOnHDgsZDwfoJWMpgPWo1DqieGeww8hmvdJ6PsCmaMIBbAHsndk75A+CgYR371
Z5lU8thiY3ID0AEfS8lQjINwBzPWgvJCUPx74baKgP3/GeibkznzAmjU04CjnWH2
Hcs7ZYA5LxWXpl9gElwqcEF+fyx6ErBMoWUvIt9zN0M06fhO95rMbcujT7rilwaB
BNwvs5k6t4SZOLDITxZINpMDA6qmp+tVKN7s2itVBZX3Le3crmisuH/5rKj6HRdA
TFRtRexn7HNemOBFUr4gk4g9hcWHOLj+/Oynvilut36EbWo25mbmzxU4Ec9NrfU1
dXCasXo3uupblk4SfXq8byd65FGbahtJMPBQB07zoqO9E24ZfgfDxC2moA/E2InP
JrsgIieC2Ef42521DRWwrlupbFzlrfodHPEr0SJuPwtW67lKypkMRoTC2av8hM5v
0RBVoz8ejoOEMqUIAFax8V0FjBFQGPmMOqN8EBz2oXBp6TqFg1rJlAwhGEd/PDYq
cwoeSK8ir/BPXpHFqeCl1jAkf07DyiTv+dilLMEbVf27ur1i9wX9bp/Uyl67Zj8p
mywtkZ/KqNjj4ZZdiSSOjeER9n5ALAuW4kNQ31zkQLfS+FX+wWzF7lZyDybOxv2m
ybTkszTjAvhYe8EixafBWuXf7R+B6o5BbrEwgzi7OjmkFMkgRTJ8gbkXOld0grV9
k1uqW0pLFyRfj5jwOgnzLV8GJe2T+RSnOyxRnw80Oe6f4Xr4pMHLqW0JDZLxWjQn
Ocqt8CBaGKeNQx3vYcG4Uav+H+mxmaA+A/wqjaNtWpWc+95uwNCNgU+ek4evgFdl
qZM0mNgevWlspcL+JiPrXUuOPUmbcRdj5na16G4+iUkmhtDFv35EZkXJg3/KW+rl
vCKOuJb2WiL+surL+e7by9bv/nyStLO4R9QdcpQgfUkcSY9VNjnbYgrV4P3+FXeZ
6ChuV9t6fiXS13OvhoOWGJMURCc0XIcAcJ6uqf641KstT2r5WR7E7VEnZOO1UFHo
CDPNtM2B23Q3mHFZCL722lj9MN8dCasnWUBjk3eHz+04gmivEYMBAX39SdxDzx7I
7/CN2VjJ4wK7vJDj+vNxkD/SisZVQgvU1ngotqrV0c4ZHHeESeDS7elK1gKgc9mt
nEhLK2mKjnfI/sHw9Edt8qKBwo6y7XL9p4fEhjK2DJnUpVbjlSB6LFTcutKwFyAv
kjtm9gBrehKVPdkssgv2gJuCY3mNE6xgXrbHAmn+a+irJV783JkYRE9aT/65bCcs
jYhP42iqjF56bSxiezyPt8NR3J9fUjCj0j1Tht4VOk4qhsKW+svaiphadvq4bZwc
gM4wO0V3BVgo7Nh9/Y4vpvYtNl4J/Y8iU1VJbMcMIkK1Hy1pXlLWz9pTUrpfCydM
HAIe0ImwQ0rIfFadWoeQ5u90+aCTSSuYJolKJJ49NruYEaHEEzJk6P7rd6ERTKTk
Jra1Qt1vsRkgmntG+6TDxfcdIfPMLXU8hvOO1VPaEsKD9MXCxGHptDWkWhit/jk/
TE5fLJ0K+qFjZUW5d95oqyjf2UTB9Y+vrGbc2FjX7dPazyxSjUl4Ja8jsYVta6/7
VHo85b8X5bdQPAvy9dk+42oiRqXudTrxThE4wBo8ew86/E6rmYkPw88L4gfIHJmf
C5hWGHgJ/PmaNTlHC1j+zLJcZAV8AZKmYNqUfl0nhXZr3t6IQu0FHRM1143ZPX9L
KkDAae68kwgpiKb1rCRIlnwTuQLesRk+m/LNRw96cyS/H1bc4NOrnpOpU00HAwTn
/CBrT+PV7VLXxoq0V/ja12wSoMXN8RunhvCloWOe2Na0mkKDDFiWlX1dTgvyv8FR
ot4dAj+ugYFauRGbVbLExtBIQHVs4Ety+NglzIZScEbPPDdIPCdAPwdd3os1jR4U
bDpxRLeSJSmXxPDgJC3q0ExL/ExE4/GVPVhovr5pa515ntWGmmIbuKRFDqkxdjqO
D7YErDStClWkfKNit/+hxfO8wrhTL8Qux6ztENzwD3Hq0oi1RYLxwvOH0ClHGSb4
R5Xdl4LNDapt0PjAQmwGaaTvVs85ZRk8PijPjbJq+cpLGuYanq2rjvdfuy4+uvUR
r4NeEspcMDp2zMJWPiBoslmAHUc/lGRT+3AZ6+LrJyfeY+mt1zfPSs7vl8MYFrex
Luy2PNM+JQPeMfqIavvW+3/wbQEuVyFyfl7MWjWeNwqlBF/ueg8BsySrEreZFzlu
PhG8NI0lEem89EMSt8v43UPQrE3li9gPt5nuwzBZOlJbGKSB1N07XHru1/5SCXke
+vK0szU1pfErIL97vNJOpF3JEMgDNVQA/dnRMsAduLS9e6wwQa2bzp/ACNPXUha+
GYjjtSjOSyrQw2vTRmXZ68Apm8n+qN7bBIf3U7hYlWdOND8Sigt7OFJ/JOXvXwLK
PpKs4DZ2Gt6oZd1xln2adymcAYGyWHAFvuLVjScJOMoGc//qP0omu1S5evLGDWZR
UOVuuklPu2h+W3u4dt97OC2IhsBp6mpp5o0SMPH5CsGpUikp3CH9XvybTd8DXlB8
TnRhzQywoYKA8Orwubu8rQod4yWZl4avh3MppqUTAbExg1ldfUPbATEokePmzSuK
wemj95uELpKouyWre7mQ+MwlNDPSSpJLJQ6sH2WcriTjWXyzxlCyVeK7Mc9mFQtK
Yq1LTWQsfBGQV7TtHkFDQ01M5c2oPm5HDt4XaV0N8ydvQ/w+1BS8RT1XVG19/zli
m9fQwtuc495M/xR1+rmV/hzLQVXfEyu8RaaDDPe01GKRqpyttR4wXtNuo9TPvYCD
nMuSvb27Cr6QdtdHLO4gklslytosOp9K6IOKYr3QfhWqUF+Nn9DJ1APo8tp77FaJ
Agxa9zfrn1RY58pBzLB+7xdmMCbTGwAS4hS3h5Hx8h+mI9o+4CderplgQUtjMAjS
EarF9dS/7C1z/p3dT43h0qZTSs+eyNDmhoyZG2HIzH5J2ELVbxUO/R2Ap9sg/IMy
yG3RdmCJKQVNCW6mSJNxktl7ingRioDy7+r7uZrmFj2eN+VoDR4JIwJ+wXBMFuOl
2EWEHHKxQtl9XFu7RfIjy5IyWZDVzHfw/mkYi4GqIcycWB6rrD59GndgQNi8noLW
0y2+4TyzhFEND17yOmxjMIU+fWdubUEoYuIqBaBt1hYoS3MtJJlr5EicsAJOz+ez
ebqLVEkr0e6hCiS4rz0k1F0CNEnRYGhrW1LwQ7QaRtKviTfW0hPdH3Qm4prjafhY
itN/b0wC+5telwunpZhh//hQQ+F8VrIYTLxb5mNnyw/3nqV3XC+bCx2oLqyA/rId
Czz4lHPQfmUJW1nMSVjOwyTMIZ4+WHd/SkIVjsLdD+aGDCQGx7UqhQwdG48vS4uC
U8qcIbUjy80QDqZ/PiSJEGX03/PMuR6np8AImYyYWihWB5xeMn6FnbSruCJJEDN7
WBR+HpAy5xiu5bPk0vzXLMhH74krsxc5k2bFpqOhvYLVh0DK4fpImz9gNE6IyAqi
+X3iBxfisZQezO27XSdBZqNtjf/x4lg9oL2yu7wIIbraW71MP76374SW4lEhHhPU
2qgMGU3kGF+/XFvM6Py2bcXfzCSbCuApXU3MlXVi30kLJkS/fN93LRFXtYTgl4Tb
NW8v//JAKKg2+UT4XjXhcY+jxuH94sxUglSorZF0txF7YHiBVrC66yriC8yKBLPw
MVkGoKBfUBSo4XVjaOxj3XYwKXbCaaoevopDCqztihPd1wEpBLN8UdaRvxidxAdi
kalSj7YOWH4pKKav1i7althCEB0Sx+KXQxhVkvEuoaq9LkWhyEhPfDva/p6GoNTL
X/UgU3+c5RAeUpYKqvFMaELuXXGWiIPKSy8WCbP+FHb+FDs3P1KVzax/FxoBH9D8
qVbEnOdVi0dFGD4h16lj5oy6ft4WWl1Udf2V2HR//MwNSBMYLctTt1V3DBelYLji
7Nq7kbhqT1H4XMLjKsyQVmIwXxkkFUM5IW63xEX1VAnLgCo1PKXj5ror499aShrJ
m1Ft08pccz2PTcOjxXMsEvNTubhc3+i1ip+We9VrgPTnizsajwjLfoz29k7Zhred
D4mJQSHjjAawlByy2JseOcgBhQ6+F8RayHrTNBujDs0hhmU+9YsdiZP9eO93z4zT
L+oR0QM1SkOkpHkXaSDOuYNYzh7+88y5fS2lvKlFhYBatoJG48CsxEK10RMgGYZw
YER9T5Dv3htM4WUdOymeojtPB1Cxnc0MmtLwnm0KtDMzEDUm4eKF3+fxI1sSlSdt
/oZ8XYJL63gpeIipmKQn/JrAnbpfGSxsXv58mCtYFH6bbkMWkbIEE1iWgTxm0SFm
56VzQMh9ulnf+bz15tI6oGAAIb1hjwYYqllyTd/u4DTS4Cw/exWzykXJk3CHZgwP
3ZY087mIS05gVLhTeWWQrttxLVtK8yadcJEa1qziG4YYbYW/HBXtX8M6cVrDN1DP
NBW6EVEdp9noeSUToU6bI5t3oJHFcl0y9U+e3BMyzj5Y4F7ji6XewRljrS8cxuPJ
RWEfGnQk0FZ01q6KE/G98xEXAvCwD9/XozwuReclIfQX82VRjmlzFqA/DKh8fgzV
CuzQUGCVkpPAeHweee6hZZ+T1IvUqNROP5gSP7d+9QrlmKmVVV5KCGj/s51KnCya
dWGSJIs+Vfjy2rZEfvzQgMZe+9map2MZPPyLcKfudwXhiOxxcOfqZABHk+JQFxKU
IQedU2tgXmuEfW+XH1GjELXzDxDP+dKc93yeulF1oS5/1VOhdPx/NbXkxa8SqSNC
2nZg4glDmMGYZF3QigGvV2+7LPyC1djh3Ix68iNyBOogilqt5dvZ0478u5Fo/ZS5
WzeJV5Pxs4MEu5ZpKcW2jB9LJhJRiujd3Ei/h6S4QTe0T54zDCTNJJ7oDgfWakI2
574CsQyjkn/9lL6VlT4bcH3ilkm3oPEvL+htiiYKVgD/fMkRBZjtM0a2SGSFxX00
YVtq1oiOF90ek72tHh2Fqo7bV1qrxi4mHGLHkZOkOtTLTHIPhL8mSpS1+Pt4Uwxb
O/QBPzmzo+YfdaNw3jjREayly24GG1xSHU9U6I+P3pWmoX2wE03C1k5RrGmjevy4
5vFDXLv3Ek0PSz2JP0yrghO1I7o19PdFrzljSFrH75kAn4wdYHPa19GiuvVxQa+P
H20Bbpv+k1bMnEPOhEjnHRHEFk71o7pg0ceaUGL1chEfNDsnPDVbHgvvQHP8kttG
MRb/OUWp037Xgym9McW4jmBjOv54C7wtpttikIe5acBZKGnG0vs1B4G4QUYmik01
1Gl/I/e/bmL21ze4UDNlztNe9G5bTUojuWuZNC2VwV+BlgfBQdR9rJQzbHEakipE
qETJVw7NMBTF6WVXLUoi3aAWChyhP/hfTQCYnCpWdYQqwt79vyghSE/mW5x03aQi
V1rVi2+a7QDodOONzVKAbzuED4JAS8UBFpUyEHWSIdOSwr0XKFiPdhDOlPOk6w/y
pcm9WDL9FZA7k6+i/ji4h6SwVXfw4sdS75UKMGXa3T8x+YwPYzjUNMCmN53Cs8W8
+ICTSiS+mOm0L5U4+QHBxAz1bOM4p/Jy8jyXhH5IctT1zfFLCrJIIGyFagwtuDwB
gEqf52ZpFzS+eDSUa33NsITUuby+DwSrubEDBP588cJYW9tD67gIz6ZhUAsMTdFx
YW4YZq9HX5wtctvxbXOSs6CHlkQn6lbvyMMXnkfsasVUHymVOGzjn6CMqaBe0EPR
Q+yQNXOkefQmfD9zT5Jg9usiHtTeiihKWpRebroMeeMrHSBpw3Cf3YvF417GEOx6
ouC41BSYt77YALQUcPqy4gqGYQy4MroKX/aEV+nCKoNPJ+cS2K/utp3j+fNmucjY
5NprPcKLSpuRSGcODHmXYdt+F9BaK8JifkVzV7DdPTiNQWBo8TcBQShSvDo6nmIf
s+AMXRXvy2nIICZApGcF3OGvZxDBg+nnAN5YCuXR2FLKf8bEfdl5tU7Uw6xUt72c
FrkDMi09mv0+xfjBjl+mjPwu03ko3tYZq5SH3StpWHoPmiGwKovZxCKjuDpGtIzW
8Inx0XL0l9ZrpHwg7sHh1k1EGX+Ii7ts1jwpcTjhunDUsQQablwaOuiiD2FJo8vt
XRcj/IoshuktBZ1pIqXG4M1eBT8WwIoxUH/7kUmjKsLbZXHrasorW1y5pWEY9drC
wUSgUAHzPyweUpQe6V0M4xR0fe5P+NGgmLgwgdCPrjLKwzgEDOHLrvPK2OJUtGTE
D2b16MyNT/sJC10PBMY3Co6Jy4EwORJ2LDfwbRAwFusqQ7QPLvh7+r/OrsCddopD
MKjxYC8Do8LlCSNaI36mL/YwoMxUEXu96P6CblkD7+STL8012xrnixCWpwfCGu30
xu8s92hSs8T0rpQBcSZXZ6qHJNhWe/kfk4HNgcdNYpCFkLTm4Zd3+o6gc2Zo0wUe
BBwzx638G39VP+tdUICmSu6d5u1tAnqjXKEPHAvuQFiMJSEkFITubV9TqhQMkAbi
ALYUJifTRuaKrnUu5KElqthHe2oHtNla47W0xlHC1f96JY/2B/Yble6Iiu+9Tmtx
YiX74BkyXKaX/CyRQgjsQWC8QjL5H3cLFjiBOHn7uESStPJTT/KNZIee+ogprJFZ
Op6IrPbRVGTaWC8i9P0pGHnM4I8Q8JEX3XoWajW5LK5Kf7B83bVHCXHg9HTuvmO2
Rl8Gmq2+0CVBYh2RsFf1hADbxbi8tNxsEhWJMoL3E8DwAbHrchJaEmRfZo0TvMVe
OOFSX1ZN6+4babIzKk+GWwV/hdC3pQ2AAoP42j1y8uQ5Yi6VH1tpLxmxH/BkW64L
e+MDHfiG5Fuh9KOSyx056EKdTNloraCYiuEZwBA1FJ9051xPeWR/YVeftknhNO0L
mP227L/YgndGQkn7vXZX2QvotGPu4Hbdo2kUZbJmWcd9Q2gq28FqkArqavo89CUY
plJ6rSTspR42fn7W+Gx4CW1dEIhoGrCJlqt4OcvH2mMlkbdXUaUokGIORLvEVP9v
hREdiLNWo5oOEDkex28TLKzrHi+OkthprijHpUrx3qc0PL2A4ziNdmlHwZZ/fwbV
jywZYvvxB/UNWQ7QL+viuHW5dskqLbWbpfyB6ognpjBUO/r+EexhdUNczINn3ULQ
Yy352/sasFkr5wLdAlLLAvmjKFclJ1tEihqDC0tGPFg45YHUvcAEh6C69r0NESTM
ofcrJ7t5c0zrQ58p7xEJG6uukWbpKszst3GkExj2CmmMnE7knnfKfGvVf+6O9nW7
lgEBpjjI5EnB1Kcy0q7LFEgOwvemUwXXpt4ggbIA0N01ATobM16se0BKRqpRchnK
RFPUkIhDVbuqI9yhMfw80IomTIg60cJlOqOc2tYAIeo3xg0RNhrRa9+pPW1/zwrw
ghjPSOPYnp1LqACOsN1OqwtosNQOq7xE7ZEmXtPsvJP9RpX5RYyq3smnXO8EK38i
WLZZ48nfPMlCt55AwBIgD3LU5fTjGvb8cLSRNzKwFeKuYIIP8AVWa55e+7+meWOv
WXAeQati6+Y6Qynxnod8X/y4NvIVF9T4q+uFXW2iLOQdGHRddICN/mH7Foc2Vwu4
LSN/SD9PNvHW7Hbvhek9+ItCSpqx8viPaMAdoBE6KOWaaRKpcs9//wh86Rs7qsx5
Tx47LkaTEcKfBCkNS8rOABatJOZ4Sw/rgkKjB30rno/xOByyxTn4AJyLdP/hSGzO
ZbzJySrG7Oj0jAL3SLyF9fYo9xqB/Quqr0b4k1e6Dr4=
`pragma protect end_protected
