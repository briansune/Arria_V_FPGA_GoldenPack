// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:20 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OEsivP9Shv47TNv99gFLAQguV8EjMvyi+MPkSjlsNq9r35oTL6AY7iDzRjVwQnCE
OpPigBUK3dUPiP1jUbxkCaJDdWxANjNTxf94wm1klX95QTNk7RMxjO30JqC9EMK2
0lCYqgLpFwr+QRS82V/43AfAIi2OUl1tPBuo+A0+1GQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
QocFWMXu/+wO0MQFMi/dUvyPDg9eabwG3liiip7Y6reiM6EmdBp5gTGkVmDMdFMj
jtWQyBo0Y/m44ryzDj+J18aYTN1LEke0lfcJ+JxSe227PmURLbyKxIg2gu74jMZJ
k9MjHMI+AVU55aOV+wI/M/+FziJLjZmHecCp3IVRFYFzRHzO5JKItZ8giBas03Fz
7AZSqaS56iLmX6ay+8bDfTmOcWU16/3Dyudix+Vv5tAkyl06rb6NcjRjs6ibjnV1
1+OvYXuizKP1PK6/qMUBJ/X968bgYh0TzaDdh+GMTvwFH1K58F8YIOVftH/ZdlCT
97OdUbkssI5rXh6QGCzgzO2WBGB3xoz8rWHAKnauAl5lVsK5vCBpPotqsCRYI1PU
lL+uwsjJ0TBvqKyFNaQ1TDid81H8bPntem+Mzy7J+JqcfobwMjBUFwRoNOAFWEpi
u51SUod4DDdGTcSJK2olEO+HSyYrpnKrFCkV7K7jcQK8Z+7yRmgoygC62kJnicK1
pG9WXdendMHJ9Rv9+mY83yFBymkB0q2w//ZazQcbDUgyM9GGF+cTXGMkfGJk8XXt
PYFzKpIFG0xTWtRH5DQ0G8fdScGrt4YHykCcEwsZdrOx+Vkg4BQiStVwR3JwGaTz
jpsIyWY0rtW9R43A0wZYxxoBhVuJMbHboUM0D6v21UlxRH8I53plswg4k2/JmrdX
0wFOwZbHT8dnqofGPv1BDeW0qIjJM+A0a6a5rvLDh3ZEE817kWjuEQepoEt5igl2
iEjLklSmJZhFoPu/nSntBG3qhECgqoAUTYRTi6TTqBtiCNjjfx7aG9R92lCbrIo5
D1Vdp7vSzpTQpP7LSBG9YB1AktIjz4yLdM+6xTg98TRlsZ6rgQBXPQ7pkvIm90I7
bSQK0IQPPAgXRlv5I5eEB/BaYfIW4d9C0WHJIzSc/MGwv3X6skFaSbS6UbvWcaI7
falYVleCCoo5R5Zfxz5rLdiMP6o5WFQX5hSrk5PhhtIJq6BA/2GUd3q8dHPWqh+7
rj/ZSdYmFcpfs5eVz90+rKKc1OcpWov9uPCnj33xdaWt7KObFj5Ou2kp4wLj0UqC
8KebU19HXyHuOZ19WYHu2P+yNb/HCvbNjdlvRSHCo+wPI4/d16oor/edrBbtqgFA
pli70jfXb72k3r6f6B8vP34adL5fJUkusRTbNNMSyC5mrwvK35Y4A2nDSbqRcQhJ
1dvEMDHoJFUL5Bs4AkrO9xL/2iEnDyDUM2fIjEk4rKXdxKsPiPIHG6bcBV9GLxJf
1Uw34REt3aj64ghB+2112V6VYAetqtSVaEbieDDPsJYPuhBy8+K8BfAPWP1i+9QE
ui9x1aXBfE1Ozj+Z/ijeI+ZFDqV3BWvOoruRw2+cA8gocDA1Mt/66HzxPpM5nSk7
cAepeK8aCULLV1C9znnp1CT+zZwFFUHqA0W42fK4VobXit2LzWSsMHbsZoUyUri+
vNohnreKAOwr7YLPk2eslVt/YfZji+W5Bflg5ojD/hvFb7SA6h+ezxDLr/Uq9Wty
IS7TW0XFm7jpIDRPV2oQ9lIX84LSMPy3WR+XK252EdW5xNoLZi3GouP4y9aKi8Fp
fWyfQNwQd6RxynvriLiRX24jgxWfdghMYe+SC66dnbSV/bwGNGVOGweVxAS6I6D/
XoQtJ842K7Z26tNXtkc5QLgK0yselX87qJ/LWO+OC+dT7Grpb6fOINJmFvu1LI+z
SH4Ufe2wsz7B/onZiaQII6aF6ObwJr7klbXoycRWLt5wFQitYWA+6MWkrtP7a4Pq
6N/VuOWk5LVHiqIyBT2nYyMo00bco0J6QGp2fomG02KsjhBNg6nOXXD+d5wXs4Sg
TPxVrf/34nOcNsff+Yl+1inN/lxVjHtNc7jd/BqZaYLl2Wgdr62SGJBMlBQ3HLkT
90d0t4r23sBM+e4d5IbbDo6zZimoAlyUOb+lYmaHicnXucTYLkvc2fgNdzDHr+xK
HKEv2SAOeBKkYHvTFHmSu3Sy8k6tFBP9otZfjFIwRItsffWOLOYKnVhKXJgwtDbk
GUrT329EkgTl9JaOFhXcDL2tfMHHjLVzXTVdwgIpBDjwC5OHl0uOoehOKlT+pbJk
XlITExkfY1GnciGgsQB208jd13wdFyTUvyfgPMKOAexYTsSBT+Xed1ysK/i1RJFl
La41OmuOsy6DkHOq5SxUaEbjI8ZmJvLz9PUH5YoFmj6ABIwBbU+M4rwjYvGlQUth
GwKUb2h281xycG6IdMlyQUdhwD7uXete621ZMCZrxLGI7PpfWsZ87TbDENJbt3yV
0zWxHtM4HJAMMMXSkoW7Ncgtn90TclFhQmxf+4gaOexaXJJaGtPBkJXJaQi8jwq2
tF/o4wtOLDBVsz3rrj3KSA3O214lowACGTD2hyHGW4u9SYMtJSKrjLj760JbxlYK
6B5C2DzuNQAnYkfmPH3h9A+btEf6ZDk8fNEznKUuxdAznOqVHFbxWlizZ57gd6R7
CqCoEymFEUG3OlOFUahmf2N+i2oq65tFBVN71s6kq3k1Vjq86nt/VGGXHxuuS0M/
Nsw1d84XicZL86+cXQKrZjCvdmqrmmrL+0NDyYNx1W+6AbBKVtZVfWjQnjNhFeBB
lmEhG6LCdkLzkn7s7yxkQwT0V2GTClFwv+j7ly8D3b8NlscAwP9Ds/c9D/z+PcfE
VlxtLPfC60/0eLatICIYbb83dFmI5tGswfISEM9mMffNqII5A6QeCPA61H7RkoTB
1GaC0HqXo++sNW0v1K+yjKTtRYUPFp4UxHG+IElsNpjxlRba5UfupRczjXBAAbp3
j23R4o5SbtPYHQ0EJC9qWXy93cCaPpz7I/5+NJxqJiSJ8rTMhcZVS4vEYNXAawzd
wFLCytbYlsItfDDBgDXdysXBBnajaFpAMUbUbDXTpKBOXkbETodKSX898ty2KmIr
N6YiLRPtZA3PfjutUyB5xv3fRmY8CbMZPrPU6qEX1iNoYzLdgI0th7rsWD2xyLJl
NJI0BE5J8fsKYABTh1U2koDpYvnseJWfb5fLEzw1BJ4m8+QyDA3cDaBjEV5m9xye
8D/gZeOPV6x4tE6lq3ssMGnBPI9AMMvVBh3cqDGIdS7r7onnKl52In0pjiRPddzr
wPCfRGHlfVKEGwc16W3AqaYHuWIu1CM347umyMPT16Lz+Td6NJ4l6q33bNNtnN4D
KW6P5vl6KiUvlPPxVxJxRv696GzpHioAAXkHfHmw82Y2jNw/G70H84oBMc3yss5T
4gTvIp/zUzknrMd77ZEDSPK1/EoPFXRQrN5v/BgvCbtsN+BfNtA+s7y3jfO2RfuP
Y6yv47HnrWkC5XWuMSYm0CSkD00xY+NsjiXf61gIkEaEYq0Rr3mHGOa5xwYEclmK
yLt6uPO6X1ITvhESN/GOvoNZXJPXwCknZMdzcz5nPpn3DDXI1VgRBXscnXhE75fg
9CBSkUZDKQbUT4utiiu/OWKauOcc7kGMyqnhPu75qNOiMSBQ1ID+hLEg60QMH1hr
/S0S5otTF8dtCFc52EAt3vtPRXBW4fvmnfjtlT2TkjTjNiUCB4S/KNKAZqe8zDBo
VWWWXWQ0XsNPYfC5c1JZ+rYFCwLE3zdkCW+whqtHJC7NKKZKSlw2EcqVtQxFKtZU
PUMM2a46YQutpr8AH7CHXnMmK7fq5/m1WGoijOhHx5e1BRI61jDb4HHQ0wy/V5x4
foHiwapXkOtP6t9uIiVwUxfOHAX04KYzERaXGKLOwS6AqVfcHHCyzt1AQ3POWP37
gdzptaVo+eY0ks82g4VBaiyP1xPLbNirr3kjNj4U/x19B4IjFxWehSBmTzcvSsNb
1OPe22IPrF99Gw6Iawk6tVJfoNCh6YlsJQRuMfmWiv6royx12qbzUpHOimLHHGv3
d1IBd/OvtjgFJqLZZh01EMfx5n8tSR3jm3XL3TPNe85OPghzKv2h3izwUr5X44dq
/eKpiTDQG7OqwV9PY+8ELOobUqbnwyami3qtjtLbAP+TRUdOcSfgMU0oYskYE3TI
LeTzQgYAOUYrtIRPAMiv+016a4IOU1LOchulVpjKZeaJaLGdg4ExevrmO7rms/h2
EUt52w9sOA830uVrZTK0dDd7zV8UE6yFan5XivvLvMaZaMvYG705HoObn03tpNFN
5x14NcBO2G4pUu733NMyKuyHqmzoM9QWYtyB7EMurDuRTJzK2+VAEIUfIItd5TJS
h24NYHeRSWZIce3nfhWQhiQaFXXXgbVnO2lgebxdGNK5ycN1uNkXkGDR2HQhaBFd
RYPKjX4jNdxJrKUnYtUQ9h06pz8nqbjdif4oViz2hZrkdSeTP8k3ksxHUJFO/WpK
r4PmcEr7PSmHaalUhrLkOS8ipy1tUjQE24B5hFzpvgq47u3ix0ffUhSEsDkjdAW3
cj3clBRHSXxqbPy5D44KSdS+mcM0hDxzwiL6tA6FhtK13xcxF2Vv0wm3qBoROIW2
/GsnkNElGRIe0wc3IELUkGtjrzNnQq5GqIs9RQpER64f9Copwmf5YbE7G0z1qLSg
6xWC48wOLfv4RpWKAV9vUQYQGGts/IxL2TYEPglz+WlfhTQlbp5P+/iSHHLbT0h1
4jwgkQWi3MZIb2QVKVeI/N2iOrnCS8y44xC1cnh/JSBrDn9bpHH8bQnZuSfVvoyF
p9nuqOqsHuElFNpTDIDz0xhloXxPvNKw0Emi1rRfQcjPqiNd16zARA3hdiI4fVSf
+0wY7NjUh25UZ7QkijwphzS5D90Rfbq0givUZDSJ99MHqsLspAcIs9qQ9+T+SVEC
8GoMxdEVrUS40fEFI4XATT35J1sdaXNtoB6PvqGXjvg0oITWy/mCd4bEtQV/wWZm
eBP7vOLZ+wRSx8KNqTFYGkFqTrrpG+lPlJw39glSSpA/nB7T2HR8KQ29UorcNjTe
WRpged1Jc1omGvX+pdSCgU6HhC1ahNbxNPyVrCqF4IlBqKaTFzhRq/g8+Vssyu3g
7ENS1utsifYqO5wfZqpQsP0fZMEapBC1R47QIeDb9m2ECBnbkmW8P4D2N71QI95l
0IwVSB5i546/V6Qhgx2STvD66k6MHvmbCu2pv6EKnUxoW9+b4kVixA4jfuz+rlUu
LBHpIlrwBQMauRuVYhxQCucLWrKrAE6eMpdTaWFn2Q/QEApXOJ1caBQ8wEU5TmqK
ozzZR9l4u9Gy9h2OlmL4xrc44pyEwJ1hQNjxbsuy+dXQBDrN+1XxYXppf/FiSc3z
gLd5hJ9rfiCamdCRwC/fScaudC/EO1JC/nDnF41dfPW0udSlt6C9x9PKyQbH3JR0
0GO5/06ayI6aMtVyTOzvKCVh5hTHJV83YVUy8VWTdLeZMJqpnypMmYGeM77PH69w
cJ2n5XLPiAz+FtO9cIvncyRzYstf5DvIgWMLPlVyL+F/sLXGsH0RuE5jV8e2Vy0J
R/gCaQj9g7aVJ2eWePgsCpsouOW8sNvdR4vfHWP1tPmLw6eb1MSaQIy5F/5jWaoK
eXNWpcNGYIhAP8/17hA1+2aolp7dU2PB/TSAcwKTyyaHUPdz6nF7gVVorgc4laLK
cdEqmOzahEc0GuSkvR9A1qJMuVF7EU+NggUL0CcP9Dg8KJMFfTQs4EZJ+v5Mrnlc
epPH2RCrW0z0opVM5/pKFqI+UcEIODyF/sjC4kYnRk5zgB9OwjGj2kUqF26YsAhi
6AUjrhWTvf04KzpC3zWHtpeEjsXmo2qhnuaDMOVbfX4P6g+CbVC2zJkSJvoFNq4c
v1PNFHc+uRD558pmCIzMy6jaIaClK3pQG4I2v8WfPIGv21cXnqKIuoHKlJFEifhb
zk/UPgqur8ldchtRJkHvsm9aKghW0o0O1UfcPgpitkZiqrPF6+Nh+e4S5ZtMfxeU
jAGqA5nVMzCv21/RrOY/yWPzDCoTUUqnu9EJN5l4RkA+yZak5hUoOPqynGDFVVeV
sgPmNNnmRwUBVHoD5vbeE5oJSSQ91sWcv+eyc1ztcneYKpzFjx8lBWzpvH8LM53J
062LEWs8//bA5FWKdwu1g2Jjiga2MXnBsGAuV5XudA9eCy0ouzV5arHqR4RqVa1j
dS61fREYiixHdlHR3NPoBKzzvQfaZyiKFYqdu1kWAjGok0GnZTDsqFT+L4+tlpbo
o50xBFrXz7YTbRynun4jR0KjOdWqQoBb0xn03PmnQlEIPfB6Zns9cuhxXxYHhXu7
kgT0r/hfaz++MzAwrrtnNmvNwGxFaBkYiKFlSxAAEnqlxNYwlWOe3UhJLSSi6oOr
fcEyh+45RBGTA1/bU1Swv3kjrCnHZjG7S4t1RotvsiXfML+1QPGpK/5BTp8y2+f6
niNsYDhaE+kE8+ZRb1+bca7tX4a6MpvPQFVxs4kctK9amWcfXqrXYllyCFbDZuE8
/HmAee8KJ+kDaMVQek/naUtBluZPsvyLGm1poRiHWyj8b/LwZPYGTp5cwPpf3+PC
sKR4J3I3Sl663dMC++IHhOjIEKGEuKELgNI47MhZl5b72qJES1dgJaaoby6VSbvm
xxejXpuhzfku0IPSFkVopSQhwFC7aglixV0w4QUmtELFXqgS9cUDcbEl06m9H8Su
pYTiRBRmh1a/oocTUqYkO24J+UUAnGKS92Oh8Ijr+rGI/LzV008C/KsFqxPBMG3W
i1IVRSFskGQVFNy9hIKere1zF6ZOUUs3NZPA+aXejyFuvZomF52Gqq96O6Ggdn9z
/Z014w18bcdgeBsoUmsNd/I7fa68bqF34S6tQzxkKrKzRZrqRwNBjWtyebTj/FtU
EtmjmQDVHYlE6vN6F+RWssZunRHlZOIOZ0LpUS3Z07BA6yNtwYTtkVxKK1mKHKUV
LQUrCIDTllQXndcDHnURkJbNWWs+Orio70mLOZwriB/+zfVoTXoXeqapaudkGmdI
+EEPD93n9DDYb6+pStJJAOcbK8vNZb3lfSDzAhZyCMC5SuGq/Iqbigid3UEAy+R2
HaQDZG5dwK/wngtGS6LdKGBr5LCw1+A3SYBUi7zWffKryvXrWSZ8WatM0WZmhoGg
vVrGmy2nHSmpBxS1/JLYe9JkZohKZ5iLNTA6YbhQRM9CF/x7ecRBNwi74cOfXZS5
sv/gN9hJX2PvTIfXeSMWsEf82RsbPaHHnDiw1MIle6dBJlMH9sNRlYS3UnLbC/ri
yiXFsl/z6T7Asmb3RR6qn9SdWawphJiMm3gnDXe9a4+YrbvYeF1bYUb1owMi5Hnx
4dCwKp2dlHlMbYUB0ZSKQNQUc7mvILlobb26wy9t6UGOGDHzbEZOrfD6IE72Oj7q
j/i0/+X7GB5Ql+GvgffR8bug9U91rBmQxwel+bKQwwFPREraON2cXhZOc9pfs6kz
emYf+IW2GwrNVFClX7k5Xpex7Xfc7WUy82XiRJrCK+xzHYK4y176BjRkdJ8qkfNc
Nl66xtuAdOVlawSkSJHkzRVxa3RzJz+hHo4PbELQdyZdhbQhtnKPi94w+jJMOWhG
o5/Z7B+4Eif830fOj5NCv/AxxxufNhcbvRknG/48opYxb41qTOqdPlOda/q79V7S
fKiKTvzKNc7BROSV+5fdzxrZvBwSwzOLi0MKavqXrMsXm4gADP6Zs8fXrtyp+Yx2
MTltr1O1mmPpyjImtVZXGKrQC1OC7c9n+8miSpJWYic2W9zYsvxyHk5APRzA5A7T
LoF2ZhbZ+0Ux+QezhEPaMLbF8nazFzFD/A0Js1Mqj1smnJV8atw8wTRAK5C3BA/U
XGodxFVApJ5XKAuS1Py32UFMDz9b+WkP64+7FcF0OGP7AMw0mkq+xjDSaTXWr7wC
cbIf3GQ8G0y5CAKBQDT/TJ87UEkeiiWLMBGucMpiuAdAhsCJTcGKTSekrwg71OMs
kTdjZEp40cB7UGEZzK+uhr3dRTqvilPRAefZJ1L4ClpRPQc8gE2rBSxTrJr+kvke
ibG8oHHfpfBhEYwHAQfxMnL2tDZeELHHXqwHzl+How15GqENOKXZZlqWs2cmdJJW
NNt1rxaWvbCECWSZRkI9PXl5Rc/eh1ryGEF3nIiqDh5u9n5chhidp1SaNdqIcEAa
NfkxrxCPBhPwXIU9vN59utjFY0Ezfu0s/oJ8hbliVwqhuRjV24Z+r99iI3448TP6
zU9gDehBfvUOvqxRA1bcat+zNN7qlAANO9EfpfvODcB3CVNmFImo3hlt+czptB4s
YI4Q/YvGheDhgN+LUmt7ZZ1u44HBbmmvvmIUp25af46lLYVbNTPCwrQKWeQd2iqR
UVDRp7zoc7CRpS2RautenOOiixvHNAXp5cVtkAVm/4K5aGnI4jI3nWA/kRMlN5yu
cqL720fKH0xOdXtKkSOV0VylxorU6XDnkgQSvPGOSiI95xsef0137QDo5Zyxd+a4
jqM0cNeAaPvjN8Vk5hY4Mokv5er1gIcOnfo/MKq64u6ttGWKB2b8plQoB2kyfHdM
itM9LZMUkEDBTUqzJaVfI0CUhHVWqCp3vFcNE09M4m0dK5R4Mdv9oGGvKNwA0obz
o5FBWZqdL1x8he8bk4DLTJd1fJ3MSWeYnPH64IgS+NAi7Z5dBb4UgQRz0VEYS3yv
xQ0IND+qMQniWG/bIqFPUUr19c3462GbUVhCQhj5MzTq7/qzvl5PSxDQ9zePdGW8
YcI5X7OcCOu61EItql8WRIEfgji8AhbZ5FvmDMjY0RFZOgBzD2bjrPMLvqqUwnol
gr1+kNnjE4lvqlT/f/9eF8/M7LaVXw0Mh/RWuHplbk42r3xY1BXm7yjgV9Ognk7V
eZONu54HnNWuErEgVgAPIfYAZY2bnMVkAxq5GOMXzjqNF5bPCWrm14spChHcjZnk
2u5dUTsDZ7RmxnoTe5k4hhshh5Mb53abCIv2f+c9D4wMjvwpYLWp4JoX5ZXJAMMt
/R1osNH3zFtLODugXPNh2JWRGyI/rLK1FVwDZhX1AhKcs2Kj3nFP6z53mAuBrI3G
TDnLsikss4yKdOe2nnDUrNN6TUV43U8grawiMgnFXANJoIMKqzezEdvHx0rxixP3
fXtEzHPn1BVjI3lv2puKImXjevQKPuIjsy4aDa3dAT1SvkXr/UVoKEsbZfG8IRRh
2KzL9b7KbBz0QlsQzgNuj8QW6SCYD8koGOQzm+xwK2uHGDiV2RpHZ7KjBzTWBTkc
8CIEUNTcknLCAMUwtU/DkqGfYBvRq2Obt+owFHRPMFMFQ9caXwahwD7RNRuJNAQa
NUM/ZMfQSrFwr0Owof5kO8cTeF6J3DeU1xguZ9ht3BNU0adTl/7a3DCgQCZsAxAP
3JN+5FfEqf6lFuxQB6JvmbebFIY2D6cZcqbXiNZpBjtU3sVXyTrxEgCdsRqbVpge
OE7CaFhSRFmWpQ2nXFVDiLUGKCNUBKPJtcO+3jD+lMJqE7U+aBWNhkhDDN79f8eX
fpEjC2D9/FTJ1ZjpZAIrcbmjYZgRnhYm8SItPRX0dJ8aenNyziGvF+NDVAEra/Im
g295hahI6Y6RueadNAh85ehuR6txhPKkh/Ab0wi9saLN3GN1seLS3FGsSM2Yjl01
eZXYLUhz0QywR/q6k3L18W0Lxd7lX0gqkJolHPzIqVzZJ8QwfrIPzIty6MBrjOYg
XjeWhaLDVYJQg7mIQzYuJ0fr/AwAUZ7NWlTZt21iAPX6N6DSPDbDyYyQEQBwWyVQ
j/+WQY4NzRybp3gDKRWF9M5Jl9nzAkuDGOZLJwz32oXXSa+IWMfVN81djhneHngd
6JrMiwt1qPONyAQc/WPzQKzkOQaDi2VfXnq8+93tvj2s/Q+x0OfCSrvcrBl23qvR
84z1sOP7LZvaq43ED/LcSQla+1ibU8lC5v3BNMkdrkp6m2V6auwPLhb4iHM5OTH3
BtIvfy2aJPEEbFmtCyiwVMg3PiKKX4hH8Be7GOV0pBGOvD2p96NMDz6/V5E0fBuC
L3VS1wJWaJEp7cq5z5kMcM6zHYEDpy4cwkDDSYL25Vp5cEs/+MYvB02DqInvhE9E
d2/RN3kXrRSG4CbrKt6yePGHSDMb9cOiyJQxFIn4j6yYn9GqbGY7GNbAmNzHsN4h
g+FF7xJf+YdkjX5SrqP/BocqYHLG0carqTt704uWdbPr933br6Fy6Ni5hIHVknAr
Fh3ZpGgpqFIEa/I2QaSF2rbhL4Eb5eKsA5j5WqY7A4Tm6cFovni56GWeV9GcF6tC
HTP3qYIEXZA+zMha38l/D8VI366ohVQtvDbKS/hka1BmTaxIwnUqPw783xs3p439
EhVeWe/1A2jlvVY7fJoBp2LoifmJEKDVTh2D1Wg06Ehfq4Y8VUs6hoP7IZ95IanL
HUNssnzCFw7MlI90zBDA7tEjT3LOW16uHh9RXA4z8n1ywLxqNT6ZmxCODjLgGepC
k+x6ZX6KS4xT9BVzFHUSK+Q+GBR6bsRJ/Vex2k201Oz0KndDRdXp85pZJG0ViELR
XJPqGmAMK3FhbDWl2yVC/4I5eIXKiUygUny8zXKXOSCaH3j568iyBEx7gtxmLR+f
G9eSyY/4/4S5qjEG2QZtG6Mwv1qsEQQ37WBbH7MrvEGuotqOoaCWsGvsaZsPd46B
t2Zr0VeX1uwS57oiLyK3Pcil+42ghfydP2kvE2WHK7+z23F5xYWcJ2fa4vX9xSD9
OQ0TaQ7JrvERQtmGxZ4NpuEfME77AvbfrhTKcSWqA9TGAfGZmfTcJ7RNg7kz5QUj
M/qTsBtzu2/0LDFSfyNIYaY9prBOFDtJvfUuFCtgrXeEaYE9kBQncTN9a/VxueJR
+zQ0TG52ESbD9jD58oT+hoZXVsqwLHae3ikjSZ04XDCTvvXtYVoni/MX6T3GgIlp
6pM8puYP643S6il8LrNY839RyqgxHHVf2z+RPACxYQzXsWGW1NcQ/3TCEKDDofyF
W0yGWomhs6XB9XLhfuTaQeJK1H18iejNZ2sXK/I40ng5oo3JI9K8lVuwIpMXgKwk
OofDFm2IUDY5m4gs1DqkI+zLYIT3aRlpdYuRNcrpC33I1cafd2uHt1aqyYkdkeuF
hKJKRtwnO/w6k1bbEro6wMNLcE90ewJdnki/+ZrD0bJcYNLJuSESx+68oLJRwV2r
nELfM9wwq9YsHslGMZLqg/gwbEFSeMtvaYbjWLbt+JB9jmQ+1NP0sTA+s09Xy1g8
atGrRLTEJ5DJJBr1AvW7yKTOKxJvtLRRNh4IUGOoqYOw4VmfHXE/U2dOFVOoF7pM
FG9up76TKE5dpODVA48GzeYCwKcmgNbmMDJDVSNMLz44kiGV7WieQg82oum8vhxs
VsResOrFCJRk80rxQNbnMmNXMrbi2pfLZwTJMor/w4zw/8QK7P5smzoEc3M39ZOG
eCfzbyIiQkodpkQqCNsZRFnKip+EaqOLVydE+SDFAGWFPqpry3lKurQi0/qH+FTp
xOEV1DpB2jpSZ2XEl7V+dGTLILThZxW4YmWyr0PEK5zSUInxd/pXMTDZN2zS11vq
TeLrtEEUs7x2HsnOoRlsgxVVYavgYrM+0hBTeB4mydFEAbNJaV92ha52AtWXczBU
1cl0RZE1ksgMi0ZJ3SA7kOtA9qei1iqdvqKj0HvzqTPzQxhLjlQ7PBzf3rWqLvDE
/c3S4ZG1uHtI6NW03Gydx0rTcXT2ewl8vvpnHNqsh0WNSZQJlIlpgSN7XJmqHpuu
NOLW/1yeUmjvfO7gQhCFriOfE6miJhSIJ1daCMWXR2VYf+nL/9SkvDeBHo0BWMPN
EUQxTmlFXyVS0TrRoqRy8VUTSOKuZBE75pdFktWWvnrlTe4SNQJw3ptmQt4ZARYh
Z0p2lXHFVoCz2aokn5w8YNPf2QriRX/Nc/Ul1d6pIw9IiO8fnuNux9mHAhjY0/vJ
Qg0OMBZOl/wXdUoWWZjmUk/y4bA2hsgdlKQ6ZwDz4OQX6mRgAbxHf9l4qBq+0RuR
OO3CN54hC1AIW6mGWV/roLG8CnUMjPcSSL9ZtpklG5k+PKR4Pg/D82/w/hgnLgpf
nYn9mLahj+xYiO234/26I5nbZNNoeo/qdYvyWwin0UULGM2wvuUf5t1JVdpvuEbU
49Z+y/IJPMyndsh2zVFSJeRuFqWgtAYnFGxAQI1xE/S9UH5eDgj9plsdVSI/Dgps
fWWUdnG704FBB45Xilp9QwycVB6AqWJCWpNyOyDNcg1ltwsMgBU+gEaAjl3/AA4y
Ba4mgDtQZ7fiCPVBjxWCxeJFn/VpKTle/r1ccjqkVovesDTeXbhv8wOTOgzZq/gX
bV3D8XmfektejnCXOSNvMF/AWhTpzFxmPdx1vHedU1Ug1j/ZkZLFvtIIhvcO67xe
V120MSOXcy8t/WQOVUAe34ruwFgk7e/460iHjIEI5OAzckE69pHfALeqb1o6t7ob
Jk1zbQGcEfR94nAjVBJo82c1AwA+8jaUANkb3+OAz+v86ws2eAwBBeu7TDWAvGon
cKBgjBt4MlodRmaUaxHSfYDIu3rL6rrOuTck2OMZeYtNJ1WeUET1OtiLZrtFUcYz
So9bCI2UWjZuWkVhiPHQvIefqs2IHQpeplprt5wGKEgcNcpj59EVSwG4EEwHuemE
8TL6isBxPwH5FwuYM5aa6f8STKTFVZ1CDYw1QsAVdqQdEfJfb681U63X1ikGn/Kh
LucCB6Uq17zHMFaVn8gOrFdI7bj+ZlJHcaKWJh+lKticDAx4hahaSLNfsLImZ/C3
UgJh+pAGS9pcx23jm/uqWYwOjXY5EZZlFu0zEu+IuGK6yhXjKX9t99e2PCxODrWc
/egRF/3S7roqm3S8C1LOhHGxkZqkA17jQhxpSpAzPg92jiO+rGYGBpbzMjAEw4cg
Hqt2W3Dq/ZtAimfBdaK1UNeWdLlGrhn71fUFnq48XweZSUhikO8Qe3XP0ieeXTGt
P/MdhhBPMHh4BqKMHZYvGF8Hstbn8XTNF3WRlFw5W0lsPauocDCl12tKnD2BvZ3n
U5R57J/1NY7wXBmdWihvfs+jhsd4vkbow8XWdI6nxMn9p2ysq6B9L/bUEfOn9zuO
RDWma5kNwk0g7UEmGN6442WEV8saxWTXjD/MTNDa43PboXNGJTJKIrYs67T7I76w
8oH5BO3zMOidjmTUSBLfsd2cJlhiL4Yb5Sy8ACQMpO0TtFDkTUMKYHkYQjMNf50F
bE3O+fhOKVBqWiAhcmbd1yguKMS4EZc17d8EwQtlF+9iD+jYpc2QsRdgpcDuS+No
o91Syr733Nfs0d7sWxOQVezzTpAL7Q3TnCHu1slhvPxdvzIN0EBQlZu3nx/tS4N+
rIlSp24PvzN8lWTsL/dYMshC2CLN1GFZLPK4Sx/2HLnmhyCQuu7JfWxgyUUorT9W
nJvAj0mKn7Rg9j2wn9lK4WDNbYtArQZBSg6QXs9Ljk7CRDvde2+BQk4cqvg8sRFY
VO4I7LujeUzW82bxaeogPbKg9g+uXIiOAtZ4KIuwrsS5s8UUbjyt+t/bRddjH/Y/
ZMenUGeT4wJ6TVv1dblW5SdnNO3Q3zDJG22I38J35tPjCPRwSdInzMG1Ck8tuCYW
oT33gcJrHqyIvkB/tCLyNAxPcBrLaC/xmdXR1B/b0YnLH1F7gCWW1dVVSMyKmn7U
LQUzZz1Qy6GNysYNo7ay0NUyilJrbg0vJq+K9QPFeATDdomxhA6l8HK3Bd02APb4
J7lRZjKcAzzcMtocOLS0vVH0+IGtiOMsp9M3XWLWvf49iF1np07LKxMjt8BG6SIy
rBIIbDypAIbci8BdarUU9UF9SRWOIkUOtG1cAo5Sxks6knnFerr4L5Rq3Gi2Hyl5
XY6Zd4QuL1yisbCPQroyOCAQysdfpaYwe0MViDISjWLoBs5c3ZrlI166kneecD/2
U1TBvllwiMz6zMi6G871+1kXIae7bT4rhmWukczEP2UgdTOZBuhwwBML8YL0uQK4
5haKfmxFEDIeX5h/tf7fuil6ZkQoJeF6pkt1c4ATL19Q9fhU9KghU34HBwCguME0
nzRpST3HyGdnK2TWUZr5c3VmLVSKN6vjg4/JDlW/HICMN1V+ez30sQuyvHDohak2
C3E4ZTk5OcXZCX3O+L5izGLQyZEln5F0S4Qrn6d/7DhM+bVbO0EczdW57GBhgkzm
j9DJ3JP90WR+r019e7umPlNJsVdi/AhSbBV47a1Yvc8+mK43tdzBj+zrUfEGMm0L
sbhAB7hUaAEIbWxfCSAH6g1qd8jBDozluMNfg/dZsJ7g7535yBNfAEhK8JgcslZF
R5D8n/J7z3e75Setxi2p+8z0Ck4NxDWNj5vpGY/oX0YG2yNS8NgdSuc5W08PfG+r
cdogJr7iUiS7BTcR4V9gW6JiiNgE3MKwZBEe73P53V7S+jy0SPEvXAPtsTY28BlM
XG3QMgS4zQzUUyT+XTOSYXAPRn8CxlkvJ80k535ysFYZIFHcm/iIfBY8uh013Aqa
Afia0F/z1xHRfaARt9xiiy/YQfgyj5MDz+MmOYinsD6qWmiJemlqzFfANGDwqerC
jugYu/BVUI8pTE4R0Pnr9rFJL0XEyijLNq4auOyOz1BCFrNOmJms1RuIbmiUyv3j
UfqI/eju/cA2V1MXtCqJ3wJBj5eBtKzG9HXBhRWc4hXhMip3fhwqcSKFMBAcdH4c
ctTtbCrQdrCSf4uLSDlxHrbGtjbCAXYtUZET/Cx7ArDzNtq5PA4evn+AsiwDm/H+
EygWAfpNxln3GI5mEB5E+IadbPaqEYj0wlgMTKxpMq+6jhj9Fp5F18FfxJy9WE1R
qYjdbd1YqLFM8UV5UYkM7Lli4ylHfRSYvS+joUFhSnNTun0eVpGLGgTcggfq8X+w
F66LhRcytiHY+1EghVaW3xlsEfVKNwzupjEfmEJ1jZUmLkZVr/lAoZVEE/weBfrF
B/JTTs+TXV88G9qlYtiNqVqTHBpNu0KU8/0up2I9xLYLZ4/aJCCcB/uc0+WFm7DG
b6IKDN7/WaBlBko+VNBOOy9w5BBsf+fqHCMi+TXwAdhyVCwjYO3012RWyzICRJa+
J1RIg53oWa1u21QHRgHb0KzGtCRfSe1r8wy0WK7MU9OhCHMnPx0IS9D8wdv/Mx4T
yo4DMfMqROcIvx9sfPQ9v44//1GHr0FIdA/WMfBmLjQ12JKL2oTh9pT2rjy3sjel
Y6f5ZIma4XC/S1E3tqoGpoxuchoq4Be1JuUZPSvFI1mkCK/e2L4Lm8qGOcNsp/vL
rC/JPqcQuMvQp61G7Hu+Bqe00ioSITILFjS5N7qWbZd8aFP24jvXY3yVLvQO2HVb
UckjgZfsQWADThk3vg3JT42TPgy9C4VC1UZouMa/nQe4YMtggw6DOmF8w8pYUfwp
C21A5YHVCRS91z9pa/rBYn4Ns/NmvPk0I/MLr6PcRNPiig7l/ipkxTu5ncazQcDc
v9kP/kvTNHjQsq2szKwXVhJqdpU4ijtxMJXzUWF/iZoCBgNl9iK3SJsM/0rdzZBZ
n5G7OC8rGcKl0UZeWm4xAMoTGSmHnkhUFWjikuTdjBBJpBofEBHCs0Lx8jRJKq1t
9YE8cjwFyoPDpqOXPaGURdjthAY42nGRhEyvUocgWpTgGC5wvG39+0GtLT2HkeWh
+xzlb5t+46Bm/+1feFS4gnTNfQANNwRBnB+G9Ox3lt9rKathTc6/Cj5oM7ttHNCP
uXIMLmRBp7qOHS+EoTpQEal3MakQ1x88dgTwBCFZdYJ7zBJcrWwGvGagjnZz4do4
BIggncr272dUIiZAthMQhATg8+I+/svLRRxVVlmhmm0fbrWb3Pntm3MyWhM2o390
YMKQe88g6+F3pJ1jBFhRnYkFrxdrvATGCGhPSMQtnM0sXEwPDXjya0DYdu3Q7ZC9
YsYCpbnO0v+AFrwfO1ByazxoXHhyBVdWnsBMEdMz4bXpCijPJ+DQBi4mwKe42I6Y
wIKtB4j7OrSFhmTxW/BgZWvyywTjzN6jrBfCzu42HWMhMwaKLkx+MgXhJ09d5cZC
SWg7zAP/mj7dMocbsc8ALzu4dW6HxYGNIfbsMiQFmPNYXipiLl0CGrR5mKPzIYZn
NmXoFO3zXz9vEbbOAWhsVLcOIZ2zOe6VkWbHdJmY91YwqwYWdrHbrBiDiX3qSFWF
5FeHwe9DicvMg5hqjC5C1ER0ZWkfK9akDA3inazU2TSO/nOOEI96BrNPLuK2xaCV
kY/jlsz4OeA2+jV7HJ82+TYWL66Htt/nDnnvPg60+bcIXhkySS1PF6Ukbe2KKufQ
hGfwDThx3pgWTrVjiuP6WxYhd6OfERUwMbmbKYvxBeouHJkoP+vQwv+aJhpvPge7
A29ARozcXz2//yS/rCJ9IMaLuoLI8Grv/BprJzHiAanEb2+uEfgVQ+fW/Pv2w3+O
czZWtgOMNuTSMsedplFyQW6E3aeJPsvYJsbK9ZKVPh305CzvjxEjiNrTdGb/IW9G
9/XOCN6/El0UfrrxKQ/IF4ZnJ7AwfQTEk38Z5rHF0vpXgH3Vv77jNN928Ax9LElC
00EkIK7DVmLgyn1l2KqiBe6XJf9xHpok2m2y254E6VkPTQ9R1XlFqglEVv2K34xo
bpAQhigfXoRWpGrlMXPD7hWJiFPGu4cKr21qHGjN45I+MFntjyvLOup8dzLc9aRs
`pragma protect end_protected
