// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:53 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dmLWjTyfGxCVXOxJ7UUyahs0GMGtb8lxrDAr6/rR1rdNGikobgglL9i4gTbGzCXO
3ZfvHLl8gXPKFHzgIY+7u1StErFC+xo7YOJnsoPo0O6X/8LRj8v7Ny9gAnJlyn2U
ujQn5ZHM9h7UemxsZHY0fHHt3QUVJikFQQSQgc5JRDo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5280)
x7QvDkzbmp/ixFUgwubddNeuwsGaCxPK3MEH8FwqlXH2bARRk/YUl2JeLcD7QWkl
/3Q9jy3MN1wvnnf6h4S0IrHGx2KlZvbv95gETs/qg00hwmfXgtq2HqQLDqbX3OBx
efwSe0Wwx5Cg8b/DlA49J0XK2qdZ/AKXfJ8n/W7Sr57Pl/sUf9jtM/KL2ZqBajNM
I4YiqdrqbZNdDNbXX23fs5WzpINUvoiRHWx3c5RdMLVvf5DViVNz7jGnsEuAiAus
KdxTf7N8/WSF8tM4OLqZPpEWKBfEJz0qHYRE313sdnFjQPXKjnkySGDb5UOH2wij
ADjrndgSi7rdzYY+EtDJZnmOOFD+K+oLfHOms+j6fP7gH/bV8uRPC92OZfd7FVo5
a2wtG11CWNolN12d5HcGcOH5gHKqGGpMPioYT7gNfMsjgFE5UEV+S4monKLr2zbA
Nt9MdNGpMAfZB6VIJiWr2cLB/iMihfY1Jf6YMgqER+w5D+t3nUdgl/lAPGfOv7Z2
rCnVL2jqSGHigpid6jq3fVyhH6vQ8Rqnl4eDescF4ooyZOwc5giG6bo8NpZbSEpD
AiOWJ3dOAhRtiVvRI2i8r8qaw6R6A486MdsoMLUK1qF5yZgIpigsBArxl3kJqDal
Zu3CqbJfVDSJHEmvdYmynP7fIslJuXYDVAyd1qJngR8TRoIf5xRMRQo/09qup4Nx
ElZZZbCTT7jROn6rkPumM/VRe/lxXbZTzp3S+r00Ts+lk1O5eFpEkdbkdzwjehuN
8rP3OOG3rOaaInr69GblhQrmeg7xKWbzF69Kwp1rLzTAcSxit6JqlfVYy1Evz/z+
XnGzSS0bZcTdDuEgbIQHdeIYoQ4shvtv2YUj/KkusazgSXZ1Doiqdeptdc22/pqv
WZ2osdbZHwuMVlTK9IR0hNyZC5ZS8x7lF3kvNqGUEt8MSAN2y0M0YlOdwrCLphPe
Ufh0HzDp/Evz54CaKLYhy6MFFvj9vePNMm1yPf8uPvMKIrmebD3MiN9qLqmpDAQO
Vxy3JvOmVsAvcusOq2oz1BKgt3Jydl/s2zPLmGaUvNoTD+ooWReFivP3zY3ebJki
5L8WXv1kXMPVuTOqGS6AmerBWq15OfZegLkN+TPFTd4cUfsWnXFBEX7vkryv/x2s
myOhxindzLrx7hj/V/rh0kWNd1DOAcJI9IGC3eB2POG5Qs9Qv9Uth7RzriJU/Wv2
vWOEjS75z8NxqFbmG628jdyrtrFodQoYaGGDOv8gcfkCHyub3sFA8dsJXu12DDku
h+gNOrVZLoOB2tdffg/q0+DDMxFGeq6qu6IWuEOdri9bWojnWlpmFpYV2OQ8lG9P
QK7hWV1p/a9uiPGROHF5ebskPfEmdopt+51Od0wEbhQVHJSZDc2MVKX2auArBqA2
jUJgQe8yrYx2rgwrrVk/StveJkB1c53XLbr1OSslAc6j97OzrsaPgTobhpM7j1TX
0e6DItZ0kg8p1oV5IoQgSsj4LLRXRKhG/Z3t5QEsYuueCQxCrCwn8n2JZTGisVKV
vHOd/oVkqiikcwl8KLjP7gWYd9MxGNURSiJj7acA3BNmRbfOUIJVbZKTk+Squ/tx
lE9/T+eWXjdjFI+gBWEUbSADaSAFZNGoNntu+7tBqqM/bjE9d073SsGmSHjlCWlE
BC/LcgQyvwf0I8ioSMjaSDqL+KZ7+737G8mv24bFn22XwgTFTGrfM02I4mM+I/Nh
W/FMTwM9oqgWYULN4OUgKFIwzbJRtToQFY3lphgVkqK714oKLeBdtOaZvLhMmdFp
7UZMwUpRjqdknqrrLeo9dCOugGbjE8pIGQE+k9cBz7lfIK61eqmSMFl/fetdVlue
0vMEd1586nAJeaLviiyU0UjdPsm/y9iXh7lGjRgOKJ3K0h/pV3cmu036BPi+J0O7
ruZTnNMV1aOVEw+eVowzBUPG5GdokU6qOcKmUednnoLfnUHfpV4u+uBhCS+ZCtx1
RJZzVcvYhQmwg8upgfj1Okt4C+T+0WTlQF9DgS/HA8gOVy4xmAxqlvGJDZBX8aoB
b8VnVCd/2jkZ03YY6aPMBDK67MiTdVdxr2hkiOz8N28IVbtcj6NCXAH4TmEKFSl6
gqtCYEwVXQ32mg5TiIRT3tUWa7cx0P4HB8QTeQAUFQuCpPBEcsFBhxsOu+hmYZsK
2amXCfEGmj0MoEyhVH0ytlqMqlycox6xhgOhm7zddKgx5X9czdBiEz0+awJk4qf+
BB5OAyXz5WEH3s9iVoP/1u7OXluLJwobRk5THr9/Lbu4aDeCqp1y66GtV1MdYew2
sflbEP01O+mtYC+6HOHGpOiSLpdNcIt/PTUaSdjN9P3GZWt5VDCPxZBOjGtB43ZZ
BKKe/wccMxSLjqrWVBon9DXbTdyfJ8qAm/t702EXVK2bepJlq5IDoC+VBZKvjUGm
daetXEdnEe7gdH/KWEOYTrlyFYjHc5fgQ8kxEi9WnKuiRJdJjt2QjmoZ5UZSluGa
EZq+c02i2OI+Zivr4vOjDlta+Yt0b5b+kTWRUK0TCeXsLwNQorYBcMnT4oWo6Mf8
kt6XwczSHhiiB220eHYNZnmLIL5YH43gPsGgQ0H8toQYo4eHCuJ2NzqvVn6ibCaZ
l8NCWuEeSR1UDA9dd7VSSH5H1VFu9QPOzzZVwRLbcfw7wNVO1vNfIqNzx0lvFX33
bGuIt40rfJAesSgS5F2C3Rav4biUlSMUvhpQ1HfhBnqJBqQ78fn2ur/l/t5VNxBY
bqJagjY1JVGiXwu/LyONs2kZHT7BmMy08c6GNHVxFHS5K7vaonnF3TcSgr1N33qW
YNyRqAhhKWatDj596wh7Hz2ll1H5jgCeRFV9NXSz73jiOZn5Q17m55GmTSLCo4/S
0cMMMGC5Zn9q53+wMmKGl9Vk06F+JW0C7AbC3MeuUfcBMG63dSLmVu0RXaC47RfB
VgFj8Xi2tDX0gLQmuBUH/rWPMwDGyu1twtUiUZkGrTDY8ptPYl07dGZb49YXT5mZ
uaSDvQ8a62+lZ9qXEgh+V+g8AacZvLDz4oXUv50Ys7rkEqHDG4F1bnkqUVAJWXCr
qpiWnZXw9cwFmONiJqob9XWoS85kNAGizPBYgHqm1NS/3g6gFBjhwZCTrx7OBwpt
O5mhexqSST1j03+cUNf0HfoH/FT01XUsV8qbR2rtSRxedi6XRBT7WyKG170f4ZYx
2LYNirL8MY62X7cEmUaQJ99Sc1F1guiiiEu4y5iDkVV5OtN6leHYt21QKFmCOn2D
X3UjyNXzp0gkj+groR+5jBkxSUb1WL8aR3bjUCNRwELO1Ah/8f53SP6e0apvsNgr
PCc5iq6kgFCN9qNWdfnhB284TpM64vVg8fVDn8PpsGXZm6bTMc1/neA3o3aP7Qgs
KrN03nrA+QKTdQqNf0lN+3Gd4XP3j0lGMrMgaos6OaxnqkoLoi2YKZq8j+wC1GFP
PjcNkxphXQZRL1bapaBt5W7UmGGZvdmvZgIsobgdYdj4naQJNBu00jS+t5Uk8bRZ
81f4NuZhhxAjBE0H3VkLonFjxLBEPIj7X+KBkgMglBNHOkRJlOuGduGBtayxGMl2
ueaQ5B+BQXymrGajSOLEWKpeY6pKq7eWq4XjVDJQTAFw/Q0hQCeubsevLcgH6a2T
bbDkF34jUWpFYP7Y9x5f/UX+iGNZONA//xjM2A/okYQ9G+CNpo1VdovrEQPzfge7
jcH5BQJJM7gb1Ra1i3aELpJ8TcX0WzJ2LQxYmnC9MN7GHIjA1ZrPpQQ+04DVA3qw
ULov0YdsyzfvQJqY8UyXggYvOy2+rc16j47xN1fhHQAMVcACWDsHdKMarvtFKqCf
5iS5Dj3A0FcyiwFv2YNBgO8OYsj/YFBnX3UYnF4XUkYj2HgOvHBMbkl7AUyCZ3Cd
8+GO6LQ5rK71WSDmfc7eCy6rcdUuRqsoNRN9F0TEE5eYdpl/Ak0VthjrV/Vbx324
RupXviE/4SqDL5wYCNIuDkdLW/Zgt+W4TmSmF+5xVE7nA133araVn2dA7QQuPFef
NvNnjXFvrWd3ImOHUeGlCmiF1BFBT4VoYs3f+kj1VvgEM70lZrXlf/ZCJGgU+JDY
Rix/8WdA8gtvJsfUNU64At+gietAW6XAda3FV3sdV424ZiPpq9LEANkgVlZ70Etw
k0oifenbTlmnDkHqIovFKo7/S3UK9xuyDzZodOmyrtLxLFNylzjxoJf8++KD2Wh3
IdbfEe3UTrT0BFl6lAatQLbWx47KyV5teBQOzaBKAcOiovXgJ3Q60d4b7M+IuwJR
On0eu1LeQ0tlewgM3sVVT0ptcjoYwvNQr0Pa6oJDrwZctjnb5i2cjIf69s1atcpi
4yI4ySp38y2M5REmNVjBaEpjmS16ZHNNZJAO2e6oxcEMT1d0MXFkdjTGhx1IVmAX
/kA+T9DDXrlf+zdbrAl2D2RKZy02xI0Lf5Y4LUO1ZYI+bLxY3ra5HnUYBWg5v6du
ANVX+hRWGznCUYmSAQFskYp044rSvTKECKAJ6XuKldiAYqN3ePLc4sjf+CaY3J+G
g0/alS7IzqUSwmH7FfdUGop2I5fWsjX8jagkfNZBeucXaQxS+zFbVNFyVGndbxhc
69as71UUqVUdOZDnhclGm9qhOVkC/h//9sG/iio8g9ANVGoCyAUZ1ihfeHFAuGxJ
YlN8OOF2VOFzO1qmAUjmqyahiRoGa10u22jak/tWorsShkUGzipqnOCqtF7Fn92G
vjEC1Km7PKHbcqoMQ0RApRE43zOX3Kja+xieWIIKLI5dM8N0zusof0e2UkkwoPzF
XgvVY/npXRsfyh6jQO9bkaCik2dtUiXyC8yuasI2pHhSh3vRDuCuNlvidyVDIfLV
Riv0EqYIlOj2GiyH0YtqKDwyACwkv6Ohz54CzgU7eT2OchumeewFIOZ/xyXhLtaJ
scUPFQPRZbkATBa1vN/Kiy2hbbWQiOIa0waGTs7/Jzt7Fn/UB31eQiIYNZz54Ntb
rTeMbNM9iyXMhlhmWoOGJxrlWqBS1UCdCFVTl8Sb3DldD5pB/Rq5EKiKffum/rE6
8HCgDdfaf74EhdqCJ9go6vJWDAyRkv9Qn6P7IUBWMg3FxTe8u6Y8pvlKmVuPnrgg
uV1/wW6QzjDLSl86auhZyqvE27nQc7FgPHwifoUsc0PTo+YNZq6vjzpep+yY3m1S
mixuU0oGZhzcq5BtSpheC/rC71B43gHgp9ZvTXIoBNrs5YRda91pCbI4MEmhCybg
9OCrZYdf9ICuvDcJOma0RF88QHHg/HNfkbnc6WOEtciE4wECyThWtBX88wclGXQ2
W9zTqwpr6HEy+NGzQvXtpGcYGY7TgnrkFtD6JkyCEwljTLHd/oGyO5MWqTFKr+6y
+AaJkU5xrqsNYSUisT3WkOBmVfRgDLCCKVe6oB21uBBPbOse24MKM2SXvbjKDrkJ
7wjUaIzNNytZ4Ja8riKK0yIeCCuO10Y3MyvIYxGnUQZvj1hSjZd8G9vykzsCQ7k7
ZTBacdhxo+3V8OVnVk2vbGRGYhg7ECcbd8cMlIW5zrDK5gVaLV8ebaTUwmSFSlsI
qcn58b5rjOZf9pJKLzPJ6JHjRiAN+aSNgR1KK1Imbdj0kqZzFASVZQ92NJU6mYTZ
U+tTQXQnJra1HF7tUlQjWaiA+swbrfRrZDaRy0/8pW0vgVIaqVfX/ta0prQ8yq82
TG/abP5renzzIlX9jTPbvgLOaPwIpMDuB/CRhu3k3MB04HYZAaDfreWpBhWD+OIF
iLTyvS8K+dAt2CZJTuB/g1JCY1T1CGFP+Axae8DNBMdTnOFaNuoDymmyUZ3V23s3
J1eiPhmfk7w5PyPq7Fx6hJe1dRN1jL3VWhC6ClnJfRjGzMCgLmZn0gYfdJFMIUfW
0FA/rLadb/Bvfb2OxTAx98yuFjorBFD6XAts/5qKfd1rcuXeltCEWagYvPqE2oLA
g/f43ABtSfby/RXIKd2vr0MvN23bc6343e+RJULWsik3u9xeICF0vXycmyqoRSIH
9kLzo75f9IKMsp4e7vdgxLrZ2K/sEhIwQtEC7gIL+Px/onjQSIaIrZQrGdFDhlQw
PFE/EetUqyhK7cBBaQeX5LTwOZrr/eInXH3MmuBG2ug3wfJXDgEHzsr5CNAksyRa
Iw7HBwuFwqacRnOJHo1/dALayZHBC+bHJGnOn7GXuHDjqL6l1JX3tgM6Nh9Dc70k
nrNC1GduQLr4Bbpa/PCqMxXNWOMgJUllUSjQVs6Z8vdOmhyOxVWKm2FmDItohK3F
Dtoyi0k6YH+SeVLO8ZhjiudTBfkva1h1cfXYcjie5HLKnKnacjqadxZA4fQoCOqD
J6Xcf4d/gJGCC0cfGL7VciDg6+yYlNzF4uJIMpp/gSmUFXQOoUjednHxp3hAuIRP
xakDGSCIZTJAof5aylfXpoanKCAtApWNOy/+TU3F2REEUjN2SvGQ9MEhDfouMXfe
Df/QahhtsZAd9QIrAlEg1fyFrvlbUp2kXaqGncvEVcN27ukZMZX4KMmXl+MAHFAD
b6ot/yvG3/r3zyUA/R5a7ICD2pjw6MDzSzQymSzWXA3L4xmrt/radMKBz8yFJehA
AhVf/3DagqKcN8JpqS/M5gXdUhJDkQzlL4XJWRiFadjleII9L2Sx2M/vpMVmMHxJ
j4t/qEcsmLljKExtdr0t/qQbzVIV+PDEqdVcqbuwJaKXoGY55S0Os4LB1DvNYDTy
zJoneUIE8/SyDw6af+EY3U7hIiHZ1vmSJOujC7Lfh8qZ8KgSH4OSdam/Ua/kNXOD
w5AxDs52fRvLjyG0MLdUZBrNMQTWYHJ6ipkrGSYp7hKSOmQm3bdFRZYp7jZn8TQ9
AmWwZvCUV4Hf1GMtszZkLDL1HW/+aUGv/GG0iNVei3eL+BPTfPpXcJ2dx0ojwMF3
xhXcoBl4S8qf1lPNhZOW36zdPesXu+Bpkm4aQY+EuRVCqrxEmTyUdZkwGpHL/IEz
OMIFnUIQnFOR3YxpCXR2sWtIOuf7JpcIKE6YgfU2FQgxZ9AmKZVKqHchDXaCl5Xe
`pragma protect end_protected
