// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
XK1Hc1SMg2YmhhzhbWyGn39Hd4Gu+Qgh/tgX68v4GOBdmghEM0GQeKl6+L2zM6fQuSAUCqJNQyAo
vzDIIzL6eFAZWxKMhnIFIWCymq7pZnSt8VZWkhnY6Zj8jnkQO1FIwQMoGmn/8micRDd0S7KI2T0e
r/+7rWHre3+ZABRUGvjsE8yS7p8GvK2oHWGjxYQIrtEtMWKaMtHnRjO6BgvymlS75ic7BjXgHZKK
msN9TF77HzRQQxCaVItSFdVXSUddzKetzZwgkWhqNXl4EiGHJbYnkzeFsaM0SwtLTGghxVkn1Euk
wjAKMPMyAgF47vG5+I1bQXjUs4e4tycHrjRpcA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 26320)
lGyDZGMhW0Aq2V0aAcTyckEbjluuAM5e3/xk4xQ94P23JKTgoC8ZaNkIFLvSg8PeNPtmfg4mgz/Q
HFCGTPollMFg4PNlIfUtLn5jQhw15AGUE4MdOY40sLWcmeYP0GCnoCY858/6WLvC8kvOcTYwyA56
cJAmcqzKxHKzOxf8QK+e/pN8Xtm68qyCP6WRs33Yw1Jf5xgc/GTodSLwWqXMu1Y3sOEw78Qg8z7m
l93R+1QMirMcLia58A8aatnTDa9OhSXAJRiVjth6DWKWsJwrY5u87J6VlaCWG8RX1hdJgSUJmK+z
457xfFB+Sg9FCA3R26wd0gqnehqJ8yZK89V1fKOHpco6shaVktccLvPUOr37nT8hz/afvl0dZqJd
mY0lyH1hZi8wPdJpqF/ubMrQuOJNS9+XSkX/EiY0yYwrtk03gj5yMXBZbJljqCM8nAGdPiVQBgUr
Ol212TS1TJs3V3mUTm4XChMabxcrCrh5BRO+jTWnFEBmz2gAcf7kGVo7nJ+t5aInocXYzAKVygW/
Lt5sSZG3brc+bIJ9uzNNd4nzUu7+MPp3RdL3Xs3+TuxOgvzqO/dH5fXqpO5h3pWoB3evFgu+17Vx
sRqNs3yGZCtDwb15ANgkypKF3moKIuFLiUIgB7+OCldLGaAUAvTgBf3WjZ36TKIPcapHtvRw6F0/
O1vz0CrNxJlJfRQ78hWbzyEn2j1KX8OxxoWLLz3puB2G+tLP1IWl5N15qChc2+vR2u+sss0Dn5b4
nOeNfnCTfJL1Y+KY05AJhbSwCAm1h7YRDa+mrWIg2UV8V3gw7+Ajx9U5YHYSneIdEAEx0VwBIHIr
bmnbx6cwloYzR2b6SUTfq894G77J1sFuO682DHD+2EkQGig4Hz2ZnZprzqVGNBaYGHKzPlr4DZTp
VPzJVzn+XI0/SuhPRmlCLZ922tVKDCRRV8xQypZXDr9aZDT3wdGbhoeFy5Ds4YI/XnvXbFydcWmL
8+FjixGgK7VdfEa9m2pvdNBd+tIiMSdC4TvwhAzDN5iNuSHNS9g/dLRbdbMMxWNCqd1o3cBJlqLE
te4b2huAvLv/XQ6/uQUT7UExJU3ByRC6WhmaQXq6e9w7dS4Ymm6IGFgF3vzMWO9sj6/MqshGzhB4
L26uvjsotc/k8YymyyO3W2dEcYEy1t3Oriec6XCr34YAzg8Q6z7mtLW86rJ9kTyz2JQ3pJ69R4Hn
y1Wz5Y6tFTsPT379RnAHrGKV9QBNa4LyIrQKlIvQz/1LhR0pnRbbjXcPysKqd99nHeBuSFaF9Ecv
MSRu6T0l2CvUJyW4dMjrhA+J4gzvXMTEdYZj/JpYHagNZsfReMtLh4lbhC8NyBHnBUwWdeJPvkHL
0JwXf/vUnRsY5NJ+p7LiBeA8dg3woYVPt0P4UJmHNEUx7vvDJHPKxXZyPTvMcOIkQ037+W1tiIZD
jZf+9GwRFNeG6PrsetgE8cwV0cQylGX71AR2zQN4nEfWR0Mi7ehGPgAc+qiyn3cw9CuJ3K5KBf1L
KGKkwU4mlJJsqRrfWivkXwGQEHoNENpNXJlhFQLlGoKhhbn8ZO2CCscOi9gTbGfx5OSxHsnToS1M
7QF9UODbmUaXOLL+gM2xhQrSQu9FbfLfhmBBYyoGxMnjVh47j/xvPgLiuuYU2W7JVWhFqZVs0q/L
Dmt9VeBbG3YDf2uPbeg18WypsxkQG5UFyRYCm6/HcfKjVLvf7SzRu/1gIaEwDov4yfWbL4AhIdDn
a7mB9K6Dud8fFJgB07Xe+I/010ryQBzWPaNRG03uJknaO0WMLBQOfsvW189Uyo+j+TrYH9omrVOt
2M1Pw+Ou4/RAqeFgmK32FIA1wKByeUoHTJyAONFfWnkmjAyRUp//sLP2q9yB4vGIpOz/0hW2XCQS
WJdg7nIEK0+QjEa1JJx5l5oC0z0ZBRfAXGjMjPka/LjdfDwwM6TuScP1r8aPef6Sl0elfkDbqRJ4
cHlRNM4DPGQ5oSZyphpaSqx56ee4ZZ6Tyb7J10F54TmrXO++jhhrzdCPaTqtaQYDcBz5ewt5gjLR
FEbaaLJ3yurPEcXpJvbzdqDA5UfU5Cs086KRyx0DmA9wZAmU+nprvGteu8+mThV9bekPWPW3eytP
9JQDNeGVhyBB0cBounA87wMzyXe0rVee7YeY+SZhOVpT1LJPfm071B0Jvix8mb9CZ8o0g1wt99zh
i5TBbdSYXH0FC7aIf5eB0SAeV861pQ55oi5zMm5FZpeA26gtJDNaNt51DVq+ZH+r6d1L3K4CQ0NF
9JVqOcab0XyyoxBHvM1bKRsAX37zZZEbt2BiPHS7vLlCye5v/4xQ837ALk6/8TbrvFlout3GLr5H
+1NX8KLv4sfSMryM3UaD4JXJ6vvTV5ubVzur+shdiJPfG1fvOeFHvRgZiH/2fgD5Zg5E8et4+TBT
4jAgjf9SyETDTM+ZPAHxc/qB3pEoTAkQeiOET1SzTJvBe47rYcCma2i1NKLaGwilrEm7SYZTqu5J
HHV2hSj+JBrMNFAgw7IHmkGMG7NSZ6vky4GYs5y6paNNF1bpwRIxhqhe4nOQPVqYXdvvbp5Zs2dB
PuVF9ck4gZVgodzYtg4O8USZist1xbo8vibO8vKqMeBfaWjYW5tSAcSunOVcdZ4SSDafpOTbzixT
KI2xt4C+SJ9HJAfBQKr7LNWJCJDpoUqmxdSyjICWzSmr9uW2nN17+nWnUyyyDCNh4K7qNGufM9tW
6ZYlaDtvOR8YKmm2T/H5bnmzKJ1mxSLEc7/sYrIBLMw+agmNAracd/QXif0pl9dUE91ZpKCSCw72
qvOdvJhW3Bx1Ia9R9QFXWdq/6RIBvFxUcLCs3VKqcDlysNNUKWrkb6YWk+ldbfnGrKNu2Iyvwhda
V/PndvN297NjEVI2aglmwFgDUtzMx4e9NR8HqV+dnTxGR5Vltmru1+CxGR+OmXkAO3qqyTAheKd4
FMpORg6yUQRL3OiwobQijkhSof8GdqK9eWfBANUAGJobIJYvlkN/JdNuR9qIRjl08WRe/Fag3aCv
LniUBKvcbZNan4vNKY0xFLfhbYbARumeCIOD+SaWHuoTCB4eYIM4BHbihWXiO8ubyrd9LouKB6xY
KAqdpUJahvyAzT9vUoVBqGet4gB+3oAMZ1i7J2PrnGtkyfWYe0PZG2IHLPDEiYXkrn5NlMIBHD2+
35AsV5F0jNMenvCqqkAHLv5G7EUj459PKU1lOhVThD684Q1MhPPLTeq5WHT5bd2PCIShWDPs8Oa4
CVzxLtgNRH94fQC/6jlcEloSbcHzom6w4ZYE+Ili7hNypWhX4t1FFOuG8FOqvN0VJbW7lmlj84do
U4AYkTmhoa54OKvwkfcqB3bPQH0B+cpsRDrFpOVqH9I+LPqotkQ0nyLinOKNuEUahscxFVS9SNDT
tUGpWwIF8MGFMaB8hKj5zSTZMTdPWTJPE8uPb7vUrMYGM05KZT8VYRuN44PfCUzC6rXsBf/kn+tl
j0y1LUoV6ALxvnctu7AOtzMTBHoOX+bNzU7LsOACZSC7fCPt8qYU70nnola/apOfl+tb0Bg75KSO
9UnL9R4+LII5m7Y9IVyiPOWjttqKho5qApAaUpEMNhJXc163cmNNyg9W6rAHyH/JMuye9ygU8xYg
9pVgZskujxPrvhFzyAqkYmhjkLbiX94RmVonTcsZhiPfdPraphmXVmqR4zpIqdKpaJPT925rZWXk
OTd+01lei3lUelOGHX5T7822vg1YhJLEHHTAc4yOtpR4iX53xJ/2df59svdtz84Mq9myXfRCxxXB
TvzwYNRH8wKTH4bK5BnMpD9AeRPM7jIC+3YEMm106lZ1VPrHv3ZsA52Hp8wRXCMJaV9Z95krw+EB
F+JUZCoHNrEXMVk9xsJoSEiAhOw+cfjacjeBjfpvcxqF19Kha1dnmVhWIuhfiXHP4e/VTOxNFBU2
2J8dztKRxuyRJuI8r37a7Kak2VhGdOdeD+x7EciWr2XcK1cDgvfVB4J7mKwnjBVfCgxo7yGhKFME
jl4dgsdqslhw6ctwohDyNPnokFd8BpKw++YGJSJzp6TKBsEGpAZzzgOQrLHe9PYcVZbiQoZtXn89
T0L5Xcrk23YYHjm0UsTfeg03S9x/Mno0mQ371OJQg3TYydH+xXllfYx/pOOTTQlyqvx4qorFCTUM
eEVfT32DyImvSxr6I4guZpZry9jGGc//Cfjh/lfVJ4cLPkPGeQNqfJsZyNGcTogEC2wSG2I2UVOB
Ht/237eaaYJX3pjsq9Uql6g7fwlYh2WpCjSE9aRE+FNHEYyL9AwkTuoWLpDD/TYNfpvKvpbbceV4
kdal9a7EMIgKT9Ql6wRfsW8+nsA6zzJXY4hBjV5b86y2k+LN4T7GrWkmTfcJ+oevMvFVR7384M9o
OkGEGoEpx9t5Il8ZmRUzv80Dqd+iCpvO+oP3DPBSacmOMF5mzcsGN6KkxlaSPxQFNhDMLCLpjIT+
SXkAbZ7Bw83+3q5WzyXMolc4KiNACL0d6SP9MB1MBb1TRDxeaMMh/9xykx7L26j7hX0j9+ZLllzV
1gfKTe2eXSUt+Wl8UBB0RyXMyg40jdEXhwhkmor5UtJBXmDEqFI6wtPpNbfCSKXe3IXumbbp+ulV
L/jCMFRpk5furYqd9X7DdbNdRhJyEi7UY7sTzsp61PK7/K/pB7hIsOBh1tqYS8tqzN/DoHPJldmA
docG1hXW211H9oEiaNda81cOP6nBgJ+ajRlHdeNXXEg9oQGvKmTSfLOoKpYfFVoGl+BhGtQCeEM/
DEUtz/AkNntjC4pZdXzNkHAqpLeaJZXmqB7ozzs/yudWyD22tXUkDy7BtH8EQf03k1ned4lILiEN
S9r7qVSNQ/U4OjyAeFtUIEvZiQ7IlrFRaDTZJxJiKxdQ6GNoB/nHmNn359p6+JUJQ1n1lhQSYJDX
73tSpevWSHcZYinUIeabEb8G6lQCD3VyDOKdwzCJtzZCqqDrvRftawQdiWeQI/87naDgzveoqYaH
8VTIuAd+ZXKGfjwMHryYgbpHUAD5exh8sCp5MSr05g5aG7xDaGNem2MxinSlcIX0zfFl+ovJ9y6I
7kle15fnSg++eZHX7+x+v5G4BGJJGJClyh55MB+Bn2ePjS5Vfd3eRv1KKKN3TV5T3w7BYLZapveT
uM6DygQJIqSIByEs4SCfXyadss8uUStmdjlzMpcBboxDrtLh6AePIkuz6cWQP4WnWlXTLDPhIdPj
jiOV/SaoMV5RmwMfLIXi/JjLzDPktjpWnuNSjDJpSo6t/wqglAuijntvY2KK4i9Sn8JbdKOfdcPL
2E6aiRby6o/Lh7u77PN7R2Z/ilkWAPmrnCujJZdku7tjTPwFz7T3S2t+orINJ4eRvfKbqT21SQhR
qprNDBdOzbDEZFtcNO1ZVSp74BWjQLPvtpUCHG0UzhE6pdL7oy1/0O79oOve+AyQkNlt5NOYy8vh
bgefRzseTzEfojIP6/E5vWcuNdELVL+zgHKC9Rw+ENJQ1ZBbsmhz6VO3rne6yjbsrKpFg2bLFyTB
aj+jV832zijU9WCnCxoyDvUnmhRR/JbR415/28yFXpGBMF1/NOo6kDSRYNDXNOk9g1vkgQkg5Ymn
A6YHdMtjjCDx2ZtQ9C9rrfLFWZpTg2y0v+S6iOElnAgj4+Ll0enPpYh60j7E89lgvmyMuaD+N1hg
PvdbA48utSC3w+8xxOQsHklFo4pghZmY4YfLgYgWuOhj7LEQYJ1XH6b1G/kxixdAIYc8nzzBYJvw
q+R6ZBtomt8TxRS///Y1QIyt+TaMaov1TVtgtjSnJUdcSqIYmNJb7Y1HdO8al7tx9jALoou2Qr+d
WrvOLVvlmsvAL/QLH0DtDHwgxEJCYypqfslyHflQVL991+DZL/4Z7XWSCjf9wTsLejUlpCbWDEuv
Ag4WAvaXhrjxLUtbJr6MPXk3ZxoIl+dqJMrMTyhhKmvFnyT7v4YCyfYdHvTbVZH7e76SB1a5d/kU
ZTy7MNjXhvmfsWQwoAHLqZTsUbveJvxw1p2SVmQHsxz2Ep3MtqHUMT71j7uINNbfQ8KOP9xZIc8w
n3R25Lj6c5/0xWljjvQrihB1eZcyjuSLTnqtBO/PlvObpPkiQi1JFg6ayHA1IyEVEM3ID7UC0miU
R8lVCw0q96ld+TnAuB1KE7xM/V0IDSYbBtvI1gbB81QG7B60D3vmTA1LbY8M2diElyRdLMwC49XG
0zpikNHJdqQe5vI+auQ/GDluiSFM+ilV36Emb/XM+W25tIfiF+WtjY+ya8f4aa1Uz9wvb9cltesm
+aWEXcsr2fEhkKPb/hlku68onoMc8zIorajHnqKrmqvH1XiapSC2g/gearDbEmgLbMRQiKgWe7H7
li9JLxZmxswjSsL97cxvSteoJQucZ+CrOkKI5/8aD1jkwWlRL4OKZthxo457Y50M2y0eHRxulfhk
Gu8d8XLFbQ3fvx7eXSRJjHLlfPYTwyUGTgPUyUMoCB5nCVmCzK5w1StW3mjBhrLl2tFrDWDdF+5u
a3PEVC5gF+9gPMWV7ygjxGgAGwbmEi+RVj7jljChUTqhpnvddCz1iFiMh0MiXiLAB4fRMYaQVLhz
4FTbf6jUaTbUliR+Cm0YVOUTL2cWei2ICGjfogLvILQKMGpqkTVGNTgpdKJVpJfAyJz8dsGwSrag
5HsZyoc0AQ9BpHLdejVLpaiDVjMtT/0RQz8x7uk+H3Wuv6gGmkB+nJBvWB+Uk8xX46Ka8mPm5oEZ
QZK/HNbGsbMBoCvv+VTkIJs4Uu6+yteY3yqoRWkpuFx4y+8NiyFeWCUqBR9n8ZkPgiNhNh1r1HXN
sot2niLQ4U/gbDdqEukO6+hpkjfYMUSUr2iSD0R6PuCrmSIfPKnPh2L6RpNxos7G9PaZCSk5MWoB
kR/kVYkmqKZZYmlqolQckZCCK/vXbyCx0H3qxPty7bzlCZDbBcVZizBEc4tkmONEoML0mq/b5U6c
AbC5ArFfQP0ikLyhj03w7Hv0iOkrSQ/JszlDdtIkq8EMZTLmQE1d99C9KkUuyuJTSRXEhwMJxOri
LtvkAawIybH9Dk1zwX/lVSqV/i/YyKOX7FFfhD6U/V/OuS9Zn+nneE10+960wmrV3oYCCQCw5Xbr
qGorDKsXyLGB5oXiRm+e63WA+ZavpLdwsbUuV1Fc8qcZp93NOeIcPkAHuoCfwvien+PJxyiZDwum
b+m8OvdV6fhACQJsfL8AaL29QFcNwizcb9n8YNHT7HLJWjmyXddLF/ic5RSX383eCemQl09AG1hz
nsDJFAGbF6rmbFT+clDM4B90ez4tMKqmTJ5ooQwqlLHRJRlgOoQRkV5NROnul6bS9BMx/f0OPj82
7+v0X6HNhLBigxAKP62bObYXAYpqKTMywjAltDCwL+rTIW2g4K3EvaK2QhWiPqVT4Shd84GmU/u1
LBcx/nVoBrYqyvpjzEA71NXvHPkRSnj4Ez8KfVsckT0NucfkyMYJ8evLjs3j9Gew4tNPmYeL3ZkP
fbEVcBkTdRXu16s49JfKn+IW/5B/0yyyAxJl2Llw3IA/T0KTIoMIMGw6KQlpCh/6puobcM8aCnjW
xKWeDlAUuJ67HqZKil43f7H/mfCgmVAe+UlCv28I5/aOXq98MHsRigGBXUlWY/8TBUMddLpdtv7L
p/MkDBRBB0ysL9uNYOZBlxJxDtmlDGOX15lIsuaNaoSzS9qTc3cooGmouM01ya669IdSLmb93lVJ
cgVJb56eJbsdMyueuf0f4mQJ9LRgfbxgEvWdcGW1eCbN2EFn9bp96Gdy5kV8+3/TGaXu4GYkwNoA
3q9yszbtE5UuvoITk9tgME67q29vRoN0fchsV4+L2ZVyDG8+TyhI4StFPWQ7k1bypdZaFPi1nsrz
uiFrtX31iPPgZ50/uGSHzkfvlyrWCQPMYJFzMA5zXVcxaf/CAmHQi+x67YS2neII5ph8kWTi3uML
GfO4sn7MHYhdglFqeS98zlZFUmoBWAHWwAFShZZ9e7qSosDPZXPF+Tko8Qw2M5aRB2kKbKPmNkpR
uZxxIrwABb7NDgunRyJI7lHBZ7etpPHEzO1YhST6rml2lfxj5cHGhqGLStIRjHFKp4jKr9DUG6WJ
N1Xmne2fbWDuId4LBBvk8+j+6Qcbx73MbeKOntPZMD7WWmBRhuoGPhi6JrKwcLyrz/uQx0hB7kJi
InX/VevTGvygmfOJgEdVtbw1bIUwQ6NMOkw7ZdWIyHK225NmGsDqlNDqYsJ+PvJGBtyvXBAX+E7i
OBMlzaYjizy87u1whlbC7e0qfx5mEy7Rq2dQDB9Z3z7fSnNnmJFKiUUUG1rB7MwvucuYejj/hbsx
+iHv9rhfRSQK6v/TBEHwiG1uR16ewulbi7UiF1uk3A6D1dwqqQfeGDSB3f6udcr/Ae1z+ktiP0p5
WsxUb7DnqLN6QkVbHXmR0txXMHnpEUR3EtBnPqLyGJvMMP/rq2qv3LGDKb9hfvaZUrZMSWZU3UM+
cYhxiuOFtugX2c709ozffipuBTguaLOliw17Vq5nYAcf9mgZl+Ek/vNEwK+dFocP3zFTHLBz755r
qlh+hU7cAeT56Pcnuza0vmhZKJtpfFNlJDmPqOIULRa29VNvYc6yUN5D2sWhRKhshDD2H3otqe7b
QzmIPN9UDOePRv+iLKc5Oy3v4pjLM6eIR2iCWrp5be8Nk7+BghSiDaeHYOOQzWNk9UdNJylW4DZl
GyKC850XsjhIYWTKlJcHwTodZrJh4gmfRDCJQUknn6KgGwwxSdPKbq7RcoSCtgVdFHg6ChBGCVA/
HsfazuL9s+NvYcit3vUJR7IkTmdfDMJBTlfFvLoNVONH24N2WKeY+HB2OOdXjD9OWdE/MFTlkyNu
1tzvCA76c4GEobPnaZT5KT2ghvY6Ill+h2qX3LXc2VjLoWP6aBaxqNjsOkiuBTrmsb6sX0yPRVoN
bg67ZLFF6Qd7R/HderIOUO+ProBoBD2orp1fuXNIzeEl7K2aocJ9dP/Kv0P40FIqgtCVj1Z3Z6cc
+DYHzeCazqkiaNyA8aOk1RlqYy+uYRXkr9zkJHALpoBwkhh744yQ4TH8c3TE9q4V7x62cCSt89fs
cwyWJ6riSHwbwVOGq4shm0NxJTEH2tL1Mjs3/ROaTGiY/cfZbhfQaJmGrMU9xXLWYdt82zFpPl06
RLQF4vH1Hs0aBHPY1zNNoHBHQaCTW5gk5xfw0QSEoTJdWvsAOOtG4tGajE9b6VdU2vhSg60uTvJK
Yk/r7GZEqa5ZiGsBsOUXQE/cH6niThIfsXwcpTl6/uVp3iaDycZ0ySvNCvfMC09Y0aY558W8BFx2
zPRXkv2QRCVsx9gku6V5/JgeFj1+kviH1s2r0N+zttXBl1AGX1u4ah/Sl3a6zqKY8ZkRKqOfhBJ9
mTvUWnzoTR3m9uE3koKDIUsYeehIMeSv/Yr9yaeeGpnePyeqdZoo2bABHKbKcqClDTqrpMj2qx21
fQUy8q4g0XnJvU/v+NnTV4lFvY9qf0qv26xJvxybfBbP3LRQNvficOA7ZLOHx70EOdJEI2qdliEb
hW9ckVG2+LPEoAASzyEDlUO5axwVUNuRgcP8Lg62HJX/KSBOkcvQTxgSa/u+BXriYAPGL2k1tOSU
DscaQQ/L3LU6XsMIBlNFxr8coc5PvqjESzsAeiIDtwwVOa63zRgaW73NK6zYrhXnxL/ca51YB+Jj
BNBsvZgp3VQuhivPnFXhOP/kuNeFvCpNvZ1VBm+Onb3i3wXcP7DZBuBy3Sf6ZC6E0UcUOJXj8IO5
dKe/XPzTSqGxKfEZz+SJQVJBfPTQSM3Npv39GABEfTzn7j0Uc95P/z9I6gTCPS2uMU0Y9w0StC5d
jUMZnF+oXZPqYxeeMIB9X1ZtScvSPRsTy0l/hhSl8HuBvYvOVyIvSu6W2JmZGVfVrFYTFQ1ySQ+H
N+QFkL5XYi/04wFa967CcqgX6o7BxoNnJ+SL/Hyo7/nzpvkqBMjszgMWAVAYSBXETLXE/Lc/iWR2
cJaPPDMumh8ehexFEGQrM+G1KZOEdkUTz3v3kC6wMDI6AVbZKqGFwEsaI/Zy9XClJA/1Txmdw/sZ
eK16pYUv7HvUMs+6w20YNIHX0iz/dRIFefx+MIP3DLvlRGclOmftejMSgeAF2WkvoV3SIYjzMsEd
NzCbG/pILjUmdRlAlG7JSbdwam4DL9vN+1Q0DZ/M0qsrIfo1mNmctUTi18WLJ2HOgU7Xc4iWQKxS
73cj19Gwf7jHMneoD/aO2FFA5HgnEgmgnD3G/V8YIqT+iAnZ25Uy2Ht8+yaOuA13RiyaBjaN6arI
TIkvsLUFkZDN8FnCu3s2TjGB2PksMT4WeLs3s4lGvMX6FC235ZaYm2GK2OvIvONY/n0k6pFsSzTE
LdtHUDfuJBw/XyyreRxuFCRuqyKTLY3qFUzh23BYDMSz+psG+RhOpMx3tPyfK5Z8rVodzLugBWmd
xofc8Wi4hh2KQTAa9Tdxc2OgZ8hYAWyduxmn0OPU2mR6Kqizm+RB6kTvMOH3nJhgwDCeWDir0QDJ
6tj2ofVN5nyNp1PM46zZxAdjbskjzoIeViUnbB7m8hiDUZWkqIi77o4LkfjQyazCSrZTsS38+VBN
nSlU5B4PRw47e4LQ5md/qrm3s3MBXq81eXOwTxLCqi35Dt4f5iodfLhKmIUSqsN1qtnRZL5l3U54
Zsmgs9SncAnyiXfgsZ/jRJyv1PmgZlFfDd3kf9I+i8D5zCRqaF6jz3pD1LmiKKwgaoptlGo2m6mz
TwjYypCjZQ8o1ncKE+HWPewLFBquFcES7IaEIWa1W7Bw+rnXd+bhVIZIHTeTb7xO2eOtpU/qM9/+
6osDYO7Z2fFMvGyfzTBqi0xAyuYQab+t7ezZ7veYY3MHNiOJuDlbqJfcQT+VoFO1OwhFxujZvLui
k+CS7clXST8BZ7SL25GirViDSA7qDV9Ba6sJQydh9ilyjBtgU5HyddWrBHTltbILJyazNSNUh0l0
ovFpcuHtFK7CdrPFclaEgq7kYS0IPC7+salX9T6wwH+gHfBINiOn4nzQzRuP36rzao5pP6ur83oI
mPZCKyISfMgcvxTeGEK0JLUh/GgVd6dkurcUrs7T1ZqiP2HYixFucI5PRMc/aWHIYo5vMr7DW8L4
g4935IhSsiNNaU4NlY6z83+pQ5aJHajqPdYHEAX2uVaBg1WXHA3P9T0j6MYWFfg1fFxoy9L+7v14
eqaLUhbuxoCgicirp42xABXhjCgMDWy0/Hyh6aoJ+oEbWtssnY5qujkjNyI5YdvDHs8bd/QXlgi/
3STn4ts1UsQSg9HtWDTWOoq41jTFjwpIxZpQoZFpNc1gNiWv66YCCn48GR/MT0pWLw4LOu+w6SOK
H7iLp7fraUebHuA3BjeJIjmp41Dp3NKCYmhVbMyJ4qi6sIaZ+i/USBpoTsvniLU0DwIuX8Z9JpLh
UwQASU/+/gI443EaY7wY243fWWIAYQH4WKrCosl4w/Q10ZgmNstY2SsCvcKKdAUKGqrB0EwkCM/9
U0sykkxrU70885fOBvSq/9jgYqHEVTOgHiYcBzSjBW2b6Ini1tJ8C0OIu0n4SbissQzGULld4Sih
oztDgdd83U3fzyYj9h3ajt7NUQNcq31UjLTc5ERwdRCGDGQjzTPmUdZR0mQZcdCsKlCBPJhARw2x
CzGtZ+0L0AcWJ+q0YoFUN7hys86niCKAQ4klnXPAovPGIcVjgMV/ixYwrmTKjuBCqQKUI3V3UnpC
LCkBsKzz1xmXMfGipXJEKNfFdS3gloJ+tFHTTLG55uoxMx0MvyETKiG+mGCIcXdA0psAkIlCo00z
xnkPqCRF1VTmPN0vutJJxhjUSLvKoN+hCh0QVXbrR+h8SBLXcAnkmd+e6wM5hFDmJtrePfdKPh/J
q+J0LpFjgslrZUNUxRpogtRjbmfsqzw40Wiyqk/+BER8PVnmt3/EYIQVqc87Fzms82N7yeHZ0u92
FB8K7rynnYnse6du0OX7ENwYf2hpVj/Ls6yjvgk+VN5MUNcyguxRi92lfB9XJBz6Tr9lKNBfHWPZ
OacbombziN+pENhjxvN+7jSgwRBb0ebp9YI+wFu2G5XFANrSPoq6O3nf/52bJ/ZS9ozH2LMszs4X
jGns+jxEZcnOriEPyiI/JsoZ46WhUryM1R4Hf60KQHxEUyH7Jz//jwPxN24j4vspwNaAQjRVMDiv
362jdJe89dMUgRBgR0gf3NNuevidwPW4KTWvbVN1gp+he5Xa0FF3SKfv7O5zyTLO2XezjpqPXgLV
f4bimlEI4Eik73IASbi0njuyNecrgbSC3q4RiiqRP6qxRQ4vKPwVtzKoZ4qtdm9hBHVVLYMMdQiJ
WDRuLrc17fo832keJSSkCzObjUtNwjT2MLtZeqiS1dXd0pU31ASiKhSlcQw83kbwjHB9l0cw7IKZ
9+ot06DUf9fDvyfeGVNh/CeU5bv03TOaUXN/b+e/eqNKbS1VyiJITiULSLzvWD3Os9+JwZLqFY3j
xt0t+l+XN0n2MvbFDMMMU5u/CdeN+FF5GGhlDflXnTalGlp1tD0OJ2C8Z88grN3pGDnjp8MFTAUJ
LWJJcu2HFSri/aCVvlSrNYus1h+gdYoeTyAen40mfaisvzXA48ZnEvaonBcJ8mweVMgqpRhuomq9
YWckRHNzMgGwpOroHAyQADIzdkCKCu3jJonxWhJA2MKah9CU44Ra5DWrnbfRRyzXsvQv6tDPFroP
3NIoeA5uzVW+cTvZjHlnF+K6ouSWr1BCz23t/Med8UJ7DSPNuAl23aom9fHjL0afKPe6nObItO3a
HDqvegf2ocuJ4x0Lz/+XzXespNEZsIYLUt2A666RsEs33ePzCFjoLs9zlXu47hLSPHCOp/E9wzlt
GdSSkEjXs3XGYFzj3cc35+lcwh3qhOeBmqMB+ZJgurnVB169MCHfS182cElf+xLrX5PVL1n67VO9
2CNLxgOqqxrdjOUXNAzmKB11neSftSvWgukpSVn+/xTI+pFehkdQWlAEn0Ot07q50k0zQJVaqBhs
Jr3UPhykcZreuNLUkw45dEAvXg8/4E5/L7NwjhWHn3rmuU7ArVZNQywLPAtJZNtomqz/ziCMNzH3
eIOpCg8dCW0Z2zonTNKPuZHxJ6XaTf7DDbgnKi2u3PrMyKnL1TvjN8BsN8um3aenkIwzhQdAKnxV
pCGZQMUP/r6ClvsCK4KGVcfxq0+7lHGFXhzgofDFxoFYKflK1kf/zauCp046jSitPGJk+QuwAw1x
ThxZsGSVyWsb3sR6kO9FYqLxEhtkKYg67iqg6GvNbzGTAv8MM+XMMc4MkLGWoFWV90M7oBGrzXkL
enEI+rVuwLbRcRyNthHPWpoyJ9gwSOhHjAYNkrcCmuQV0WHnlRjOHMUPtFWFBOCv5MCrv/OqTcLu
2Y2rQCwUYPdxsJVsJIglNV0yvAxvzEuBv60nUJ+lWfWxRSndbQIVpnIjvWad3NRvPuHmn5CT5iK5
In4/tc27mfRJ1KtvRlAntHR3RjOD84EgV7rDYP17Q6FjhZYQ2pzXMZ7xkHxuk8YSV6B8m7z233hi
uEUwzAC3dFmBfsA6As7eJhosQqf6HgajnfWhDP2OKvMUoo3m3Bm1cWWHfCU3diloNK9xqmeGanRu
/WuWHJuFZZ6nGSLG6f7T4w8X/Fapb5zV6+BNZkWXmE4SjY+J8QN7uS8/MQmSMaPbptGb8JQZGdPM
dL824vEAo1IYdEnQZtVAjPQ4ndAq3ysKT6jEA9H7eNmez/B6ml3jNm6PH5rSfugCUJgsKAaVvBYP
dDogV+VxX4tNhopVRVds9UY6rtwxYDXux3fdLBIpSeJMcNlTZmgoLbEngi4avCL5giFmcKwNw0jV
m4Wr83TpyRdrT6uVExigZQi2Cmr0sOwl6INZZAMrPGOB12nTyvv7oZTeXabpf1UmfamXjBUGu9PZ
OH1/PrAvNKF1T2YycJ5vrAXdSjOksXp71zCXZUjmHZxbHDkbQCPcmah8804EiCdSmV+50n6bvGlO
0nQTTdSODQJt5dxrDsv0RQDxHwvdH+Umwl4ovRw5Adk5LD+vR/XmjlVlei1msdymSDKKHblMXnze
/KHu1Zn4SRIi+1bCUD+3s7oTFsZhW0rebWfxhuOURHQokkuJ/Kug359ya4kTpejT8TpiXVC0x3ZR
8XBMCekz1cVLuvfCfVQV2/MAxoX2ALW0mQdQqdjQR37CS34hZy8ooTym8CGfkcEY0ffyXstgcl0I
IvOTFrnJ5AR8V/6M1YGThsUIh4csHlXey4izh7F2H19yryfaT4TDcBFn+KTa9yE7rXjHDTuiKGC2
HFKU4iRhSlKGFchxHLCp8e10a7OuJ4a3E+B919vvb1btwrrWfYiqKBPFwaRKS6gbK+0+CaH0U0Tp
nXnpxCshQpcQ3eF7o/JvwA9/HE2IF8h8M8R5sH+5dR50m/yzEhycma5uQ1c8mi5uKXAH5d9awix9
CQkZ5bpnCI6+rLZ8fvqYJSrAv1LAv+8ESkSX92VT4lNuYMIOFX2dwZFZ35upYmOotoWiU6fRpGt6
pQkleRjydgHUrMKrRJd+AycNqVxC80M4JuQoxb9ROE0p220TzAZtg74Fw2lrIny7D6nSJNdiFmwB
1gM3Lq/KC/VQpw2P1CcHk/Zy8savs3q22kB29cKZTG+Oel7LHdxBFD9piKGRKlXRlYf7DB9vsa23
nPAIQJ157dq/BAe+afPBywvLHIhxJBlErCHQk73Msy+KACt+8J0l1pSXez1PeliHjxMvKsaeoN9k
SG1/pBJ3c+OzGeFfT8ZlSjB5dhcaMx8fBQ66999/05IkJvz/2MFcG65DdsAR/5rFLtNhLFKQL67W
L9+uJhhmgG5/erI3WiUXYKCzBIwOGqdLTxkdKmrz7JVMDXHRvTmPn/LClXHVrzYTVjkRo85E2QUQ
6ZoksecRgOydkmEfqkCSS/ufyC82rwUsZ2n5EzsIupnnhfEmiQ5sVo8ql6e4uoTT35qWInd77ayx
+PXKBEfh32Qi8B+ALVCKGxmD+Pz4Cc/g908ClLltm/cdvKWqOavMRKzHuP63iCU0X7Kv2sv4avkm
DK707fCmSer54sIgyKZwJ7evhVBudYwe9S4vToVkz3rs0giwCGxw+R8fLEX63zYd0sKi9vMDHNfF
8QgsKhxY2EqzsPzZMLC1Lre1iQvdUPsTqUXvYEadT7CfZJhJXSuMB78eopk+ae4XIuoRvn4pn0if
OncD2EyJlLHFFQmV70YmF3l6V8ALk2iq7z7ZYO5aZhQSlIxn+VyCGrvINQVnczN1j7k6HoAckXb6
JSdfLHGQmgZYksFq2D06CjyPVSKSTGNK9EKnpb9UdXQN442jUtFoLgaY006T++Z6JCIppYMLVkb5
B+vRWN/bc3X4s7k4QxUB2TmFOZpykfx8iAd2250DDb29UnPoPGMRsbHouRNpBvYmg05RaGSvYq4U
+bIosVEKcd9Q2J4taPJlz8Im/mgL617832EhtY3cmUu+9drCrFgSCtIdl+/4eghqSi630LL5winh
3d3PTBJOAz/jYSrUwSeZ4ynyY777kTr2gOcQDKw9Y3tJHkyS1r1eLEqFtmWsDswwIskGYbJyo9PK
1jh7Ceb08O2PN+UWfRBipe2SAqw3dHQHk+mLdLwjAhMSOwOcV+fZmjO7Vd7tqSMefIHIXoS5mh8y
stZ9ez5wNUk/jGkabPVzLtp9DbvAZqP0gL/IYKbjaZa2pHzpeEx+WNsCva5PV3zhWevYeGssqwYi
Nl2Y98jd0pZ0cRbXlknGrg/9/RkPfmlyVOir/YC+uLhSNGwsHrxdCe827E/xlGtxseFksU7AuC+C
FBAVOLjcJfN/KMT9k+sTXH9YEhMfWV9mdgNnENB7UA+XRpUcN2zJxX69kYOHNRuHIzKZW2rTa1jL
K96opramASlBq/Jp3NCyLYyV5HKcCCoum7ipSt4qc5tacu9iWSvttKz7yIhauXNyjUDyHdNlzzeV
N0LdDu3mOOIWY0Lydj6ZgFqHi/boZOJfS1qReEasHZReQ3wIxylb2eMXEuSCeIyskqfgntwml4U4
JWAieXQnImbrXPXAN8W7jcHXL1NIY60P5E0tcitVDckAD3xTO9fSam3sxAyWeR2EQG3myXhiz1j2
G3cHKgxaZYmM4lrwxx9yj2zAeU33UtTeTKjO0yAzfrNdiiJx5mwCg+JSH69krtXQe20Bqr9mSOla
aZ7DRcBhLUbD5ubCsXJEqfUCOGO9AkxtrA/eqYXMjAG3xeuuSk1B6HpVq8cut2R/FvJuCbyddTFy
FM9nEHNKn0brrPdsPyRIMaGZdzra9O4+lc3uUWfgoruC8nl9rni6qU2C78MwNHHnNIc8kQI8+JQ4
JAaxF0e3EyjM5loVktZWBRVtQzyJpld9bqyCVMckrAlHmGApv3fOCZ4vtD0KMhE9JiXHFZn6sMG1
7zeXXv7f8NkbdigXh8T27GI/t/jKhY7cQd2K/4z6Ns+3wHJaRBiva7Rt8Iluxtbv6TdvpQXMHBpM
M6HyufuR6Gtj/lRY94IBuSvbR/fUxpAZNA8bgkW57aLRY/uXShNu8c2tAgzJZitITEJrMI8aRTU6
wTlpS/htuRpQGljbkL3GBjVEUga4b0FXMFcPnG5QAoHNpAI+s0/4j02N6HkEiJ4k/kY3wlXQiefV
o2o9tEdTll1TCOH5XRYyAw6qJdAbST30DpHZlzSV9NS/xjB0GaNH3QeblpXeFjBdqWMsT/rSehFz
uHhgP9TMpDBTx2Ne2cKO3piOJ1AIjWYvw+2q35UJjpPEC/l0j0KfAyPV6NJQlthfjiOTHwQ+zBQY
lqF+id3iQFwMPnnVGI0X7dtEf/NKdq0QYtXG39rxUH9GNkcibzKOgUHSZ/T1Hen37aIgadXg3DHT
hKkscOnTgZurD5m+ax6UnODW4GFfmzzVEmIVClrMNKJpbfWyrYXpXn/qgSEb9fzceazAcAf75AkP
1nZUDIrt8AttZBoeIid0CoUIVc8YQPYvScrOeLwXRLIxr6xhZsnk5MVU2J2/G2kKkBcDRq4KSnPS
Crr2ZaJkHiDBdCfyxQ4PicEOuCQwGn8xyNW2IWy2epH5sA1AQtJ1I9cMX5hOF1cm+BU7k5FOc8eY
1s9e4MoIwEMGysrCJrM3FapjMqvk89Um1WBS8QGpp53X1m4y8evNgf2ZNLjTqCfpLuFM9W4rLpgB
GdHcNBej8qhjUqey2Z4MbSNgiJK0Y8HNJzCgMn0+G7JvdE9jb+kzaDicZuLWJKJVIvJxU4cE4xE3
gudI/pE+5Q3a+tlZ0kbDeraC6vbkCyh8uT+yFyKptfMLyHRwxprLi7tyDzgI0v6basFdqWtao2b6
Vhy5A8FVrO2slGI60LcSwCzIiRNeJtUFEH1REaFcpAvkuXeIlAoS/WOa8J07Ad9kK3Ywsb7rbt2M
JhfVCoPbzCSQMBPbp5DH336axHGu7+Luu6YzakOUTsL2gaJCzXLV23nVVkCcD+KnSmzcoy6wInne
DZ3xFBYgKN7tIu/QMcuf6c+jqgF8nqcKSsllVyGpoe8xU2mRMCMZz3J/LqyHQeT6gvSZta+civ6j
84nUvyZTX5Q7uaU1FtuRzQ0FAp6e3PmI0NQifMTIx183NfIvfn7ukNPcf8kpmECdFlKFhefYrSyT
DW6uqq2s5zxwDKEm5HeQVUM6ADeLNdsTeR9O1bse4vRS41cCuDabl7ePuT2KT+eHzxcl++4dWfzI
zyLayfGuOQzEtqLda4d2eVb/+khEexilRcfeNOsD9n5A8U/ALWTrxdZD5hKZEO21yyv9frBcO/9D
fE+uvCchNEuvz7kGULSNe/JO6lCZFFlYsOu/C+WtMbuFXc2RXsWT0XZ8tFn9XHfIDnVkLiMmCi+T
lbMDOakjHwcgoVPUSY3EsaQezZycWHb+X7y1WLQrqfO6NGMvrzvYjEY7GDSt1jR/Shv3dil53n9i
tzoPtwvD6Nase6EnWyiPk7SVMDDr2pe1PwGp6JX0ca19AaU9hoayXKyOyfqYm4fBjl9whV9DeFlv
qNSIU5ARIby+GjZqCIBeSsfTxRYu8dyMiXluBqyxk7LVmIYamE4buJ+Ehw6y9VhASWacjg92v+jl
MlF6Yadq8DkvyVP320PdkJOmUi3RXv1OHpevXsPioetCAUgfPw3NO0Li72/nNiMc52tMt0YpGdme
UgI10ynrrvzZzCPUMDXLYqH9CUERPvNh5I68rl47QWPtoXF9CRMhebLAzcPt8DTcvvTIWRreGXwN
kT7TGnTDGrsdNLHrFqoGd5f2jE6Ypl97HcF9OiJEu7GnuGmFFTuYTbDupD3pUTufmyA8MGo6O4bV
xzVt/M2KRRBTkIdUO4I92c9cM/0mjAReVDHTftmod/FTWaVV8xkV6KIsp3TOqeh5ny2dvrRFirU/
xIuarbMh0Z5vdetLp/jrfRlXRUx3EyGf2BJX6e9442TaR5OXOW6tp61QySppRKzhUcYguIQS5kiL
uQ+D6vkM3g5tu1vaiBmUGnSSuxwLYpf4mohwPSEyAKn85GfRtP48fYumNqDt+8/Hw1dU7E0deUK6
Kuaf7KCZey3Pmy9B76P8ysyITTPo+B4tHQ+52zHO1MWehGt8IUo75ltSKVrC9bofxlXgTHUyUAX8
wk6B4Atll0USMMmyZHREAk11841YzlQpbr3HXKSitEE3o6oW6Atj09Bfu0tUIbh3zuHwUOhEll/h
BKjald6DP10NV6kozcE6f6Jq0WpjIswoZ+h9EkDwOqCBHK3eg8wW/zAyRyM5EaVS4a38mm1We6UA
PBbeK1bgGyZHtdXJk/p7gQ8SmGOmbbIMgC4eFSlGp8cfPDaUDCGGJcNv9bR+wblCflRfX6PyH+yr
nCVm0cSMa5EsR67tWrDdl6QSA0iwHbY1JxgH8Rzot0vv/BZ15sY7yBj2OwZCjKEK9CWxdQ+oFLh8
T1pZzqyMJ9b5FDPtJLIC6Assooth8DrjbD9H771BZybuKZislNTiWXc3b6JjU02gdqc+h6Mhm4bM
kiuS/zDoi4nTQv7yrxRJx0PeGMu+uhXzqDCXK8Me9qiQQzNVG6sLuHNptJMZvvc2Ogt7vJFBfbgb
I3jPsyO0mBrWJwnYOXVTQwjFQmicAy7Y76QNkHzsNfTv+OMQEG1HzQgD69Oh6G0gfBlqM2acMfiN
xktUXz9JOsV9/3SvOrPfF2O9BBQoQaaoMMdHgdLacbG6os5wWQm3zc8z/m/DUDQ6IOzv/dHD7QHN
oqwDXj/9SqaGkXHF2ayH5jNEQhWOK9m80YJSxakauhHhVj6QIkhwxqO05a0AsysptgOGOgV5nv84
b8eiaDA7YzCd1OC0WgBk+osqlf2kKenyX5gYMAk1YucZWecT9oB0zqfPLOvHOl1X48Z39HSSKbUG
tXmU6wlZnSFHYlUvM5nJhXPGPq3oGzwDEtcXrfhhGmGzZdBZG0M3P+0gp00pK7pq64Vvnf9M7a52
wsa84ed0d/3WI0cxLq08hTrlALZ1CnHPUCcnwnZiMIYrrabIEA8j0MwC9sh7/2sblV6F2aEH055R
8SQKkW65TAUjGQJ+kW8LfdUK7gHgMNMss5+9MMDv0+l7hLYZZjbKTKxhHErAzGNps8fpNwOQR7u0
lg2EtuCfdG4wgdFzGFjlL8KP1ijZotjZvePxmbSSoHhXomSOiiI4kHFUB3Z+q4uKhNuRiSG3pB5L
zNf9RSvKDGPUadkYHwgUe9CJI8pJ3sb/CBSAomxzz5ag8hF6jfTxYLUP0D3WYHQadFQBMMyMs7V6
dZejIL4pBBHub1n8TPyrYubPJYPrUhB6GDWdn8Hq8j2sIQDO2nNIexaI/yWCMYuZTFIcy+fFXtc2
yE5ZHcJfSoY6YiIsY4AisU9j5JN6H0OB+WVqqd0DWYRjI6goh9Wuh1uSrIlprkLwXKG+gveqJZIv
bcblNC7MzgauIIGTAhbWYVgo1vBhUQIoANe33krbpZMwWm/kaMOZXF58Xr3R3hu3OWPFHs7bq1DO
WktF3DgqvDH4Gl5YbwU4nshnJ2afQmXFuLw37SmI0fkpBZ+7wCIpkX+Zj1maVwKjO/lLPAx/gvDB
yS8t384OZAZ2FmZkP/7mFdhv6PfsGE3pSrwc/ET/lW2/gNmtX/ljcpNpDTAX+6ukItGldBS6K2sq
SmUupyciwy1iXcJV4LQtZktAFwLeinRgbWjCHgqt1S8YAB6z6elugDDqrHcns08UMAOyfS5VkeiN
LTXi4kicWGS6IbADBde9E0uD2W2dQ6gdiR3WrZvHx+e5NRa0r3+Ys2wI8php+Hl1GY3KcgR3G+BA
hQRKek52bvQrmzrMWqAVi8DxuPXXFKKH7Oiuixr2y1xWHkekxLkCdkeR6SjK8RqFY4qrr1yRxwmk
EU0/I5ZLT09Axcf2Noes0n6J41s5TFH4Zo29PFJCr3ahw1ai5RzC3Ig4ByrXEzs5n5c2zShJ33ta
Qs6oA9Ad/L5wPIKXxL/3UXwO1tR1JfMx3ROUfPGSV3rvEzBXfFB5BdpyqtdFn+aL088EdrH1exgp
Fp8cdRCoQokY/paqe9WC5HNlGFZBayNTYaknNSz6pyKFOiqe1PB8DmDeC1c6w7BYw5SAuWCNBDeD
lc7xrQ+24xjUJlEai99BEbU2tVw0N+pBv6vtXZMfNC2nXpMfmWTaGgRrdgk8P94igO37ORto+xEu
qAuRXnQehNWmG6VeJvWFkQWrgbLZSn2pHVpbrQdA53hgUefrBjrqjJGNlBNBKZhiKvnZ5AszSwpi
L5RolGtqe6jQs2Y6FZSdJTXR78SMycIChxTiS7o/6o6Op4CKs1H++yu4nfraBt/uRy5F0x4Hr9lb
dBesqNy2j4s7Iotv2xZGa6tkSLGV3IrCOhCQgb2NLHnoxKNKbOA99DGLtxY0+WL+tnIRyjZlD4W5
GuGvK8/wSe1Dhg0NXnnUiKVYDk9JrzoViRsMPC3SK4+QTAGyEdTwqqeSkriJwIjoEYAWNZsIYqGo
Z1sY9itzVwnXI9Oby05AV6cyUdrDbHZ+oty06Rt3EOXvH8SuvP1z6kfMNqzkWVq5J6eqnMWpmOA0
aLktIZUFXNtfgwSTi4bhYtqWvOxel6UwJJ9ztKy2uDm+eLEvDMtOWpuYNPGlW2KDfQxRLBeIbhtS
+ahIiobbDWlryJA6mL2v7thgJLZbq2qKmMMwIMs1HAHOcx2KNPDtvXFCHbop/22/heSP0fYwE5Nj
oyTSARTiTQSdW56FPKILLDGSW4gv8ZPy96qCuuEBNOyVz0636nlKrQ4jSbLIkdmzs/AXI3nDpKcq
1xKCKq0NLqZwzUsq7aVgj4hq67YFTabg/xh4o3wScSq1rn+31xiPlAURnWUbnagq+w2VZhpRVm8s
+OB6vXje3BwHAqGK2KHO7LPWqsYPPiQrtDhKT9tgoM5pHhPUG8sNL2VgvaWCx3Q2JnnU6CQ+eFz4
RkRYa/9DxyaQyKUl3A3ae/pKuMIYzz8r1JimayE/OVcjQUigmDeKI6J1y/2njtH/UAzdZsRXU184
6iO2Naz3xT21oDdopDLrNr84pCUTId4jwQ0qEhX0tiwC3kKm4VohmNK6xKuuJwQDvsBf9jwlIP90
7p2jfyJin23S0EEORUUVcm+TTUCJJPon71YJesRFHuiF+X94YPb09AZtjAfaHHqViEgtDO6v17DR
+vqBzPEdn970YBKRS7Y1MX9M6CjECBQ+528dI7xUZU20Tamv4D/6YdJyACdY4ld3ZoVyFiDNn5Hq
pibL/nBTf/y4vrFlQcSA3pxVKFg6fe5LhgJIGSo8pRyaCB5wD72UqdOn3USk4PCJyf6Rh4uQo/uo
QtAyNzM0PleN3hp6vFWaMAhw5NhxDkTwAL6w0r0OaHBbUutZ5JGJmQMs86o7/gQjHWmTeUT18X6d
Ayshxse2Eiu3F+kV5i3tupI4ssGqU1NPu2LxbvQp9tuWg080YQjJsjeFv/0wF/sT78TXUZLXBlat
2/XhLiP87O9RQc4+Iwv346n4VHby+37IfvWTCeK2GxC79C6pDBDkUVWj6hQkRtpMOsylOmtE9k0V
LgQ75LJ1bTFn5Xh8vTz6Ng2MmD8XNzz9GMFyaXGQpDyadDQ3FerbFvQf2Ygo2RBEnl515E7+Ok6N
prIUtVT8FhGL5Tp3QxyCIJNZuib1a0LEjUb3ksVBa0Px94xKrSAC29SoeHvy6QGkjMFB5XX8TkC4
+J+1LFmsBDyViRMMPZaAyq7evzwAXnozJmEiX35MGj45HraZkDo1RlwWWt5/0DGaT/B4WZy9MHhb
4p/vkYGyu8akB81zkDfWIujb1mfynY1yiUHGlVWv8SvibVGrLAWNrJ/W7QQC1ZzBQ/M/CrjqXXno
DkjFU/zZwAz0GOFCMNkzTiAcpXJsxPlNN9elVxdyet3waYd0L3+3fufkyaVKtqPDxvEf2+nR4mYL
Fqt4kQ46n/VtF7vQD9DBj/u//vXSO7gGxVX2EoBH/7KLAXrvtsT5NyBYlt5xoi80wVyTxBevQRNi
bK2TzlBQCcNdJc4Dhp6a/KaSMEVJxyI+/LJ+078d+TMkjzSVJeQb0BT8Nge0duICj+ot/aFTK7VT
XQSOAtCnMweKxh0ssacCCmn5Y4WR6J4gsA2HCXqml/QiYQju4nkPyquI0RKXMaoEvostW7qNNUqD
5A352l5ZFOHOsv1HSd4Qg5nf3gc4+NwahEpJOVObx4WokluVMglX43+4d05oF2xNcn1RyRU7Dpxr
P+rUoUM2q0sQgGWMseaKHLtOSFYcX5PnLcnCoZKLj5xpXk0aXJrLGtVMRoh2tsqGoJUxidkRP7Hh
aYV+U3xdbjD06QAuPDimOxw7qImcJaJvf6ssvEBKlKFpeb4rm7H3VdpN1NW4LggBX3Vkgqub23q+
eAP85FtDUXiu2Xfo+dfnaxNNl5B4E4f8yWKT/aBt2qh31r4OzUJNJFFEc1cQ47AyiEn2aIyeZSwl
AKPI2BS2pWOwZLt72dC8QB0jOAg2vevqJkUKsxn9uTdy93zhsaYFJc8PbVrK1ssn/ggU6pg/d63n
84HPh4epBfe5gS+btFToNQLFas6yZf8h8BXYOeCez62/E8I6vJKky+9hdF6Ly9LiYnH6WO0EM2e7
NmwZAfeXwskYS2X6vZcrSyWCcD5OMSJLfK31umwjE6gpaiKL87mQfRS3qeqlV+TSPhdsdcE4Uzms
Dsd+ZUe+VVzVAoYkd1fJ4LE2XMdSMcughPHk48Wc7Otmzx/q0EOOybjl1RvULiHKhGjO3zWSvYKm
fXslkpz+fPgMqhGXmYUx3HxqVzdxN/EX0ChofrPg9YsGDtSxVp4P5NwiilsnrlJZlLymT7ZCiiIW
duVqOQA05AZu3t2vnTGddmdw6UEY+zPjrRfEwggmZA7UPFbb4z24sW4YTLsvYFykJem6VvhmV9BR
MOwz6Oz06VOI0WiLIqQFExRwbeUc3mOHg2CAbHa/qtVBODrHjXOcMhRXHeZlutuGMblGGNv+6cDP
/J/NjlTMTfqedTg8tVYVsPpGa5O3f3WnqFUAtBz8Tr4M/lQKCTSBKkiRN1rkrWa1QaMdVZR/oSac
6/GYqbN6wc9Bzfq9iINOazLBV94qFbdOwJJle9oVKv5mcdITDTUDckk2VxsC0nWDsJmsG6iAFNQF
NooLO/LCnYHeZdSJwc2qoLqA74SQcv7XSM3q2O+dxPUhuuIH7OWFC6OLiQ1NpkA/a8xlUQ0c+FUx
JFaFbXAlmWv1GlFcrr2vj0/WXNwWFRKy4V89IBnIxSpcv3f3G+Kf+9XfH3tTprfQvI6tFosjM5ui
Y8buj1hfQUP5JNICbW1tQdSq5LF08jX79Qg4R69gprWAQasJ7AeqDqovPlGCRL9BM0HIr7oNl0Ao
i4quUlh6HESC0nb0KHT8Mhf3IxIvrAX4JP55BKGYoxKJ8i4p4nQqZoyzlsXSFmQUBO3hU35axr23
82m65Rcpr2LmPViHeV6p1aTZQ+m89dQvJeWSr25q4w9aIsXFhJDGcwu4zCZiC9nuxxm4FBcA0M4z
TYgMd9NHTu0azHWVe+c94+C5IA3MCpnIkBsrl/B0tIRR63Gnj5mSX7stmuZZGVMthGjMwMjcRAZE
d+ZCFRNQx7MPR6Gs7L7iUs88d/W4r0YRzcDfWNC185AJnp8Mr2EsT3BOtS/RlwonRud5GIjNGNU1
xEah3hqR4N+ojCOuiJ1FvGUuv0xE19N/AOd8uQptDKr33bcJ4wzAxGzBjNc1vipd2pOkwfs1qSaY
4wZ2uc0ho/Y9Twio/x6UhNpsWy3N7GUMe5a+M/+NVLhaSSonRQqlng9lM+OLyaRNzQgH529SDoAW
6m1eyLIGZ+DbLhFfady8qMOGEcQuwEP0i1VEmstROEiBvJ7jPYjt9MAjOs/ucexVhro1cwWqjTHi
MHEOt1RFLUV5LpmrBQVhn8zDTOriFSvYu1u5K5MIXtYF8nbGDGt4rTWqbKOSPMvVCSv4siuaXLah
HTJ44dmXb62+eaCX8uA1p/PT1YloXg878ohiVFSRzUo1QtGdidFiAO4Z5HEFQ6xJYoTHK8482NqM
cPvYSg+EBC8bheULxJZZ8eF2TPT1K/gkhzsOMbNnGxrWX7vWdB1xmfZhhx8FskD4cDyrPCqyCQtY
LGbZxK6zHok4dGcFjDnDKtFudyL3OrCn9MOeVS/LQJCp9L+patQkPmbTbDCpXAKBM4dOcgAI2BUO
ig8Ss+D9GUNffglroKMKKksZoREotiZjKFHlNuLknZLfT04hom7JYMiy6P8ixAM+gYZqq7lu7mBa
hechVeWVgGwKj4M0X1JMx18yoBTPZesOK+GAP7XXizkgo97o+VRU8I4sw8ioRMNeaiYshZsG6L+v
2957q8c3T49KhKsSKnWbaExD3XdMi84kABP3KiXibv3VBiRdsXPS3fnyCMMXzIOeD1+LQbF00sei
EEp0KEZ2aA8Cp6jBaWkWJ14HOcTeS/3g4KNJOxSDaEt0nRQsKyTkqNNmIOZcJgcR5KmFtKOvj4AA
mkRcnh/bmrKVGHi539fmyT85sF/mTY2CWw6RaT/Q05AomtX7HywQwF4tyiVfDPHV3wFi8qcHxxgU
D6gbm1W6QIqnKTCMXWirddRvlp9in7PpvDWvQyCmYWCE1trQgau2QGCYiJk1BljmxgaiVJ3qcKed
lAcaf+bj+yDUHEsBjPbXkdd2E0PYu2pS8ZOhsoBOksg8iLXLOHxc43fx5QfTSe3GxZrxn1NZNP/6
yUtRviIFv+QLyksm6lXwzfhLlNsZ2hLP0jvff81MRTFcroYgfldjK4cxqosq6RRT9ck92CBc01N2
vyhplCm0LZE4xanb0CHSIZmkt1U5zAoC9+FDL27nB8LsAHy01fB7YMjwmt7uepEP9LzYns51kWPN
DM3J7YdSnWydhuHbJ2zOxqUPgDx39MPrAYCgdoBdnDpRf6pAUmf2MVRV1BqNtVKZvFHk37X+WNZA
+MQruBdZKzZfOwglf4gUiziwuKNk5c9anDWkmAxl5q4CXgsdJM1g7qFniy0yC5gz8WyLA9MUt2C6
vZEXD2SGk9J+qezfC/kagfUkOzPPrnt1eYu1semvhrOBOhDM0p/lLD02KRqqJYgMaVBs/p8mG6Xw
tdU4rerNo4+X9EWh/flyJtk5oxK1MvfH7K4/A83GpjyCv9zGbaovEo1mTE63gV3c8yGHLLONQ1ET
REc9EUxviD6dF+YwD4MuYQ9r/Cy5dW16X0hgEk+O+4B5mqbjocFLcDFQ7r9KRreAATLN1QVVtInk
5kIMV8twQYF9IDdWj1AOIuvsM8cXTtLE8VnWu0rtgrXscdMlfJeuT/t+T+QKqr/0fbLBgxTRL08j
E2XBRSzdxEOqkOTph3u77bk88qe+n7UP8FNIqLLjyzmwIpuNdtbZm8XTmLx2F+tOT1h/P3+8s5Cw
uT/IWMRploQ+ixqf8NQAL+98gL/gv9j8MteeWte9TdklvRn3h60osPpnNBJT2scLHLk6zUflXeAd
YsL011oIazCYZGzboFI45blP0gwFe+aEVeFoNfmJktogf9ccagodVV0wW9TlqllT++LZuAl6ZmSM
2s5EW8rl25BbdfTtX+g8nqAofXpKNvKiJ7kcqa3udCg4Lzj1SR6mR4gFHY8XIh0vFnKMCuLiIuia
ZgZytuf5H4nIVPv7NwAUnHy72SZ3Fwax1RXn159e6ehFYz5F+qKvrsDY6bFTQktIa058KCr6dzGG
SwUfJ+yIs80X6k80B+Md/95z6siPFxH4U3cUrzF6045GVMjicdXfYDl/iYMbfQrsdWxc/DZ0oTMK
4K5DYTccrUqjs9UHlV3OLZEMqCHf920vGAXUtrJuBqNyUiUYAVo8yzeqEvwDiUQpgMhGJQBtJg6+
aXAR1pJ7nSJ3qPa6toSceGfPl1YQIoGhtXYPTajmPoGE8KszVw7UI/EMW0z2bqTfYnwk9DinWBK4
d4hW4Zoafm3vMMuE/mhVjjQ9g3DexMqpuF438LyG121Z/+Jj+CEOlrceROATkuo9O9MqfN0QAlx8
67Uf6SxipfOMFxmpsC0fL4r7az16pWajxBMU0/AmXvT5wMPKz8P5IjBK63S0LAFAjBT8epreYpAH
IwbM7U/ZPWSCxpcbid3yRmFRWoQ05sT4fxlXIaUKmpMBIk0kE8WB8Fkf7nsoyVbMnIWI/GousPBT
OQLKXIcdIK9HsVb1jQkWKKbmG2QOgkWSy+vIegWmQbEeoof7WO4UBE3MDaOr31aA1uwTjqNHieiL
tTdiQPB2oTlIb3aEc4Fd2kJYgqFuKnF5qcETHsbPOhb9JsPsUyfJxCgTUqnGdybW++1FOiAmj3ks
0QOXYVg9ls41/OTeyJVj/PsX2j0Xd02I2//D8k0UpzSWeg9NvRDkAaOhYQB3OS4sQwLiVFA8GR4A
fz9x37UYSxcPbc/tKB5gq9i6AEjIN9CLi8JY007lT6RkMSAWdUpwzh6S/JR1knBK/CZl4CyKxN2a
xv7QeYHUBM1zIDN2sgW2lIisZ6RXDkEktXJJ0gaw/b3ias++HMBongGCGu16h0CrphVoi7JV5d3J
N6oo5s9edXauzVObiFL7e6BDPub9v6Z/DLzL2+4bSdMoV49uFq+oubvAm/AmP+kS+b638OXsNBKd
dHrldKfNF1VMDTiqoduQEWZJQke2r9LWT71/kXOzoH7X7Zc7JG1/hNds1fPxTHvKkpJvF8dfi44c
+jydRzve69ik/kmFWPhMs7EW/qH/J7MELgsZZ9YRkSn0fDasDO7FXfL7mlZpcSeOWXnbD5DSj6GO
bkzejGGKh7z8LmmDbTwKxxS77UXqMNswF5CJSiysp642G5KKR+QgUVDSO+gUUuZZmLy9lHheOqBe
/EwICtgZqa1aYau87askOoedbIEvNO56lpBDCIQ0HcEDikK0PmfxXqPNBDhtQ9c3e+gwfy4FiksH
7GXGf/ap0Z1pM25c1eJsFeA6KC8dgRjwJXDMU81a36ilhOgGrVj6yL6LHPtGTJXj0YrW9PP0kAWJ
SsPBr28RvzNiaTM9AwOVJu3G7dMDwOVgc8jsB1FSgeeVFYkIa3IEu8ZJqech43oEZiJ8my6eKvjo
DxP7hKUgt0BzvUJmlNfSXMyHgNw/g7PIiD+xaUPpnZpIyX36XRtuSec8Rpi28LQEbWjWOsa+yapR
a8fBOdO3cRDCOz63c0F5hI+kv2XMESoNcvIXykaqbe1DfHA2ebZN3BLoyGnZbGxnaXrRAgAgSWKV
LUZwNhBa78FQ3hIj1JjXk4pfzVJN0Hx2zSxKnxYE5IHK0FoKn37v8JF4GUKYvBtF0PEpUUNv/dnL
Bj/8yZR6zuPQWWFeK/3O5KoX6cKIDq5hJQaWN+CV3DuqSWJ7U8T3jyQjIqxxKLqVkbG4rirmfwcS
OzRMoSHi9+sMI0ISKUL7CnVxXEZ7MsLZHW9PU1UP6JEpCUuyIwzoSwCjQuE4ocWRqx2C4cwEyhqA
BsS3OOQBLjFmXaXEQq3+9D51WljbOaqfBobD6X0KrQC/u6MiUJFsNWI2Q9fUCZzMyhuSRKb3a0pz
bBQoQZRPjaeykhLVV3YmtoJOOwyvgsx5v/CmgrrVkZt8Re+BIswLFC1xRQVs/a68DQLk6SCYB9ut
7xUt5s1VDBYlvS8Zs83rJuWaek6n3KMKIEmbLfNcbnfnbiPXc28V9ZpQuzYmIm6XUwwlKoFY+RWU
LAjhVWCZiESqTjYaGluQyHq4WOOCgV+lHd4YS7wpTh8MNLdQkOe/5O6kHa1Xt5q5+P8XDlj0CS/Y
KzgFDZpoxxiXQI12yf+AY/A/RGbKVZkiGAkDXdb7cb0AktqULaEqNnAOQZeqtK2nh/wwTv4l0zIu
pxmtqWaXom9AO9qc3YFbslnE9FcKRIYz8QTyFdefey6rERywYn5JjRfYxZ6U2P13pMSbDxUKJtr5
KddibEXDpIP7m6XtwHN+hb95ucNnFpu1nGQsK5yMPbjXtAOvAiZoGUIQAm37dk4pw1FDg3aTUm10
ySTPgBrT7UiqbusA6ejJkZ5iD59yUi7R9s9cJSlRNnUEAhoTa7Ts3f0UdH776reBr2Jhn49f5fqH
OPm/yWc45YCba/CxSN5MxP7TQFaHI1u1EU07Ebe7KaA3Dfb8y5i1BZEwvhH5PWAj9ObzrxWqwbt5
+7yKQHNpx1vQNo6kg4aJiXYNPG6WIh20AMsMfs1tjW/ok17kMsPJ29beEcPmtxBIz8WsHwz5xFn4
JUcFA+Gmu9LSmLUYxlTocr5SJ+SBthOnOptmVsB4ELej3bgTi+JmIuM8HT/4/SmZIbe7ohOKvKyk
GRhpzrItqw311srD9edD75/wrtgIzRZNEEN/G8Na3I38W84RQ4JCETdipuC+czvN/LZjGMIG+Igy
JnrYFHF42e7osYFciDiZyaQd1vDS/lTpYsJIfTCQJalk3e81nPDAMKkXzOSIVQ3LJ14lAGKSBEHH
JTtIJ8oLVyWB76O2Q1jruNLYDHS7iU740/iihU0QQhl7YpAIcGwLFF7mZi41t0ktIh64pN6BPMYu
WFVE5nK30FOEaZBlS05rUMmzJDlpoE5r2smgJDdMa0EoH3WO6LywHBlCJRkfrc/dEgbREi6m1nbd
WGy17r1S4y1TMx0d6Xoq6KQk2l3o3hotEgvJ9hkZRHMx54pfe1PR3zoZceIuRxCxw+oj67gkR7GM
97LGs1NY7qgd+FbYVqTOLKn7/MzlyqFZnFtjSkJcMmkQgcHEt7y01qo6NuPjy8DXCcTCvm4Y87WZ
Kwoh6C9u30DVUOikQTtl52z0BmoY1F9QDMalAHfgyoE0YM7lLkK+AxqAkvKnad3xQKVaFoHDIgWe
YTuhDuIYJ75dlw9YmmjGKR1bUWvzfKcQ2BcKHironDfmh/ZnhLxWdLB5beQSstf64J1y9khaWSje
4cc8gdaJhKfkWvJ+P/Xt9WC10xCjYxqLp9MD9oXA5twoh9hgLIVOgeFWjIAquC2WSA7txaQYW3De
J8iq/wT+4n6ykCADIcT6FjCvhM4Y58fuM4Q7+3bKNdHlNqdLojnyH3jbrz2z1jtXv1zbkDTnFHhs
IguEWAvYJKvEMEgMJg2bFJy69AGfct/xNx1yclgDbnIw7AMEyYyN/SFVkC/gHRvk0CC1TLF9Igyj
x/89wdLdoI5wj/HFmPQm8fFIh1/i/cLYwhaFyrFcyPSg13KLeBm0XQV+FUDCFHywdjl3k8SKFSCr
CRpoG6WhePRmQY2X/Ah6r6QoPs7VyfY/8SAYnqvufdq6KgcumuCINrCqeqNpACeAzpy7DZjyH5gS
SZXkt4i8aylvZMDzwyTUA7AnE679+HaH+vrIabmP4/wLeAfXX3L0M8tUBVCAW6OgsYIPtO5Kjll8
WBoFAYhN61FiL9AIKr+0R1sL8L0fdcBBd3D8Tb5R1DWj4SuQF1rpf2EKt0XayqXETOtLfgdI7hVZ
cFxqYF1lQWrRCFde5k04LdfubBDb05hwZ63eXfiRO6eRsu5d+ThEIsl5x8wAlJej98D811bhPlvz
VcxqMBuL4KHi7WDNbuGq1ga6tH77ydurh/RDvwh7/UUwzVPbW6sZA4g88AevAX9/93fP7+a9jjYs
Ac5Hr3RfZ8sxe80pWZ2/YLHDIhE9IhreMDFhmMypYWJlmll9rec3Q/+pGyn+rp9H8XplSdi+eSOx
UBG47cVVitz8sJaOpZ9Tv+7TYyH2Q+0CAubsNN/qVWTQUgYC1RbEZAEtlzrIXJMYPm7WyTvB4qA2
dY5yHMaMIudaUWk5eS+1HUGo+KIYwz7pXg0n/djGR4MkZRYaTj7it8IPSyVryWEOu50KSHgHx7rO
HsdKAL0nw30o+pFL9am2e9x5aZoVFKSHV68C1nGt4c2za6ecByXzkYKig/1kQMHsMA7K3fGW9HVb
uYTx1fySJd1s2MIhbGF5LjihC4kZ7WzgoLwIg9aDgZqujkk+CcPc6ESBVKBosSAP4AdPNMA+THNH
obzo0mnJ18lFEMe1TlqeBLB+OdS0E1nr9mWFLVsDEFwgbZBkZfgWo7TMmh9ERWndtqIer4kwBfWN
wgC35zJny3XFl8V7oaji7pqAxLtb/a3mULB80IpGfdpSq/ZGAdv6RJk10LN9YyDcJVQ8XjhfpzXX
zgK37cryyauXUnaHKbPJDAwrbHm29nmNwIa7OvNFzCObtZ4t9N/BpXDcxdsK4jM8S+9EF3cFquOJ
sR0USUdUQgG2oaTPO/7c6KOvA7kCOaHhMhLhDrV3Kz9vgWYV7yUZIVO+UUhnYZ1dEhJAS+TvkMMK
hzQI+vnN+bzj6Gi7pb8VeR+tcgzDuffkCWRtCebfyGdgmdhu3bBrWs4eNnEOMl9xvWIitBZ48uPn
0/LbpcEpyCXgqHo688gESMW52Lj5LmF6alddTGC6drJb7HfGWcnfp3O4k6Z2jPkjSejse5RzHwMw
Gg5QsiihE7gJDcTcyHRRQshjYEfzDxzORoFfQEHRHBkswTgEFKvR3iVTw13EUZ+ie5PBar6mD23V
aIaplTcCi1rvrq5LvvE4LSBKz+LuF7VXSskkKH9vBCztv04dM6o/cdmLq0E56y4se5ymSHfyxpkj
YdAwzzb+3SE07XJck4Pv9EZ9gutNrVWyKN2EuFxnRfz7YmJjl/kJso9pDi+ZnRbH3TkABuYh4NW4
FBTNGHWxozI3aSgHH8EqkuzZc8IbYZUTP2yFzsj75T7oR4nj688TCn+XzodBK3g5Xa0ciIUAc8vQ
4F7OqAcO5yBx0P+LVFsqHg/KOHLEI5IMoKPNg9AgYpZO/MT01QiGtQ/N9ZAezc7ki3hIZB+N531y
wX40enc0ZveSG1VXFb9NaYvAanBYBTudgJRyVGm6dKVF2CyWXZMy19TP1PpofLI8cFQZDUjWfv0s
S51H963FqZz6T86j88TVp4TM05s5iZzvQYNYSuGa55XNkNVf1kv3sqz93l3ZsC1kMoVFIONwrcXV
k5qwzpRVtZFzBNn/Vj/vvuscXGzxfKCwW5ABVWlGMRPiQIBmyUXlqRuwVJ4bBEogXiehy1kKHsZ4
x57iXA24vPRS7sShHKZmjLLDHabQ9alrhshUdFhF916V1uU0POrgi0h0GtyNX1AB2+UBjSSJJneQ
pCo//GuK6Cq4wPDP/cfPl25XdAjmB//wc3LIKe4l+SJokw5wcl9K4fBeHtAQRHdUaS5ah1+TquKl
oGTKYYf6UmVzasaLMKOT4JgTYEfmZuKOQGWWBnSfqEv9e5UszUNctZ4HQdZ45qq8LAlJGFIQj3SV
XPCwDZ30Z4LEL6EaxhET4cfsp04NjJpRFwq+13PVrcSezXCJD7LlrYa1PCOA1XAxNEzBIDeGXzbE
xdzhJ2nHjERzdpURKt04x3H+h2+x4Mls7OUOypU6B5T4/KO50aTQR5thCscJzmxHZ1XRgnh3TDG6
GQxxwy4wvEGzgUG/UF7zeYhi2rzIbvo82AvQhHQy8x1a3ErNf5t9Y1syqMxiLuoeI5nIpn05PGue
HUwQW1fWMWKP3/j44emgRg5rZQFjbobypUL9pOtmA0s99i9A5lBqd+K1sqxd/CAnRDwwkpYOHljl
SyAMiv3Hi7bMUcrDr0fz8r2zskeqQ+THyAZAj+4ggy0jhi/0HoGSKoBCRoOG45+ffB2hbEJxru79
8UG9lwGhGZw78gt4AxiDCcO/T+EYgMhVA9DleZKTaNBm2Vl4zZvAMe88kTIDsyUR2TnKMvaBwThr
A7F5bJcburg4PJUfyYGRGWv44mUoQHaUIN979Z6QBYPFWWgwmYTfPDHCaLgGZHeejMOMjL4U5CqA
tUh0VuDgBA1Jvn0WTYl0BZi4HZI5YOB/xogtb8Qfbdw3x9A5+GFVuhZJqHJecqit1Ikyj2lz9Vt8
dyn/ixDQDz1dkit7rnlPEs2IqjgjudN4XPsAub9wXUT42cimi2l+sZvcRtOhnFzZ95xkDfEcr3JS
aodFO+vA9DbJE9+EVlhQKNrET8+T/fD9gZBgie2eG2z4zbNyKt3FuU5Yf/2LmpZwv6q9PK8dzP/C
E5Zxf+THJZucM7YMG0ujzAo++8AoHFyhX9/3NEvYEKEFamRFF/DmXwQzv6hOD4ogzbfbzyO1smy3
pQrt4Rsw/PRCUnFZzbMGESkZnnNZ2zsJcnzuEpvR3OP2nRy4/eG3jwDXQgdHBTlGM/dCZVcTClyx
+MiaggByeNl1y207vmLtuIgII/ZQwNGiYow0ApiPZ5g7bSUtOkkjDaT4OY920sbxQaqvnea117GA
+HsZXHZS4AQdrTvpnCzBOmjFlZP4DkL0q8VDmRaLzX4B2CWBZoeWNuTfk6EAUmkeCDvj4JI9o692
nZXzcNjCc+uDR9Lck7CFQ+WulFMacaYSKvbXrdjJjbAsy5SvnHP9xCFUzApp9fxwN715zeM3WN4t
y473TwDxZzVk4ps6AnHeDO6WrBfs/SSb0TLd2vJmxOhB8zoHq1OCmdSpdfvYLHzz7vtixpEwd8i7
PReEtYMLdcsEtWrYKY+4kF1psxkGcxoWub4xVIFF/NQul4yXFY+P3qeIXySBFdugV37uqPG96Ffp
GaodJ1raoh3SG4aeGvlat6LOdPGbrgpf8byxbWd8myHfhlV25BIIXCDkN/XO/8YVsFYay30N7HJd
yF+Dx9hVWV5V+v05fsxK4ezvdnGMm5zxnJAOcfchGthGDh9qCe8DYmyo8/BxwMiKanebH7JN2fSW
FnlPB8H35g6VpkduxQ3NfvoyjTuS9Ofxc3cdtWDicf8L5Wrw3hCdHxlcwbfJi84swjZskrKv7ARy
FUVVgIwv0/iSF21TbN+jJ3ODAiQnPfNC2tcOKaWS2TBGDigd0wd938ZNsXwkPJd5Zn0q/M6RLqLO
qR63ICpLmGnoHgk4Au/2BIf5hOu2oIvKFeTLLXHyz4CsC4k/u5g7pGl8b42KWW8alZ7FORiGyIYv
TUuK95PhOE6q/LMSLVWXU3bKHKTWcPuEMEVRXkv4t8loZLcw3EUbRPJuiUaZI3NLR+En+txhbzA8
bakdcm4evit1mFRc0cqDEpg4ImxwlxswPb0+sjLOiC4INZHLOhA2fVUQyaG53FfuNFIk6dnobUEx
cxZmOQvoqDfYoTv0YKGE5naqxF4X2kSjlVo3LUbOqBkq2kzFln7Tl8B4eHT/ukqx33P0Ez0wF2tz
8jcCOXeLUCOBrfHNR+a1KZdPhAjHwbdj+V3ZXAq3y2HiRb7hboltiTVyNZckL5vP3gCyvG/RxZ8U
pG39KywUmMS2330lDEOjBGn/ew8dpmn04+G1GZ/ovZS7kaHY2gSo+1R8vpTcuMFJUHGbBxoK8AiZ
wo5sHYlj+D1wJtRoNR8jWiymYe8JRd8sAvPDOVA1/sXUsP7n9J5Nwdf7HlfL6Qrv2Oiap2SAizLO
kzqYZMj1QHjp7DoM4s+vK/hnk7v139y1ebTC2bpFJVnbDQEasu/828ktqTQNAeaQwY2cCtslsUxd
GnvpJdxtq/BBfBclpF8fiJcqNbc0hU3PeNiapVYlUeTEhYpE+cAShRvqhSO7UdNO2uaORza7d+SL
HcJCDAIB3GmvGznjQZ2u3/niKtiPuH36iCxtxXs+wPxhZFgjM8AIrcw1/GYHASoeG+g/BVyLKfu7
c9LPdXYJkiubSNHX3yAn9QQwZdmLFQNUGPZRZRpoKgyIZWa0r7oBYJOFiieaqhe/tULgS7+ZwxYr
vvP2RAvQNj6f6y4wX5PszqauBFMeSIRFdCkxBnI+DzPnWxgFifSSJT7kP/z8lduO1DR6MrrADrnp
Vn/W8WOwFbZLtgJ0SQZf3SJaQo+j8yujeR/ODONGmM+GZ9w374qCUDviH51vTMp3gR58jmkPEgrL
HXAkX/UrsNCZevi8Dyr4xJEnc67Os8WCLls75MgLpUeg2qrgit8kWmOV57VOYBdDgWQ+38hlUrE0
vDkoyhHKC/Hy7EIjpEnsrc4EFGx8b5OmJte4BqAsEF6jBbJr26iPubOcVq6lWEQnzfsQihQY1lHI
iWPFoCGwFKdk+eACtODq+Skle9rZFY4EBYZ/NZv71RvF0LVe6cQeAPKiDLCYXnvE8T+abtYurgAg
isRh2RzcewL2IpaDEHY8mt7ClB3r8CZ6ioQrHL88RmkpRiYDy7ek2w/LufaaPeVSINMH2xW6OA3Z
n2TZMUyIAwWwgVt8kRaqK1ouirIjVPIzBtcIbX3/8ixlFdxi7ol3xTp9O4xSDfrExZ+RgaEuvYr3
Pk4VSXg/ENOBBpAq7oaGGyFOcM2gsFj+cUJ/WcPOFykzUu2jheJv8r8vdUiZsGFDQxk3DM/bvl7l
4xXWnCDMOkxBBM9Dk4AecAn8CW+XhrrTKljwpQ5GKS3KwoANklT6wGEcQcFGC0iCj7AAyKYjv8f9
haSIYvHufnUHSyRRB97dGrl8XpABJajwF6WcTRrmaUJArb8u0dIatBhv/APEw3MBu3rNMDZHbEKT
GnzeuhwmGwJWjQ3NK6Jt6v+3jSyEcCmThO0QL0jzaPah32kfXTIpDm37UQ==
`pragma protect end_protected
