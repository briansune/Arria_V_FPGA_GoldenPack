// low_latency_10g_1ch.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module low_latency_10g_1ch (
		output wire       alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy, // alt_xcvr_reconfig_0_reconfig_busy.reconfig_busy
		input  wire       clk_50_clk,                                      //                            clk_50.clk
		input  wire       clk_50_reset_reset_n,                            //                      clk_50_reset.reset_n
		output wire       pll_0_locked_export,                             //                      pll_0_locked.export
		input  wire       refclk_in_clk,                                   //                         refclk_in.clk
		input  wire       refclk_reset_reset_n,                            //                      refclk_reset.reset_n
		output wire [0:0] xcvr_custom_phy_0_pll_locked_export,             //      xcvr_custom_phy_0_pll_locked.export
		output wire       xcvr_custom_phy_0_rx_ready_export,               //        xcvr_custom_phy_0_rx_ready.export
		input  wire [1:0] xcvr_custom_phy_0_rx_serial_data_export,         //  xcvr_custom_phy_0_rx_serial_data.export
		output wire       xcvr_custom_phy_0_tx_ready_export,               //        xcvr_custom_phy_0_tx_ready.export
		output wire [1:0] xcvr_custom_phy_0_tx_serial_data_export          //  xcvr_custom_phy_0_tx_serial_data.export
	);

	wire          timing_adapter_sfp_a_rx_out_valid;                               // timing_adapter_SFP_A_rx:out_valid -> data_pattern_check_SFP_A:asi_valid
	wire   [39:0] timing_adapter_sfp_a_rx_out_data;                                // timing_adapter_SFP_A_rx:out_data -> data_pattern_check_SFP_A:asi_data
	wire          timing_adapter_sfp_a_rx_out_ready;                               // data_pattern_check_SFP_A:asi_ready -> timing_adapter_SFP_A_rx:out_ready
	wire          timing_adapter_sfp_b_rx_out_valid;                               // timing_adapter_SFP_B_rx:out_valid -> data_pattern_check_SFP_B:asi_valid
	wire   [39:0] timing_adapter_sfp_b_rx_out_data;                                // timing_adapter_SFP_B_rx:out_data -> data_pattern_check_SFP_B:asi_data
	wire          timing_adapter_sfp_b_rx_out_ready;                               // data_pattern_check_SFP_B:asi_ready -> timing_adapter_SFP_B_rx:out_ready
	wire   [39:0] timing_adapter_sfp_a_tx_out_data;                                // timing_adapter_SFP_A_tx:out_data -> xcvr_custom_phy_0:tx_parallel_data0
	wire   [39:0] timing_adapter_sfp_b_tx_out_data;                                // timing_adapter_SFP_B_tx:out_data -> xcvr_custom_phy_0:tx_parallel_data1
	wire          data_pattern_gen_sfp_a_pattern_out_valid;                        // data_pattern_gen_SFP_A:aso_valid -> timing_adapter_SFP_A_tx:in_valid
	wire   [39:0] data_pattern_gen_sfp_a_pattern_out_data;                         // data_pattern_gen_SFP_A:aso_data -> timing_adapter_SFP_A_tx:in_data
	wire          data_pattern_gen_sfp_a_pattern_out_ready;                        // timing_adapter_SFP_A_tx:in_ready -> data_pattern_gen_SFP_A:aso_ready
	wire          data_pattern_gen_sfp_b_pattern_out_valid;                        // data_pattern_gen_SFP_B:aso_valid -> timing_adapter_SFP_B_tx:in_valid
	wire   [39:0] data_pattern_gen_sfp_b_pattern_out_data;                         // data_pattern_gen_SFP_B:aso_data -> timing_adapter_SFP_B_tx:in_data
	wire          data_pattern_gen_sfp_b_pattern_out_ready;                        // timing_adapter_SFP_B_tx:in_ready -> data_pattern_gen_SFP_B:aso_ready
	wire   [39:0] xcvr_custom_phy_0_rx_parallel_data0_data;                        // xcvr_custom_phy_0:rx_parallel_data0 -> timing_adapter_SFP_A_rx:in_data
	wire   [39:0] xcvr_custom_phy_0_rx_parallel_data1_data;                        // xcvr_custom_phy_0:rx_parallel_data1 -> timing_adapter_SFP_B_rx:in_data
	wire          pll_0_outclk0_clk;                                               // pll_0:outclk_0 -> [alt_xcvr_reconfig_0:mgmt_clk_clk, data_pattern_check_SFP_A:csr_clk_clk, data_pattern_check_SFP_B:csr_clk_clk, data_pattern_gen_SFP_A:csr_clk_clk, data_pattern_gen_SFP_B:csr_clk_clk, master_0:clk_clk, mm_interconnect_0:pll_0_outclk0_clk, rst_controller:clk, xcvr_custom_phy_0:phy_mgmt_clk]
	wire          xcvr_custom_phy_0_rx_clkout0_clk;                                // xcvr_custom_phy_0:rx_clkout0 -> [data_pattern_check_SFP_A:pattern_in_clk_clk, rst_controller_001:clk, timing_adapter_SFP_A_rx:clk]
	wire          xcvr_custom_phy_0_rx_clkout1_clk;                                // xcvr_custom_phy_0:rx_clkout1 -> [data_pattern_check_SFP_B:pattern_in_clk_clk, rst_controller_003:clk, timing_adapter_SFP_B_rx:clk]
	wire          xcvr_custom_phy_0_tx_clkout0_clk;                                // xcvr_custom_phy_0:tx_clkout0 -> [data_pattern_gen_SFP_A:pattern_out_clk_clk, rst_controller_002:clk, timing_adapter_SFP_A_tx:clk]
	wire          xcvr_custom_phy_0_tx_clkout1_clk;                                // xcvr_custom_phy_0:tx_clkout1 -> [data_pattern_gen_SFP_B:pattern_out_clk_clk, rst_controller_004:clk, timing_adapter_SFP_B_tx:clk]
	wire  [183:0] xcvr_custom_phy_0_reconfig_from_xcvr_reconfig_from_xcvr;         // xcvr_custom_phy_0:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire  [279:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr;           // alt_xcvr_reconfig_0:reconfig_to_xcvr -> xcvr_custom_phy_0:reconfig_to_xcvr
	wire   [31:0] master_0_master_readdata;                                        // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire          master_0_master_waitrequest;                                     // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire   [31:0] master_0_master_address;                                         // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire          master_0_master_read;                                            // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire    [3:0] master_0_master_byteenable;                                      // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire          master_0_master_readdatavalid;                                   // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire          master_0_master_write;                                           // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire   [31:0] master_0_master_writedata;                                       // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire   [31:0] mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_readdata;   // data_pattern_check_SFP_A:csr_slave_readdata -> mm_interconnect_0:data_pattern_check_SFP_A_csr_slave_readdata
	wire    [2:0] mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_address;    // mm_interconnect_0:data_pattern_check_SFP_A_csr_slave_address -> data_pattern_check_SFP_A:csr_slave_address
	wire          mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_read;       // mm_interconnect_0:data_pattern_check_SFP_A_csr_slave_read -> data_pattern_check_SFP_A:csr_slave_read
	wire    [3:0] mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_byteenable; // mm_interconnect_0:data_pattern_check_SFP_A_csr_slave_byteenable -> data_pattern_check_SFP_A:csr_slave_byteenable
	wire          mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_write;      // mm_interconnect_0:data_pattern_check_SFP_A_csr_slave_write -> data_pattern_check_SFP_A:csr_slave_write
	wire   [31:0] mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_writedata;  // mm_interconnect_0:data_pattern_check_SFP_A_csr_slave_writedata -> data_pattern_check_SFP_A:csr_slave_writedata
	wire   [31:0] mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_readdata;   // data_pattern_check_SFP_B:csr_slave_readdata -> mm_interconnect_0:data_pattern_check_SFP_B_csr_slave_readdata
	wire    [2:0] mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_address;    // mm_interconnect_0:data_pattern_check_SFP_B_csr_slave_address -> data_pattern_check_SFP_B:csr_slave_address
	wire          mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_read;       // mm_interconnect_0:data_pattern_check_SFP_B_csr_slave_read -> data_pattern_check_SFP_B:csr_slave_read
	wire    [3:0] mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_byteenable; // mm_interconnect_0:data_pattern_check_SFP_B_csr_slave_byteenable -> data_pattern_check_SFP_B:csr_slave_byteenable
	wire          mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_write;      // mm_interconnect_0:data_pattern_check_SFP_B_csr_slave_write -> data_pattern_check_SFP_B:csr_slave_write
	wire   [31:0] mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_writedata;  // mm_interconnect_0:data_pattern_check_SFP_B_csr_slave_writedata -> data_pattern_check_SFP_B:csr_slave_writedata
	wire   [31:0] mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_readdata;     // data_pattern_gen_SFP_A:csr_slave_readdata -> mm_interconnect_0:data_pattern_gen_SFP_A_csr_slave_readdata
	wire    [2:0] mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_address;      // mm_interconnect_0:data_pattern_gen_SFP_A_csr_slave_address -> data_pattern_gen_SFP_A:csr_slave_address
	wire          mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_read;         // mm_interconnect_0:data_pattern_gen_SFP_A_csr_slave_read -> data_pattern_gen_SFP_A:csr_slave_read
	wire    [3:0] mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_byteenable;   // mm_interconnect_0:data_pattern_gen_SFP_A_csr_slave_byteenable -> data_pattern_gen_SFP_A:csr_slave_byteenable
	wire          mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_write;        // mm_interconnect_0:data_pattern_gen_SFP_A_csr_slave_write -> data_pattern_gen_SFP_A:csr_slave_write
	wire   [31:0] mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_writedata;    // mm_interconnect_0:data_pattern_gen_SFP_A_csr_slave_writedata -> data_pattern_gen_SFP_A:csr_slave_writedata
	wire   [31:0] mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_readdata;     // data_pattern_gen_SFP_B:csr_slave_readdata -> mm_interconnect_0:data_pattern_gen_SFP_B_csr_slave_readdata
	wire    [2:0] mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_address;      // mm_interconnect_0:data_pattern_gen_SFP_B_csr_slave_address -> data_pattern_gen_SFP_B:csr_slave_address
	wire          mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_read;         // mm_interconnect_0:data_pattern_gen_SFP_B_csr_slave_read -> data_pattern_gen_SFP_B:csr_slave_read
	wire    [3:0] mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_byteenable;   // mm_interconnect_0:data_pattern_gen_SFP_B_csr_slave_byteenable -> data_pattern_gen_SFP_B:csr_slave_byteenable
	wire          mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_write;        // mm_interconnect_0:data_pattern_gen_SFP_B_csr_slave_write -> data_pattern_gen_SFP_B:csr_slave_write
	wire   [31:0] mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_writedata;    // mm_interconnect_0:data_pattern_gen_SFP_B_csr_slave_writedata -> data_pattern_gen_SFP_B:csr_slave_writedata
	wire   [31:0] mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_readdata;           // xcvr_custom_phy_0:phy_mgmt_readdata -> mm_interconnect_0:xcvr_custom_phy_0_phy_mgmt_readdata
	wire          mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_waitrequest;        // xcvr_custom_phy_0:phy_mgmt_waitrequest -> mm_interconnect_0:xcvr_custom_phy_0_phy_mgmt_waitrequest
	wire    [8:0] mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_address;            // mm_interconnect_0:xcvr_custom_phy_0_phy_mgmt_address -> xcvr_custom_phy_0:phy_mgmt_address
	wire          mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_read;               // mm_interconnect_0:xcvr_custom_phy_0_phy_mgmt_read -> xcvr_custom_phy_0:phy_mgmt_read
	wire          mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_write;              // mm_interconnect_0:xcvr_custom_phy_0_phy_mgmt_write -> xcvr_custom_phy_0:phy_mgmt_write
	wire   [31:0] mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_writedata;          // mm_interconnect_0:xcvr_custom_phy_0_phy_mgmt_writedata -> xcvr_custom_phy_0:phy_mgmt_writedata
	wire   [31:0] mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_readdata;    // alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> mm_interconnect_0:alt_xcvr_reconfig_0_reconfig_mgmt_readdata
	wire          mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest; // alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> mm_interconnect_0:alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest
	wire    [6:0] mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_address;     // mm_interconnect_0:alt_xcvr_reconfig_0_reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	wire          mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_read;        // mm_interconnect_0:alt_xcvr_reconfig_0_reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	wire          mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_write;       // mm_interconnect_0:alt_xcvr_reconfig_0_reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	wire   [31:0] mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_writedata;   // mm_interconnect_0:alt_xcvr_reconfig_0_reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	wire          rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, data_pattern_check_SFP_A:reset_reset, data_pattern_check_SFP_B:reset_reset, data_pattern_gen_SFP_A:reset_reset, data_pattern_gen_SFP_B:reset_reset, mm_interconnect_0:data_pattern_check_SFP_A_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, xcvr_custom_phy_0:phy_mgmt_clk_reset]
	wire          rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> timing_adapter_SFP_A_rx:reset_n
	wire          rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> timing_adapter_SFP_A_tx:reset_n
	wire          rst_controller_003_reset_out_reset;                              // rst_controller_003:reset_out -> timing_adapter_SFP_B_rx:reset_n
	wire          rst_controller_004_reset_out_reset;                              // rst_controller_004:reset_out -> timing_adapter_SFP_B_tx:reset_n
	wire    [1:0] xcvr_custom_phy_0_tx_clkout;                                     // port fragment
	wire   [79:0] xcvr_custom_phy_0_rx_parallel_data;                              // port fragment
	wire    [1:0] xcvr_custom_phy_0_rx_clkout;                                     // port fragment

	alt_xcvr_reconfig #(
		.device_family                 ("Arria V"),
		.number_of_reconfig_interfaces (4),
		.enable_offset                 (1),
		.enable_lc                     (0),
		.enable_dcd                    (1),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (1),
		.enable_ber                    (0),
		.enable_dfe                    (1),
		.enable_adce                   (1),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),                 //      reconfig_busy.reconfig_busy
		.cal_busy_in               (),                                                                //        cal_busy_in.cal_busy_in
		.mgmt_clk_clk              (pll_0_outclk0_clk),                                               //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                                  //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_address),     //      reconfig_mgmt.address
		.reconfig_mgmt_read        (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_read),        //                   .read
		.reconfig_mgmt_readdata    (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_readdata),    //                   .readdata
		.reconfig_mgmt_waitrequest (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest), //                   .waitrequest
		.reconfig_mgmt_write       (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_write),       //                   .write
		.reconfig_mgmt_writedata   (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_writedata),   //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),           //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (xcvr_custom_phy_0_reconfig_from_xcvr_reconfig_from_xcvr),         // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                                //        (terminated)
		.rx_cal_busy               (),                                                                //        (terminated)
		.reconfig_mif_address      (),                                                                //        (terminated)
		.reconfig_mif_read         (),                                                                //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                            //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                             //        (terminated)
	);

	low_latency_10g_1ch_data_pattern_check_SFP_A #(
		.ST_DATA_W            (40),
		.NUM_CYCLES_FOR_LOCK  (40),
		.BYPASS_ENABLED       (0),
		.AVALON_ENABLED       (1),
		.FREQ_CNTER_ENABLED   (0),
		.CROSS_CLK_SYNC_DEPTH (2)
	) data_pattern_check_sfp_a (
		.csr_clk_clk          (pll_0_outclk0_clk),                                               //        csr_clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                                  //          reset.reset
		.csr_slave_address    (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_address),    //      csr_slave.address
		.csr_slave_write      (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_write),      //               .write
		.csr_slave_read       (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_read),       //               .read
		.csr_slave_byteenable (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_byteenable), //               .byteenable
		.csr_slave_writedata  (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_writedata),  //               .writedata
		.csr_slave_readdata   (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_readdata),   //               .readdata
		.pattern_in_clk_clk   (xcvr_custom_phy_0_rx_clkout0_clk),                                // pattern_in_clk.clk
		.asi_valid            (timing_adapter_sfp_a_rx_out_valid),                               //     pattern_in.valid
		.asi_ready            (timing_adapter_sfp_a_rx_out_ready),                               //               .ready
		.asi_data             (timing_adapter_sfp_a_rx_out_data)                                 //               .data
	);

	low_latency_10g_1ch_data_pattern_check_SFP_A #(
		.ST_DATA_W            (40),
		.NUM_CYCLES_FOR_LOCK  (40),
		.BYPASS_ENABLED       (0),
		.AVALON_ENABLED       (1),
		.FREQ_CNTER_ENABLED   (0),
		.CROSS_CLK_SYNC_DEPTH (2)
	) data_pattern_check_sfp_b (
		.csr_clk_clk          (pll_0_outclk0_clk),                                               //        csr_clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                                  //          reset.reset
		.csr_slave_address    (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_address),    //      csr_slave.address
		.csr_slave_write      (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_write),      //               .write
		.csr_slave_read       (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_read),       //               .read
		.csr_slave_byteenable (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_byteenable), //               .byteenable
		.csr_slave_writedata  (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_writedata),  //               .writedata
		.csr_slave_readdata   (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_readdata),   //               .readdata
		.pattern_in_clk_clk   (xcvr_custom_phy_0_rx_clkout1_clk),                                // pattern_in_clk.clk
		.asi_valid            (timing_adapter_sfp_b_rx_out_valid),                               //     pattern_in.valid
		.asi_ready            (timing_adapter_sfp_b_rx_out_ready),                               //               .ready
		.asi_data             (timing_adapter_sfp_b_rx_out_data)                                 //               .data
	);

	low_latency_10g_1ch_data_pattern_gen_SFP_A #(
		.ST_DATA_W            (40),
		.BYPASS_ENABLED       (0),
		.AVALON_ENABLED       (1),
		.CROSS_CLK_SYNC_DEPTH (2)
	) data_pattern_gen_sfp_a (
		.csr_clk_clk          (pll_0_outclk0_clk),                                             //         csr_clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                                //           reset.reset
		.csr_slave_address    (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_address),    //       csr_slave.address
		.csr_slave_write      (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_write),      //                .write
		.csr_slave_read       (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_read),       //                .read
		.csr_slave_byteenable (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_byteenable), //                .byteenable
		.csr_slave_writedata  (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_writedata),  //                .writedata
		.csr_slave_readdata   (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_readdata),   //                .readdata
		.pattern_out_clk_clk  (xcvr_custom_phy_0_tx_clkout0_clk),                              // pattern_out_clk.clk
		.aso_valid            (data_pattern_gen_sfp_a_pattern_out_valid),                      //     pattern_out.valid
		.aso_ready            (data_pattern_gen_sfp_a_pattern_out_ready),                      //                .ready
		.aso_data             (data_pattern_gen_sfp_a_pattern_out_data)                        //                .data
	);

	low_latency_10g_1ch_data_pattern_gen_SFP_A #(
		.ST_DATA_W            (40),
		.BYPASS_ENABLED       (0),
		.AVALON_ENABLED       (1),
		.CROSS_CLK_SYNC_DEPTH (2)
	) data_pattern_gen_sfp_b (
		.csr_clk_clk          (pll_0_outclk0_clk),                                             //         csr_clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                                //           reset.reset
		.csr_slave_address    (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_address),    //       csr_slave.address
		.csr_slave_write      (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_write),      //                .write
		.csr_slave_read       (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_read),       //                .read
		.csr_slave_byteenable (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_byteenable), //                .byteenable
		.csr_slave_writedata  (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_writedata),  //                .writedata
		.csr_slave_readdata   (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_readdata),   //                .readdata
		.pattern_out_clk_clk  (xcvr_custom_phy_0_tx_clkout1_clk),                              // pattern_out_clk.clk
		.aso_valid            (data_pattern_gen_sfp_b_pattern_out_valid),                      //     pattern_out.valid
		.aso_ready            (data_pattern_gen_sfp_b_pattern_out_ready),                      //                .ready
		.aso_data             (data_pattern_gen_sfp_b_pattern_out_data)                        //                .data
	);

	low_latency_10g_1ch_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (pll_0_outclk0_clk),             //          clk.clk
		.clk_reset_reset      (~clk_50_reset_reset_n),         //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	low_latency_10g_1ch_pll_0 pll_0 (
		.refclk   (clk_50_clk),            //  refclk.clk
		.rst      (~clk_50_reset_reset_n), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),     // outclk0.clk
		.locked   (pll_0_locked_export)    //  locked.export
	);

	low_latency_10g_1ch_timing_adapter_SFP_A_rx timing_adapter_sfp_a_rx (
		.clk       (xcvr_custom_phy_0_rx_clkout0_clk),         //   clk.clk
		.reset_n   (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.in_data   (xcvr_custom_phy_0_rx_parallel_data0_data), //    in.data
		.out_data  (timing_adapter_sfp_a_rx_out_data),         //   out.data
		.out_valid (timing_adapter_sfp_a_rx_out_valid),        //      .valid
		.out_ready (timing_adapter_sfp_a_rx_out_ready)         //      .ready
	);

	low_latency_10g_1ch_timing_adapter_SFP_A_tx timing_adapter_sfp_a_tx (
		.clk      (xcvr_custom_phy_0_tx_clkout0_clk),         //   clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.in_data  (data_pattern_gen_sfp_a_pattern_out_data),  //    in.data
		.in_valid (data_pattern_gen_sfp_a_pattern_out_valid), //      .valid
		.in_ready (data_pattern_gen_sfp_a_pattern_out_ready), //      .ready
		.out_data (timing_adapter_sfp_a_tx_out_data)          //   out.data
	);

	low_latency_10g_1ch_timing_adapter_SFP_A_rx timing_adapter_sfp_b_rx (
		.clk       (xcvr_custom_phy_0_rx_clkout1_clk),         //   clk.clk
		.reset_n   (~rst_controller_003_reset_out_reset),      // reset.reset_n
		.in_data   (xcvr_custom_phy_0_rx_parallel_data1_data), //    in.data
		.out_data  (timing_adapter_sfp_b_rx_out_data),         //   out.data
		.out_valid (timing_adapter_sfp_b_rx_out_valid),        //      .valid
		.out_ready (timing_adapter_sfp_b_rx_out_ready)         //      .ready
	);

	low_latency_10g_1ch_timing_adapter_SFP_A_tx timing_adapter_sfp_b_tx (
		.clk      (xcvr_custom_phy_0_tx_clkout1_clk),         //   clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),      // reset.reset_n
		.in_data  (data_pattern_gen_sfp_b_pattern_out_data),  //    in.data
		.in_valid (data_pattern_gen_sfp_b_pattern_out_valid), //      .valid
		.in_ready (data_pattern_gen_sfp_b_pattern_out_ready), //      .ready
		.out_data (timing_adapter_sfp_b_tx_out_data)          //   out.data
	);

	altera_xcvr_custom #(
		.device_family                         ("Arria V"),
		.protocol_hint                         ("basic"),
		.operation_mode                        ("Duplex"),
		.lanes                                 (2),
		.bonded_group_size                     (1),
		.bonded_mode                           ("xN"),
		.pma_bonding_mode                      ("x1"),
		.pcs_pma_width                         (20),
		.ser_base_factor                       (10),
		.ser_words                             (4),
		.data_rate                             ("6250Mbps"),
		.base_data_rate                        ("6250 Mbps"),
		.en_synce_support                      (0),
		.tx_bitslip_enable                     ("false"),
		.rx_use_coreclk                        ("false"),
		.tx_use_coreclk                        ("false"),
		.use_8b10b                             ("false"),
		.use_8b10b_manual_control              ("false"),
		.std_tx_pcfifo_mode                    ("low_latency"),
		.std_rx_pcfifo_mode                    ("low_latency"),
		.word_aligner_mode                     ("manual"),
		.word_aligner_state_machine_datacnt    (1),
		.word_aligner_state_machine_errcnt     (1),
		.word_aligner_state_machine_patterncnt (10),
		.word_aligner_pattern_length           (20),
		.word_align_pattern                    ("11111001111111111010"),
		.run_length_violation_checking         (40),
		.use_rate_match_fifo                   (0),
		.rate_match_pattern1                   ("11010000111010000011"),
		.rate_match_pattern2                   ("00101111000101111100"),
		.byte_order_mode                       ("none"),
		.byte_order_pattern                    ("111111011"),
		.byte_order_pad_pattern                ("000000000"),
		.coreclk_0ppm_enable                   ("false"),
		.pll_refclk_cnt                        (1),
		.pll_refclk_freq                       ("156.25 MHz"),
		.pll_refclk_select                     ("0"),
		.cdr_refclk_select                     (0),
		.plls                                  (1),
		.pll_type                              ("CMU"),
		.pll_select                            (0),
		.pll_reconfig                          (0),
		.pll_external_enable                   (0),
		.gxb_analog_power                      ("AUTO"),
		.pll_lock_speed                        ("AUTO"),
		.tx_analog_power                       ("AUTO"),
		.tx_slew_rate                          ("OFF"),
		.tx_termination                        ("OCT_100_OHMS"),
		.tx_use_external_termination           ("false"),
		.tx_preemp_pretap                      (0),
		.tx_preemp_pretap_inv                  ("false"),
		.tx_preemp_tap_1                       (0),
		.tx_preemp_tap_2                       (0),
		.tx_preemp_tap_2_inv                   ("false"),
		.tx_vod_selection                      (2),
		.tx_common_mode                        ("0.65V"),
		.rx_pll_lock_speed                     ("AUTO"),
		.rx_common_mode                        ("0.82V"),
		.rx_termination                        ("OCT_100_OHMS"),
		.rx_use_external_termination           ("false"),
		.rx_eq_dc_gain                         (1),
		.rx_eq_ctrl                            (16),
		.mgmt_clk_in_mhz                       (250),
		.embedded_reset                        (1),
		.channel_interface                     (0)
	) xcvr_custom_phy_0 (
		.phy_mgmt_clk                (pll_0_outclk0_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //       phy_mgmt_clk.clk
		.phy_mgmt_clk_reset          (rst_controller_reset_out_reset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // phy_mgmt_clk_reset.reset
		.phy_mgmt_address            (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           phy_mgmt.address
		.phy_mgmt_read               (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .read
		.phy_mgmt_readdata           (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .readdata
		.phy_mgmt_waitrequest        (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .waitrequest
		.phy_mgmt_write              (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .write
		.phy_mgmt_writedata          (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .writedata
		.tx_ready                    (xcvr_custom_phy_0_tx_ready_export),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //           tx_ready.export
		.rx_ready                    (xcvr_custom_phy_0_rx_ready_export),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //           rx_ready.export
		.pll_ref_clk                 (refclk_in_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        pll_ref_clk.clk
		.tx_serial_data              (xcvr_custom_phy_0_tx_serial_data_export),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //     tx_serial_data.export
		.pll_locked                  (xcvr_custom_phy_0_pll_locked_export),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //         pll_locked.export
		.rx_serial_data              (xcvr_custom_phy_0_rx_serial_data_export),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //     rx_serial_data.export
		.tx_clkout                   ({xcvr_custom_phy_0_tx_clkout[1],xcvr_custom_phy_0_tx_clkout[0]}),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //         tx_clkout0.clk
		.rx_clkout                   ({xcvr_custom_phy_0_rx_clkout[1],xcvr_custom_phy_0_rx_clkout[0]}),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //         rx_clkout0.clk
		.tx_parallel_data            ({timing_adapter_sfp_b_tx_out_data[0],timing_adapter_sfp_b_tx_out_data[1],timing_adapter_sfp_b_tx_out_data[2],timing_adapter_sfp_b_tx_out_data[3],timing_adapter_sfp_b_tx_out_data[4],timing_adapter_sfp_b_tx_out_data[5],timing_adapter_sfp_b_tx_out_data[6],timing_adapter_sfp_b_tx_out_data[7],timing_adapter_sfp_b_tx_out_data[8],timing_adapter_sfp_b_tx_out_data[9],timing_adapter_sfp_b_tx_out_data[10],timing_adapter_sfp_b_tx_out_data[11],timing_adapter_sfp_b_tx_out_data[12],timing_adapter_sfp_b_tx_out_data[13],timing_adapter_sfp_b_tx_out_data[14],timing_adapter_sfp_b_tx_out_data[15],timing_adapter_sfp_b_tx_out_data[16],timing_adapter_sfp_b_tx_out_data[17],timing_adapter_sfp_b_tx_out_data[18],timing_adapter_sfp_b_tx_out_data[19],timing_adapter_sfp_b_tx_out_data[20],timing_adapter_sfp_b_tx_out_data[21],timing_adapter_sfp_b_tx_out_data[22],timing_adapter_sfp_b_tx_out_data[23],timing_adapter_sfp_b_tx_out_data[24],timing_adapter_sfp_b_tx_out_data[25],timing_adapter_sfp_b_tx_out_data[26],timing_adapter_sfp_b_tx_out_data[27],timing_adapter_sfp_b_tx_out_data[28],timing_adapter_sfp_b_tx_out_data[29],timing_adapter_sfp_b_tx_out_data[30],timing_adapter_sfp_b_tx_out_data[31],timing_adapter_sfp_b_tx_out_data[32],timing_adapter_sfp_b_tx_out_data[33],timing_adapter_sfp_b_tx_out_data[34],timing_adapter_sfp_b_tx_out_data[35],timing_adapter_sfp_b_tx_out_data[36],timing_adapter_sfp_b_tx_out_data[37],timing_adapter_sfp_b_tx_out_data[38],timing_adapter_sfp_b_tx_out_data[39],timing_adapter_sfp_a_tx_out_data[0],timing_adapter_sfp_a_tx_out_data[1],timing_adapter_sfp_a_tx_out_data[2],timing_adapter_sfp_a_tx_out_data[3],timing_adapter_sfp_a_tx_out_data[4],timing_adapter_sfp_a_tx_out_data[5],timing_adapter_sfp_a_tx_out_data[6],timing_adapter_sfp_a_tx_out_data[7],timing_adapter_sfp_a_tx_out_data[8],timing_adapter_sfp_a_tx_out_data[9],timing_adapter_sfp_a_tx_out_data[10],timing_adapter_sfp_a_tx_out_data[11],timing_adapter_sfp_a_tx_out_data[12],timing_adapter_sfp_a_tx_out_data[13],timing_adapter_sfp_a_tx_out_data[14],timing_adapter_sfp_a_tx_out_data[15],timing_adapter_sfp_a_tx_out_data[16],timing_adapter_sfp_a_tx_out_data[17],timing_adapter_sfp_a_tx_out_data[18],timing_adapter_sfp_a_tx_out_data[19],timing_adapter_sfp_a_tx_out_data[20],timing_adapter_sfp_a_tx_out_data[21],timing_adapter_sfp_a_tx_out_data[22],timing_adapter_sfp_a_tx_out_data[23],timing_adapter_sfp_a_tx_out_data[24],timing_adapter_sfp_a_tx_out_data[25],timing_adapter_sfp_a_tx_out_data[26],timing_adapter_sfp_a_tx_out_data[27],timing_adapter_sfp_a_tx_out_data[28],timing_adapter_sfp_a_tx_out_data[29],timing_adapter_sfp_a_tx_out_data[30],timing_adapter_sfp_a_tx_out_data[31],timing_adapter_sfp_a_tx_out_data[32],timing_adapter_sfp_a_tx_out_data[33],timing_adapter_sfp_a_tx_out_data[34],timing_adapter_sfp_a_tx_out_data[35],timing_adapter_sfp_a_tx_out_data[36],timing_adapter_sfp_a_tx_out_data[37],timing_adapter_sfp_a_tx_out_data[38],timing_adapter_sfp_a_tx_out_data[39]}),                                                                                                                                                                           //  tx_parallel_data0.data
		.rx_parallel_data            ({xcvr_custom_phy_0_rx_parallel_data[79],xcvr_custom_phy_0_rx_parallel_data[78],xcvr_custom_phy_0_rx_parallel_data[77],xcvr_custom_phy_0_rx_parallel_data[76],xcvr_custom_phy_0_rx_parallel_data[75],xcvr_custom_phy_0_rx_parallel_data[74],xcvr_custom_phy_0_rx_parallel_data[73],xcvr_custom_phy_0_rx_parallel_data[72],xcvr_custom_phy_0_rx_parallel_data[71],xcvr_custom_phy_0_rx_parallel_data[70],xcvr_custom_phy_0_rx_parallel_data[69],xcvr_custom_phy_0_rx_parallel_data[68],xcvr_custom_phy_0_rx_parallel_data[67],xcvr_custom_phy_0_rx_parallel_data[66],xcvr_custom_phy_0_rx_parallel_data[65],xcvr_custom_phy_0_rx_parallel_data[64],xcvr_custom_phy_0_rx_parallel_data[63],xcvr_custom_phy_0_rx_parallel_data[62],xcvr_custom_phy_0_rx_parallel_data[61],xcvr_custom_phy_0_rx_parallel_data[60],xcvr_custom_phy_0_rx_parallel_data[59],xcvr_custom_phy_0_rx_parallel_data[58],xcvr_custom_phy_0_rx_parallel_data[57],xcvr_custom_phy_0_rx_parallel_data[56],xcvr_custom_phy_0_rx_parallel_data[55],xcvr_custom_phy_0_rx_parallel_data[54],xcvr_custom_phy_0_rx_parallel_data[53],xcvr_custom_phy_0_rx_parallel_data[52],xcvr_custom_phy_0_rx_parallel_data[51],xcvr_custom_phy_0_rx_parallel_data[50],xcvr_custom_phy_0_rx_parallel_data[49],xcvr_custom_phy_0_rx_parallel_data[48],xcvr_custom_phy_0_rx_parallel_data[47],xcvr_custom_phy_0_rx_parallel_data[46],xcvr_custom_phy_0_rx_parallel_data[45],xcvr_custom_phy_0_rx_parallel_data[44],xcvr_custom_phy_0_rx_parallel_data[43],xcvr_custom_phy_0_rx_parallel_data[42],xcvr_custom_phy_0_rx_parallel_data[41],xcvr_custom_phy_0_rx_parallel_data[40],xcvr_custom_phy_0_rx_parallel_data[39],xcvr_custom_phy_0_rx_parallel_data[38],xcvr_custom_phy_0_rx_parallel_data[37],xcvr_custom_phy_0_rx_parallel_data[36],xcvr_custom_phy_0_rx_parallel_data[35],xcvr_custom_phy_0_rx_parallel_data[34],xcvr_custom_phy_0_rx_parallel_data[33],xcvr_custom_phy_0_rx_parallel_data[32],xcvr_custom_phy_0_rx_parallel_data[31],xcvr_custom_phy_0_rx_parallel_data[30],xcvr_custom_phy_0_rx_parallel_data[29],xcvr_custom_phy_0_rx_parallel_data[28],xcvr_custom_phy_0_rx_parallel_data[27],xcvr_custom_phy_0_rx_parallel_data[26],xcvr_custom_phy_0_rx_parallel_data[25],xcvr_custom_phy_0_rx_parallel_data[24],xcvr_custom_phy_0_rx_parallel_data[23],xcvr_custom_phy_0_rx_parallel_data[22],xcvr_custom_phy_0_rx_parallel_data[21],xcvr_custom_phy_0_rx_parallel_data[20],xcvr_custom_phy_0_rx_parallel_data[19],xcvr_custom_phy_0_rx_parallel_data[18],xcvr_custom_phy_0_rx_parallel_data[17],xcvr_custom_phy_0_rx_parallel_data[16],xcvr_custom_phy_0_rx_parallel_data[15],xcvr_custom_phy_0_rx_parallel_data[14],xcvr_custom_phy_0_rx_parallel_data[13],xcvr_custom_phy_0_rx_parallel_data[12],xcvr_custom_phy_0_rx_parallel_data[11],xcvr_custom_phy_0_rx_parallel_data[10],xcvr_custom_phy_0_rx_parallel_data[9],xcvr_custom_phy_0_rx_parallel_data[8],xcvr_custom_phy_0_rx_parallel_data[7],xcvr_custom_phy_0_rx_parallel_data[6],xcvr_custom_phy_0_rx_parallel_data[5],xcvr_custom_phy_0_rx_parallel_data[4],xcvr_custom_phy_0_rx_parallel_data[3],xcvr_custom_phy_0_rx_parallel_data[2],xcvr_custom_phy_0_rx_parallel_data[1],xcvr_custom_phy_0_rx_parallel_data[0]}), //  rx_parallel_data0.data
		.reconfig_from_xcvr          (xcvr_custom_phy_0_reconfig_from_xcvr_reconfig_from_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 // reconfig_from_xcvr.reconfig_from_xcvr
		.reconfig_to_xcvr            (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //   reconfig_to_xcvr.reconfig_to_xcvr
		.tx_forceelecidle            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.tx_bitslipboundaryselect    (10'b0000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
		.rx_runningdisp              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_disperr                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_errdetect                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_is_lockedtoref           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_is_lockedtodata          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_signaldetect             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_patterndetect            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_syncstatus               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_bitslipboundaryselectout (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_enabyteord               (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.rx_bitslip                  (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.rx_rmfifodatainserted       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_rmfifodatadeleted        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_rlv                      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_byteordflag              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.tx_coreclkin                (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.rx_coreclkin                (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.rx_recovered_clk            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.cdr_ref_clk                 (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //        (terminated)
		.tx_datak                    (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //        (terminated)
		.tx_dispval                  (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //        (terminated)
		.tx_forcedisp                (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //        (terminated)
		.rx_datak                    (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.pll_powerdown               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //        (terminated)
		.tx_digitalreset             (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.tx_analogreset              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.tx_cal_busy                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.rx_digitalreset             (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.rx_analogreset              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //        (terminated)
		.rx_cal_busy                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.ext_pll_clk                 (2'b00)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //        (terminated)
	);

	low_latency_10g_1ch_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                                          (pll_0_outclk0_clk),                                               //                                        pll_0_outclk0.clk
		.data_pattern_check_SFP_A_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                  // data_pattern_check_SFP_A_reset_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                  //             master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_address                                    (master_0_master_address),                                         //                                      master_0_master.address
		.master_0_master_waitrequest                                (master_0_master_waitrequest),                                     //                                                     .waitrequest
		.master_0_master_byteenable                                 (master_0_master_byteenable),                                      //                                                     .byteenable
		.master_0_master_read                                       (master_0_master_read),                                            //                                                     .read
		.master_0_master_readdata                                   (master_0_master_readdata),                                        //                                                     .readdata
		.master_0_master_readdatavalid                              (master_0_master_readdatavalid),                                   //                                                     .readdatavalid
		.master_0_master_write                                      (master_0_master_write),                                           //                                                     .write
		.master_0_master_writedata                                  (master_0_master_writedata),                                       //                                                     .writedata
		.alt_xcvr_reconfig_0_reconfig_mgmt_address                  (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_address),     //                    alt_xcvr_reconfig_0_reconfig_mgmt.address
		.alt_xcvr_reconfig_0_reconfig_mgmt_write                    (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_write),       //                                                     .write
		.alt_xcvr_reconfig_0_reconfig_mgmt_read                     (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_read),        //                                                     .read
		.alt_xcvr_reconfig_0_reconfig_mgmt_readdata                 (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_readdata),    //                                                     .readdata
		.alt_xcvr_reconfig_0_reconfig_mgmt_writedata                (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_writedata),   //                                                     .writedata
		.alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest              (mm_interconnect_0_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest), //                                                     .waitrequest
		.data_pattern_check_SFP_A_csr_slave_address                 (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_address),    //                   data_pattern_check_SFP_A_csr_slave.address
		.data_pattern_check_SFP_A_csr_slave_write                   (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_write),      //                                                     .write
		.data_pattern_check_SFP_A_csr_slave_read                    (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_read),       //                                                     .read
		.data_pattern_check_SFP_A_csr_slave_readdata                (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_readdata),   //                                                     .readdata
		.data_pattern_check_SFP_A_csr_slave_writedata               (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_writedata),  //                                                     .writedata
		.data_pattern_check_SFP_A_csr_slave_byteenable              (mm_interconnect_0_data_pattern_check_sfp_a_csr_slave_byteenable), //                                                     .byteenable
		.data_pattern_check_SFP_B_csr_slave_address                 (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_address),    //                   data_pattern_check_SFP_B_csr_slave.address
		.data_pattern_check_SFP_B_csr_slave_write                   (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_write),      //                                                     .write
		.data_pattern_check_SFP_B_csr_slave_read                    (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_read),       //                                                     .read
		.data_pattern_check_SFP_B_csr_slave_readdata                (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_readdata),   //                                                     .readdata
		.data_pattern_check_SFP_B_csr_slave_writedata               (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_writedata),  //                                                     .writedata
		.data_pattern_check_SFP_B_csr_slave_byteenable              (mm_interconnect_0_data_pattern_check_sfp_b_csr_slave_byteenable), //                                                     .byteenable
		.data_pattern_gen_SFP_A_csr_slave_address                   (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_address),      //                     data_pattern_gen_SFP_A_csr_slave.address
		.data_pattern_gen_SFP_A_csr_slave_write                     (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_write),        //                                                     .write
		.data_pattern_gen_SFP_A_csr_slave_read                      (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_read),         //                                                     .read
		.data_pattern_gen_SFP_A_csr_slave_readdata                  (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_readdata),     //                                                     .readdata
		.data_pattern_gen_SFP_A_csr_slave_writedata                 (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_writedata),    //                                                     .writedata
		.data_pattern_gen_SFP_A_csr_slave_byteenable                (mm_interconnect_0_data_pattern_gen_sfp_a_csr_slave_byteenable),   //                                                     .byteenable
		.data_pattern_gen_SFP_B_csr_slave_address                   (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_address),      //                     data_pattern_gen_SFP_B_csr_slave.address
		.data_pattern_gen_SFP_B_csr_slave_write                     (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_write),        //                                                     .write
		.data_pattern_gen_SFP_B_csr_slave_read                      (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_read),         //                                                     .read
		.data_pattern_gen_SFP_B_csr_slave_readdata                  (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_readdata),     //                                                     .readdata
		.data_pattern_gen_SFP_B_csr_slave_writedata                 (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_writedata),    //                                                     .writedata
		.data_pattern_gen_SFP_B_csr_slave_byteenable                (mm_interconnect_0_data_pattern_gen_sfp_b_csr_slave_byteenable),   //                                                     .byteenable
		.xcvr_custom_phy_0_phy_mgmt_address                         (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_address),            //                           xcvr_custom_phy_0_phy_mgmt.address
		.xcvr_custom_phy_0_phy_mgmt_write                           (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_write),              //                                                     .write
		.xcvr_custom_phy_0_phy_mgmt_read                            (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_read),               //                                                     .read
		.xcvr_custom_phy_0_phy_mgmt_readdata                        (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_readdata),           //                                                     .readdata
		.xcvr_custom_phy_0_phy_mgmt_writedata                       (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_writedata),          //                                                     .writedata
		.xcvr_custom_phy_0_phy_mgmt_waitrequest                     (mm_interconnect_0_xcvr_custom_phy_0_phy_mgmt_waitrequest)         //                                                     .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clk_50_reset_reset_n),          // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~clk_50_reset_reset_n),              // reset_in0.reset
		.clk            (xcvr_custom_phy_0_rx_clkout0_clk),   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~clk_50_reset_reset_n),              // reset_in0.reset
		.clk            (xcvr_custom_phy_0_tx_clkout0_clk),   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~clk_50_reset_reset_n),              // reset_in0.reset
		.clk            (xcvr_custom_phy_0_rx_clkout1_clk),   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~clk_50_reset_reset_n),              // reset_in0.reset
		.clk            (xcvr_custom_phy_0_tx_clkout1_clk),   //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign xcvr_custom_phy_0_rx_parallel_data0_data = { xcvr_custom_phy_0_rx_parallel_data[0], xcvr_custom_phy_0_rx_parallel_data[1], xcvr_custom_phy_0_rx_parallel_data[2], xcvr_custom_phy_0_rx_parallel_data[3], xcvr_custom_phy_0_rx_parallel_data[4], xcvr_custom_phy_0_rx_parallel_data[5], xcvr_custom_phy_0_rx_parallel_data[6], xcvr_custom_phy_0_rx_parallel_data[7], xcvr_custom_phy_0_rx_parallel_data[8], xcvr_custom_phy_0_rx_parallel_data[9], xcvr_custom_phy_0_rx_parallel_data[10], xcvr_custom_phy_0_rx_parallel_data[11], xcvr_custom_phy_0_rx_parallel_data[12], xcvr_custom_phy_0_rx_parallel_data[13], xcvr_custom_phy_0_rx_parallel_data[14], xcvr_custom_phy_0_rx_parallel_data[15], xcvr_custom_phy_0_rx_parallel_data[16], xcvr_custom_phy_0_rx_parallel_data[17], xcvr_custom_phy_0_rx_parallel_data[18], xcvr_custom_phy_0_rx_parallel_data[19], xcvr_custom_phy_0_rx_parallel_data[20], xcvr_custom_phy_0_rx_parallel_data[21], xcvr_custom_phy_0_rx_parallel_data[22], xcvr_custom_phy_0_rx_parallel_data[23], xcvr_custom_phy_0_rx_parallel_data[24], xcvr_custom_phy_0_rx_parallel_data[25], xcvr_custom_phy_0_rx_parallel_data[26], xcvr_custom_phy_0_rx_parallel_data[27], xcvr_custom_phy_0_rx_parallel_data[28], xcvr_custom_phy_0_rx_parallel_data[29], xcvr_custom_phy_0_rx_parallel_data[30], xcvr_custom_phy_0_rx_parallel_data[31], xcvr_custom_phy_0_rx_parallel_data[32], xcvr_custom_phy_0_rx_parallel_data[33], xcvr_custom_phy_0_rx_parallel_data[34], xcvr_custom_phy_0_rx_parallel_data[35], xcvr_custom_phy_0_rx_parallel_data[36], xcvr_custom_phy_0_rx_parallel_data[37], xcvr_custom_phy_0_rx_parallel_data[38], xcvr_custom_phy_0_rx_parallel_data[39] };

	assign xcvr_custom_phy_0_rx_parallel_data1_data = { xcvr_custom_phy_0_rx_parallel_data[40], xcvr_custom_phy_0_rx_parallel_data[41], xcvr_custom_phy_0_rx_parallel_data[42], xcvr_custom_phy_0_rx_parallel_data[43], xcvr_custom_phy_0_rx_parallel_data[44], xcvr_custom_phy_0_rx_parallel_data[45], xcvr_custom_phy_0_rx_parallel_data[46], xcvr_custom_phy_0_rx_parallel_data[47], xcvr_custom_phy_0_rx_parallel_data[48], xcvr_custom_phy_0_rx_parallel_data[49], xcvr_custom_phy_0_rx_parallel_data[50], xcvr_custom_phy_0_rx_parallel_data[51], xcvr_custom_phy_0_rx_parallel_data[52], xcvr_custom_phy_0_rx_parallel_data[53], xcvr_custom_phy_0_rx_parallel_data[54], xcvr_custom_phy_0_rx_parallel_data[55], xcvr_custom_phy_0_rx_parallel_data[56], xcvr_custom_phy_0_rx_parallel_data[57], xcvr_custom_phy_0_rx_parallel_data[58], xcvr_custom_phy_0_rx_parallel_data[59], xcvr_custom_phy_0_rx_parallel_data[60], xcvr_custom_phy_0_rx_parallel_data[61], xcvr_custom_phy_0_rx_parallel_data[62], xcvr_custom_phy_0_rx_parallel_data[63], xcvr_custom_phy_0_rx_parallel_data[64], xcvr_custom_phy_0_rx_parallel_data[65], xcvr_custom_phy_0_rx_parallel_data[66], xcvr_custom_phy_0_rx_parallel_data[67], xcvr_custom_phy_0_rx_parallel_data[68], xcvr_custom_phy_0_rx_parallel_data[69], xcvr_custom_phy_0_rx_parallel_data[70], xcvr_custom_phy_0_rx_parallel_data[71], xcvr_custom_phy_0_rx_parallel_data[72], xcvr_custom_phy_0_rx_parallel_data[73], xcvr_custom_phy_0_rx_parallel_data[74], xcvr_custom_phy_0_rx_parallel_data[75], xcvr_custom_phy_0_rx_parallel_data[76], xcvr_custom_phy_0_rx_parallel_data[77], xcvr_custom_phy_0_rx_parallel_data[78], xcvr_custom_phy_0_rx_parallel_data[79] };

	assign xcvr_custom_phy_0_rx_clkout0_clk = { xcvr_custom_phy_0_rx_clkout[0] };

	assign xcvr_custom_phy_0_rx_clkout1_clk = { xcvr_custom_phy_0_rx_clkout[1] };

	assign xcvr_custom_phy_0_tx_clkout0_clk = { xcvr_custom_phy_0_tx_clkout[0] };

	assign xcvr_custom_phy_0_tx_clkout1_clk = { xcvr_custom_phy_0_tx_clkout[1] };

endmodule
