// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
wtiDDxfEZ1g3/BrRw0nQDwGWPcXYdIA7huBrSQfKSEF8XyaeRIRmdWgXOWro2nF2NJW+gbB+P6Zm
vIanCRpESIbFBJMrAIhrSfl8SbR3F5CqJmc/wtTSnEXcFHCxSFBaHrfeiifUyGg7KijWkyzeFD/M
tQDIiyeOtoXY/FUpV1Vqzj+WhRnieu5ATL7/gYSvqbviDyK6OKB1rClGJnmRx4mW+T8hUZc1AOG2
Dg8DpfLTCjckiqOCq+NooveeyIOs40unQpsqBVp0aIaB3IWz6V3xO3ZCtIoscmnZIK2jrFOpJNRK
6Ihql6WBy/+xbXIpM3zZdPQ48nOL4XKH8Y3/Tg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
02u1cKZ9Qzjg2AMakDRuxW0r96KZHmivWiviv5/1QqPVhzg2OtL1+W3k9rFXmQRGNnEoghRU2aUf
0kAZcVhzHJlBOB15x339c4DfWb4We/cN/5luAjk360iIkaiJASyw2dxByaTabYGMaoZVxS0znsdC
Is1tXK+0emB4VYltFcax8bKzvki4IXECx12KqEGFInJz1B3SoD3EkSJ9y1iG+kPhg2lRdwDZyW5g
+giyR9HbpSp+m/oUNPaOeMBhnJYh3buCXayu4mthGYWcqR5zS2Ctk7qsBbD4LJY2bwvelQFqIgJ+
gfXYW2AW1cXA9Y/XHP5LRbMRwIotLSaxBdixX74V51WsEGZuB4RURxVxNvuTpwSTaHWnC5euwzVs
a1zmp8hntH9Ojss18iXDzftc9/70jjUTOZvymBFJXxpAUu1GJyGzQbJGbg9rD354YZFtw21yBBd4
iWMsgCAbKSM9kEmKWqgNoPQk1kLgKsVX5hg+Olye68c7Ac3yW+sDM1+hG9PhKsdCyLkBEuC5YnGH
7sZ/dzN+g2buWLsAFqhSVPP9or5Pb4ekizQQv2Jx+rOpagzcAUqG2T5xOFv0ZthM2p10G77efbeu
AYsfV0YT7vkyvhaOTeDygEyze6KcjaHgtlPkbeldHcLiB7ni5RVC42h1Xy8h2qyrIc0Pd3/Y2vCl
QXgt665Hn8BnBjatiZ6q84KzisXJiHVScUUVPhawclQiIdzzzk1PXlHEh2Fo0IgwpmbtaWjXVvR7
RMkJ4e0W/rlR343CjPUJqOuoQo47Hri23oMrkwYzguuO5o0Wk9lkD5fw8r+OZ0ZPJRUTg50pXkyT
l5GqkqHy+1kTiHrBBY9mw2bWPRc7MLnBtOGck2Mgg7hhtzN3wNjOX5QpV7OsW6dCxk5A4V8NieNA
ZguV7y+856Uu25mNMqWZRuu1mzeAxyzlZFyseT+wJS1hspsR9UvZ1wW5i3GrMD1O3/ng/GiqGZF1
vqpimA9YzwqM5oVmP1xMcX5lw6gFIKj74qNy2LDVRlg78C5LoHri2WFUZEwRW2NHhJjfLk4jZ9uh
aQSzo3Z3Skpg7b1TWR7cZiTFllcGpXU55I1i4vQYj69rcykvWmRGSEwf5kMZ3Kz1Bv2N2o118D9Z
zPdc9NxyBPYLlzmOCAl5/krvJIA6XKSOo3xenxVvlaegN8V7ZcG3cz2spQJ+CyqPBHWIzGQIGEwB
MGK1DUE5Mk77ovRj/HU0n0/yYLQg+/U6Zf3nepgeR4ZDEOEOBlfiEsCgzcwZz/ZvTzTZLbwX/mZs
/UBa+Dq5IwCnGEP+cu/LpU9bpt8qLpLQlPwmIFPtT9YYUrhK9+2Q54BugwskHrEAGxeC4fzct58q
T4mi1KX38BkV0a3QN/a5lLEHRyUWDLACTlP4fvfugJRe3sQdxjtYxPhPzRA0RdSYOoeITw6aP6m5
EJoReGZBvOa9HHRkbM6sxpIUXJvMEZvmEgNZqTI6yyTYpL+byQirbB/wNtHVvUXI+Oxo2wdS34Ng
36E8lq2ijkR/xHanmbWTt3GYu8payKpsNkiqiIze1O5bhmcSjzxDmNQCTu8GIEfnAOuTKI+XmSgz
ZfwVRsExvZK2y0VYVgih5SilUj3zVat20eOdtqRz/6w27N4b+Rc7nPl3J2WKaLLfyAnxIkOYWSjH
Hv/2MC5kmCl5Dr9bRj6e1PlKfe85oLY9Vb6inQONvw0OJBzpk7FL7yGR/+UOZ325PonLILNtRwNk
yVAOCAwEDkHhd8snbk/vvE7Y2KQVI6/Uv+wFw+aJDnbJ7n8mNvHwbsXAU4pPtmvZjVkQWyRaVM2C
l2wkMwM9z/r8ArNT4p9m3/Ans+FocIim6LTStXb0hvqIM37sapKcizh40vGhH7spn6QIF3yoauPD
KndK9Q1FAGZdoYqU5ITTe6woFHMJvX5S0pSDYjBm3icrLTQUluD9N5TAY2VBuVCnnWjTHPhzB+z+
LV7r2TIQQ+W93vLpCJm3lM+7Zl4suf+1DGAijKPPQP/j+VmlR93poKX42RUdIbOnGxOK+ihG/+U9
ro8RKpTfplzjrxhE6/VhSYp1ZH4y2qQOqEh80XjY3g2wVOEhYdjEzQwyvO9vbvP0nhRCKqby5pd+
rUoKBxTrNQFb7wPvZytYhD0fD0sQ6940gv58nCtiYcfMb3JKWj/lShJybRZ9ViewAeFcLxlRYxri
oHGe85s16g370sWoPmQUhoehP8e3fubnqsfRlIMQCxXp/by1xmD/QSJlsNCb8nzXyzf5YZFq+H1s
o3yhg1epdWMRAitrL7MBb18OebMC5dI0vo4DlWkQOVj/Qp/7q9wyDqWyUAEkS4Gk0koJxx1bUeVA
V5hRBKiva7flgrcl66L8gzBihj+dSG8ZzBh7Vc7vDnUHYpaEy4iq2SqLM0w0TxdPfgQJhmwsVCsg
qWZtFkSHa0dHTr0PYTrcxHKlPITtcpeylZFKwMRKpSbvRFe8nd5lSOELHxycE7VjqQ1D49cmPGy7
ny9XaqE94O0b1N4c4PSjwrRTxF4YZXuyArz+B06r/jFbAovwYq5FZnpl1vMtFtVZrPyz25vPQmy4
PTFwEBlEn4oPW1eEfxcHZWb8klrxDZtENZNKc9TyRLaOdb1yfmSRLg83D71s7bzU23zGQCZXorBS
cE+unZazemhC3vOoFp13LhybAQZF9xXDi0pP551Uv+bH1G4/QTeXGml6pJb0mIdDiMc/z6xBNYOu
c7gymlrzn2CwdushiowhjP7pWcx9HuH1j2/0V84M7jz/erJGR5YfZmCsODdKp6YAGBVjF0QGQBCT
ycgyWGRKiQa8oDr+Q9qTWBxwtb/dsde5rgl31ZpzLB1GWbuw+FZM/oQve+u+NnK6xN+iVmaXfsY6
XBdHC+i1eL9hyfQd/RQmRS85tY2ORNWpI7vZjsqGFhwDAVMznLVHpdhMXHjJKWhKvmlp4pHSQI7x
w4hTOVsxu6U45oZJ06gX7uF05sU9dW6kBDFXhPXoVJkdCkpYbwA8PPCRcgsXKcPGnxGtK4fppb2J
NVYNsmS6yNj0b7bJXz5fwOEFuNihcbM5gkA/cSjX7ILhPNE36wbHQqhAkHTnU0gUrisaJuRQvWzA
4TulJWq/W7T6XZq01CCNxXQkidm1JjlbU52GrmYnr9RzSllk5ctNEc6AAaJSbus4dQ3wT4xWNkwU
Kbdk1XmbMeBizpNpFpycAK3sMMpHB1Q4ZlTb+wHWiXVNGe3GlqRtH3lAsL1LyPMnEW5DJlckJLkk
a9g8EVfxZ8aTaJQNIDrJ/WkEzcAruMIXGVjZR3szlc90ACfKIyyv8pwCl/AqnvlFG7yqVThc1o0K
ZdMfKrayUfzvMAPK8Mcus9qooyjZaanS2FgOMHeU4G2MNUv0OwAB5II0k6OM4dHLwV8ykS1e5ma0
jhRiosnaXR4C/p8NDsK1bOI5BSaWUxbhjjk0sj/lg4YNJiAEv6aHg9ifkxCGEolT7P/XU2qOro0V
lB4JZJuvCLGkPXOwSz/MMpuif11ZpDiFAw/Oz0gcwDQ0s6PiY/CTVwH0f58ki46XzYv0b49OCXvq
IFc4pkn2+4r0sEJyXjAsv/cScWQcra/pAbX3mk3JcSwB0AlTf7iFs6l2RkKDCJa4YOTtS4RPcRSX
wrD4/RfqTl2WOh6/fqIlP7cPA5Mnrd96Xawozom76/dmxnGalMQKoeQK48HBrdhA+9YDHhe5ZSRa
DYOw3wE+owtlVA0/l7cSCwcQXVH+TjX6AHPIsPUShLE5/BgvaUf9CoXJ5HjPt0E7LIaGUoq0DYAY
f/+Rg4qXrIv7Oa63vM6ijuN7FNy2cjx9mApE4BArVNf2g/nKKE7Jf7Z8arfWBu0aJgDuThYkEMvp
ZVSSWueq6NtE4QU+IXSm3y16q1Tsnugfgl0rV/8Y35/OekgsWu5Unjk6GKb3DjhzyiiScc0SciMO
FqTtLGHNKh33aasN5WvdC/hvhV5xcWlALg+bGIAdD7Kwjuzz7+2s74ZE7+dFgkzbuthdBdZWE0Om
vyvAMzww7T3H1QPLNNgVN/4Vzglz8K0Zh8TWdCKOVKMVuatoFq4rLvqYFYFZABeC8iiDk0ZGPjtJ
kmFVDSriQV4/8x5yrmOONqqO55H2WG2QGjOOt6Qpb7TuDD+Fh/h7xDIEuwYq3CaXpAcv3AsIP2fB
G37ZJvznTyqY5mCfpB/YIdBq7jkEUYhVEXylHmEF+u28SK5e1qSABf094pUzqUZU/YkUmAawCZ1U
gDZVSKR/el1XKFGmrvgLdYEV9SOmlzRBeDmM/B3KNTsFqEjffTMEvVF/xL1QIJburHYHUcuZtVbf
1z9CXXLzJVMMi3+Guu8zoG70F/Fv6WpTCY/b67ek9wRw5QAjUwTPqP1NLJNtdvDELKBZmew19Q2A
qc6nhdWKFyJQELWhCBtsnrr8cUk/7PSI/awxFovNk4GNfRbhcPMrqml01/T9oB1JjYwApvEiv+7n
EFsKaW/rWqolaUxpFf9KjrVPaq11haDYG/akglQd1GCh/mlgdV08nX5mNzq/HX9uWPTbg+qrIDwb
FzRo/k5v8mWlLcRx/tmJ9oPTqwGAn3g++8C5s//UwaVxwo17uQN4wOOOQORlb6qOHqYPZUuTuPnQ
G1CcWkNXOoDw36EyrZZSfCCblS7CjNA6KVxMSwtxvxKp/++yCdVI5xwWmQzfSRUFjU5baWkXtFPY
JFq/p1tK2gelE0L1o2Jm87FhH1GJUPLE1Qo5KcE6tMdc0W/qXCR3a5CKV2KDf+yuHqFwgdiYgFrV
AAoTyLHjFbpINHGqcxDMIdMkHrWq2yX8zXFfzYMvcCedf2fs7907A4d7J8bpNElM/4LCIshxFvF3
0yR2RtIPaEJ+/dRx6+eUS6V2ThbmOafgtSiAao62M+eJuI5MVDb9UEFhvt+ukLS4uJLlYF/nSwHP
YN5TthrCY78zsnmGctt8Ai9OAt983Qo6BjYPwQNcKEevaC0hBHzvl7OLnDgLVRJ4Z81UYjyEBJJV
QrosFpj795xcOjmqzXk4tI2yYj+sLZoPVI+bKLuTFBaWeH7Ngxcs8nPKmvbpEBpNjlrvg5b6mTF8
F11wDaAAqnBYDDOnLF/4rUqLe+DKhtr58U6JEu0KiEYnzF2NeOshSD08drRBvr0SgoFdMKIh6DhI
+tE97wBX0TNiIRiD7nvZdvuFjuM7urEBYFNtb/VRG1SBV2lXid/1HGSIsYGdLyUi0D+aaynu/5Gg
UwrtoJGvEt7F8kGC4iQm9fIras/d/0y5jLDjV5KdRXOyBZ73KdscAubpfmwN+SBImvW0ldhHGsRe
gFBb3VXX40B8rjdeJAoyDyNmHO+N0/4csaT1ju0EokcAHd+9Lx7F5Jz8gD2eUvQbFMh6tzVYU9Nu
dqkgOdqqsBkEBSMYFpsIAz+DWiUirlsv7CwIhkqhzyJcY/VPcgb6thU/9LGAZ2IcD3YTOnqzCEs8
JvoQqWn+u9raUn+TWg5ZdHL8Vjku5blXifRCg4zOLPgqEe/lGkiMv6sUsG4EdzXuZpTqtsdc9PoU
BvsW4RmbuzNDDcokBtRAaUW/Degn3SErFgKjTUeQoI+ymFlfZEBhrlgMGK7ZesYsonUvAEzBNAzX
vJmpqUAsDD5HtxN95cAgGo+so5+wH9GlTD2kx2AuiZZVA8VLeWpKqorVpa7d20/X6AmUPC121U7T
RoJ3qGTogAxuWf5/xaN2Re6hkGlXy5pegD/xAP9iiFR1Z8s/1g2IU35vmEJEFxqBw1qKm6YpB35h
ncclpB4Gwa8RgLSkYW5LPubv7YOBhsJm0UyErjPBtvQCpur5xJx5h/Af4ELT7h+IfWMO6QRfpAi7
fT/d9xblQNQ5l8uaPFRWobo5yIK9k8Eh1zoOR2A0fq/+69ilVQnibzX4O3TC57bT4HeFTEXcLyEd
e0hhsdyt0K5tccNJJp3ERUnoSjZml7xuM39KV+GqaU6sNGJnbDTgwyX+/VQCvJLspmlQNQhgI1zZ
2SySXSB+2DJQxnBtUAnsLPQ1LJW4tvd/YrcugUE9xRhKsZLGQdW/yckB206cbOpLHxfK7CgtSJW6
SjH/8yABK+A4X+jukRde58Qey2IDw1uHOiKHNNFP7MYZQCJmWslA9AceHt6N7yLXr8wio1wbMJP9
/cNei1pv+T0TLtxSKiDjCuLxPlaXbM4r+/7elsLcstpfgyH0Ox7d7g6sHq+ZeR6NwQz8pL4VnBxl
7+Y9QHTBLehQiHZ5xLJreVC+cobQOS6FUioee8uuSwIoKyUPkpVndXztPSURLW1GFHwIHEnsYNJF
X/Zf/+krqebRYnQbIjBn/IcVSDtfvCoB32WcfruQUz9DHe3HaBOD8kkF+SMjTVZS8O2cV8YWcK+j
OjvR1hJsmxBY6G1XBnZK2moIn7nE4as8i7L3SBlVg6VsqkUgYaR8rOkBJwUcNUwUgNsgDmmCwSAw
fl2jFF5LDREVJQ/zg35iigQ70WMiab5zCD4pRmZkAiDLhOTzfQIaFOTe4qxarnvCOWJCGzyiemDf
lDQcwWOKNyaF+J4G4b9JTrUO2lP5QB2lJCaRaufiU2zVVSrf9NAtamcWSrfJK086aqeJkqpkWdBL
B1jsC4777BD63cXXjrxl/xhvPqZDGzy5KP6Q0PP1l8+3a4Cwp+7YnB9tKmC/wA5hWo42Ne3myKCh
gmfwiaaSPShYdY2sLMPoMoeBkqXZ5fh55TRO8W8svGDpBnCCbTt+P+hXNqoxE0A7H5JxOBbSSXk1
GZR03cKqtwSwl9qrWuJN7HrKjxorvNEZBEeyWgWChNm/7OFdIowWVNLevfENmEXlPzFaSUD5M+Kz
mosLOmWHbr1lsMhP5x74dVbvuvRZ7WO6mLblndFcE+Grd3scf6VMGi231HTv4tbMlgY82LfVweK1
WQFXcphc8l+xAYYrstTz/rCCyxpn/k/hFAJoTd+n31sAx7fhAjBIsevNoNZvY/OJQ9TarVHwzJCK
oel47sxJI5M6RZXUuOqVr+3xtNhxtqy5StW/xeQNlw0UFvT0xtEKSAnfZGG7OqdgaDholDF7wCCh
Z6vYmklhgmX4bgmmDhR16/CI0RBwDpUDUCSbMLoJg1+93tPJxJk4D3oF0DnsXMfbxEOuOYABgIOQ
8ACBEQKyF82rsVN7F64gKda7+SHsPTazNPHyACC3y159dlD9MUzNDKvIA/Wy4mZV79NXgRoipJyT
t/2rI0b58BnYOFUYKZ4zFGEnQD8vWeyCU0EU/HFGFsxvDH5buXsm96NfPLV1ShUrjo2/XLbHOCM1
+DbVAJHlzCau2P3kBUKdi0LETVhY49VtiMI5z/VDik3ZoW5wa2BaKBcZpjGpcYDMBQ6Uwt+dOkfd
AYV0g90y3HJiWiFw5Qi274g1lxC4yjo7k208QGSQx0FqQcxI76wAYYPuEqJ8oJBkzlnpNfCzQC2K
2kHRfTPqrHdpGdBmtWtydWgBvy02gza7mH004W9gJon/I/9RzasJRt1ftteCe7ovVwyKP+Ld/Oox
8V+oL7fCXcntQyz1I8MCggDio+rHsQoGtumkSljenfDGKBwiGvEHOHaPU4oGp1BZ4LPnRiKyjCiQ
RLy5W87/0bdaI3nanRGAjQvej93Rhkroba3/NzXSXdP2aW41gQj0VC4ZCzxOCUMFWEDlGPrcEtXW
Fh/T
`pragma protect end_protected
