// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:27:26 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WwgKO+hEO+1CPt65kTcHqLzwvpJiDXr4XciVKs6GDF+Yrhzj9focF8IVxVwf5Gsn
fb5330DiyVeO2IBaIm1mVVl9td9i/lY8AqEr65pRwGQayb9T05vLhjjUNu8jdVZj
GoXFxv4qWM02PyRge+I/kmt1W7wuA+JN9eyfh3F//MA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8000)
oy/VaXFLlaJyoH1dXVyLxRvh0eV4nL5vehmta5/qnIzQfdujqd2WsFxLdQoZPeNu
MYUzKhtg55PAaUsowkoHZO32GMO13vV+r7p23chkU/pV75ewB086B4gWzNRnLM8Y
DeN8PlWiJS8+6wxGbZ27no1K3ItCkEAKyCYVgMOREHp31IDatLu1GvwEixDAp6wK
3lGU3bHx4nhWBtDbiIRHonuRwvSBJ0LDSddyNWgYUoJoC10Ms0M6RNImSG+4OLUS
1ocL6D86uHWXp6HS2d7DF0HQchduA3dhnRYVJ7BJcFFQEPpgOja50fnGwkY3z6dA
xx0P+ZMxu1yCcRRKdYo1K6Od/fXs89q1y5KZYJEgMGpyqtO7y+Qy91uWzSMSL5Or
/Awu2Ib6TjMw51U6Ho43rhJJkL05fHOdCtjsRkwiSymjw2rTU8cYRgRFSaBzBOj9
CGcAdO1Ux74Sx6/TdImcgMAsPRdwmWUg5dWNt3vr57BG2o959a4LjxJfRFJCZpH7
TFxJiylBbsE8NBs+2u7puIm6FCcg77ENyA9TWkBVAjBaFG6uPilTINxAeuC7j6AL
WOiJu5Zwc2P5DkEzdRGMhqBkLFXhbLOxsrg11LY22aXoFKwN6ywlW22sb6v9tyom
/j+7HsuZ/6LL55nI8Tf7AXqVl9E240u39VKM7l9FTR7zU3X3tDu2CESpSKuMn9K6
qBnNCs78LMkfCrrCrmSHHSqc+KuH/3ht0srIpbU92exZpvNaM7xN7d0NJ45qy8Uq
eYX7WYAXRJy30sZvKa42JFDZYYlNZ4JTWZzhtsz+M7f9aFqqxO6tl6gAEt7a+xZs
ykGpu3oLDdMDbLRdAxgmhUDPHERU2smdbdkQT1qbSkySxnb1YW5Q2QtJMHGn0vZp
Pa4Izqfi6EGBcSpeA0RsvnN8nAJ16c0dlJ2skZ/SYGBwVvgVGbs9M93ERlv24BIe
6fb7gYp6i/628pda2EXfg8i3yPTcBAGpCAJQFKaChlglmLK/5iiGdJqN/UDQPNBA
A7m146Agxu5B/BcGYeigifrbXGDPSbGUIkYf/0Fh67AFHVQqh6tgZQOSUuMucm6b
d2YKCWmXCPYreaQfvCgbVAEfDWIPFeqRfY3VDam4rceoNBov1HrEcaureN9yCUpz
8HRSXeEuaLhs+dpOHFg8J7t4E+edjr65aId48y0VCN1cEzm1RiE+Hb6pKNZ59+zk
nXEl6MhyHrTs7Pqp0RZNOTRU127qqPYYLe73xig6pvda9JYh07ERvhhVk9ODX9QA
maq5e6y9/rn04rhEfqNYnKJJRYB5OPkcl0KgSZZHA+FlC9dPIT7qzVqgaOE84BE0
8shA85J8yNA0of2DGnlApXvlEXL7dsGlPVCUVCD3vHzCaz9XvVPAKD0tzSUPT0+u
1ulB0UgFB+e4Qwhro1sIn9KwAxX6uJLx3nYwLxCENukqVkPJwR23+Ktr4NVl8NGT
1rkO7DbfjrFAphB1F7g4LtBSH+vPUAkB+C0Is1reQqg3oddcnbVzGeLUTCCkdOMA
hB8ZJXTX9DXdHg2e39gDV6cH0Knwrp2rcLymNk7i1zQdp6DzQa+S/TQEy53E2a6d
inUwu3wlcNXSPwKPOyFi8kvfhb+jLYBbFgWJ6+AZWz4n2O5jcI3t99c/oRQxBk5x
5Z6aTYQr2KGR4/WFd74lP2C7zL43D83SLqoWLL34hi4CFl35eJxpReJxiMR5crtV
5cm2CCq/FsiRRrJLCCspGpuyXmhUrICzT2AUvP5XD01mn9TwyKKDWt6hvPIacq9X
2Du8aNTtMCeLLZzvDHP3ChHxsRKXCq0PrDbI1ldOFQuPvWaRNg1QQKnWx0r8Flvx
B1rztVwB5ZW7PLjlyl6J9tSiuEDLIZgeZFoYuNXnERtrpXF6HdBHrGmMTDFOkbCY
giXFQejrIvAZPFFtIEqv8FarQJkx3WbuqFgKE15i0777LrgoKYf6YuF779Zq8b6e
X13k5yPYNfjdm/af3JaWMFwF29usYW/8AXEGoDvAD3GoLtczKXXgpxQphSh01l7b
wPn9I26LfKv48WAtMx7GdR46swfCEAMTb0AOcEXGcN9/CD0sSCBMiNkX0/Y8Obtk
BbNR7A8g5BUlmyuHlxRn3q8ZA3GpDRKJ4Jg31d3R8oBzBatc8yE2dthMTtQZ6Kve
FdA2RR85w8223qQXHR/NlefdhZRcnyQbh6hT4FSTUXvNa/IR6x5QCWXeL73wNFvZ
Lt6RaXh2aObXQMNLb+JtDUIurGVbkazBv41sB++vgMct0kYXbD0XPLS0DWU8K6jh
5CalzonnEQ+32kajFXo4D4gcjsij6XMahfrpDYPXWGNwpcZPJItkk8yHxehadK7r
E5ScquUCnsNm6Vw4TOGY6j+4ElP56mtBqpjEDIsilCDeqiwjWDBrSNBKQ6Vv1Lon
mxuzFnuJyirTN6S7sz2YwNd/rhmD4c2V35yp0GdGP1efFxBKPYLSejHqTslXJjoZ
kQ78S64fEdmSMm2KfqD18IFdbp0uB9aHB+r+9ADKsDhOi1ng+9D+X5tSeOAzTt6c
kb4ZGNuM05/Q1G2+mIvBmy6MKNnsP9xzqUv6bVmVBkC/OwXap646S1nKHDys11ej
hacy/FS7DdU6Wi7gpmbCkQsGYiB8ueRikllJYiRTf9M04wmeJlT+vo9Xh+E7toWM
h2h+vgmbzlirmbv1FxhuFvgZGaPQ6dlpxgyp2tiA7VV2JJVFQe+L5CtFnMR5Vwpc
3FLQu1Ts/ttAUZK5yIAaham4hrzoMh5msiGyLtjo0VyGXLoEquJfg2OnUpZoz5+y
Y+d5lXTha0W9FSGHmfni8D1n9NtYD6ZNNsjL6V7hFgL34uZNjK2xVtGUgDJvKztS
yvbh++Co4ZYzsvUcY4rcY6K0EdFbDsCiCtL+F6IAWY1Dnf/XRs9/fNtRLLvV5F9B
QA+pMz5SPMhXNw0OvaF81R14dAL5nxTgFWL25oUV4A/fmh59v96zNKpge3ryl1ZH
g4mhEAwWv8VC9CXNHz/QDJkn4Y//+qr8EvUmc6PnpbTGbs40+E6Ni5rvB2F6tIUI
og/PsxxXgFgCUrh2knN4f8CzJOIwNti3vvKrwdRQHfiX6mioqFrQi+WRY5VD88E0
TK+dtKPy4KqadlgoIIYXfnNlpboqaaozRXIcIz3SQnDRor8LfvHNhp4aoy40G6IV
33zohXaEzuWPXzWPYR3Nru0v69PdxzutexE4aD8ISu4yX9O7B++TqGSspJnxB5P0
SAMtYiIFxMIT6S8jCGq5dvMQGcDKE/Uhxrlq53IYYU+KZ7peqU/LKss4ZJjHYcX4
FIBGMyLekD+s9Rwv3x1wIXXuHEw1MMJlPy0ma3SuMHMT/yaTmDnHTkLp/cW30kgn
TVBJJrSqObW/IAtvDKqt91nfThBdffkmWbhhcK8o2cv2NRAGIzW/+nYUBbItTsSu
zPNrq8CSCWSld7lo2xXdQvv27ymAlS2ndzKO7mGEZKUaDt9MAh4L7QbBDkoDQjrA
O2wzCqMY8m/IMWqvjto3zbRC74rOpI6qMdW7gKF39VzB1cyv38+ws6EkITy6l6SQ
PK6Z8kso4QgzzX//YQ33MUdjpQp9X+Gk397+Yq2i4toRGwN3LAihp+tydR/gKS0F
09vNUgUVWXRAYtJlGLXMZS3VRiO/chonO6Zh6vJwoONxGuGL+Obdo2musWhyhY5A
1gX+srBSrj7zdz4ULQgJHxzpBVtaB0Bc6q/3fYKpvlFDCCyxV6XcgeyaZZqc5JG2
dsrBkqktZVW6qOmGya34pwTmsjGeaAEkiSom34IYTgw1TBo0iRIKd7tsTKvVDBOA
P+1cXRy13BxerU66hB6yQ1Xo7XAoZewNpnarvC0aviRk+RIbCTokOxmFSNZxVnBt
3u3X/CKraC0oeqL+XWMy2Oc1D8PljxkCWKLawwElOCe5LgRjWj0n/dYVooPe5BF6
rq/OTFrpxxYN36Bz3pDpgDhdZScDfXJfPV/S7Joigj2lhukllFoYLFY76ywsLVXF
D2rdSjyEyktthvfjT1rSt8dKdlxyfptPIjjLG2o3Npe5lZ9w/fi8uCwbboW6pbXb
lsjIpiviDGpdOLNPLPHWE4Sl0FrWAP97rb1YpfmnvbFajUsmC7IAZan8aZmaZtKW
alP+mR1zMWxWycdUnuj9jufTIZVEueEbrF4sdNx1E5+vyyL8yTmQQJajgIIaTDzq
fqliI7KizETO5zeqZPNT+o8YVbWOwh3W94AFYahL5mZTa8YQDUmLIo9TShZGeCim
zINVXhbUHR/waQy4bUJyOSAC2b+YsZ8BivKpMdYvWqnDV+jNK+KbXJqUKen9cfRL
uqHOxoBiNxAykJLUZzmaDvBJ1QTnQy0o1wDJHyYMJPpx100uDi8H517fP0L1o4Rb
L5HUFpulGsUUbLbt07+jqGx4aGOShdXbENkXOgS+YYDGpoB23yzPIhvwuyC2m33A
Lj4KGYkkc9yPwpZ0LxILO8MeCF/Ht8iBCtB+3J2EaKgQ6kWnu9cpFge20VD17WAE
AtqHqgh2NY9U8Yguy6nqRb1zoqprKctvhWwhahSUeUNFJSR6NiRHUkjz/wt3Hrse
pn4GlwkgkEtwiiN/DirFv2JssI+/mX5G0V11k1Uo7pcHEZPX/cfrysslGWYqP2lP
+69EdSQWkZNx903ns2jp+hufrfTe+ElAXZdhAh/97RmnrhOb8R++Zm6O0P7XYj3F
Adb9/G22ySXbbQGkPW0vBnCPunT0vrkaJjTBnQS2tMxDX+IYDe0n13U0bfK8dP3O
mR0rIfczpiVNQ0HQn4aTx5jrOjd96HmxTdaBUZIhRWTFRblRdWz6rNo8yz0bT8EK
IO+46yJ66PIPT1Xm0n3/U2oFlKXsg6HHI/aazpSN+18Uu78c05QgyUl/Oq3oOl3J
318y4Pa3luZzPM/rDWcOadufMDCKxwGdi9qPDxCqvD+OtazzyiR+sI/L16Ddpciw
/jxh5FK3XVi3r4TqNgMnVzU5SN1w1msGyf7qdr5aKjKwq5uocIYeyQTY/WA1QCXd
BGWI9g1hEE2N47Uq4WyKWCWatszwHy2RxJssQwc+Mned0RBZSIM9oYWSNdPUtj8i
Vkk+jTungnb98R099JiOM3CDmMKAnbbWjO7XSGQ3XgBNkUJwBVe4htN9gkK3JavR
g4oUszh8CSJtq5zqecwAavle4+Bn1kZieew7KJM6S9RRfLmWZuGnO8cHNV8Yprq8
LxZTsoPpmxCqb3qBGnHcHnGgEjPjtR0S3hA0jvwA8eFHMXq+46cqlkecy0qVMc31
idVOiG9woqT0Pr80qlyngmz8xiGt/OLcOfFU3whG2dkP5ZntW72yKSIMIxM0EVBQ
f/6fREn61PeFkcGBcaCDdb4/pSMeDcDSmdY+fAg1DFmuh45ReEMc2MyOe0m5xIEr
ohkmi4x/p2eWHkndWJPv8kIqsMHhs6X6sSVQD/gsjqkZfVbwZcGI2eWyrE9ZOR1J
kMx6Jgc95Lzu09S4PudU7HgmKCs7zbo/o3Q72d+HgKF4Z2ChG31eJZycdjD5N+oH
RCP19+FqR1OhauHkjod8k0SvFfCNV3nEOCsv129wYToblVtPDLVB+6EV3zdsuCQw
Ak1zPqH5o9bFnsDldUIwYIotsbKOpOlI1aSbRI/88+MSLHEfRdutsWA5Vq6ioY6/
CPN8t2OOwyA3NYkB6Rx1RCKsgVeaj+vfpmF9UyDMfmiOBimyTkEPswRS4r9foU/m
1KNhW4vrg0pY+3Vuz8IQtm20xHh6F4dTMpjZf3eEhEhnx4RrZ+3E6Ym67QiD9PwY
8m5Tyi0b6datSNczgkQKROOjDH61idw92EViRfwGlXp/rufgDMQEmuFhAQd/Ros+
nz3EKMLi2Db0ztQctN79GFGDsW4PJEAIB/PlBM/QgxxYdSsezht31sxNtCq3HOsF
fruCKKAvPjk8rosZlzBkKtb++m2VnNk6+jBmAADvHsYCw9ie5pnVRlEBzWScppfu
LGJEgE/u+hnrmWKzLqRqVdWxGTWDoNvUI0Nnb4BGjO/+zfWuAlvH3jL4Dte1RenS
tX+O8szqJKtn1c1RiQzSeTXMyrH/hiGTnlTb1IvOQh7V7P2ejUAF7UADMeAKmO64
x8tour0M/zHPmLRUqdedli1jrdXu/8dhP8PW2MQK0Bq4rcsmcs6kXotm5tfZeNQo
+IV1476t5+Fzl7RuII3t7CSIcUQVxOjL7+VHIaq2SWDqTEIUS3S/SIzXmsztyGzg
SEzGsiGbwn3LkvkSjM9/Y0RrfqQLr0zgPp19uYV51wGqfAjc5ftew7EZiRxyMqzN
8Sg+zHNGUui6VxQBZa/P7PYGolaHI/JIleFaAyKkyVyj/P/mp4wbbfcOQPWRrIyG
UKlkIzfaMFavskOzbx0HMp3BuInCguG7XKmi5KHQZENeSZ8xmtzSwRm5hDuTAyQM
mzSGTKL4a1t/f216rSP+bltbUiZexuyPqgWAx8cVYWBWPWsWl6m1OGNNg/BtQolg
yui8VhzqxfckgRlBgaFQ8xxRcRNMYmiPhSO1nnaj34baB1XtRzgnw8IF8+fda6Gg
ZW15y4JktyICKppb1b0RfsHFXzNiKLMSxCdSB7eoUDjVYeVDH8pyyKa2Te9n7oo+
5qqwg3vIEoytKA755ToIqmNSL0EOTDgz7YC9umZlAAhzUOZJHbXoceanssh7D1Qn
HdghFJBXjebcZR3PmTvrWhC5CDR0444g+fTii7LxGwHLntd3D/+UPzz+D387SUnO
FSSx0nP/Fokcd2lPf/FZs73KIfvRm5bnzcTXKIZQ3itW9Gf2HBUo94d978tv8NIl
ZL8maKt5Yb/doOYqosyvglCHfuhzHtSp4kiv6KRHGMJfNayB5qMC3SB0LOsssV/l
guGonoYCA9Ia9tIarJdAwJCnGQNtZjovFA5+qyhv87Psz/8aawYG/teX+/OxCrK2
yQz8kqp1VgJlbiOymlOfJ+jcJPpPF3/POxaGSps2e3VUyp16w/VhqKJl69jjtaVU
fdHmH28phz/kK0/eTwJrB10nmN2W0OtnJoDQnHbxngqVCyIRZTPWSxqwnkzmecjC
zORrBRlmMGyV3RL2TRCXQNHVvi3KVUhHRrKFtvwUOYZ7etMEkQ7Ai44aVtnwcG0e
kzUeswZ8MKMxBW0VYQIc4Bm0jCJ2qCB+rm+0dqCPjg2UZMq0IgYhw1C9PjDVoLOH
XZLPRX44iQbqn/PicdrSD+l9kdD1qwNrVeXZAxk14WctlEpRkJpkY43fdsv6ZqRm
u+M0ZtGd/9KTLhvE8tW6KBj+vG3V9LSr8FsN6teZZVa7uCd05ytIc5joMz+zF4rl
UORht4lc7HD1J8y0p8Erlx0jnrzX1nSkWBaQFGPpGvhJIZSHGbg6O2YCGCma5g/K
1GEBaYBTiv4W9soWFHDb1ZmgB4NQ04bdD6kJylSewewlo0De5WbDPGWVRmXCtbm+
nwmsRiYgdWbc2ZGnhx58mEQoPXtadAs/nz4BzSMAlduAJrkfp3wVjYvBClXLEDL2
3AUuDYcniELTpMJO3z+bAzKRfYkEAHH1klKYUg+2/i2Rn8kRVAuqYuGOHtXEFhi+
jnbK3fFZKGr5cUUQY6mdUutJt6TChleeherAm5l+SqvkyV30yAoE4tIYL/gukTQb
JQ3pLjH6NmB1M9/no3tKDLf7T94jzml1e7GE1fPTj0M1LSiEiLSYXeL/e93sVAwx
1QX/fGM3l2ImsNAMkkbpBqrKOBj0LTNMusL/TCUXL7g7QcDAurg4fYXmKUPIXfvw
gr51QYhwsbuDaEttoT055N1nRZDWLITzop1ob/n6EIeZeSNAzwDpebiUzdTpeSb+
Lt5NVJbWFQzhuHQww4BpH+WxZkxQQjGVd278Np/di4+fuTm+UDF1BBbFL1Dt16Pq
HPc0/NY0lmdRPGhHLNJPh2GX9tC3cqYSVGNQVyvauAFrSbpcChYX7yvEwbI2Fpwj
UChfoyWrsXLijZg5I3+2D4L95VEN4NhumVSkbENvmP3rR6RxxZASXrpblNDfqz+z
XJquJNb3BI1GWPiCLwVvuZAW8xZPeJziKJ1oTp3ymrSIED11d50c+dw0YiLVkK+3
0QxLGFqOITxhPvYD6KKQcaNw/QTe0mvxSWEhaZC/+r5i06bPXVNU4PFYmOyhE6KJ
tCW4wKsIIONbPvjO9V+wZX3xAKuueMc8UWn+HDPe3kNKeL4i0+mmIAeEsofmB8Sb
k6KQ2fMalbF171k0c2AZTcMMm+y9FC1bqdPqCHGeF2976y/ydcwBZtPudDtn9xO0
hxNJCcJTbqPkBAsHkZcNB56Cy7aikyJvqKfylVudZjc/CPCx7aTrGmKcTf7tye7x
ffxL61tDE9gh3NscGqG02lauQgaQu6U5h1sURoxHIcmJF+ZPFOiuISF4GgnomPLq
OSnnNQ/wZOU3drfH/TMZeZz39EIUG+i64z/uNqc8EjgIlr3/K5oM+9GlHgj+69NL
PgMHQFTx2fo4dUFYNu8+ZJnc6VIm2wHp/QvC8yUeouWhs8Vnbs399xtaGxt1pFg1
yojQ6ykGWgQ73SvbWwpIXeb92rZilC2C87WVhFviHaekCSr8WT4dX7P9p7cFZQal
rAzvOpS3vcuFq9SskLC9DMKqUTH8SK/N+EKyCDUXRzQPIZVmBh9iBsa2oLeSJkDo
DDoeNX33VoTo20ikPKsHwhdYZqzmd9kBwlVPn1sf3jFkEWuqfP3lyxJnVf7RnAvp
IDdbABnRp9oJtc98S+vvK2AMkVx4GQxruIP8L+skR//uii+1pKiceU7qq23UWZX7
cqMZLXYmvZDeHH2vdLVs42ZElWAqOhNsIWlBc+jBzjaAJtjJsK5Bg2/4x+ZKe3Pj
VSs+lmuYKvXIULFFwdx/3m1Zwk0Ge0g8XCftdgcu86+AFxqTixbG/Le+x7KB+WOo
PtSxNStyQ6hzcZ3+s27aaj8Pcz+68oIQiZlQdOeT9pgQjHiXuy2KaYz6+MFVjuXB
kLijwL5t3S3c7rZXA05aOMhlgGIsM+br2p3el+MdDNV1u6TnxZCVw9+0gAc83MKH
CErQdMVsNEJCZ7vHpgQWjuyr4+63cMQZe91h3KotK5ZkVss3z4qGh6iz7IGd6tsZ
yF9iuAjqiY2NkRbTxRGrR4eSjF2HM7oEbGEHmDaSR7tUpeP33TJx+cI1pISdMP7Y
cP5H7QjvFUJeDQ6pW9MyfD2uhzPycfyPTcoaS920gSFiBP9DhLPHn/jiGZJnntzZ
UkZexzlOP28E2neonrf5WmSoVXsGgY77/84olmTtGDqUAoMnw4T5suWQtNB4fZ85
qbnEm8wrChm92crkqH+54pkRFJ6mt9ediJKRBTsygI+wzrx4CkF5Hwjz0HLkp3ah
zgQsVuKOjdqHrnBkH51L2J6+vR47Qt7ZvZy7qC20zOnQ/fOZ8pAXa7xKmviDTZaH
zCPVtQRywbbH9t4IJZy+nn6Pz+ivYfWRiYC4PWXtl8NcQyASAiSVZpR6NP2v1V4T
UpP7q/xCylGhV85vKUW+oylRzX34jG7xH2TW7FMW0wMGzJiKWdpjK28FJww6o6V9
awCoNRxADHaQPKsEhiNg1rTZzkrMO7ZDzN41a4dQjGUya7QXkjJvpn5SDrarQSh5
81gxxCQUwqmcsTYg2zgUwypdisx2NUUHaYnUCF3AmplUFm9RKpnhhKjzTG3N9+CH
JlbevnGy2gJA2eT/zLN3/HVLi6/K0OBpDE/NtGdmyJ9ETczwl/Kvjk4017ebbXjI
3gEReS4zIsACr1ISCHNfbsjvP83PllQa93ww3qKRtX5re5BPLC3006y7ebu25/o0
ULgtDunYsXDJ9VW/zUbkrAXO7349BMuVSLPH1tWgc/Oqa+Oit2YixUVtKX94kMXL
JJOPjXB81OLDxv7hbVdFHP+s3p9cBPu/0EdUiuE5EJL8V9MQo5KcCtJ4IzAKHXu2
mxsrUANv3auSBb7MZ7MJsdM0GyDuxSmBDAbbFvOz8EKzzkVBYE5D87UOeQxOonm/
2T3cJRfyql3uqnNAaDCwWHxs2YDT1iUslGV4g9Z1SyAuAiVGFO9gXxt2B97La3xX
rEaXs/gnKU1vCnzx0Al8t17FcaAtJU0nBvSpGkU0momDpE2tABlyT+LzsJr6wKhM
gSLBvOz3x3h/vq3G3giZ1BItevF/AdmAmIDBTGAllkZbeDIp+G8NwAYVrQPTHtzQ
YIaJ1akZYXsyr8C8SzxA4tFC5yweiKydbTrL2MauArQU6m1EheB0kIq9yT6GuyYW
4UV7nZXSinJTBpYbVMLeQ+fdjMMx7OxIqPTPKP8sbQQKLgzIyx7rIG4S4dQNyDik
ngR22jOi6KepyYAiMvTDwb+F5S6BcI3arqmevDX1hw6r1VwZeVmpnWQwTnPrTwQM
tLZqptQp8UJCiOAhMSA5bFAg/vZX38dmHtYpYt2F2Z0lhBtErd6SxNq8lgogdSy7
n/d2Y6+qB+lT8pmarGX8Ax6P7tr/e7cF89PEiCBY4LfK5i+BlevWcMS5ow6f8v4M
vEr3uGMZllGrmdRNl1kb3A+71+EnBawF2CdCKPEFsAFjZta89fzYoATun5Rsn4OI
oag9E6Qcsl5iNOWrlkv9HdpMXhqoiydTyyTUxtamatY=
`pragma protect end_protected
