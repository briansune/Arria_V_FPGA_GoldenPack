��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O�Ä��/����f&4<LY�^P@Fx�)}��QF�I*Po&�p-��s���p�����,,Q�x�LH��o�}�����I��HX�	�hc�S�1�5%�ؼ�y0BqD��.�
���
f�۫i��_�A��ڞ���`�y��Z���9,JxG�k_��(ڊd�����$|#�C�ɖ��q�C^
�����X�F"��uO�#%����4�k�@CO���"� �C[��ĩ�Ю��A|,/\_����N��h`����H8n�!�7��V$��R�0�O��U^[�)R�n�c2�4�8�Ibu>)��\�"FGK��VC�^R޸��x;������r9.���l�dRQ���%���/70��2�^�[gR8D^�,��oܐ*�J�lM̌�xy�h0�F��pJ0�5��gi- F�b����8�"��r7�T�_���!Z�1�'�e�؍�ʾ�Ҟƒ��}
�I�Ix�_��6d�ϥ��
��E����♂��Sa��!�ms;�A�/������_-���?��g��F��<&���_&�W�5�p�!� �pY�SdP�d��N��%��D�|Sm�	��ȸ-��P2ϸ��/�>m��d�ș��9��$?����]����'a&�'�o�A"��E� ��c������U� �z����iB�~�4�񹹃G����[����
��DZo��QÆ����ֱ���ڍ��ʛx�\$��
�A���~�$?�΄$`"~T����N���8�:�L�{��S�]�����!��s8�7{6g+��E,�[w��x(���@@��JR"�FU�༶i����]XM}�]w��c��OxEO�))Uދ3���m�g���%���&��.���8`�#Z��;��޹r�.,�}�.�ZP ���g����l���e~{�nb��"��t�*(c<Es���˱q!�H�����a��^ì���Ͷ���9T�3(�e��-��břPٱ	�7kJ�6X��!�>�sjA�*��I�^�6@�n�\�C����A{(J$��d�	a�VMX]Yf�R����u�/�G6U4`|�����G����0�!.��#��t�b��~#��y���z�/�&4��F/��tn޺�|�-�$�5���"o��Xʘ��Sz�6=� 1ݭR8)v�}�����0�#���E���Ӊ��k��E*Q�)���1�P��bg�;'CK��@q��6�b3)ʁ����c��fQ�~R��'��XP�
�)h�'�r�Q�sd�|[����t?��\Mq})yr�%�./BTi�y��<��a�HY���QR��nQX+���>;�D�f(�|�$��x���W��}N�Y=����]l�ܠ�Դ�g��4d��҂���ƌɝ�w�qMec���&Y��ܕ��ԧ6�����X/�ݪ��T�oS� ��Ax�p���.h��	)T���g��|7$<9ȭRC��{�!��*�� d�q����U!�����������)��A�p	E齠+C�l5�c�}���g���8<� l��߁��W������|B<W# A�s2$���ø�ef1P\�e�ݰ��{ �Y���u�׉z� ���n�:	�3�1����M�%3a�5
r��U�9���^p���^Vg��o$��P��̾��x ��m�/G+- �*ɤʻ�{uج�o�� ���غ}��r��L����}�0��{���T�i���������JMk�.�|:����=:���'Ë�ʳ�5
���WJq	�]/�~[����J��������X�+�2�����x9A#j
y�1z_�D����8�}���G��Ϯb��u���lg�G�`M�6�ӑ�_(B��~����N����hy8/�F_��|���Np����dLG5y��j���6F����Z�}D
��ǒ�h�rm��h��?�9��J��F��-���fuT�� ����0�>�����>�y@/��g^q��.�+C���0 b?����8�9_�1�u��.X��"Fz�������$�r�������!�n��O��k*v���`>��,jrм!n��ߛȬ��z�;��CH/��w����vm�����ˌ@�\�,f|�ӎ�(�?N ���Q�1�^�������ݞ'�%��鸂ej�ΨKIT�]tG���Gi����{��7�Z<}��9_']������s�$r?�������ImQ�t���ZF�:����o��F�WR�z�K���d?��ܴQ�z�g��+�/�O�H.�D�@۞��_�=�P���F��9պ�C�Gz�]sME^�ǰp���%{��� ?�3.K�zčO�QKș��њ�9l��^N�� hO�@u�֧���6R���'V���?�r:���%""�]5�Y�v���|�x_��S.�E��(�K�5���������')��>%U,�7�=>�w�W9�!�,�q��ݙ���D�E4���\����ǳ����x�7I�E���z���c2��z�U/���ݷ��>ݝㇻ��~��E F����ǂ�#���R�,4���rM2B�Sk����d��7��E[h4Gт�°`��:|R�s���}r)v,^�E�CZws�ڶ�6B>N����{�b7�v����'/*�oG���m�n�� 7oQ�5�*��:��4���o˖5|����&ja���f�ƋO����5fm��Zʲfv����O�"v��_��4��+�`�8�c�=O���hZwDjr���?#���L�x�����&h.��~\T{�F�Ǜ4$�a/o:$���#R3�p�E��:�4r��0O�F	*��T�%�>���@�˻O�9������n�q ����6넇.�OzH~��r���s���_܃ ����
�"���Mѩ�PAY� }C �6Tm�����'�P��N|5u*��k��o�W�@� ��V$��z�=�t��=_<1W�x&�񾕺�"7�Յ�Tf�"���zz�G�4]Z���cA�쐌{��q�9-��� �󓦕ذ��y���L>�l�-�&w�����uS�[��s���#��D���-�H�7?Ww���h��*�J��x�O1fe�z�����6_� #=H9(������v�M��ꪾWv��P?8�����-]G+n�FǊG�j�8�S]�p� �.b�Ä�1l�>HeKm�%.���C��Kg�P�t���JZqG� �Ͼ�9e���]I����eY��Hl���		2t�T@���Lv�i)�����2�e�n�_���H.<�2�z���g3��T(�@ٵ\�?n�n�7tG'�=�y�y$/j���Ѱ-��*���{�$[ 7��ҵfՑ���bD"����2�.�Bҵ�;����s���o��3a����D�O1a�2h8�$�OA�X��IƮ8ڣ�������ئ���;�'v�{��=(5�/�ڣM����e��a�)�ʁ"��<�N�'�a�^�qlv}K8} &���' �aG�D��[�i�OV�g�!0z� 2�F�����5���w��X�U�@�!�"�QE1L\V�O:�:��p�P��X��l�̬��£2�щ�n�x'�L����F�9��k�M0��k�S*[?�<�f|��+'6M��y���Xz��O������/+Rz��y���P��ٹ�
+�T��d^Ԋa�� ��D�T�e�ݝ2iap��ݧ		}��JY��*90?��i^��n�\��'d�i��J�=�EK��X\�DL8we���	�6ڢ!VW�N *��>x����3#U��+b�wp��
��[�O��4���@�7�(�,L�M��tYB%/����+�BK�k|7��N�(@��u�����Hua5�D�����/T�p�}9���"��2�'�F|�2�
@bT�������듼/�|��B�g�F���W>i	9�ȭpÚ��P;V�2vx�qh1��b�W��<�YA���CeNhg���Kp`[�L�=?{��ϝ"��z9�� Pi���yZ�MKDS�c��0VyFu��m,����{ʨ�/�1Ō��eG)c}F��M!�O
��%Q�"u⮺R�8�k����l�R'=��	�R�7�N��-�������z�vl_�ȷ�1��漖Җ�H�X���d�3������`��:���>O&�p�wF'6p�\�ZnP����{�II���I�y`�� �*ue�pX��F���B$H>�J��F��t��oP���& v(_���ao��[U�7Pה(�RNg<��w�RYw��u�aY�SѴ��M����O^s�'G_ϻY}��V\M�g	�2���P��W\��P�5�Yԃ�v��/���be�������n#IN[
%���/����<�XCnt,���̔�3��QgQ�A�e0v$�M+��7Z]I�[���2c�gN�	 �<�(�۵xiՌ����0��Z����l �m?�b]`�.��9�La*FF��:*���.�1�6*n-�������x�]�̒�Wt�y��� ��\؜�y��%��#� ^u�G���	�]�C1��~1�Ш&"�9������N� ��r�F�`V�+/�;;��-�G�Q�Ţ�!������.�F�W�������S����0Z������C�P&��Ct����P�;1"��MؾKp�p@�P�՝�>�+��t��KV���Li��Q�m���i��	�����z�̌���b$��>�4���-6����X�Ľ����)���+�C��o�(!O�[J8�O�t�����[��E�Ɏo�I�J3M�9��I}. �Rr��i
�?�������f��E��$�7�z�@��<���ve[? d�\ք�ۭ�ϰzH#S=�Գ�P��&�>�' ��eb(�ʂ���R��a}2z�cnw�ap�s�:"���9ҍ� N��G7�����i�D��7rU!�@��ԭ�i;�yK\�c��S��}����k�l����ҐT�}�:�b��0�|w�+����1��r1߇�;��N�%���\y��?N9���j������j�˕��4�$��/�\��7i��˺�E�n9��� .���0�i�mU@�:��P�E�֚�E����5՟GP�n� q�~��5px��ʼו�}n�s�?Bv���P�&�(y$���8h�at�B�k{CB�e� Ovs��r��"�5���K��`}����^H���%�C�/9�(�
M������0����I���/5Rgq�"�`V�'M�W�5��%�[˴�8�����p��~�m	�tR���䁪=^�&�u⅀���W�ɰ��m"��	�*n�l?%P��tqTa�b}��{�.|��S���
䃏�I�;v!��N+��s�@�i�6����S�"3_ł���E8�%vV�+{*���0���s�H�ϑ��s�خN^��V&��L9�+흏�|g
��ٔ�����FfT� ]�8E���$��ؿR�Sl��t4_��E�Y��Ɲ$��cù�GZ��{&9� C�9�4
ۣ	) �ϵ�`��Jif�8�HX���ؖqS�G����_�-Px�x��)?����r;ְ�#��j}��RBt�������O�4^
�ގ��fT_�[�n�#��-�n�΀�g�+�/h��.���۽�&��YN��N�;0%����c][8�~Y��
'�sD��Q����6h�����| 9)���:깿:L��l~P���B�{�$lz������"Ms�8A��҃�e�������!o��9X$z�f~M�娌|���l>m�v�_�l#�|��#g��:��0�a�J$0�t���:R8����7�TǶ��G_��5)��Ȭ�"Լ��{ �<�<��+�um��X�1�2MK)�j�<oW��f=�R"�rX_W@��	y�;�_ˉ��?�*ܧS����eId����W:N�W<��P�7z4`�RZ�>C���Y4�bi��������3y{�-�ȃRVc�,���y<��AJ*e"m���W"ߦ�e�4��;~Vb�+8dt�^��Z,�Q�@������w�F��Vs�f�z��� 苘7뒣I=� !�͑��9ǒ��E�VU����^X�����㴞�\���`Oq$9D�[�V,Η���ɵ���G໕&�DN����pIt���4�!{@P������j�i�9��3ۧ�d�z������3���/�8�$�|r�G��L���/mk������م��� �w9r�1sȡ^�n���2v�ޘ�RTu�dFT��zb��ҳ���#��,4��%�8Mqm�����`�
��`O���T�w�[�4K*i+1��Mͣ�������]�����t0���Öӭ��
,V�����iv؍FQ�z3e-xQHM,�o�)�S[�U{ێ��[� �[�RcGH��D���
�:Hڎ��<ݧ�[�"�i���-%D�pwx�ƛ�G��V[C�ψ���%��{��$�����2FC_�=F���l�쭟��p׋�~�|����Ҏ\&������I�M��ͯ���@l�Xm�6���4z�)�@O�]��/�ϙ%C���$��� A����C�,n���y[�X_z����Ѐ�(��5���Th�<V�Y�
���w�C���x�n4_}2���	��'P:�p��R��U[V��)�b�#�f?��0B���m3��ұc�ʮ�T�@��Oq�p���ӵ�]:<JͿ��Mw���NN�	g�ϱ��7���"�
�h���C#r*���?O�%��JeHÁ����D68�����h�P���t�Q4�q2\��ɝ�u&\���YC!]R�*��
��cKȗz�F�G�����k��֝wb��+,�vP�������0'�`=*�f������t�0�f��B�}U@;�3ʵ���*!�VzKVb]?_`��<Ꮕf����>�&Ōl����a:I�!%�y�z����w�BqT�b@�B��!�߱���?�2��[�5;Yh���i$�`��AgD��>�#D��ʯi{ߵ$��C�a��j �ڣjp�@����٭��2����7WZ���PJ�����WlNSrF���x4��J��ʝ(C�Bj,��s�G���(���S/����4�B��y��V)=���ղ9#��P/��l��˸�� �(]{���VJR�)��V\��)Λ38AϏ���xO�<��r����G���������:kbF�F��ןߋ�ݮ.�qOFe�
�4�n�%27k����(��i0gi�f�L.��~1Q����O�JF�Vd�Rhtk��a����S�6��Rw\�kUB%h�������H���k���ݻ6��{�EO5��N�j(���~�N��y�S��}��(�q]?�z���I�S6�(�;��jW��/�p���"cx���<�ZǏ@*��K���3۲P��ȿ��CF)�b� �������<�t/�3#��#�����*�lM���4�j��H�l,��I���������#֏n�ݤ��Ƕ'0�_��w���K���#zA雿s�	@7}��n'B�:�rb�����rdxŊJR�T���:�7S��x�wY%X�`�ʊ�`)̒�S.x82��!?rY^�[�~��,[��p'i��GG�48��)�����Ô2����2{'�Җ凭�j~:.���lH��Xbǚ7d�18�{=vx�9#D-�۰�jM��ĞV��&� �J�	��<0��L�w`�;��)�����HD��!����V=@<�b�?��9�x���ȉ�����w՚mP��i�2���w{&��ϰ�s��o6dP�L�dT�
KV�Q�)!��(lׇ�u:�*aa�Q?@��S[ZլmK�ڏ�Q[l�R³P�	�҂]q�~KIR������t�K�&��Sd����
}�CJ����S�Ex)�*N٩�Ų�}-�6c���9&.��Q��Ȑ��2�a���� ��O��.�����������Bcr�\�|S�[M:1��I�:�7�	ž������0��g,��"�;o=� ��GQ	�㍻+������~�a���S�n���-��V��i5���F���2j�]J�4��v��R�7�evMP���6z�-�)��B{,Kdf��"gx���a�/L��P��ǃ�c֚ʈ#��U�D}z��!mL6!U}�ÄTոR�.V�)�/u_6�����������^�����ɚK�ݸ��B�)l\�$�&�o �<�ӎ�h.�e穮�i��V(�_�rd�@u_���$]	v؏��3�D�\ G4[��BdT:�X7�og�aY�=s}pܹEA�f�{�����v�ǒ�~�+�R�Iq_~^o���eS:�
�K�X<"�˪�b����h>}�R!���uC8б�>z&%O�ƜfN�S��B,�|�����0�ֶ`	t�h��f���#6#�*�i><j�Z�"2E<[����cfKC�*JL��B�\
Pc�S�ߧ-���F"O~���68pq����|�.]�<����ќF���ؓUwS�;׀�^���m�jX8ܲ&X��c�T�0u��`n��'Ao����@2�w�����:ZW��t� ����T�aj�o���������q(²ă(B��T�Ā��1F*�}�Dݽ#j���_+'� �}A�� Z�����6��C�`�p��]\�l`����u�V7x���bo#�u��1ׯ�!7�@�vU
�s��"�N�Cޱ��v�u�)NH:���8a&�ir���Cག9ga��?@����j[}.Zl�f��{~_������Sͤq�R�~U��t��&Ri��CO�r�|�r�g`�sb���Г���z3�zH�J�r/�1�&}�)5b�`�C4U���-qn�����s}�E	8�Y��y�1�8�	1��y_���?��u�����.��uX��f���\��<�<n0��� �)G;��@%1.㌢��g<w'U{l_'k}Ό.o���CjJ�IR�! �#ϼ��ZQ��ʽ���qr;��u���h�o��N.�)�H)]�)
���\���M�����&�6��&2<��[L�w}��9s�X����[#eV������M5��P����T��v�����by[�`���q�&@%�)���r6���4:etp�kn/���GƅӒ���a�.o���{Y��x�[m V��mȷx3Y�����}P�b���c���]l���hܯ]���(6��)��ka�I�a�]E��^�2ũNf�|���68!j��-��QUƺImk$����a�z����Qp?e(z����~Pl$�E��mX)�w@��벽���2ړl⡴>���2�>���q75�a� �dSe36ܽ�46���U. 6S�A�,�1��0'�����.8��_X6��%Qoz�c3�V�M��	�����mF���A5��������y����j�[
G䰳[�����{�39�<��tLa?t�/�O�C�.q��̳c=�v����O��bq�g,�o����Fϔ��xZ䍙����0�^�@��Ӽ�{P..�(X[��:@g+ƮAT���f�snP#�M/�����歋X��y��bK���<:V?��0��v��};lW��;F9*���"���,����J���"�0W&�kn��s��_OA�������G�4���#$�8s.�� b�҂���/�#��b.��%: �>z��i�SWP����f}���e��,g�J(�c�QYd�~��xC t�!�ڝ}:&��&�%䙙�FeE��95���:�)�~���6p��u�L�Z�Ys��2�a�}���<_�ls9-���c7�Ky��+7���]F�P ���p��������$�3��U*xn��^���.DnL8l`��AꟜ}9��A��n\�K��#���~�!�|��"��'	#��=o��4C�A�Mj�7��n5lS}wI�+� *�9�%tb+=^ŵ+5�fί�3��n��>�����+
�=��?�����I̤�ګw_>�vf��On��V�W/�Oa�Q���nLzU-Í��iy����<\� X$!a��Tp�kz
�m����
�W�b�=3�o��wΏ�rl��,�Q�|�0!����&	փ+!>�X�4r�����&�9�b8o2��v�<��/u�{�Ϝ&�*b�v���L��Ӗ�2D�g��9<�L��D�qH˘R�����q��^1��lT��9G��sŁ���ڊ��ڽ*�"���5>���6�+�?h�ݮ��	�b� ��Z����\q�Ԛ�v�*�W�2��W+A�A]Y�B��|���0�T����y�@L.}�̺+����i�����#�uh�;�=���G��Y�����7���{{�o�نXwS��8nbX"�ONs���q��7O����)n{���x�ǘ�lӣ5����z
�$�렯���#&+�Y�g{p!BRȦm7쯜lT�a�@Ha��s]؆i�s"A�?%�H,�=�	%� @�q
0v[�ǭCw���y.���q�M6ড়l�~PQPlp�f5�u<I\6ȃ�4�[��-�D�֦�h*�B3�����ل���#3ΕNi�c��1=z��"�F6vK~E�6����銯[��Ǭ�=x�z�&~�c�7�G�����Oϔ����yT��X�IDä���Ç�(|���Cr	ﭷ�T���4��%A����M나�'��D���b�Z�:i����+�l����/ϲ�յ	�~�j8��OWψ��w��YocL%Xtf��&Y�"k Ҏ����c9�������N�����Nδ��7����X�
�PO�3<]@bQ޶�%P�?sU%R�NZ޷���=�z�vJ��*����Wwl'�2�`s���,R2GW�i�0�g�o_
p�h�i^寔,^�������C�</�q�yHn16�I�ԙ���Աri��m.%P��"`3 ���zX!�$,c�_��$��E(z|9b'�̪��Hm��
l7%��mNwɇ�r�jT�Ձ+�/ߑ�݉^{t&
�t?o��*��
��{�/j�Ӱux�,���d9�M�RO�7��<�@�^��t0�6 �UC5o#j^8Y7Z4��b
�T��]�Xd��sm�?��<�C����fƱ� �2c���x� ��_�����-��f�'ު�V�CȚ����GS�<����k�QϥR�E�8-Tȱ��W��e��c�A��FI�b��&����֚tqr(�kBM��x
��%�	�Q�Fsu۫wV�/�U!f=��1w! �	�7�HB~��| �fB&�K��aU��ȇ�ls��)S��~(bnb���$z����r�EmraA⥴���o9xB�����F��pJ[�t�o�Q��ݘP���_�c�
R���i�%a��8u��U_}��ڂ�x�ڀ
1����l]��e��D*�>d�'߀D4"�]T�21ӗ�W�#��@�?d�o^,��sqO+��s���$Ě~ ܗv�зVDT������6b_�I8���|j9�&�!���@�xͼ[?���|�j��� /������ĸy�Im�t.�"
���:��an,�O�@�����`�k�;Ҥm���K�� �l�8�t.$O�l6o��cb����*0ϥɩם�z
�˜�=z�L:s��M��C^�X)�-�%�f%�ܴs�|�9=�7&�vQo^W#dڸk�i>EO�\��	�.���6�w��;��B�oċ訯�<���:��?t���h���x�&�!0�,�΂u�Y�3ˡf	�󄟱S{��с�#�/�wE�do�TܯaOV�q�5��%4�U�"�2E�E�����y�L�;�D�J������y��B��j�L=��p�ٮKjV6|��
[�3b������4�Y�Q����V �O�J43K�a��*�T��ml:S��f%�1o`*�,)��s�U3��RY�WȔ<ĩӯٕ��qQ�z���u*o���#T�s.hs��b�^�%׍�T,U
^x�6��3��T�������얨��W�Q�w�觥h�<��w�I��0Ӻ���1�����m�rT�g�5!�v����8n爷�s[}�����ϴzjo�Jf�=�6�����ի���?����z'�%����ZZ��-=N��˷�E���&P�8����J��B׺����m� 7�9���0���#-��惯E��oF�;(�c�c~��Ur ����#�
)��2+g�+���她co�7ѶXl&��ߦ.���&�t�U^�K�C�[|4��3�/���\�}S���������
�˚2�x�5�x�ߊ{l,+�=@_3I�Nj�����>� �1��_L*a'����uoO9J�Wia@��
�i�汝�<���͉���W���xd�D&i�`�DY�.��PG����F�Җ��2�'$ѵM�h��~E�z��9�������y响�T����m�^�p�f~�|�40�4��:��}�Z(�?�y_��&�*��v���Ӕ5��e��{���߬7�V�Ą�Ż�Z���⏚�z��j���Y~A��jA_�7b�$4L����D�e��4�8[aڬy��4�g>Z�Y(A��~��-1´ǩ��ޤ�8^�}��q��nb�&�D����I�PL��B7�F�16��7� A{F.��y(;i:��,�H!a.�5 �&U�M�tI����-�lv�f���`��*5l+32MXp|܆����q��P8ڼb���I�4){��Z@3&��?�
gR��҈r`;�^�#�1sK���S=e��2��l������ �z&�E0E]dd�;J��� U�d� :B�!��K��l�x�j����>��\�
��ՠ����L��HG�:��b�a:����f��("��]X۫Ĝ��O[�_�g(�AF��@<��QF�!�[�I�4?���������z�����������|=���"�ٞ��C�7��Z�&��8��Ї)BW�V)�J�ID�kƛ0|�����å�3ɹ�r�o�Q���9?�.+��`���9�6&��M��M���D���z%�*, ���+��5骎k�+q;Y.&cL9�ߚu}n����*A�cJI�9_��%?�;-�F�AjFR&��o����͜g��vUzkڃa+�:����pz&���L
PwAW��W���ؑd^��
k7ƒ������{�H\�]T�%]X�����XXu|�j-����a��b��37SuGybݥ3�܅��G��g �����\nP ����h�Z�����L�Tm��Lf����S`h!��ܻF��e�Qa����6r��O�H"!�Ֆc�_ڒ��Yy9�l�$�FCB&s��8#���`GM��&t��9�H֘`���c76��E�_ſ:��D�%mN���[ə��t�D@���`�	�"�=h%-��nN�f���s7�f�WC�M��jc�?l���]���}T���7�������2�ђƾX\Q�3���O
��!��TO�Z��
�F�R�m�j��n��KX_��%��rW�nTy�,u�����P���X\����g�O���ޮy����.��ߟ�z�M<�J2ZY l}>n��L&����')IZ���l��#eD�e�-j�7m.n(��|�E��#fț�Y.L��%�E�	���C��.ɉ�N�9�q���6���z�}[5��^�G�N�L� h�8	=�ƿ?�H�>�g�袽k<�@z�aL��N���x�Ҷ/�W\BǇ�����X'.���x��>P��:�]-�<�M�2��檳��C-'�ͮ���2���W|00����3(D�o괔�S��C�*&�_���-8�
tuo��K��jc�I��NZ��,}r�O1Bߖ�,A���.c[��.Ű�V���������&�v6����]������Zڼ�t$�-9��ߦ���q+r~_���s�����O.��@�ʌ�ER�ޤ�;����7}{g�IJL��T���c$,OK�?��d`�OĸH��vR���4�80�m�Qz#�Ff��U�)��?����f�I$��'������_�R�/��ύ�[��u���'�ʄɱѿ_lW�/�:_>LC��MҖ�f�ج�Ŕ��t��'��4�^I����ӋE�it�W�fh~�-eq�I��ə�5)bj��>��DeK���'{Z��GAZ
&�,��d����خ�:���q[����@�_Br�C���.q�)۔R���>�Z�c�Q �C\�o���Ξ�4����5x׈�yԵ����8_�)�e�����7YGY��,��V��C�"�Q�����pA���#�`QW����~�̀��<�-?����Eƹv��d�d�?� ��>+��'�n�n;8��C����6�H.���4o�9�҂���	�d�'�Z]��%�?�I_�S�X0lr>�fg�V���s�:��E�R��Mb� ��a�;p�^.�46����LV�q�R*�0�@ʦ�w�+_EU<+��T0�O�ԊޠL����,'8}y�~��'.<`��BG�I(E(���_��<�#��,��Z�a�����\���'������x���+�<������%�6��Kg��H� �z�zl��B{â���S:��p�%�<%�1*ԡ,xYZ�O����.P��1w\~eX�?si�N��,k��x��5f��?�ࢅ�^]䧙�P'M<��p��{�Q�Dy m��,����J`������g���H-R�5r�a���9��ed��5������,B�N�y=�j=x�J���8�i)�M���Ձ�I��}�ˣo�kl��v$ET�u�p�����3�(��JC@����#ooz}�B4����0���kz)�����?�7��)�ccBC���p��?rS�[��8*ԻR�-�}JV4S�:��s��|:��ۥ�S�v��s}�
�^??n��j���rx}�,\ws��|6�JN�_�L�r-ڻ�|	�M�BLJ]�Q�uA����^�����^Fu������a���ֆǇ_$kb�F��i�x�� ė��R���l��jB_�r�ٖ���/W����'�2n��]��:m��a�P�3��j�r�0_�K�Ÿ0��H�3�;�y�hlY{� ��==�>��)���������ל^�]j*c,����(�֫�#�����q�BJ�=��_8��3ޮ�L���m'5��������mP��v='T�nA�fv;���f�Aφ?�Ɯ���^+��b��"�>c��Y�PYV N��`��Ȩ�� ���S=�d���
,��xە�����5{�/���欎X�k�d���=+Z��u-
b�V�>���j�]�b�����-�2��4���R=�Č��~ϡ��m��g�w���*4�k�Nlb~�����o�!��2�YG,qSi@ƨe�(X��G{��lSih0z��3O��{�r�s�E����X:3���+Ȥ�n�&��Y�)��b�G=;�~�nL�T��!{s����u���R�������`���?O=��w�2�!g��*��E>�\��k�F�G^2��aD̓h�Y�*�b��O\O�FV�3_槄7��%�x@�w�[���%V��QSV#���C/���x�B�Oޗ�ۖvO�6��=�ҲgBq�v��ԡ��z�v��֯�LH�L��"�գ��As�9�YA%�〦Z�}ǵ���ͅO��5;�0�a�e��Ѻ������ӆU?�c2r�<�H����+E�2��vo
,}��X�͓�)$F�9�T7w,8��?�E-*nV0V}��Ŧ]a$�hye?����+��N��"������1Ya*hBc��V�7ι�7T���}Z¤ї����d*m*�F"0��������ژ��)�S#W��G낆�'��W����RmO
����k��YĞ����\���r0�k7����?���d"���S�؇��T��X�+S��kkL��h��Dn��"B����L�fV���[��-�kʱ6%��T���]g��0�a���%݋��d��pTYt���^D�N��P�ceS�Q�j�4�W�� �Ö��f��h.�%�ov�^�ߘ�`b!Kޕǥt��_ H$�����[Zv|��"R&�ޚ�1O���N�����llrИ�Q�'Gd�ʑ}�A��	�7 M]����Z���F�S�5͡3%Sd�Z������(:��Ǯ�)�:�S��e���$YuF�� ��C�}VS����E�Dحw�d^��!)�hȪ���M)޾r�4X�5�	���(z�����e����_��
��K�T�K��?��8k�3Z�">g�\{���*x�n�E�e�q���c�ki����拵�~�u���O��w���`�W�X���:xM�	�ە��˹Xd�*�d����tjYw�)�"8@��AJ�SD���8�ⱖ|5���X0��YH��n���0�S����X�� ��]�i�)�E��f.���~�0�@G��l:п�E���rX���������r��!����n���4l�)M�#eq:����;C�	�j5���,o�zF�q��c�v����%O��FQ��i�і	O9�+�'Vw�r�,�;$��Mn٦�X3r�����!g-(�C�g�X#]�� �(j/ir��*B,an7[g�gJ�&�ϫ*���{��/;�WdğfvH�R�<�:BZ�������Fc�I)W� ���N���cg@[y�*G������Cm��w>��K ��j=AK1^��+C���ر�y� @��v2]�N|9��@�1��;�D6��jq�,$�{L�faF�M
�L�������RR#��s�?Z,A��O��I,%�t3��]�g��ׁ'��w�Gp	t�<��-�[����2e���F���p0�S����ȁ�l��Ȍ�T<9~±<d �S���F!]��PYC��:W�s	�f�n)�#<�N��+�}jVc{�Cڿuق�(��zޑ ���lT�(���i�8��\>���|����!����2׊���W����Y��5��y�)t&���ut�L)?Q�� ��{>\o��۰�N���@����d����Mz�ρ�#ؒq A K"�Vͱd���[�J-P#bd��ɇzD���eU��"���G�7e��-�fc��Ƙ
.S���`,�C�"ZAs�ytJ-��S���Ι�d�I��+[�q��]�?5���ђu>�TV�Z0XP��e'�р�A�J]>x�EcM���`�b@�vhiE"��79��ڪ(�	�>�>q��7�w㥔�	��a_�D�JeP����py�B����j�2^��`�9����~�
4<�e�7�����2� @���&����9`#�#��u�s'����^���ǘ:Y�gy�;��`NTz�/�)]\i,mY��ѽ�����h�w~�d��t�W=����/�E#��$��ڝ���m��%V���R~�<<�	��sS"�v�`D׽��7��WBx�T}��&�p�Iv��Cgٴwܕ�?�G�Ȓ��0-ynP�U0rS�m,�-���J��>��gB`ʴf��P��;��ӮZ֖�"Or^P�T ���抢�ֲ%�OI Z��9±�TA��	���"N��F��A��o]�R��
3d/�規V��OA���,�S����U�,��>g����.�w��!j�^96Xc �o�Жp�����p�Ԛ[��P+.^%���Jɮ�e�Ϻ�햾qÍ��*fy��M�Ӌ�9�U6.���f�L�
Pj��>�[�d=��m�<���!�6f���F��ϣ���Fx䷰�%r�����-��0X+������ k����� ss�5z��N�o�䯗�����N�<�c�~��1}Gy��Kц���ӄ��/��i�|ޫC�C_���t�n�`nL����Ϗ$Ѱy^Ҋ����jR��5:[�:A��VKʙO%�h�M�K���rƁ��ῤ
�55�2��u��l]��I�g	�P�/�#�{�ᦳV/'QE"���o�I�CN?����������j-��;6�A	SF�)pb`�z���y�C9��ʟ��Z-��:�:�z���9.t:ͥ����j|�.أ�]Wb�6��F�*���ձ����Ī*g�_Q�Ss���f�:�3~g��L�|���e�m��7~��O����=����n�BD#�e�^J:6%9�3��hj1��a*�Hh�Q�q��ā�J�7:yG7?X	�����ˢ�ñ��'�s1�Db�_^�F+G���S�mDF��r�JI]?��F?�����{c�j��s�k���@��`P��#s�F[����Hv%�E�L3 �Z���z<�.��+�Gj�G���$Vx��TZɽ�1�&r	�d��x���F�uuf��%H�L D@x����*.������Qs�KO�E�Z�T���}�A�c�h��P=b����lޟ:�h�pA����9�������s�1Q
��\a~:UZu�Y�Trx�E���4�-4aTzRp@2��k��S��iX?�6XF�4(��>!��uh[�����=��qU�U[��S���ԣ;�/�o	�W�>U��S��o`�5a�މ�B6e�i+t�� �q�hl���ӫ�ɣmd���M|��5u� ���l��˹�s��]򹡓����"��a�#Y�z�4m�s!jݫ
Ĥ�q�oR��TJऀe�W����$M݀�ݳ�e!�t����8R�|�v�
r����;�g����>���G�]a�jaP�� ���EEBp� +[���L���t��VnYXmN,���h�t���3Y�ɘ���dC��HBJ���V�9+c7��?�aZ����N��(�$yfȨ�����'��z��x8�D,�J�k��q�8�������K2�x]���y�6,sja�󠏙.��.R��'�O�3	s��#�v�%8��ɶ������`������$�Y�D����G��gs(�AS�d3d��n��^;��� ��<L�lyi`2s���ȅ��ӯ|�����A�b��2A<��G"�:	��p#��]��`�L�.��+s�w����+0f���;KYb��u��K�<�jL�a;dG%WSh�OlO�I�t�u��w��meg_3d�W��ĐX��$}H",�o�I���ws�@�7Vv�^Rˁ=Y�z��䙩��%e�~���$T���O��[]�US>�ޖ�
���b������f|S��W~M|Y��_�dkd
�p��*p�C%ʠ�h$�~p\�ˤ���d33����Y����C�=H:������B=@�A줜�͕�r<zY0�o�*��+D�TAvK��򨣬z�2���a�%���Ly�x��G�H`�-��R���AQ+@���W��/��n���+D����ʊ� TE���yw��b�������I������f��m���F�u����֢�H�149T��]q }���7�[����k_sS<f����*��a+(�����9	��2ǂj撢���";� :���k�5�:�{<J�8�/�h:ny���4Pר )9��e|b����ׄ��$
'�+Ԓ��ֳ�g�����"Y�i�U믶������ol:��pTRF�j��j���1�g�;���T�g�����xٴE�9�`���-"ۊb�t��[������2�����$�xZ��~u�P*4����D_@kpu�Ml4���K�iC���m[�Y������A���:��­_ǲOe��k`(p9'y��~
k�L��9�l����/A����"	�\��&�4�N��o����v��4x�Ѯ1�S�x!�W:������7@�E��ɓf��.�����zKT���/���\�䟯Ə���	(=��0�A�qC(���[űV2N��M�/Y�7�E@����GJ���
���nn�(Xv���س�Si�΅\ܞ�o��W�:�B���V�\1,#y��i�x�����=�ȎØ`Gl1M�����y���Й�E�<7R]^�fӝ��gBM�M�,tA�-�p|�����7�<�����#I��_W�j�#��J��)�:hy��*�ij����MS���_&��Y&]F�V���n��}��f)iTҰi�5Y��+l<U�P�(K!��G[����������fe
��f��OP��Fs���Xb9����x�k��.�\���NR	w-�x���ދ��?�D#���扽�w����7�/oGFc�.0{�([&|3���X�����'�����M�����(��Ϋ��_�ێ�(�,CS��*2�>�^6/�P�-�����#���ز �z�{�dj<��5�~~k:2��V�K_A�C��"��@����q�X
��P�4j:�@�ni~�����ȹW��	1�4)k/�*���㊞X��5����|�H}���|�����%����ى�d5=2��`29#l^2�!̽����Au��͈];A�u3��fSަ��r(w�*ewm�桲��_�_##�i.S�_�`z��=%��3�i�`I&[+VU��f(M%���V�eX�f���cr��(�(0\�Ц��j�9�cD���m�� �s�s�/� ��Z���]ʠNk
]���*4F�cb�b�����P�ǐ����pK4�,��| �%��5.]-��~�A��I���=KL5_�ڑ�~	Q�=�ݾ��TM��:�|�k��S�>��b`D�5�F���"��s�9ԍ`^�W�3x=�cg1$?�p�d��ʦ����O�R�ﻗ��my:ݟ��r���4����hU>����ٙ��&���ظ��a�lyDbGi��H`��L�B��s{xf ���/��~&>p�rB�l��;жMw����a�.��������V��k�NT�p�]3P������ꟼ����o��D�Q8�0�c��EO���M��A�(�#�SB�o���I\��������X5\�j}L���܎Ƴ�y�����E��=�qQ�\�?�Ϯmc	5�+t�2x�c�Sr��1S�l�P�l�+�.��ܶțG��B�%�ѦE��4-M,��ȕL��;�;1�.RN�#s�._�5���>O�;A�܎�;2#\ްxT��-�ڭ�}(�#�h��y�@�l�:#����@���
 ��;��X�?妥v��Ľ��&	ec��ҳ}�C��w�S�h��>	j�dx�L��cV�8�new��idW�Z�f�y�C�(��? *NnJJ�
Z�wrW���.a��Q�s����:M�!FQ[=�p����<S�9�,��U_7!��-Z/�7�����78�?X�J�ǥ��ְ�=�o���^�a5�֐�1�U�et��~hÀ�O�ta�G�l���jd�+��
�����(h���])󳗓�č�Б;Ќ��)2��9���d�G� 
��շ�vY��+���t���ro�]�#����W�[�d��Օ�c-(s��ߧ�loKޡ{U�K��#M1���axqN/Mg��ꨍ��(�Kc�!�Z�9s�,"6:����L����aԝ^�7�&5e������܉��}e,>�&7�!:W������S�6�RjZE�˾��-mf�r�KCw��&�\gQ�b��/!�w23��3�c���:�7O�y?E�Ђ�#�'�.�U3X-�sUamvܔ���6?T�R�o2P�q�_݀x�����"}�"�#�$<M���-�.\���y`s�gb@��"f�O��@�L9���f�+��ATxh�.����%*]��QjK���D�iQm-Qm����R@Xn�����2��H��,��D��C��t�a`B?AI��@3���Ył�u �0�P�]�d�Ž �\O48�֚܃Ǌ�
�9es�eJ5��j���Pلɢ���ҴRd��Ko�=��&�FQ Oٙt�'�C�x�Z�6���ew�/BToD̀���ޜ7��Ir{ė�ꭍ&Q6BN���}C��6hI�@��q���5���U