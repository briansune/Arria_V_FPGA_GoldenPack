��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)���vG4��NB*v�^%��_�rG�v�2�H!�W��m�e��
�H��2������6:ǘ�>Moy�ձ5Ċ���������U����3-�lP�FQݪ�2�fU�B�QZ�.�Q�'��2Ɏ�im����I=҅���6�i��mMv�����K���3"�(FU�_~�fW��VlִJ������6.� 2�B����9�T�H�� �ä� �<K�˗C:�b��u���W�ǉ�Ɩ�8KO�����4X�ְZk�_�2����J��� }��=�f|%H���3Oh*ң�qe5B�{���s��!��Lk���""� �
���["�Y~�)\2k�cvJQ8p��&'p��[.P%wk����//�?=�hpǿ�5��]�x�Bޜ���r�VD�.�1/��y����ۣ�|� Hk7� �����U$=!b3ByC�S�i�_H2'��!���F0����3�d�(w*�vLX���-v��`j�w��`8qP��ݑ|G��d���ԫה7 �k{v�X��=�^ �q)�Tk#�1o��O;�D#^*"���W��n(�B5XSy}K�F���mlE��;n���#���v8�{�1�k>��Ѩ0��\�wC�[t�:���/H '��Q�\W���M�r!�P�CHOH/1o������)�O������:͎�t7wkt���[<R3C�赻� p��I���6$p�����Y��^*�R|����-��q�QS���n�T1i��,Gnȑ�G1H��]�5�z�#$�C6�K�*�UPx��E�m�����ɞs�o��!�{��r�W�c���]Զ@��,X'f�b�K���TB��5��-�-��`�� y�� !"����w���y��2݃���|��/zp��u���s�ƶy���~)��k+���I���,�-qJA[�D6�����уe�1�old�\�4W]J�0���(Ɯ �%���8DX�!�xDF�Kbi�W�ᒋ���+���1� ���N ˥��ֵ�-�9+x�ۛ�/h�j�o�@�+ի��%bF����A��q�ӎ�yrJv�H�ܠ�\?�Be���
�z��S��J�|�'���8����'k�]�-H��f@]CA#s�橶�H��FsB�bٯyM�1P	��o��X۞(>h� G����G�#�l��4��qy�RGAu�c�����wZ�M����IB·p&ҷ��Ȇ98��@Ae��4����,��3XmT��D%���E��y7�9*TZ�i��!n��b���p1��3I�\���n�����?�Ӛ�S����'�.�tc��Z��'C�o� F��z��O6��ڱ�<�]^�|�onaBz�Cš���I|�#pAU�9N��DV�P����f[���'�(0��Yu�N�$�{�=��~��3l���b�R���͍�5�>R���{x��� �^ے��4���R	�
	�ܕH1��_-�E��K��=�ĕ��=���7��š	蠸�q�(��Uo��u�(v��e�dᅠh?3T�j�+�㯅��y�y��e��]�$��Z�--��/@��z	����6��h$��J�"u~u���]�l��1p ���){�c�%��^��A��&���v<+�����Ǒ?_N.�����eRh�@�p�O�f�����~L�&f��P�A˶SK�!��i<8��?o��ڒ#)��)u��ely��-�p�,ce��P��I.�C�����)���q�����+�j�~��ל
?C�e���e�?x>4IaCS:�����8#D@�i��y]����3Hl�N�sGC��]����3.��0��Μ&Q���W����1�%+����r&w6q��GS@�`�5&�6��H��-��l�ّ��d	��l�n�� �L���M�N�K6�&�����`�o�h0ۉicY��d��2�$OFu��������Ұ�!v%g�9S�d�e���;a�>��2##�r�����r.O�ւ�b>�'�!��PL����5	�8���K��Q4�&� a�;�,�I�呂��nk�Ⱥ�y`�P=��I˸R�ߪuL/�
���㠂�J�N��1$�*��Da�c���͋�F �2m:�!u(�N���D�������S䵖�ى"/܂O{��zpM�Jg>��F��O��b��F�i���e$ŕ��O1	�f"��p����-��~���OU�9�*���}V�)��ם0�9F�-���E���h ����g�r΋G9l}��<z��zr���� Y��(l��-0�����n{�0� M��|m���Y���M1��!�/��N��~)��=�7��*X�Q���_P5W��Ez�#���^=U�b�E�Ŏ/�ǐ�o���
єCJ�3^�p����բ�;W'�z�i�'5�~�ܾ���\�4D��ԛ���>��bX;/F�l�%��rp|%T��xm?��rA���2h�$o�h>�.��&���\ه'TOk��e�6&Lo⑟d�Y��H���C������I�f�l�}��a�>�+�ڡ�~hZ�-���'���N�̜��/{4��WQ���-o��	-2�(�����f��
Z�_�f�"�
��l��}�]�q_�w���&���4������Y���Wf˝�~���lx��8��9�ΐ��}<������̉�c�~�3����J�-X���T{X���ﻰ��b��ɹ�6�?�8�Æ�`5�uT�Բ	���V65��a˫qe�U��w�<��\��+ Q~|�O`��\�Q����+�65����h���:��e�6�*��Î_�c-�Ï��D�g���0��Z=�1s�]<�����1��o�b%�����VM��+f_���\1!�K�e9+�\����\�%1:�^s(]�L9ih��+�j�N���%5즑�>�Bu0u�d��b�L]��U�
�)���?�<��.*�/���wU��*�E�>�4X�t���]�cl� T�F�1
��ƿ8�p�f��u ���Mn�>��ֲf^-���C�,���7ͰR�w�Xe��Oq�Ō�x����AF�P�Է:�4߻!�Y��g_�)Ka��3��X�p�~Q�=���bY�~?i,�tA���d�W�AK����T�O��E9D�[�\���ߢ�u(��q�)X��/�����O4�`����P'o|��۩̟`ө^1��t���P@j��W�<�����r�E���&n2��:eB�G�X7."c��uRp�s�J+i��!�ɇ���)kH�%4�/F)RF����v��<�jvǹ���̭,�|ތ������ ���q�óc�uc��;n� &^��d���������[j�����F8�8Ð�pTI�Zj�����8p�a���R�Ӻw��_�F�5)9u�|��W��l�����*6�����XG���&t_n�Ǡ�x0�Y]�A|v)EKn��=����!�F����E���'��R��7��d<x�]@'e�Y.�kxܮ��)j9�ʗJ�k �x��ͬȧ�e?����j^������휪��e�"%����&�'G?�Mx3�`~�~�"�o�}4�-�7�������9�$i��S!�
��H���S����WiH@7�P5�Zx�b�H�ɟ�7+�A�w�B�y^+�t,f^�ԏI���捸��FH�a�4ff<p]�����i�L��2�㝬3�'V�+�/����Ґ�jj�&��Ъ��զ{��|�)�6�u�+�=��1=�Q��d��8�
_�'�x[#ᶤv�"�����,��.��O����.>���S�D,r��g�+��X�Pj���1T�;x����Y���)�� �Uq�x7}�1��5�lG�㧅�F���V����IP������(a�1lBƳ��[L��"+m*f[ڇmǧ7�m�,�K��R�9�C���ѕ��B�+�Z��LL�`�wK�W]H�i��`*�L�WZ��_^ ����f}�(/�A{:��u���E�OÇ�8�R��c�)6���^e1~�d�"с�"픉X��kqyɶ�r��uB "O�Q�e9|y�r$_s�5�K߶�)�t�z��$���-C����o��v0����r}��xu���M��Y'9�H��s˜fzv.:n�A���<�\ǟ[�k�ZK��ON�IZ6	e�`�A�LE�HM��܎��¡����f�}�D��
��j��Ϭ\H�F�-����NKp��dex�N�^߮�<_�[f�ضn�J���#ꈎ��7���T��5Q0c1���r���a%�Zyz��l������6�l,�u�">�����U��e2�g���6��Ov�{ʆo��L:9J���>�8Ŏ��Nf�*-�h�Eċb'F��$��r�MI�ŝ!��T�т,)��4�����)w�Շ6�bx�x���i�����T?߈�(��`�^�K�gm�od�^:9&��<��<����MeE���D�ry�!F|&龖<l�i2�t�8��\�=��5��N��ev`�U��h�.!)����#^��eװM�I��#E�c+x���`�&�+,v��[s��6�@Y���Ļ隡j�uO �C�YJ��&P��i��Գ�tB��1 /8N�/�������J�J�l��uhT*}�]i�Q�f���'Rn�>"d��"�o���Xҋ͞x��m���$�؈�?��2^<G�}G7�ۯ�N�3z��-l�A$��z����Õ����P-Fn�%��-XG!O��S/�\<dc�g�U�+�i��~��A|#��8��S]���>7�	Z�F��ǯ�m�h!��9C1�b����dܛ��S��_��vm5\�*�!��^\ᰅ�������$+7�<p���@�Y�c���2�_^[�7�1-�MYk��Tm��T^.��5�;ȑ�e���17z�8W�{�����&+cd�W!d=��+�	v�We)�N�nN�%�]�\���4������~U�g�4+��h����sA5�ejw�q���B�Z��U�ަ��h�t�l��(��J�j
�����,�1���)�P-���>�2�_P"�[:� 
� �aH��nk��FG �f�g������/؀dO���|r��s��7�(KXV�c�2ێ`��V��i�z��u*Lf��3PbK3}Rk�U��^���P"
H��s_Ђ�q��%0v!�$��y�UCV�p>4{Ǯ�a�Q����Q�v�u($��_�P/8J9 ��HH�D��K��45�{���jqw�>�D�Wx;N�!SP_�(ˢ�l��w�q�?4�:½k���Br�
��qj�þ�鿀���m�% ����{3B���DL�H���_M��.s]�9{�-x��y'���
��lf)$�@����(37C����ޞ�[�1�B�d��Y���m���޲(����].�%�̗Ƭ��� ��AY���tZ
�$��m&+)u��]��/�ԨI ޳��ɸ��_FKB��ފgs^��@�1jg��w^D��x72���먛"R���kd~5���81F�9��Xta�����j�ür��pִ���%Ɍ���6�8�bQ��r���5^�]i�H�īt)��]�J88[YN�#D�F�@䅂bNu�r�'�������b��r�x;��v�~uA\"�:��̀
ŧ��#i���'����C�]�O �)Q#��	�~��������A�n(Kƙ�`z]��?�����bJ8��Kҁ���W��\Zm�I��(�>�kv�$oÕ?p5�+b��R>p$�$t�|j;���@��lX��J&�%$fއ׆����� ���U�{.��/��p���Z
�>��)WS��$6nuu�|	g��u6�U#.��VU�~���پ&4+d:��e���P%����9�H�H2�wTӨ�`��v�8V�i~zT&G��D3���	��cV%��C�������X/���e��֡��!=Fi7�'	�_�����SB&7�P���Gz�xs������,%ܒ	J"��_�3#cl�e�+�g#F���#�v��Ҙ?;��Sx�L:n�.c,�n;*��W�"6���/��zԤY��VN���Л��s�^���9(~-yd&�x�7�u,f kK������p��*2n�cTi��8Vrv��/��θ�6��x�l�U��K�M�}�:@�嵓O��=���]q�_���?��`��y����\�m�P�Ӌ�4V�b��J�RU���=����m��fn�/��V
����I�CW��-����i�J��C
�C_�T)��B�8r�Q�!�8���9V��%
��v;�R��c������J~�'.�2����3Fq_�?%?L�Vr$���"fxl1�'�g ��:�#4)x�2�n�ո/�_#d�E��!�3�!`(�9�=���4���@�z��Ph탓�4�y�뭌v39��9)�����\�̙`��ڠ,;����V$��j��-e\���K��3��F���u�n��^a�0��q���%����u�n^�Ԭ�tX"��
^�=����t��ss9)/9�ŷ�ejne�N��/C7���`ܦ3�Fgə��`���]�e�zҤ/ɲ�� �� t/��/�3<�M48�tX�^��\E h�7f���w�P�0�'|�I&�U�-�1�?�n��c��_��-�9�F����rHB��������$H}=�Z`����/�Q��hA\���l�gG�����*>e���9M�f�m���\\����׸E�8Hn��	_V�Ҋ�o�ɜ5X0����. u�@=/C�@%U�f�����v�J%6�}��L���ZwD^M������Yw}��"�&z��v�Xѕx�c:�˓��T���TC�#�T��\"����`�0���D�7����Գ
S�A��*鱈)r�z~�b������ǁ�/Ǹ�(��H�x=���\[��is��O��w�n:���u���a�`\$ޑ}@ϸ����C�xMđ� k������|\C}~U�+�ܩ�M�A��<~ST3p���[���!cP�5\?�~$�A��0:\��osՄ�>����\�+&$�䆴�J��#�+�W����O�Ȁ2r��|�Z�r����hNo��))�,c��?rU��CAJ���U���R`V�NH�����\�rJ"Ǭ7�}-T�-��徜Ȅ��q��CL�{ՄN��s����A��9��������?�Y�#E�:q=f�9��	� �Ve�������-�	h���}On�#���� ���I�x���ykrC�U�������e;?�#�08t�6�q�N�I�ZV��Ne�( ������x忀�qՑ0��L�b-��n��۠5�����j�|	-ߴ���]�H{c�j�b�;�5��B?i�N�\��sn�>2�p�'�0B��s���7hэ�b�z*Ŏ�v['�)DZ ����s�v}Z|��|������"�Y�b��"I�� ���b���T��L�U
�4�" d�V��hʱ]�雇��*�@a#dB��~.m�I�u�-�W�d��n����?�zF��sW�Q����f��|���Ҫ}9�\��T��5t'a������sj+b�P5q��?� 1%������:���\WvL�"��Y�54�5�r�(o=�I�Zn\L�^$w;�TYF�8@]��f#�P���$��C�Ճ��J�r���<�2��s��;r����)�����+��+_��T*&^נ���?�;�4����4�#$���s�\4?�����n�̢�X�����:�|��U�:w�����_9�����{:�5�#}Z���bu=[��R�}gd�7�aXu���K8X��G����a�V��������s�cU"������ܺ�vn�������m�߫ԟΔ��^w��[��o�[�c�p��|r�.{�B�� =@�s�E�@�7��Ykj��D}�"*���>b=��4���9�m_��)«O�9���0�8��������o)Ӊ.���z�d�?�0��/��y���-�"t��L	m���	#ذ�>����r2y}��SdӠ=��0��"���	1��2�^c;O���zs��Y�����I�j�:4"�!���a9#�uO�����av  �p���[�{C��Q��W-n2˚a��"���Q,�I�H0�櫈��YV�k���Ke�|����\�"Z�"��ͫk�Us�����ca[��.\ڪz@�K#! �;�(��S��&_�3��MT[�-���L�<�_�9x�(��j> @�{�)H�*uTk6�"xFl�`AC<_/�b�q�9-�_���N��e��`��ΛJ�C2�ڣJ�FVc��K��"L�.�/g�����)P<��Y]��"��͠�zƻ8!�8z\�	�T,�G� c7�O`š��������g@
�/ ����T�3����6�O�G�	�T���(����\��uL����Y�G(��O�����c�-�|DZ��*���taaOio<4�(_E�$"��O�es$F�c;x�k��<,tP�܌���-)��ϛ ʥ-gL61}ZP�Z�#|�	 U��� �\�:r�Ü������������f�YV�_#��\��R"�aԺ<_N�)s�b+��<��1*��.p���E��T��N�"���W�A.XV"G¢t�%36���������AR�z���8���pI'��O]�R_ގ��g~@7OHt�y��Х}Q^�5�WabC�feRp��s���t%����S��.�+hF�����6h�25UEOi���P}��G�f��vA�gyd��9�ױ�e�i[��Wa|{]_���'��|򕱙KO�-�a.�~�4;�viG�PR�T���<m��zA�>�xl�!����P*AL�Fs��J��z�.y= �m�
n��k�#�x�o(��-�)�$����,D������|�.>��aܯ��n��&N5�>��m�2�j�:���,H���(]ߌ+vVP����OA��\l���	�o%�ՇH��ߜ�c&�⇓��8�t��k|3�A�`�L��G�ҭ���	D��c��� OpX������|w�����-����5p���3
/,h?�:���di�T����Ѩ��k���j ��3��#&gA����[���C�:�j�O,c^?}��lJfh:?kv�f�`�
��ˁ�YQ�ͮ�9�q�.M�	h�C3`���w� M|��1IA�t�^B3��pSk.�zt��.����Y��4�"�m�98Di��*��Y��p���7����1I���*L9*{���GV����4�bԟ7�j�\
in�Z��;�����U���dY�}^�:Ѿ��	��?Y�,�#�(�l��6G�|E��aT���șS�3�ið�>��u��9@9ۍ��U�Ak��_Ծi_�P�u�H+W��])�G�xg�����y�4r�l���GT��L�5؆m���u��t��d¼#.0����P���@/��� �^J��ż��3�;'@W�5(�$>���d��p�6[�1|�N=���K`[��fǦ]m�:�l� e�F��͵[fO�'��5rt�wF��Qy���(�zyU�l=eT�p�(Qf�#�XqS߿-��zN=yZH`��*UY�v]�Y�M�c%i��R��j��'k�j�gW��+G9q��5\�%���s4��	�5e=4y"K�}R��x��tV� 0��p�w+�T	�U.�5;�H�x�:���9�^+�Ɖ��g����{ ��v�E�-����%��Q��/t��l&T"�z�-fظ>�����E!A̘-��ٓғ>��}˯Ԃ�L�s�X�7�C�=�BlAQ/G�af1!�0���oИc�O#n*Y�&(Fx���v�����7&4Z8Py��\�Ttb�aG�m��3t[����'
4��b��Q=Z�	Mc�09�i`J$t��l}V�d���g�td���N��H
W�ǅ�dE��`M�5)��r��Bʁ��}Өǌ�D���ٺN��_� ���)@�0��5Q�E]��[Tq��6��ߖ㱎��e�������}�ˢ@��
�K�@�i���$�9F!b�m�n:��n~@�T&4���;�e�������1S�wt�R���f�O��*[�*A9��y��[sj�k3�m�Y��錗�:-!Yn�;�\��`�ð}'���J��ڞE�t{���9��S��B���w��ܾ��T�A3�OAv������L$� �V�v-�)ں)�פ*[�mޗ��88��a�.���U��A��<cYm�7AaQ�ϻ�����=���7J������T!�K;�����\(�Af��h���Qm'E���D�I�ٽscͳj�]o��	�}o���OĒ~��J�ې��o�����B�����3:�����fS�}$�v��Ȕp�JJxiO�߀������Pp���961[B~�rI�M!uc����h8����X�23t�e:�f*� ���H��3Va'�&N��l�t�V!1Xg�le0Q�Ѩ	I���*�T^�PY8_���B"B�GEV;1���UGZtn�"�>F���#��֯!�:@�,�}�	���K���/��_W1qo���������֋�<
�)v}.���?��z%1������A)=�t��a���yD�c�Ti+**i� ��h�c��b|�o����s,�@�4w�%^i��*Ű!jX��nD.�j��k�?��z����
����^nr��>��ꈝewk%70d��&g'�D�i��`�)��x�hyt��m��*G���G��Ko\	}�����o����	>����ejH8��}d�G`�{�Ϫ�?�*м��F%�(#W�R�Ԕ{�r���/F�5W�	������'H�eL�9�X�ۏ�7���XÑ�6B�$I��Q�}�� �i�0�;u�:pe}���?��2�Y<.�J'	)��Un�D8h}`�\�����\�X�m���r�r_&K�ף�h}���B ^wK�mhZ�'�;��S��P�LL�v�� fx�f�/^�,c��kQE>ba�$������m�,��md!#��$U� ��cŝ�KI�}���'���n7�&������u�&�O��o��Tfl^IZ)j�h^ss,4{��G�%�'9}�����<gA
�e�CF�S�]uB[�aH�Ffc�S��a���p�i%,o�V���,�u���{*&Z�F���Jg>��Y#�K�
�^İ}�f`����F��ߖ����Ua�oI;�\ W�/,�ߐ�nu���]�D��%U��b24V�pw�w�;�6P�N
)����ܷ�z�צ2�� x��Ɯۻ������i4 ��Q���d6��3Z�'�E�a �)R� �5Y19ݔZ�<��z����Ā,A�CC�����C}�;�-��$.iu���5�yګ@�.L��@�{��C^�Dv�)}��k�.�c�g���$�B�S��c�'4#B�߬�=�8t�ͻ�>��dF���*��`�����f�~��E��F3k��E� ��.�7��ߨ���u<���d��W�:���<�6s7\��D�Df�c�cK����\j�� �XI_A���b�3_pߓ�<�켛�d�o: 3�1p�A :�m��H8#���l�D�}���~j+� ʱ�pc��nu][�8xL��S���T��C�*]�x��zd �d9�_Y���>L��!��Y0U��Π�rTZ�Ԝup�R�>A��G���5O�u�m�WZ��T��μy,A�,�c+\;pCtx�|3�E:�:E��Q{2�X�D�!�i;��e�Dc�^wͦ��U�s @q�d�� �/!�B ���}�\�2nցiD��cm��,��6��bw��@D1e�)�ﲆI�k9�g �r"�Z��u�W��a[���L�$tV|^?�qEtܻ�tFs��d64g��z��!�w4��>G�p�����U�٨z[�\�w�@pPW^߉}2�;��t��G�����)�b��YOZ�Wx%�w�kL��?�-��j�����-���bq#��<h���3��{�rz3����t"--�iu�JMɅ]�dg���J����o�t-%�8�����u��c]D�)UD4��W�����u1�xY�B�0��ҩ�m��!��A�m{�f~�E$��?Mi+mxI���z]�o��K�d,Wbښj�C���)���������@��/g!�]��ޗ<*����:3�FQSܺ�dSQy�;�����!��!�XD��@�z�ɍ�5�$~�� ����$mL'�"��9ݒQG�T�лz �ǽ�
�,L>��S�e�sp,1җ�,A�e��1��\'���Yy!`��'⠌F8��+�P�D5a�?Y�>�Ʝ���=�ʒA8�"����.�gl���q��K����$6�	��h���s)�9㲱!	��?Xg�3)F�%����dJI�ǡ��0-�Q����jsܗ���>L�����*��,g���^o�)�/-�s䭪��`��-퉌�"�(��M�G��=<�ۻ:�����x�c�����FA��{�,�6�%�mo�a�S�}�5���:�)f���jMRtF�k��.�v��E�Y�\�%��a0$�ű���O	��I�돈��Ք9p��d��W��$����_���2��{�d ����9:��2�Z��^���o�D�I��6h�;��?B/
�� xlQ���c�,�)�@fXm�Q헆�.G'Z�TzSއ��Ǧ��/̼U�W�쩗�>���b"�����s:gP3w��,��3K���u�a�����n���ކ���n����BRp]�h�4�wr�Q��f���� ��������8��>a�|��VuA��H��,[�'^���MK�{_YK?}��n���<�=�����=��Ήu��I���t���uGin���U:��֢�޶�$�k�����"��!�؁��CrɊ[�d#O��C��, m��_~«"q��)��ma�tPVi�l����:������ f��x�����[�m�����$a_1��� �Z�� z#��E)���þ�Lm��HM�_!��RÄ
9V�����w�* 1��]����n�-mA9�\�N�m���F���Oس~�) ��3�W��o�0�{Sِ��OV�x�<�L�t�X�TJyP�'�f��Qn�W7G�u>�b���)݃���|��]ǰ�-�~�dH�.7s#]�a�~]��V��
�%>����F2z�=�(��)��[�1�C�)nre�,#�c�&Aj@�SQ)������P���M�d�	���*P��*����`�I�~�ծ�5ܛ�g��� xc�BK2ޤЮ��Z����3O8��k(|�)~�4��������;�C�p&�`+�W�&�Y�V]�ک�f���E�	�K�}v�:��6+-���NϨ}�ib�TI�Nj����[�)Wȴ��؆�̩�>z���'�
洼������2����T�j��^���ޢKU��Q	���L&�6(S}����5q��J�Aا��Xp�=�PP���C~������B��� �zZK�i�Ŏ��u-�/%b����T�Q�Z�eJb��n�&�A&H�E���!-lK��ta����e(I���4�K��ި�7K��Y��;@z�6$�6���6R#	���8�96䃞�,�|�q=�2^�Ң�C��K��3���8QW��7���vb5n�lY�7y�O��FIߟݢ��I*������	}/e�w�xyR}�y_܈@V�$0����1���m����Y��K6y[،4���K�ظ,@�;����=fP2��
U6]b�4���O�A2�l�!�XD�T"<V���2W�0�)_�
�cB�Z����Y�M��#�K=�/�b���;��f��|%IAJ��~����r8��F�kx�Rb��HNZ�E��p��GOa��'{ض��@�Q��Z`c�T�}��K��|�_C�?'#�x��N	l��;(��ȧ�6�1��֯���;N�G��0���P��ftn'�J��.t�z͘�H�4�i�'Qr�s�y���7��Q��:�xa�:�(ѣ��c�LfD
-#�O�u�آ;!��ks�uiw�>k`�Gu�`/���xIL5C𻴎V��@��w��Eq�wX+��2�L
XH{*^(W�"�N9�cʁ�:��%�cS���{q�c��ǿIk�#֭�t�d�ʹm����kqt
�4l�Pv�G��h��ut�̑z��z��]���4��%�.x@��o�Ԍ�7e�qp�T� �Y��E�I�^��4y^J�3�#��^(.�I������i���aVS����Q�9�o����7�,��tp:v��<����a@��Sx+��X��0�GeL�s�g�5�Q5E�;qsnF,9,	����on�*��WCO���}�������)/#���5	u0��M�gA{���Ps �e �8����ܜ�����`�>�k�xxgtn��R�W����o�;WDU�wL^$�S�-�s��l�	dX�'��HT�L0�:¡�e�[V;W�����g����Zs��7
y�w�ԥ[Yе�����<¾��X3��)�g��Ƚ�����DFv�:���������;t3E���P�j����I��	D?M��N���)	�āe�����)~��12������̙p(,�(Q�'4a#P�P�.�ŝO�r�|y16�I��L ��N��ۙL��qj���[��){�oH�N��~Ғ�[@�:��yZ���`�6{NY�Z�a#��|�"�8��7'`�|=�Qb������i��m�>�t�%����H���lF�vt��sx�#��������u\���P�[��g7�{�����yN�"Sb	p96�t�5&�U�T��L�I	HD��kJ����GՍ��JxpQ��z1L��9>Α�G��r��A�d�|<h����	'>��+�抹}|�
������$l�p3,����t^�O��Svt{d;���(�.v+B��ϔ��y��D�Tm��`0��'O1ʏ���pm��f��b|d�=���6��I�q�Po��nq8E\?
�J�L����F��=bke&���^ܝd�@��h`� �q���?���V��S��R>�(��Is o�#��|xԢ����Hyr�1�i#���E�I�!Q�����}��m�	�e����������-5���l�X��5"uҘ�sTݫ5�q���Iʗ�M�^q$%����㽮-�߬'�A�ʢ�u��_2���o) ���=m���xwm^�x�����O�U��c�jeh������E*���(.��שđ�1�h�4UN{�����re�
��Z2�,NMd�t�������]��Y�ksN(��=�TN��$��`�m(�h�9D]��.wi��)�v�h�г)Y�ӷ���T�j�R���CBU�}�ʳ쀊
C$F��FQ�տ�����k�R�/p��ݛN6{�6F�~��-RY,�ozM��(TI�_)�$`9�ʷFx���K��"aπ�C�����v
�e��o7�0>u�-Cp��i"��if*�]���B��qs]��2l�5����U.�6u"=o�d�s�~��{39&]��#�9�[r��^�O��]֒L EL���y.��%������kO��pR4���A���`�G`d����䏳H�/���d8��nt��M�V[K_a�Jw�����Zх�ܢ�9}�-EuQDN��	,��?h�����X���m�S� �����+3;-����}T]f�˅�2=����8�oƈ��_TM8�k��e'd���iVh7��21�kk�7�?�$�MO}�X��b�(���B�	� ��`�H\|�P��(��J-j�LC/1�R��]�k�:��	��[8��L4~@�bx��2er������,�J�:	U.8��U���+ొus��(�Uz��0��	�R�dr;��:��uhB�Q{���i��tx�i���XH<���ۦ�8�9����ǐ��y���6h�ej�0�GO��%���2m�uY��{6 B;s���:� �-G0~��8.�j�<��vc&����_0jq��b�?����RK�Y�3��~���H:��p8�g)`u~բ��Q�!$�X��%�<��*�&��{Μ��u%&���jו��龜�jZP1e�|v���I��xR}��z�O��]!�8���|��՚1�.�?˗}[Ǿ}+I<�R���+XZ^��������Wy�$�$2�J�y�}500YLr�<[@4(J�Qo䝕J5-�S�!p�âww��~߻>�x��F����`;Z��Za珱���غ�Oh��� v�=���<G��M���c��ӭN'\�v�����M��Y�h�Nâ�W	�{Z����o+��bS۱�n��Ӧ���5rZgP�y�+3�y��_Ȝ�ΈWE�c���E��W�h�ϧ0$�"΅���o�m|8��E�\����k���B�Q�u��Ȫ��3��eP�s7����9�h	��Lî2D#�:ٯA�q��AA��']���	WW���:��\3�U���N&�U�`�u�9�� 9�j-l>if+3��Z1��E`�9�Z��bB"�ڱ�x*�Ĭ�s���9�{4��uk�l�	�� ��b,�q?��4��T4���W��y
vj�0�>��o{@���@��fP���~��[4�(��~�S�5�N$g?��'��ZK�,vk���p�%?o��n�#f���*OcZG�I�X�+n�d��EXH9��lMI>I�r��S�z������A����'��6C ����X��q��!�d��P�oݞ� 0�>��!74�H��B �X����8@�G�|�`?6�rJ/D�aK��7�T�x$����Ж,;>�����h},6=��������(�8��``l	��KL�[Z�ʤ��]R�aY\�!���ݫ{�xl-yKQ���x��Og�a�~*���j�΃�l?���x���
F��ĥ��_�^Ft`ݽ��s��y���]^�P�tn�$�WҨ�S�Hb�i~W�Y����P�:3$�$O��it���8��.��Zf��� ������8K���&G�|Ǽ	���������q+�ˀ=��潸Rc�uOd�%D��Uw8�~�j�"8��c�3�� �͂*��àm�d�=ﳣ���2AU��Ӱ�R6ʗ���n�����~�/�#�ʃ��̀L��t��<���9���r�#ml\�K���| �����\w@�U>��dV���KS�s ߇����-�Ɲqf
��~���zd�K�w؂j����{�R���zހ����� [�\��S�_i1��"2�&���8����1�I�h	��_��{����v�9l'	���x�[���r��a��}��ބ(�Gխ^\�����v�4����t��4#��&ǎ��,��Y��J%I@~�E�!����u��ǑXAh'�X���EPX��y��Z~�.�[�I�~6�n�>.RoA�ћ@�Dx�f�1r��z=�l����4Z�4Z5�q�9�Y����M�@�$���걋��*�G�A&�D�GZ�2�;�3����"��a�t��1]������5��D���GR��$���*�˓��{q8�{j��X�uG ��!�-zɠ�v��ѥ2�G*v6�Y�2w28F?bF5uKN�/�<�؛���Zl�&���~�6`��:��ަ�H���+f��rW��q�st�i�LP]���A�>�DD�u�"e�_���� V�q�Njn�k����.�
��דv6�F)��nfBt����]�d��Ì9D3���k���B富������to�}��(Am�ԫ0���Ѐ���o������eޣ�-Lpj����G�wb�M�1���y���
��+2�M�b g(������{́0�L�q=�hm�G��i�"Y4��?^��ٍ��Xo���[Y` ��K�������j�]�{�,��_n�����J̹W�����f��a�J�S����7�^v���Rx6PW�VK��7��-憇��B��������0�i���͞�����%22�h�=��Y���/�Vk�ORӫ\�k�c��N����U��HD��kKP�	�qJ2J��SE���?�B�֛���D���%��&m4���L�� LM4���;B��}��SQ�S�Ũ��l�G��}���b�ak�7���85"t���s,ŏ�5B�E��/C�@�=�*ug���&�B��7��wg��S$�qE"����R@ ���ۋr��@��ڤ!q��K�˟5)j��Q��q�B�x5O��/u69ddio��˻,������?"4�@�K:���.�C�񺧁��άx����h3V/|L�noQ!l�R�Ҕ�ﺱ�'���J���,���g���N��*���jy���[��h��*ұ��"*�1�E=XJ0h�q[�^��8^_��O��G�k�Ra��ܳw�z9�jRG��le�pbNrk�(�{ɡ`|�|bdm(��܇>��Vt�pX�WJ�eX|��7yz ��K��+�-��ѰU��M�=k��!k��p�;
%V�GC�1��]�h��M�����A�Q��N��瓆@Z�OQ��ͽhLE�ω~���,�|D�������mv����y�(���j�9���^_�X�8�+��R���4�"8< �$�.��?���ۂ/T��9:�Z�v>L�{M&B�x�t�Y ,n�?�)��/XlU\�-75E�Q�
H�UV��R_���pj�ɧF~����"U�����d7��[-`��R'I��z���XY��Lx�q0m��`������=m�v1\xAF�/�\`��J��P�њ���Ttzo�6��>���Fe�Fok�eI�z�Lp���U�T�>�Z�;ԓ������#7,�� �iΕ��P�}�.B�3�U��W�����?�b�E��J�HVZf�e�U]s۽\�w*��uaB)���r�t�̔dˑ>��sC������x��-<E�%���x&2LB����95Ib}�cF��uE�#�ǭ�U�FzgS]�t�I� 5X򚇄*H0b9I����'��@E�,ӷ3e����#=��g��)RQ�Z�L�E��]�u�pPr��KN�Q�al-;��m��U)}�&tv���vc�n;"at��,��ns�H��|j�C�Q�]���6T�q�HM:��Ѫ��$4���.��+�xǌ��t�c���}D��u#ƌq��� MU����T2m�1���.2��	�6�[��![� �jW%�U��d��Qa����ڹ�~@����c�ڙ�zH��� z�ql7.�����޺� ~f�|~_�8>�Lzy�JC��� �23�k"DV��o�%���O�Ӥz�Xx]�<<[.i���[����B��i-!鋵�>`I�\(먠�mD!i�e�4���L���<8�z��rg�Ws�ߧo$OP�����ӫ�,ƶ�:�<�{���.�H D�K�5��P K�>bT{g�74H'�Y�ĉM٘V+id-̜�YĲ� l��C6�q|��&;�+:�Y����0�8t���6봴�,�[x-/3=��,Sj}P|�/�f
ɖ4(I(��G����G��g`���	7�ѫ4�E��$��՚�݀�0�蟓v�7�"ˇ��-[羟��*u��5֘+Q�u��y�n||��U%�y��mt��=yf�2�\Z(�)��;���F�s9���'��V2�ח��H�l�1�����p_�E��KW�$tzt��a�-L��{u	V��3�x�"���d�p&�"
b�@�se�uM����m�31����Z�x�ܣgQ��+���!�1�[��7�kJ3�N�N���e��њ�`��X�Y�A��1Ȍ ?M���W�گY�q)��Ê�ө�*(��>)���'{����x���1�[n�a��F@�)�`���l��ү�|?_d�:�����	�֘t`(Q@��T��N�o�$k/��e�.�F��6ևg�QXr�)+�;]�z���ͬ�siu�s#џE\���An�U'H��$�
�1q&]&F|:;N��dr�gbM�{(ǔ`B��ŀ�3�4f�)ά����u�H��X3��Q; O�|In`��H�3?���B|\���U��ɪzK��8�PŔ���U͈q�S�os�z�9�@� ����0�T;������?�a�$�=�L]g>�,��ID�!y���y)Ů��G��k��%�2�I�G�gk#H}x�фo#�M��Ȓ-ܫF�J���]6�QZj ����d$��{��B���юZl���N��쪸��K� ��
!o��M��p�7��M�E�H��B�T`A�q�;©��Z�rgM�����8��1M�/��g�nQY|^�Í���!����q�-dD}H�B���>d���ʗ�����ιڡ��B�G�8b)E׮P�\��e
.�s���"P�#��G$��⵨��I��,�S��0�|�'z��P� }����ϝ@�k1`|"�,�����Ag��-|"����#$�e
n9��>}��3[w��
��z�����%��6n�[�ah�7���!�LC�=#XQ�Kʜ͔�D���2-Bu����o��a5�**C=�6�G$������WC~�����j�X
F���]�A�� ZΌ�X:}[j��0��뼫�V��P��c���/� �=o����:!�
.�pm�zh�Aa;~C�d��?="�IJL*�]���U���8�����Gt$��~�9�F�gGߵ�Tij�኿����¾^݈��͜x�J�?a��L]�ؓ�U��A�V�k��g�8�{���ӻ5sHo�:��;��N�,�hhc##�/�69Ѹ0Z0����l$��
�\�4î��N��,D�`�$�NS&lE@&G�� ;v�Kni����ϟ��Vu�`�����,��u�*���P�+O(��T���n�CGIR��8��ټ�~�}B��%j��:*	�B��7�����΂_�~>����7'�y�q8������!3�4�U5�wܦ�͓�˶W�����&�}:Ɵ@h�fՈ�b�n\��e���q�͜�?�+��>�:/��o ��:r���7)'�gJ	.v������s���n,�T�"^�&�!�K��΍
��cM��&ȝ5)�#����nှ�L_PH)����i�=K��
�����%�Ɖ��
��R��X���|�
���H[p\�RL��b���}���э��|)m�[�	9}�8!��*Ɯ(Te�La��y�$G��D�m��B��7�Bo_���ŵMB���[���zy��UNR�}�`���g�;�@��d'�c�U(�?"N�<�����4���7n�:JVn��ߑ��H����:�,OGe�7 H�\	��'Vp��M�����Y���Z���|�H����}K��]�D���|9��raO�.��쫺�o䏏���ih�V�s:�-�ʘ���AIw��_�[r�L��l���������r��������_�s��������m����� c�@��3<�q'e끞Y�G��UL���v�q�:IW�&�1-+q�$g��i���a���٤m���+J�����/\��*ۨR��;e�*!"�����i{LT��O�?|-�$/uyK.�������R��<G%��,amy�Ғ�Ys��{�C��n�#��01�<�BݬA�m��WP�����KĞs�C����P�Ɨ�
��ӓYǝ0��v�n�U�X�A��mzg�  )�4��������ތ�� �DHta〧�3��np;����r��_��W��a�3|��L��}�6$jr_��}jÓ����58��^bBu���<�8�񎁴�]����Jʆ��Ӱ
���UT7?g��A�r&ӻNÙ(v�@��<�C��I�vu�i�M{��I�G�\�TE�\���ZdX��T
���SL�9L���.���*k|�z��ǔ����]���s0c&�0�0A?�T�9�A�nˤ�>.t+�ҹ2�֬����u��?d	]{*����2��OsO�ʡ����@A?tv�[o����//�1�Ж���Y��$�[��W.9>�Fc�>�����#�^}�L[��k�?1۳��n&��c�#��O��G)|��Oxi�*�(\���;uH���Ⱦl�V�1��b����A~_yH^C��:A- ���V��܀cG�p�Dvr)�Ei-},�*=b��i$�r�:���?��`A�1'�z5^�ك��-�ʭ4KF��i�t�J
�lg.U�k%�P�,-~�	�������HK6�O�����>�^�K���da��"�Yϔ�������$	%�S��g=I���]�G�������N��N��q���"�� �xDk߭h|��<Q�U,�ɔj�����3�� ��jřt�.G�~6�c���	L��q1.����E��ACbH�|bJٍ�\�-p?8�n�ɜ5D��w ���Pu8��!!��8^�30�̄x+R:(f7���J���t'�Hd�0i�]�`;�'��y �lǹ��{[��8�0xpw�l}@��<��w}/D��m�E������'H������W�������i�2E����]	"����HE�,X��n�F#e�e:�Q��S0�S�~x?Z/�_�,#\�ep�D�y�Lzv	D����,�Ӯ�X���F����XC��H�L�(
�JZ�$���^�FX-Wo�Iz �E� M��&}����47s9�fZ1��D��x�+|���siog�P+�C�zx��۵QN�$ҕ�&/�HVJ�r�ݛ^���O3+e!Bs���~j�j���;�'>	ya׹��!��5�Z��{�>8����* q@�:�4���tFI;NR��v�2)2�"��oOq��$�5P�#��,!�sڠF}�N���#����UBD�q)D�p����@��\��/�P-�/����C�:�uڔA+�O�����
ݟ�D��>��6\��7��&�+��#5���\)%��MQ[Q����A�&���i�>�A��p�+nZ���ɶA�w� ��-� �|;$P�S��Y�t��=մ�Q1��r^Z'��܋NB�9(1��x1�*�$�%�ן�%�ۃi��3G�E�B������ص�4�����#3�#��Ӟ���Z|
 "�����6�1����&	5<��*��')܎7�-!�Ѷ��u��6�A��Xx�d���2�e�<��<��ME�ԒQ9�CI�����z�qЉ��46�==n2�0���ˀV+&V��Pr+~���[�SM�� �-�\���R�ŏC$�^�s^U��4u���J��~���O���B�J'X�nn��u�����"JVf���	�c���j݆�g9��H�յ����K��N��3�q���{7��kk�A��p/��t����t4���1�$��5�#X�ǂ����k�M#��	�7/?�����ǳp�O�8]	��2!�e��Y�&$�c��RuP`���p���,�9Gf�%\�Ywsb�ڞ�U�.�@lU-s��r�B��d%���M�sy��g����2��{��� �a�tLE�U��{����,�t}���۝��|�i\\�������mWƒ������S� '�
>��8�0~�|�W;���h������l�Uqo����P:�����3��Qd
��J�/3�0x�ng2nX���Ҕ�x�Vs�Ig�jy���{���d��~��SԶ�^^�{��制D�����Y]@��t�&���4P������+�~��{��Y��$�H���"���'�_	@�P�F���y�_U��_%�X�sj�KS�!#'v�|��G��:�(<j�JJ~����6e:�>�h4���	�G��!d��o��$.XSM^�����f&��>��YC)�D^�N��3-'L����#�\�M&,�H����&k�sv4���b`��{���`΄�~0̳.��Y���eU��D�H���vc}bT[]���-��0,�eX�~>]�]~��_ġ�r���Ŀ��W�r���W]
�BT�9y3~��a��S��Y.�	��N��� ��ݵ*�2�2�r��F�T�dZ����ֈd�j���k�_��y�gx���jy�-����mw�%�]�e;��V�j�����U�7A��gF?^S�����ݶ�4�t�:�O@U`�1\ğ;�[L�W^ya�{UԈO���@���#�!#�$H"V^sgDWL�п�'�\Nv�s���*��\hL,\E�h��%�e��\��� >(�~ޭ�-(�:�״Yo�^J���KW�t�e�����!�����]�Z�[%������H�ofwm)p"ʖڛ�A��QvK�	��K
��B�l��z!�a5U#yL���G<�{�9}T*
i|8���M�D���ww��O'� �y3�u�&E �[�b�l��猍����N�G�Ir$ pѼɶ�q���Q@�at蘒��G\I�#<D4���i���?�>��z�X9н���a`��������0_�	 J�,�(q3�2u}�Zד���3���Y�^��a����α�y4��0���E��~��q�(�ޞe>����-��2�@.�^�pS(����b;���D�T"��&%P�-vJ���c�����a@(r��L}x�Uɰ���0��g��~�E�]��x�N�������6�\_�|=�T�BR-��n�;s�������G
�t�Ew�C��� ���Xa�Y�%�Uԇ�&_H�>8Q�ڥ�$FZ&��w�3k���^؅`
���aAb�w�8���O���Ƹ�\��V�:���f˅��l�ޢA�4�?�Q¬������֧:ǉy��P���~�%v�0E�D'�ּI�2Q���	Ϲ��0����hZ� K�~�]o.�IZ�P��c�-�����	#��y���v����� AzU"�ހ��Ϝ��6��?�`���)�<\q}�j0���L�>0����~U�|lԄ�
)��KqƼ�Ўd�;.3�h�1�~)�3Eb����*u��s��,�Q�Q����P��f��/�����E_��㝕��\J	P?��������U%${��#�R1�Ъ7B}��ʮ*X��dOn�	�H\GE����a�HU�JC0c��I���G����=|�z���0;g���|*Ƿ�~��Xب�!�\��R���Nwi�V�%L��������w,��q@�k����38HY����_�y����(��4���ܩ����	p��,�W���N�9[F�$R�|bK�P�O�*�C)���-ɥH��@�2��[ئ�������=���"��]0�Y7R�ʪ�Ρ��Ϭ[��$
:���IU�n��6����a(���ʫ[�)�z�4?�p��UWp[j�Di��	ZA~����W:K��ڟ���)��m'~^�_)���$�i�@�v���U­��b �-X�j.��3V?z��4�G�ܜ�����nH�G��@�'���3��%��R��_WB@�1*D��V����:h� �W��Тn��SI��K���5�2d���H� @"�+�!�ީ疮�<� CWح�W*���Zn�����-��7�SULy �\l���L;s��F�X�k�p��ݝ���dSG����gpl�%��B���`*���i�����UF��޲�x4?"/e⛳�@��Lf�A�p��ܚ_����o�Ht��	�����)�\l"��V��%�ў�??<Ku��>΃
�y)���,�GN�"�c�3W�P����E��/N?0���Vߎy=$��#0���p��#
@��5��������G�9��r��P�#�!E����b��P�Iٚ�i�p��r�ɘ[��w����nx�zܕ�ĸ���SS�y2�0�t�h�T�+w�S[*k�[��c����B�z5ږ����M��� ks�b�~1=O�V�o��=����?x���ȼȁ�W�7�)y�G���11q�fHЛ�d}�`|��+z��k�Y�ؖ~��?)n�m�l�,W����SϺe���i� Ϸ݌(X9�%R�8����Ya!Lb�>J�]��g�]�l��W7��d�ф�i�߯tl�M��I�4���.YCo��0�8C���p�[Ne��(�ng$>j8�j�1e�ZN��B�+���|�o��g���f��L3B��b�Lb�n���C��~υX ��k*�vV�(���]�lY���H�L���ǿ�t���~Ao#G���
�R���j� 8�O@�a�= �0�EA�a_��%t`B����GsOkJ%������-ߞ�oN�b��ql�E��~G�A���;�^���f�2,2�iC��Ŏ.�a1�X��{kk�. �SȯM`��',������$�3`�!SZ���,kӶ�̲��ʞ":�Ē򞃹#���}����T:��<Zn�h�$��^@��v,���d��NRՅ�N�ۧ�t��v��3�F�M����ѧϔI�;���Ysތa��Hw;�=�Py|U�v�*�-��W`��✡ɛ�oUǆ��Vd�춬t�%B?�>A��6�fQ$7Vh6�r�=i�;l?���uQI�@k�fŝ��ڻ��.XD�-��W�\o;%E�5���'����a.�Zq�N�Έ�-��8��[��A���=��A�Cv�s��=	��8Ht<�Vn����f0��1�a����u��J����XZ�Q?��I��
�K��9���j�(C5QL�c��;��s�7.�K�~�:��)y���n5��U>�̀�]���R���{��a��.�����@�M�"� �vU�vpJ�� ����Y5�C��XU֙J�(Aq�uBy 54�`�E֨2G�o�g��Kѡ���1v� bYN��v�V�o�|����-x�d�tӈy��,�?m�f"�;�=:m$�!�z�۪q��݁��Lt��sK#�Nvj|z˝m�@�<�����zúǴ�v�GO (f����k�6�S��~��.��r��da���4�]�2#��>kӟ���5�E�OJ,#K ���U����j�o�:=������4 (H�}mC�XM) ����P�͛dY���{u��us��S��CRd����(����KBi=��d���:d�AB͚�b,~ ���B�#l^�
4��*�$q��X<<o���`@a��p�� ��_y��{�S%eMKKƎ.�2i���%��!@�"���2��bQ:w� 1��U���R�r/D!�~��:P������&�.���N7Q�5b����k�^��`���C�t�N�|[��IN<��Y�!_�;��.<[�AN	{�fҁ����O�z��{�!!��0h��>��ǐ��+%�zB���9f�33p�z�QG9��"/���d����P��Jq�}e�k�bx�dW?s���N2�s}�/d�(�v���#i.x�l��ϪV�̃pM�.�¬f�D;|ѱ�EM��Sա�(%Yj�7K�>��)岞E*����h���./�qx<�AQ�͔ֈ8�z/������L�t,[�X6�3zώ�y�p��^�F�+>!+w���x?�f��.$-z���sF
�/Ycz?W(�Ka�R�h��ٽ��Ցz�t�<��q:�+c�[:))�} ]ql�n�
��Bл&c�_�$���)0M��d,h<�f�5Ol�k %a,�d$�+���\�jH���^H��G���,fv�5+uW;�zS�2u67��X�+G�кP�RL�C�_�K����ps��iC��?��k�2=���y��qY��6%�����^d�8m�Z,���=����`&�PN9WX��BW�����>z��j7;����It��E$�!i�$a �ךK5��핒9Q�� Ak*���s^a���3�R7�V;U��������B:�����Q��1�E�7�����&��z�u:�c"�G�Kj_��U����CO�!`�H/�-*�h�&l(�巺���> �a�y%�[�q��{"<����64���zBǯb�Rl��v� M��?�'���E����s��jI�O�j�d�"~�*v�{�Lx�U*��V�s�z����yY��5��L���,ʰ�*�2�+�? k��];'̀"1\h���T�9�]��{n}�F�҈ݺ_�eM91D�w;���v��4^q�R�9��ј��JM�!�ۺ'��|r�e�e�4It(�����wD�`�l����<���2
���tS\��:��^�	VTC��'j��	�
��2ڻע2�p�-�Q�p+�m4�k�� I��<��24,_�u��I3�J���#DK��`%,auM����U�T|��ŉ�� 4�K���S��ڸ��l��>�c.ұ�w��N���=;8����R����NRՙ$�D�[�ɱ.��Փ���,
�����<���]=7*����n�@�e�
|~|�(\$���Ja��M}�+��.b1�=��t�B��<��xNO����=Ojs�����-f-P�N�"?de�E����x��q�V�+�Szo�&{2��ub,r��7�����v�wD)��,UK�x]���$]����7�6uJq�����tŅp�"PɷP��|���g)��`u�t��tE��I�\�����2\�'f֐KQ'_&&l��)����~���ǐ�W�{�ԛ���G���x�Z�k��.�k��#]~@�����»ֆ�ܫp�ƞ68D�E����r��7����E�
'Zj�e�L�?����ڔ�\u��C���`#L>���l�-�2���2���LF�d�V�Gr{j�\_:P������i]�|?���1��&�W�2�iQ��H9�q՗�7���Vf&��CC'�`
|�\���<�!�x�ް�H�;��t�ԥ��ow+�#�i�#>�A�x��a��+�3����'��X�Z�r5诳7h�Ǎ�Y.B�Nɒ�a�>ιX[�֣E{<򨻁�?�,�L	'���7iD�䢙g�	�V_����z8m ���)��y�IzW��=[��<(�)��op�뢈�#�$��Bfγ2����cX�=����/dJ��*>Q+3o�_.<��1�f��N(��@�|�ک�gsZŰ�p�MB�A���8�����=��@����-q,vĠ��d�	��i���
N�^a�v������ޑ�z� �\��,�s�v���?Z�v��Ry�_H�e-w��J��+�Nհ�i2g�wQ5¿S��mL���$����t�!��ʹ5���Q`��6�Њ<�v�}���
`o�إP�����2�L4��dq��y#��<2��@����fB�ED�s�|`�ܠ�v���p���Ib��~P�y�3ݽ:$$���<9�n�%��7�UV����9U�fR~K皥���V'?�����<���t���q���ж
�;ŵ�%��]Ul6�GO�
jh"3�A?W͐:\����{0���D��S���� �Qp�22����p�����(S�zؤ�B��t�=M-��9��I�h��E�f�4Ϸ�K����Gӱ+,�F�Ef�P0��2u������sH�p�]w}z��i9��ӆ����v?Y?��-�#a.�*�����:KN*��/G��	����������`xYħ�i>ؐ�nO؀^��nV����<���p�L6�X���޾�1�����H�R��������Y0ϛL�4���i0{Z��d��f+y-�z$�	��H���+��*�(�ܗ�B>�U��!�LM���I�b;��n��y�� ��	��ˮ��h
�m��`'�B�YQ��!^BG�	��^��e�)䳳Zsc�AaK��0}������,�HΘy�n���x���$n�d�hg7�3�_�6 �iJg9�p3�*�T8��耪K�gz�U�� Q3Ċ�^2'r}�>���~-Ph�Z�LYRT~4�17�������������SN�2x�v�M}����pH
y!N��5�'�M������<�5�n�E-�Q����@=o;�AB.�%�G�%�l0r��.��)��DC�A�M��RԇG��DO�m���Ty����k_�;L^5�Y���UVah$SP1��
>�%w�B�f���E�q�]�qAF���P��#8rU�d(��wa�ӯ_�-G+���)����x�=�"2�r�f��Rɐ��Q�k�N���I<d(^�I'�ɨ��0@��E���i�����I`m��NE ��$��
��F�ۥ�2}��m��)*h�go��L�o.���s�����g0�<�����%QxWt>�gj˿�ߡzI�k�_�~�O����_7o+���~�v��6&Xq���q
�DN|a�^���ٯ#v$��D_�4$d!c�|��|T������fǩ`��6Z��}<�_	K�����o�]���b9B�k�!A�%%x��^�e�Z�^�&�m/�A�������_#�3K�_@�9:#�@�B:8,��e��xg�f�{��v]�G6K}���1n�����8���)���F���:9�N|�O�|���UZ�'38���I�Qpg��Y3Zr�'㩧��A%'���艃φ�ǣK�	@���x0\1���5;���X�a-S�	D��:NqcG�B��4FΏ�Mh��>O_�,�m�h��Dv���=9Vs$�7R��V{84cdYT������SC��#وm�ШOK70��r��O2�\wWj`ce푏#7h��0�c�x�[�hε�߲B1��]��xf"�)g���l\�"eAсlc��B���\��Mj'��t���ZU"��5��3������8�N��/3����A�>��ݼ'~���)r#D��i*�N)�C?Nc㘏{��Ո�} ����im90��e�W�Y�Z*�G
˥�"2���FwPE]��1�>��_�돀$P"B�����9
`�^nwQ�?m��OQ� p��a���㒦�ݥPQ�r�$��R�i�j8�������HVA�]�5
7*�^/e�z}z=E_s��K��-@�FYTcyF��
�bXN�fθ��\`|Q��ʓm�#y:���`}�e�g�s@���@��BC���"����U�0z��Uk�@�w������w��q0����$ҫS�ա�U>̍З�1&>�����v+Ϥ�X�Fh�6AE���.�7��,���V,@0�����x�x;-F���:	��G�4��±g���xs�6�*�18_���*CF�!��#�؆�}`���a�t�3����0:LqSYZR�Γ�.�l%�ϭ�6�T��X��"�MaD�g���ŲI����Xc�"-�z��w��- a$/7G�����p�/�X���b~���1��/�c*�J��^��V��M� 2}�A����D4�-uZ.��z���P�j�EL��8e��5P�R�m��m�݋�F�)8�(,|Ox�?\��N �m,T����z;�I
II�'�iw�(����󀁹U��|��+�Eox�3��(|{"���b[V�zLM@b�0��:�t}+���[�<�Q"�w�_�����փ��[:�d��h]���
��^{���O��Z�����u�R8�z`2�ym�Ñ�/~������������04���i�,s�:0n>m�|�b.枕�a�������G�A�fZt'���/�&��1�_?F������3�c��e�����s�c�	<@ӝp\�%^��Ĺ�G��Q�g�F6 �\Sa�BzW�/�I�yq���� N9�b��Abe5K0hiJ��[�ZCN/F�Y���Y'r5���J8�/�����0�����xz] ����蒎 ��'EC�wY�� �Ǎ������j�b|B��s��+I^nӥ3�.���O� �U���me*�xMN���l��M�9D[�ow0�\���>V��uhG���,9b���5���M������(�ւ�N y����F{���D��a�t�������mB�HkT錌�k�m�dnR�ޜY���>b��R�n9�H�~@g�
��]��a����������K�Z�$�\t��6�AM���M�}�410N`�G`}�¯ �R��.�^#���P�ΡK��IjZ��Q���TώP�.� �]G���w��ô-�u�b`s��[Y.Q'�����~�����#̑��Q?���Ynג@���#�-��+�����&_��X�@��+K̎��ԡ/�����y�'499��86�������# �w���.����#��8��iG����  ��2.�I�i���D�r	5q����޿6�OJ)��,���R����-j������n�%d"�r7o}�o�!�Lg�&�
$���ƠX +Qp��g' H(5h%�OU��Ʃ�~j�uJ�_���7�x��Ț�����L��wrܦ��VV1b�N��ƀ�+iw m�B_��)L��AyM�a���J����C�y}Bͨ|^�QN�m��)`Y��%�r�Bz�9�r�����O8�`��a|Q��5�Td���VG։Q`N	�|��X投?�o��L�ܺ��x|#���/��r���0&����KQ#�4M�	��d�T��[���7Z��)s z{��N�	����^����&�v�wW)�*
�a���"��@\j@���7%�oz�K�� �g2ٕf|��"�qx~3ص�R>�>z�ث{�HJ�۶U��yF'i>Mx�Ӆ�X8� lq�ԅ���H�����z��N���]��Z(���S��ˬ���(''������ �"z�/~8"�����GJh$�{|�A�\P�H��2Wg�Ip�K�����HEQ8�b���TeC�8����� �a�Q�ɾ��Ѳ<ߊ� ��H3֧��%���|d�q��`c�<ҜҢa�u� ���d�>!^��\�Բ�٢�Vm������
��M�Ң�7Q��Åe��h�Ӛo�?���J���/P�p�Oݝ�N� ��(�P�V\�Q�VBH�(9N���i@��Dh&s�@sذw�o���N�B\Z����N=�A�«yIY�U3û��?� h'��� v�cn��R��ޏ��tDk��%y��^�a�S��М�����H�~W�f�W e�i�n��פ����uZ��R%�F,��&T�y�2�j&F'ٜ9F�^�A.}��3�X�+~WZ�Ƕ����(@z�U�aq��g�!�,��ƺ��$ܳΌ��k)W���}�� ��y�B{�;�ZJ's���4ՈL@����5$ܛ��&/�K=M׍�n�^�I5�t�>Ǎ*퐊-2�&����-@a��B �"���$�Vy_�.�ڧ+J�>��r�[����di^��Z�J�VVǻ�*���˗�'��0�ThZ#����#}D������d�mK܂饮����פ�.��� >؛��_��J�з���U���P�~
D"���g�HRh��0��A�v��S���ϙ��Tۯ�V6�.O��*�Ӱ Q����|�0�3A�|~m#azA�����;4���d45�v����^"ы�r����a/y+�����`D6U\��?�	j����
��\mx�"LY"�$zYl�e��r����h��<>^�T��i��n�%����MN�E�4P�rsx�̇�����1Bu�$n�6u��<�\t���F�^�vJ��������(��-���f%�8K���|h�ɸ@ϲTz��_��Q��\�$v�{\o�JG���v�˵�@8���Bљw�;�c�Ӣ�q�9,x����(�ߔ�,��P"q�km>�����8�!�j��rj5m�ѥN�}�j~�%7M���OR��i�]U�S	�4<�G%��k::{�ҥf_%m�{�_e�?b�Z�S-�.�.��{��4ٿ]+�]��EU��x�i�M�?9���֓��3���h���D�5�.�����俢m���a��ћrh+ѯ #ݣ�N�����a�h��߇��I�er���'t����_Đ(�9@bZ+��;ԃ�\�n����A�}D����f�W�E��,.���������G
��uQ���QB��fXor���oGk�f���[9�Zy:MZWњ�T,��qe�?ޓr�ٟ �9��0��&���������L���%��m�og���_$����V�0�'�sAJ�M�='=����M{��Z'�������Ѝ�: H�n��A�J�H$"k�6����h:�Z�BdiSKB���(��*�����̗v�F%�r��+��g�	��һ�.z�vA�	���;i)�ɦ�j4
�O�$m��N��,�����'���0\UerEM��V<hf�[��-���Y��6`e޽���/���8�@ƞF�9���E��%[���z�h��}�k�����9���_=�͒}�������[�7��8�8`����9���)[k��g�����T����\y��ў�}�%lJT��(�rd���\�|?���Dm��{�]^/��9��r��2YO��)5i�k	|]�(�%�.TĄ�%�����y�p����^-�IA��/"*ol��9o�\�ڢ��2�JXx��QS5𢇩�M��)#D<���˶��
���5.N$K�I\��0dj��o��PFTS�^�&Wi\QS\�n��9�S��\��(H4s�#'�����R+>��P������H݁a<�!"w��}'	8E%��/N$���&�2'����̫?L�U*��f���& �5I��a��mT&�_Bf�~�Ea��st�����ʛ@�h���7��B;�ɀjP�\H�?�o��Z0���q��x���j􍘅���0���Ju1yF����n��-�D�z�fdi���9}�<�c�m�ȫdLת�n&�9+Jh:�	#o/g*�GŇ�`>KQ+4�Hr��0�m�>ަ�\��m@�j/o|�p�qq�ʻ��p��Z��I�C;u)�V����EG���f"��0�ޕ�gm�v4�ސw�ܞj�AR?Q�V�΂ cݴ^ʂ��{E�M���m9�SF�:���~z)�� w��+͍u����Y�/&��|(j&���+���q�2��6�Ϲ뷋}mX�׏;YLx��Ю��1է�]��b��/�톜
����ՙ�A)D2	��;Y>V�Ҏn#�z�6�;︝���-�N��)Ί��ރ���51'\O���b�]Zjv���*C�
��.�n�4���z���_�`30,@
F��<S������vDH`�&�>16�j޿��ُ�Bc&�˛�Zb3���g�}��.G:�?%/��s4�pZ��(�/�'�ՇZ:�j��n���FjH��ʢ'���B��`��;p�:�8��P�ZҬ2�-Ҷ��q
6���J�`׉7s��pr������D"iMkı�	����I���(��Ŗ�s�!aF4�����^Y�(d����xJ����-��`��¾��Kjη����43JL�=�c<�*j,cE�Rݓk$|��{5�'�TH��a�9�6�4��!O�ps��"���Vg��C��`�!�3{�<̭M2z��|��Q� ��7�=������_���ľ6�-���ɀ��F�J�§��(+{���bLOQE@M�,R>X�}G�ry)���]	��QNH����lG����u�y�;ٿk��,�����B������V��v͋^6ℰ4�E�q�~-|r����H�z��f��Ĺ<A��C��E��NwI4������LP�s�E�i��q�VX�]����8$��A����f�-w,��36��6~��6ӑF���A�o�(�<B�-R��R��G�.�[��)�꺏 7 �Ui@�� u���C)����T&��9C�������K��.Mۣz�Dp&<� S�ҩ{���HRe������ٰ��9��G�i�ԫw�����S�v�:�_=���SC$�I0^�+Z��$b}��n]��-�����m&��T��1��jԮ}&4&�[�nN�+{?4{^�8�9P$?L���R���׫%�-�p2s�si��mG��l�Ă^��*DyP��QAI+^#���!2�݄	x��n��E�v���"�aug��?�����sZP+�B����K���-�|!���� /�7#����':զK�����慥O!�W��i_���W�{mq�k�/�_���4�H�y2������m��4QV
���_*��Y4ϣ����   �x��3�/xΎ��x�ozO
���T����k�N Ɯ6��U�����\��(@��Mx�&��h�GD��,��G�UwN	�\��F=mX�l9��kE�c�V��N��٣ֲ���$�itt�����4M���dJ�c�ΰ�L�aC�7S��#>'�`�v�W=�Y;=��ha���ob�y�����ܬf|���!#t���޿ ܝ���R�e�j�I���+������ ��.��u�7h"�a��!���Rc
Xk;�hb�~m6�?����e��)�1�W$����`��o�a�w���:Z�4r��|��/�9EN���J>Q���:�Nn��z�5qez,Ќ)�ڸ�)�֗�%�?R灒�s���|Lc�hNnf�yn2��KDڀ5vb~o���7�eE��
z5���7�̽SF�n�>�/���)�4���\��]�(
�&�E���TA���(��\6,' ��d��p	�h�*�$��Mo���$p��n�	��!�ks��a�3�M�/�0��.d5ȱF����'��1�~�c�G'��!�L����^������$�j 4��M�c��޷�'�`�����4k�z��BX�)�4�K�X�o��k���-����4����l���u�F`�V����2,���8.��NV���� ֽ��(}��%�vSe���*ܟ�a�}4�'�K��k^�O��(�u9�V�(��:3�	��������ٍ�o�Cٟ��fsJ� FP'�Ǎ�Wkf���r�s̙Z�dk=t�Q�iE�{��n���d!�:��,߫�SaC��pB?���U4�U��2��ߡ�da��N�՛?�nz�afn��͑o?���'/h�jLIY��O�4 ��ݬ��u���)O�>�I|>A!`�^2$�>Q�ئt�¦zޣ�Ͼ�^��+94�S�����y�w^�J,[���ٮ�s�W�=�r��{4%��`6�,�4���w����Y��z�;��ɹH{컔x�
�Mgk�{�\�Ǣ��aѪ��S`�-��l��#R�� #�K��ҧ���V(��áj_����WLv��+�a�q/�dZ�uY����U���h<�KK�$�R�����#�&]�I�Ȉ�
k��?&*�٪���;(�9u����y��ȋ$w�'?��PE�W$B-<��"	��s���Q���`I�T��A�����_�3
D__;�쒢E����&���n1ʝ�Zh�M�0�ou��ư���Zŋˏ�'$ZwP�������]�� �j�ħ.��\i�BQӶ^"dH 9T�������p��X����*��⾉E�	j�dM">�N�p�XR��yh������f7y��VaA�<��~{Uo:���j�A�ֳJ���e�AC_�M���z��߆1�g����V���eT�]�]*��0�kZ�'��0�P�C&����<��N��U�b[.S�"�'g��l��f�A��g���BZӪ�[��	&�o,��.=�J>���,�=e����q�	�1�\h��O9e��r�9.7�Ah�$��8���g��`ǫ�����9mTHS�΃��ѐ]�(�=��^���KJsZI����&�1k2�~��,tb��`Vs]b��_>����R���2k����Vkk�(;հNy�2�5;��)l�O�HquoXɝ��b+1n����4�r���E��2��ps#��!��c\Ns�IW�̟����
��Ü�=VU��tn ��+�:�̧���ň�<����T8iM�V<�������,����e�R�/���!vd��FKN@�mi 2�vuC�s�8��'O�[�D���-.e�0b�i����||��ӊl���(^󄝅��)�Z�ǧ���!�|+�
�:�~�	餐�-Й�i��i�6H���Q\�WIl��f*�94E��^�I��Ck�NR�jوmsl�C#���X�>5�8C�t4d�;�S�j�־��^1V���f�N��{��8�,C�n�����vٌ
q���j0��P��GR�Ckx}C��WQ�R5�cp��ܒ���;-u���uŮ�8� �����[�P,�ӁgU{�H���_�&\�r�&n���9�S��Kw��^ �m�(%2wa����޵��_�6P�d͎�9�AvEf![$�z��� `Pp��us_����l�b��I'1����U'u�'��Z��UT ��}&��c6���,|ř�;���r�oE���c��U���1��j�A����G̟�{"����n9����C�jDL��&�ë�_� �c�c�������h�:!�mc��/���穙oDI��C�軔$��
i�KW�T��6����Q8 ��5�jw��/�	�=md+��i��.�}�w�c�m3��^ovTt�|;0�d��Y5
g���~�_�Y_�mE���#�<��)�p��Y��p���x�%��p*n��I]��y/5�,�Z�f�3;ܪ���#
�E�r�V�j�����t���/X�D���r5<�OLQߔUknyc:�2�W�<�{�B�����8�n���n�E�~���O�('?i�U'�]Jņ���ޭ޷'�r �����c������>�P��5��, ��n6ă�^sWq�	:>д�w�R5mh�ʉ{1�HR�dt,��_M��$W{�mȓ25GB-��nޮ��O� �ݳ���sqxͱ��-�<�O�㟂`
H$�zaY�
�ߠӀ�oA�
�b�o��e�c-d�%%�b҅O�LPe����i�����?�Y��o!�ZiP��J�!zJ8�/-��2�����SuDHO� ���mG���]i�j��&5�s6�8�>kԫ��`}?D�r/�\�pE�6+X�L?,G"�M����S�<�������4���l����b��S� ]������$$���(p�d��ϴ/K���bY�P�݀w?漂rǒ�)�� ?�Ns������:����Ǒ�^�\!@.qU:�]J����ɥ�wP	��;�p}/�����2��
%4�d���
Z(��*gJ{R����BG濔�դo�+&�̪�lu�M7՗�z���?R���X�BA!13�\v�밯[ζ� ���a�Q- �����\�`��R�����d&T���^y���Ӽ' =6iN�Q���0/�T�S�&;����t�zBe��	(�n�=�p���r��L���$��B�>��̱[q����S��8o���t�~��%��`�k ��'N�]��ӊ�m�q|I!6�.��ɘy��"?�6  �E�c��+iz�~�XͰWj)�,Y'���,jVp�@������R2�/0�t5���0B]���*a�JgL$S�>!O�iqX%��!�
�$�r�� ���2�`p"	Q�S���A�a�%\�O��q�&Z,��n��5��̛o�*�p�c�+�4�{3v��
UsJ��&��R�Q=��xw�P��=�u�=򲩢!|=��N}A�_w��� ��E��Aȷ�ִy1�9};�����Xx�L�N<D&1s��fr��u�>�p��">U_�2��%[�c0���/ �X����GA�V�Z�%(��_��n�����x�\��VW\��+(�M�{��d?���rմ�p}�
*pi��w]g�_�
 ��+�J� �?<��Zfa_��	��g�.
�Sי����i�z"����Av�%>����O��jWMLa�%��ըb����c��=.�iP��~�-5�MY�����Ă���0�;�Z������{�D�1���x�v�O�/������8}�_����tH-;4���"�r&V�(�ޒ�ES8'����Ʊ%��4:<�d>z���HF�be(-7|��Ij�+����?Ê��hv�<Iݻ;�DQBv2}���P,� ��[�9�y��t�+��)o�8Z��>�G4�'�Tמ�:���6�F���M����	�x<2G��"j��>D=&$���雡6�xȇ?�S��U�q}ҩ���	FQ��;G��+� $�}ot:Z]�n5SS��uLM"�e��i˩����5E�[��G}Ou<d�P���n;bG�V�/]���*��{t&��Y
�n�5h��J� m��2Xf(�<zD�\jWPb����/4-~ġ]�zr�Nc۟+������9&�u}�<�%ބ��|Õti��:�%h�PL��~�؟S�ˌ�_�9�!Ʃ���W�	�/���A[�Z��9fT[��<�Ѿ%�=�4rҎ�Ůʠ�f,�TF���5���T�#� /$&G�ܣ��*<!E��$N�̺����Sa�/��1���_��B|H�р�uk�IEMD39Ģ(������G*�g0�q!-3�����3�a\�wW<3�g�t�*��ک��4dQP���©����1��R;���v:�;��1B{f��u�jJ�%�⛊e� <�:��n"���o��Qʍm�nv�4�qw&�;�.��r=���љ�zG�'��Q�2�|6'�0c���֚b�6��bE��${���+�k[M�I�↶z��M:��� ������U�����ެ�X����sD"�2-os:Y���i{����)2�s����!�)E?�F�"rw���N֔��A�(𔶪���� �d�N��I\V�R�\:�-|���1�Hj|�㛞~0W��s=iy7?���9��T�f��3NT>sn��C1(]Й��i@�1�����?�2jk��~L���r��D����+xv���ԛ�F�E�����T���R@{��pp�[H�l��q
���%� Z�.8����Tc�� Kg�Q�1�)��� Z������U��>�;�5�t�4�#j��~� q������԰��d�,����@W����6l�R>���c|�r�#= z^O���ЯB~6@-��"1p(�s�p;!�+�ƈo'�T���}p�襤�qǬ��y�qZ�IG��Z���_=;�E��9�b����<�MO�o'$�i^~�di�0*l5[���iaT�t3���cC$��ʒEL>7��f��m^�q-�_���L��p^�=S�m�� [���F`� �w��א�B*�6�v^7���? ҟIG.M�@dE�oq,=Fq쇂��9��CO��?���vi;�&d�_!F|H�7��q?`W��m)�A�i�|�_w��4� �8��.7���J�����S�mf��c��^6`n���
Rc��������<�l۶'�M7:29�!Lż��b�s�V���U�,���̝�uʐy =��<��(	��6��;:P�~ϵҺ�@	�Y����rvݧ�Qr�t�Bf~��v�N����Q!��Z�:�2Nއb�����X�Z���9��~���.��hr��#џ�?5����$@[�2����B�q��-w7]��X�R��tt�%)��]N��[�1/*�X8M���Fi'�@H!�S':�-B�"��|脤(�Ȧ��n�hCٗ���A������&��r����E��T�>��UCQ�o�]u)��q.��54(��<d�1W�|�,8���Ș��C��v�@����NҠ�ϧ/�IǺd���%�+@Q����B���:��M�7M)��A,�
�/X�R9^��<���*|>���-�L����}�(0�XR�O��?"G������[���b��R����U�1�鰏D�"�;0�3�"�-��N���D�w[��x�����(F�`��މ�@��L�f<��3o�|�\r��٫g�C��-�p�˴�Q�\�'�!�ђ�e�@�x�2���p7`�h3I��-��J�څ��q�ߌ(����jq�i2��p�X���{P������ 8��O���(k[��sO��5����6�`�����4̡��@�v���S��yo��
����a>ς��Gw�ђ_0��g Bˋ��.������,Q�P`�	��O&�۶p����fS�Ga�RW�5_����m���u��;��
���;m��*0[\�������3����`8!ɞ�N��^�����4�U~J�0��)�����M��NǪ8�K6]}G��O�y�Z����s�V��S{o��K����lIa�`��Y-b�$^hn���W����<C՝�u�{��_?����D�?�*�m���(_P��hP�@�㕴��knA�f^!�4#�9�0-��(9�*�L:�>b�� z�.�S��&���Ԯ<a'�XN#`�2��E�=A��_��Ti���@F��.��j�����2#�t��	�n'q��#uW��KT�����+�<ܞf{�+�ߠ�dv������?�,�U�5
]���m���@ �������#�X�&Nj~^)���0Qm�Njㄸ�n��r�o��@>9�u��.���L(�ȅh6{�S�3:sk/)���#��iEi1�M���9����}-Y'��mW9�C�;8'Џ$fj�z�C�i�t.�N8�W�!5�v87�L�a����R���_�7k| +OR"'s�����/�asy�1��N��L�����u� �E�`)�23�Nإ��X�j�s3�snY>|��s�U�i���� z���aY��,Դ��paԡ4�	G��� ��,	B+��]d��D]��j����-��v��#�S�A�PBZw���N#�O�Nb�BQ%}��z��&Hdy�m���M8a���pA:�)�܎�_zR1�s����-��n9Y$�D/�K�Ć��u8d%�g6����&�ӣ�(�\��n�m/%Z]u��j��,�R����5�?B��~]@��`�
��`�����G��0 ��;yƣA��v[���h��2a[�%�S��h���h�um�
�K��6�^?���I�@r���ZF�����	�,]ҡ�������e���a����"�ʵh:�K  w��9#�A�p$��
M��p�]J�+�l�*t_.!gVeŕ���h��q�g�Ќ}���|B+�c�w���py�N�n�?M&Mj�*����,Fm<G���U�B2�OeF�P]�7����Xh5<@ċ%��W�U�]�q�{Amv�'�.Z�2Nl�M)�6ް��]�}EVթR��%J��N�t���� ��,�4��c�$��3�'1}����STSyZ�(�
PGy{I��8Qd��+�EoGP��*����vpE�_x�!C@5�m#چE��Z�U[V�Y�����%��rP�|s�S%�r��;�&�\�	��*��2�w�`�U%[('HN'awH��<f���<�n���8����Qض���0"+�O,-�J��sDn�¶0D��MezW�R�����F}�k�?S��tn*6b*���ŧ�"f���Y���Ġ�1��;kģ�x@5��R���b Z����Wx�t7H���Ve6���	��O�_�����R���PtQ,���3N��Z ��~rϦΦ@qJ�ݸN,>R��Z�dF��6�p	Nc��BEz���ƽ-����+��QǢPt
�]��S��=Z�:��x��ꯈ�Bт˚�m"YY�s	������X�����[�d9A��XZ�����%j�r1�P�%Z�{x�p�h[�ǜ�p���>ZJ�9��|x�Y/��6�Y��x8J�
Z��֊���F��9T�7F6Rb�� �O~v4�>v8������"H���|pJ���cԦX��8t�y�?����\�Y�]����϶A�	�?U�~��[h�)�����;:�xS����~�Bw_�:B����%��J�Sy���D<kP�h6���;+4�a�������#�|R4�m�)�l�V�1�-#�w��T��e�[\���a�nv�6��������@�,gG��]�V���'5�N�Y��n_��M��E�a��!S��I�
�������ˠP�}���HM>I�cW����+��[���}]�ONI���AB�sC9T"aF�A�����/��4?�TO���֒�F|��p��n���S`��bF*^��D����^�])jq�$e�PV��A���ӎ��<\
k��ғ:�G����L>U�I��$�(Xv!�E�X�)�m��ze!�*� ��":l�0Y[A�NG�YU���̟�<G?oj�b*����L�>�5T��m`�Ì���6*�ڭ�YJtu���_Pǽ1�u��0����̢�/���a�����w^�ZS�7r����\��c�hxaRh�AӡjT��޽A")�����ǘ��j9�����.⸐*�T*}��z,��HX3���r�K���_Vp����=�n��~�0���P'nPT����2��!�ٛ���)k�&F�*I���Mx�_y��:��C���?ũ�����3,�KLm:�7��ɗ���V�Kk��ijc"n�d��(w��9��J�{�Xc����@�X���?,n���9��c�8c�"Mܐ]Se�T\�>�Ga}?��d?[1�,>��.��ϴug�չqσ���L'�ُ�x0��m���&��'\2�h���Y<�{QŽ�G�
<�$�����\}u�7�s�
ˏ�f���ZC{��g����uױ��7J���G��=
g���`��V]X�1��`�O�PC���E�D�3%�����sk'�o�H���cy�kOf�L�L�A����nj���ʺLP��E`Y��	�j�����s"f�Z�b.i���,kX��"�G/"��X��R�6�!�,L8�e�rca_�z��0)_�E\7E�h�&���{
�����j�D�FFHя/�[U��[SFU!O�'�/�wo$�X�B:v�/�����[s4Hư�e�K���F��ʸ��Z�D�xp*�L_/������)E5���lu&t���X�+\��� �a`e����&t,j����SX���D#+/��@Oe�&��g��tF�f�%�x�f_	e[Uh�L<R���W��s
c�N�x?
��<\k��9R����Dx�o^1aY	��"7�`���P��bs�CoL	pw)�Ot9h�����6�61�g@)O$R����n�T���1¿��r�D_>q� d�{CB�M���]H	f��?�e!��r��=UY�2`��[+��
$P�=)�;�<C�L(�S�v^��9hԩ���
���I~!���(�6v_F_ۨc��ۇ?��e*�s;TRF����:�kwt��d�]kr�l�w%�r dAđ�e�h�j�6�J��'xƐ��)vR�gȨ|\���g!���'��~��g�1_���pI�*W	?K�Ő]�D��"���pq%Ri��`a���F��Y��c�Ɨ�v�J�,�}>�G�{|��VNϭ�quhs,Wh���`tL|�a!�}l���{���1ui��%���]�i=;�2�Ӓ�4�ǜ@��
�,���3_w(M�����M%�������Ԫģ}��ݮ7-(��w��U�f�7�=�b-DN��KWZ�N@t3C��l1�n��p�dW��N�7�I(�v9�E�:�g/�Ө�B!�����5U���y�b݉[��;�����cP���j��5w�)�pl�*�{�U���g�)$�qD��t	�-iX��Z�Eј~�$� M'�$ ��Dܪ�#�������V��t������X�� ��F��q�|��؈N&��x@5J7E�5������4L!mWoT��`3ˑ0�_-�xC�=!{�=�%r�ږ��=�����i�j��,����
Ty���XJ<D҈��	� ��z�I�/����/tW{��}ctƎuE8�w�H�E�eBd��}��׬����Sp27$!c����i�ĳC�2~��ȹɡĆ�7���]*��)V鉡�G��>�Ӷ ���!��䊋{�fEg�O�!j�1�������A(���ޤ�Z[s���dw��j�
��?��Z�(j��d.Y��*��P%j����>b�w9x�H�r��n�
ɬ�>+T�b}`Ч��j�G�e�­=�Y��G�"۬��Q�:q��\@�6E�z�����e�����V%틮�J�R�A�K|��C߃�O,�MtUܷ2E=�<Pe���o�{��u��o��oø��-�mc�r���YbN=��Ҏ�n@(�i�EXF�K��|��^O�:c���Pm�4v
����c-Bj�]T_�v;�h_�[粞~��ڡ�P�"r}��̰5c�E���~�U(r��~q���2����Ht-+D��`�E���_"n�����0�C�t�R=Ҧ�$�Bo�V�/���XJ�,��
n���s+hJ<��� -!%z	���SZ�ͦBh���{w(;),����0��_���zۮA�&�|�W=Z��vi?��q����j���
�p��|�t�̭���l!���\hB [sτP���y�ZI �8HP��5="&:��+���q�M�Y���k1(��\��_�5H�_��[��}⢌ϐF
d��o�4�v�g�z��`���u����n��4(PQ��}@#�b�"���?+����`����36���c�;b�ؓ�{�".�ˊ�<���
�2$�xx�"���t��q�75����k4]�D�@�e��Y�L�������D���j��ݻ���ҵL�?k0�Z�BԿF�b��r ��몢|�Ɯ��O\^��vv�Hk۞��qe�'҅�NEC��{4˒�v�6V��������rZ�}uDO��u�:_1,��I���<�Q��9B�Ca�&���[p��n�Ԍ*�� ��x/�J���N�gg�L���aB�L=U9�iD&Y�`��{�g�v���T��0rAz��a�b�w��!��˺�u�i����$�����p���ZJҎHȴ���W/jq�0F�ԫp<ή�� Ȝ������w��7/V�PW��)��;+�R�ȝ�@�dB�8�ϫ'd�w���H��4d�Vk���&��4�~�{�:��RcⷲQ�W�Bn^s!	�	Ѹ��"��9��amiuуfV���r�������.�����.�iS9��: .Ʃ���d� ����� ;���Кb�0����yY�a
0�nX��!~�e�t�,I�1d��lj��њ�7�ߧ?e���(VH�~��t�'�d���m����q�_{��}k�WE�m{4�����@iqv�w�3��i響j�;/���Q�|bs�]���o/28���jC F�k=�f`�����;LU9h�c��%�~��|��;� 4(|E �Ԣ�F�C��
��P}�$�a�R�N�5�v?a�}�0n	�����N�G�z��_�[�ӣ���*7lMuM�aK)��@.j�ô����RlG��*+�r*��� ���(��s��hn,S: E��;�O/�hp9��[���I��q����[�� ��Ř��x˽�zчu!�����#-Fk#]�� M�]X��{ v�ڢ�������������OF-��i��8g�K�	+�(���\W~�/�*{��H7�L�>��#;�x�x��������F�����g���M�}b�H���nt�Nffy���Jf�l�����I%�����z�g]�f�<�M��Ɉ�nn֎�-
8�	;'����H��Q���Tj��GΞ"��C��*�,
K�}������k�UG��܈��Z�����Mp�itī!4������i`���@iW��uw+�?O;�Y�RT��B�3ٕ��K����<V��4��~2�����{`���X�8��a��l^xp��>�D�U���c�FQb{s�	���=�\S�f�������P<Ͱ��x��S^o����cHCu��f�r{HC��im޽����n��iu��9�|�ҫ�ڟfdp��-�G��*iӶ\���e�/q�K&qh�|�$�Ґ�-�����{la&I/�m�א�������ӂ�%8!��yTN�1}�)�m9SVv}����w;��1��kϻr�0�649v��G�>|�|[dRs�?*��������L�G=����Ō�y ff���"r��)��N5!��fQ��a$F$*���1�L^��2P��O��X�杄B��Tt�C�e��!��R�tR3g�@1Eإ�%PlY@D���`S�t�ծ���_v0]ON��p=�>��,F�QU����ؿ8Q�j\
g3�E�N'�lcل���Hl~�N���l���҂x��d�����5����Ĥ��\��K8 �t����!���u�òFX�-FŚ.��,�g��[)V�P�5�c��^���D����%4~���e���ܑ���oJ=�j=�KM�%��)yT3����`A����� =tF�^�FD�Ӄ �s���j���֝�H֊�}QQ�G���,v%dm�j��
]�`�A���j�Frsii�;u0�U������tY5U�s�Ei�����I���O[�#��ṟ6�^rL�1&�~�����@�3~�^���k,/��A��,��vY�c@�8�W�l��O�_�����5e�ELeaKQ��k�<�f�{���3���YF/xȗK	I{ N��c�5�g��{���aV<�c��＀^�/��r��ea���\�	�����v���&��)b�e�	��A��?�v�����o^��-FO�d�Y\D����&i`0��m�����u��0nHwɷ�4�ɡ�;"�띡Ӛ`'���|�wF��=�֧X��{�&=c#�R���@�q ���Yv7@U�L�m9ާ�؅�� �O���#�:K�F[R7@�ij��W���d[����_�q�ң�H $V�� 0iAZ�>�*�C._tQ�'1jY×'��/� �mӧ���zu;s�;F�'���:)��"a,f���{�W��N:�mv�����Y
	��m��B��jU��(��Vt�Z���� �S�=D����R@p�f��B�&��
�%��j�}r��C��@O�'��>��e���²~�r�<�<��R9�f'�#�C5�)�E��u5� hS�p�]d�T�JO���Ү:���v�U��'�����;e�'x
`-~���,��a^<[��������5C�'|t��c���\Jsĩ�(�:�����
�qI9���db#���W��������՜,�d��U؃VW�Z��$��1��;z�E v3�O	h�R@���Z�t�-Bڇa4˦m�ӈ����S/�g2҃���~v���O�Wp��0f��fE�e��ߖ����H����1��+���"����q��w�vD/�اbSIu���r����?�o�kd5bR��f5G�����ߋ�3�e\�<ݤ���۹���L��ԝ�=�N%�w3�(h�^6OM���ps{���d�K(�%�Fߙ�RY��Ɏ���X�^�g�N���[x[jT��1D�#�_�C� vaY/��4���A�ψ^~į�������D0t�H%��_P�B�i@�P'�=�z����tE�|�ۇ���b�/Ҡ�%��E��tlGUm����-�-��x�j+����͠��;w׊j�����l��Qj�*�?�/_��Kˉ�<vȨ5��2؄X���[�Ƴ򘼄l͑�.J���6���ߏ��]ߞn���G���L��M��B+�>�\��n� ��쪘�;~�&4�3���.i�uG��C��; ��8�
ПP�����?IX.�̡�&��c�o�^�{�΀�~��i�;��$�"�������' ca� �Ѷ�E��$c���˵�FS�<L���s߬�ڱ��:�%�WYa H_��V��=�����Òb`:�x $1�`�jn�W�{�q,M�;Ѧ�K�`϶�sK��}����\��Z�z��L�Euq8,0�:�]���w�jN[5�t��;���r7=� ����J|�8������B~�\1ϑ��<��/��e��͢�W��*�z')�DS����OP�?D�����O�L.:�����;��~*�d������s*lG��2��A�~�`b������Q{�.�х�m������ĕ��A�W%�7m�J4�ꪆ��MFM�֛��@t�G{ɸm�5c�tq����b���� Ҕ��6�|��?���k�n�b�n��ۄ�\F���_�C��H�*�S��\��9;*��S�`z��֞�����ogJ%��Q]�N��d�3��ZAx�h�E �]��]GZ=,j(�����(�X:�'	p�LQf�3��k��%h5�eYEn�Wi[�G^�2����,&�3��I)-�]Y7O������C��Q�6gU�]�|=��⬷���cc۞?dOF ��0�T�� �z�t�D�z���ֵ��lC5TK�<˙z�X���N�F��)d�U)�M&!�;Y�U��"wc+X�]��@3�w� �Ϩ���d4��t��O��B�C�]P,T�K�?+��w٬�?~G��/;H�f�l
�5;zn[>(��ؤ:��rW$��i�ul�n�UG|�1J3]��G��ivC��`A���r�,E� �=*�����r8p�uɒU9�0(�����N����(�O�7�������AL|l=�(b��v�l�V�XIy���H��˺,ձ�+�������ti_�*�b`!�i���+m.޾�3DS����k#����Iu����W:�Y�	�~���m:���� G�ia,?<���Vu�{�/�<���݈s�	�p����5p�1N�U#<xS �N^�GYU3I�-�Y+`�]!� ���y�Xco�]rb1������?�(M�J��i�Sgv�|ڊ#����+ �J��&Q����3�A�������Æؠ���?�� ҌM��O�g�O���#��G�r����ѷ�y��������Pz���R`6^V�٘�)��F�"pG�~�h/��*[��!��?�$�6
�.��9��G����D�jRo�Zì��#+jv���R��o�ͥ:̂j��ѡLl�d�M�V�݁�p~�/��&|��ֽ�)%�Q��_�]�-�-M^[�t�2�-��P��~��:�A���s���f�A^�J�?#b��vm�ºNd7���@��9F�GrF0*�7��s����z���Vx�Xid����v~Qbm���0�C���OZ�8sf�E�J>���d��z ��8�Hh̕��#%Ϝ�m�utx�R��j����l)�j�-��./�Z���f◥EЀ������0�|��D+C+���,��*E���;L�t_Ú��U H����Պnşc"/�t�~�e���ɭٝ��rmb�F�A>޺ԆsSI�`�f
�'�<�V�|�^.�_!5��d��RF���%�e��z8�Hr����-*�d�@$�10��FܻK�_庼mm��Nݣ^
Ɇ�V#¾~�>ғ:mP����$��N"��v]�lW�7aZ*N�R9yl�������j�$6�+�B��a�&_j�Y�wB�g�'&�߽��~@^V����ҭp�V��Ȓ`���])��V0K>#��A��i
� M�R���.�'����Ҟx�ыu�M�j~����vM�����	�ҏK�������!^���I�ϟ��.)i��	%�k���G�8������-wI��-�� �@ǔ:$�˫�ѧ��"'7��H4Ewcr�#.�9�1d�q|��,3)��֎���\*�|է9��^3���H��60�3�x.�<D�c��k�UD�|s��%�3�����QX͊ݭS~Nvw�>J��E8!egG����=� ��<�(aGgδ�K"N�(~}��7�Jmᑜ]f�^ƘP���|L5�_X��U���z&r���@��g4zf],���vxB�C�8�o �2�h��k�E�.+O>
%`�)�	��n����j���T$wٜ�c�р.�r�D�#E���̧�b�L��,@�ӵ0�fYw�����?'&�gv�� ��]V�zz�s�8��F3���#:��%��+��%��79��~�&`�y����F��~�|�>��?BIv7#��E���4�c
�����e+� �I܏̰���Ɉ_�&P�p���D�mF��io���~�J¥u�v@�����K�h �\��[C/q�)��ᵂn
�a���;ɀ$�Y�f������ZiX��G�-�cJ?1`�r��el�Iu^������f,E�!?����5ioR`e��A+�9%�U��wV<��?�F3�fד{��\�n�"I���N�����]��N�׊����t��PQ��� 3U��ѭ����y�,�$k�ȵ,�=�ݗ�
y�*P9#V �m쁃0�-^�Ͳ���ٮ�"S�y��[̻d\W���N���ȉ�p��
 ^oD��+��A�<�ۂe���j��j�ev*T�ִ�N ����{��\}��YA\q���&���Iq}�T�0��k��n��c�\�q�K�Ҹ:�oю�"�T5��#"�ut5}����5z���O�b�{^ܠ���<�.���pe�R���	Q�iܻ��a\��O�3_�����vH:T`�VZ�"X���?�9E6��-�ſ�5*-�Ѐ��OM�x�74�Q�l�:6��Ǌ�ι&���ΰG�W3mi[b�Gu�����~D7��m�F��U퓖��1�|��1u�T�wY-Oկ%:a~���̠HL?�=�ry2�����c��r����g[��̓5Q N��<��$�v����\�����UɌ"����Cl���똋��nK���  ��W�D�AI�h�C{�1�����9k�j]e�9״�����ήIݼĕrX�	P�@��~�1��}��\�T�m*�Ie�}p����J+m�`�z�	�4�oQM�s,���T���=�7Cz�R�����r�C�_����H�S���Q��?��ڶC�`0��Th�gY��*�i��搗+wkܤI(�l4�r؇����k�CL����e�!٦fcZ.�v�k��G���Y8&���L�4·�C������^˪�[oAڤTԎ~4�9���~`ΔC/�������9
��⪳�ƥୃ��,m�I=���\S
�����ފ�� ƦV ,����W���}�=7���"V).�s���F�	�r��������;�VH2��5ṷ�(l;�H �mf��L��0�ʂ4<�Pe%s��KR
�>?!�Iqpԫ��������ܱM�ֈjJ\�c�\��޽�<uF�J!����~�p��1�W�o���X��[�'�-��|��rgn�{�Xy�����u���q��{����w{i�T�,�Teos�dc��i"�2��H��X!RZX��3�~�*?�8\Y�%��� J�������PBNсc�.;���&yO�ـ\���n�K��}��0��5a�dϞ�����<կ��{��'-�'93	�Y>h����ςQ";,xg?��5��Kc�����N������������H�Q]�s��^��]�����%(t�����(Y{�&���A��75��r��m�K�D�eo��1Ϊ=���:�K_Y	8�"��S��^>}z��~|%2`3�?j�R����>�Nc���L�O{3�hYDG��\.�aK�F�҅� ���
�۞7�΁�k�#`a��P�F���6�E��!��[p��g|�v��Cj՞�Z��k��kJ��J!r�5�č^��T#�ᘽݍ��3�73ppG�(��['����y6��SkJ�>%��� ������_"y�!ﻵ���"��h��/&/X�Lv��+C\�cT�H�(��$Q��/l�`N�dڪ�gZݿ��Y���X <ſa+�`8V�/eNN�&>��&BS�vz�E�����|�>�~�jB�=dD�_C��O��rg��B�ʋlZe0�d��Gq�:���R�<�I�p)D�B4Pt,O��e�dRNK�-{��aA/F�d��|6�Ug[�YFܾ桅�`�P��պ{p+R�0E(�����������^W���{p/�:P�O�
 BM���e� s>'	S�O��.�:��ѱަ!�~�i�����g�D��s6��9I�F������Ջ��g쀼�g����s�^D^�c����Ų^����kP�낆��lhY|3�]�&�c���	^�1��u3�>��u��_M�!��M�/ׯ|>`T�(�f[]�Im��ϔ�)�Sv����g�0��S}�Mm#98�jۃ��T_}JI�C-Z;��&a�����-��N���2,h��o�����h9[������P�w�ؔ4��7�uZ"��a�6��c�`M�{�n�@�A�~��
-�]z"b�l�Z�T�pa����~䴵�2��|=��0�_���
�s�]�I�#�c/��Et�LD
�j1u�Ԥ6�s��Y��wr��?��"�l�{�͋-���Z��Ÿ�i�oU��ǘ�H�(b�g�ۂ<L7�dBN/c�U����ߖ��Ǵb�b5��t��mV��F`��A1�:)�P-���y7��m~Cz���b�:v�ɑȡ�sSR�n/��aI��֭�"�yz:��tI�(��Q8>���"u���Yů����A{b�%��,=��-�Yu%��1�&�%����������zO��)��O�,�o�վ���^۔�aw��'����)����������a�.A�j0HM�QQ)��e��>�6f�l;	TI	d�á_;|tZ���Ӊ��`
x�h���p�!<G2��Q	a2j�ftf���E=DX�t�B��g��,ˀ:k,�k����3�Dx�n�S�=���h�f�,��)Qh��yR�uY�����:3��?�H���A�\�2-��8���4ђ��ݞ���&!��z�9~�������41������*Q���:݉�_��g�26��({��
!���v+����'�$�ly#�A�ZUZwP$iiy���XU���b�P+��8 ±}�����{��Բ%��Ԅ҆���`���I�X��#�P���l�=��cG}d��t�Dz�qV�Uh��ZG֮p߻E����[�^���D��.���3�~��0O" �2�)q�� 1y�k]�-q �%6��d4�: q)��e�AD���,P�u��W!�%�[�3w 9��Dr���� �$�Kي�⭁��L�;����`u�V����#�p��6��ņ}��1v}~�����!��3%GZ���b鹊a���
�n�*i� ���u/5�1�W�h��������C� �+F:P��*�~Z�f�o�LZv��Q��2�U_|�|R����r�k+����Nx�.�t��-'�/��iI��5�����o����-�ԋ��U򎑪O�.K��)� ?�n�O���-�Z;��=��
E��A.�1�y}�6ն]F*E�[a�p��F
�Ҡ�ܑ�������\����|/����{�>UҶ�T�҇X���a��ʓ��su0�al0��V�