// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:21 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PCmmuAGK8+fsMAim6A223sbuLNd3L6bpjxZh03LfmtBwS/cqmb/zvJmwl2X7JHcC
JMBIfGCH+gxPx4aZsK565VoZlLWCQwWZ31j3ha2BhM67WT/ZJND8DECs9Aj3oCHo
i1hmoz7tSlDg42dJFYrqldrv2Es0hHHolAStAbcotiM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5552)
dmY25DSwQlEA0pYm2l4MIjrcDyiS0Flc/wIVf6wKushJk8Xy2fDnUNce3JigxZNB
5og/LQTyimRJC57z3ndYMl5Cq1ttzzE+Mj9BnYCnwdU/1tR3Eq1LQaBHnjn7rxA/
2GNHW3wFiWqs79roveTuJRqE6jzDM1MgVA9+B5YzkEUh8NSXeqLOUwOpf4yW+h09
mrBwj6fNYA8/pnSqsMMCgkyhoqfBtY0HmOPPmkeZx4k9amns9ozv+wH0TruEqWxi
cVOMbGTaHOG8EhPbI9iei5F1/iSlDtc4HWrqs4qm3IjPDyG1OWwFUr0ZFRCoz7mj
JbENeUdewOdlPth9kCEYFJPWFND8vXROErz+dX85P/y+9DsVLpx+n78XoxsOz7es
vYEHuwj8Fu226ogC04FcsssKSujL4QSn5NPgpsLsGIVOXMWJV7ZaqQ5YetsW3XFU
QZIqh9vFB7YcdN/ZJcLcmL90qlQ109OyKTUPxTCjBQE65EYTnLxqAaJ5E+yfRJuX
X18GK7/gJ5KUDlE3T01Ke8xzqSgdE+hKXwlADd4zgkvMy2lEXEU9YWxcR1pX1TOk
vb0PQmYNYiIVh0OQtWcRbvVlUtcK7wQ5iSSjpATO7ii7r2712fBJTswmOhYUvf57
TraDRGUp2pdNTi6CmPTp6dXxcMdfPFRWqYGGT/c+kflYnQKEkvgnLkDZhQExQE2c
LdAJ0n2Lqqrm+Tijw9Rg1MHlBsQENInw0uha0ZgYYpHAeh+rEfIz1zBrwGbOkdT3
3fkk2nGGdp7I4HQnq3AhyGIPJnfZQee/sxEFQztPDnXW4wvzSYZXfXpwI+64q69F
BsEby7NT97yEka+zZqB233/SuIsm/FTUKE1p+xCUIkG+jBl1/ykJy0Jcx9dC0IvS
aYGKbdgaY2zDOBtLgPurAvZVidq3zZ7pccHd88EDR5HLGTMTeq/Hj9+yRxvC+T/D
o9Ihll7yssrz0MnoqwvgEW9WhqBMhYhb7KN0NvC2jnB1P6oMAbLpd0b1Qfsel2JQ
laREfnoHjNpgBfdGAqpKEjZ8I0NB1Y6sCZumxTrXIKwthZkYdzY+1m9rLSFdhnmf
wPAIZ9kjhxP3PQDkQ6XFPyjb7OYukTd6zlsdCDPGsW8akRFrCsvWOdqOx4laB0Zt
WyeDbnFWJDbjAger6lG0SLE9qNoudpSMCnv4cCrjIyZnDpBuXtvvuqv67e600AjA
q0sqnfaPrdGzRHQz5Hfc4gNvhS2Fpp74ISHJDU/7xywdQFocmJBqARSR+5p24jM/
EhNalWD2nKoDGrefn4xzHiRuMJEwOvZ9TJercr5/qo7OzuFklPxnHj6pYk7565TN
7AE2Fs9ozbk4sxmvi/eJSKvWZ5/qKmEDSlyn6XCLeJjluba+Vpa1pdgwjUjl4tU9
yMq3vu9vmBISHyLglS4JaSFAnI+eCIceraSg9nDsY2JN1yZ0pPVXviINIACoMZ25
NJTQgtSajpedE97CwHWAy4qwHKBGSsXzh4ltMPs7qV6QCovm1tqeS29OnRzDZ1be
GOSHDpwY//rTL2f8NpM0mmAWs7Rt90B7uwRwrHGemVtYubx9v7SHHvVTPLJXUIVX
jg7T8MVdS6URx/lQ198mwNe9+rIhXlvO6fHJotzP/G7jmXFeUTFyVFNamwFgq5EJ
2pzKgE6h9UQPImoVq2gxZreUeDfr8rkg/Sy+kXiqD8PkH/VqI62PZkl5viWnPhym
O9J3FIzC5om26FF8fPHAqC3Mh/PXHjmqmeO5EbELnGpVFgjt8mcs0rXbisgz9pu+
cGZKPIhynJos+CNsC/jnxz0X8MAWP0LbXexw9KLOy2+wfuE7RX9r+4AxVXnhzwPF
7NpeJmTdQ2SD9bytSmzNBrHsciiPum0IcK8vXMisO7OvNefdst2J9tpW7awq49Zc
5WX25BiGTdQYxgvV38quEnzfyfaBudzAzxc4QkrF7bwi8JeimPPssFl41trJ2zV3
3fNZJP4/UOVxf3clXXxooq4DjCGKgXZQn9dNrqvDs6/Q2w20tx30cMAPbs/2a5dB
OL6k7rZ0qv0Ci6JWVuWuOZyMG5mmeMWgiESF4v0GAMZdfIMBJeuOuYsH6JZc4Ukl
fMKldIl/oIus0bC7ADN4UCqGG7HynOs8WXqyfaTh7ePBz0450wt7dXwx+hgSk6R2
f8QlrjKF/SITmsqanLTvZsQqTN5JuurpZHG2eBq6qaNh1Hh/2EtF20rdOb+VoYIK
L5etMqb2KJJW/kGxCQYNx9nyfWWKUUbW0SE+m9+yuTk0QB6btfUeol9SXzKoWDOT
fHIJxhPFNeVdCWbismQC92ez25CYZoQRK6CVpcY8HKiH/Z88cWbOXBs56HfwzEqo
iD8Z2NqcftXgpSHNhk38WYXCCx+eIQXaY/Vd+z3KWyrb1ekR5MEs/ydKDODEcvj9
FQMmeZKwIXnnoOU3TZfDdTHGiB5AeHjOpRuAi1gnEd3rVV3qG4E+BD8cmnp1xAsT
eq0m+VnTp/1YUadACUAOMeg/zmxirHUYewu+BEWQWRXsyz3lyorjA6wUZpGM0z3E
7RkCQSNi0FUF3+nSgfuVE5ZB+MC6rROxV2V4MJpt2YqZvtZUe30Mw9ubt7w6G/Uz
Oxsg97EbSp13grcpQfy7XkPvQCEAiugw6hLSPQObH0/VO8IWHC+UycuyeD3PKK+8
zyUkX9N4rA7n0NBAJNdva/5slp75dqKLDFnDOkNykN2+zAiiTis87Ry5vjw80fo6
iLKxEfQClQ3bnbAa5UTBhjoM2UpVHRfpPlYjOP9yI+Sb2NzF0vf/uE3WEZJyak8b
VXWLBcuBz780/SVrQgrk3EmB9I62cKekV6BlErPQSdub175P0aUgCfpzoWvMfJvP
oBwJkkaCqVF2J6XVMOo/tt9r+Pw/R+yz3+TeoeROAs/C7zSHn7NdsbQS3+t3g8Bp
jk1jCytosGT/f6O2YXU3bQ7xG0qBIO9i0kx2raIDOM8ygX/txkVcwQjbxZzrfMKw
snY2ytzQjuZdcuaNsMTOIa/jI1qviWrfgl6gT+7Gx61AI0NaX757pOZGvCzZJRxK
gETnsPjImLOpz3osS/OnluAOOn9LZQdPOJEVUFvR5rirBbwIx0msZV1tc44X1Eq+
rzJpwwy8UWv6u2hcWJLWa+LO+xjUDLTlSKT4VAYLsFMqJZG6/o+vjeAy9+XPMmvG
VbmfsFZ6v8/m5kTXhanXteNjfZ+mg/x0TnlmorqO+Xd01m7NKbftNl2KA3DI+fj+
DPiZ3nA9Xzb5Rm80kZevlyz76pmKhIG1ngZqnlfksKBp4V50hPfqx55xwJB4USX/
7wmHvTMSCqoANcMPcVlqM/TbCMdJeASUqaoYoN2NTmkokWtrIyDkQBLmRTh9uyHf
k5fgXi5uftXNn9cELbtkF3nd0PLdEEJkVss5aF8PR5UnlrvcBfn7eTtJeD1In0HB
38SjCT0baSViMjVDeMaunz7jPcJL0NzPsYKFodq6GjnBR1srG1Me+LHSWF31v2hM
zFESFOVslqERUnyvmCziTKE0DWQlus+iZmB3kguwNwEsmJknYnwNww6ec+k2ZrQY
bM8hrtNEBqcHDuCGzqnmlPtZaEh++h6r2il3jI39UtsC3Rvv52RC6RYJuIePRUCX
3v4M520gbGX6MOA9A+uRP6ga/AQMN+0XOYuQcjn4OKhqJ8Oqf/MjC5zu49fxReuN
Y+y+I8+ApSvo0dS90qUNOwCp4LpDhVJbIDDS4u1pdLHh17jmuxUXs/ZCUp5lHmcf
LNlNpCDuWTAR0mLM7z5nIs/S4eqWjBf6rIxecNbXxzww9DmtnlyU2Qy13gZPhOEe
bBuvDZf2+AUj0UtjpVdWgwAQVD5b+z2QC2Rn0HJXDXEbCE5B4gjKbJwYN/sjWG3s
51Ec05ycA97ZnKkI/a9WSZs9K5AbEpza8x51Av8HvuPsiqQ8sD05FEh2bXbim66O
OfQF0i0iJ597JQ9DBt6v+KKp1qfinw3t4eApo794LmXP+KkC0ETIaHTOQm5OXqOM
RoKZrOqDVhXIVVYickLcTC82rl76sX22K/vgu0Ij7gSz33d7IJxUiT/mYcz2DapF
hIXatUF+4x1IVCx8qToPxilqIV6uTw6LewBu5W5CKtLiZ9tUZ4CIehyNDgGMYLor
MPPLdNlrVdVJvt9IFTJjqfR7eI+ioDmevLnHspENJRPz3//rfz36Yb63khoJx7Vv
vyCC6kQoBSWipdIzDahl9MO/VG8n8uIID9FXxk5NLhklK6nsBoJ3ztuK7TpfsVJ7
mdN2lHi+Nz/pVK8fqG2p+tzqFKo9yqtNXWmLm71PFl1oReTWXH2ZgA2uYii/WOdq
kLTehypzRQRIiPysWSpsqofrSsEXgYWBxPyJOpSdGVdDN8W6/hzde9VjR2KUEB2P
nmCMgVrrpW+AZwSV9QlV0O39impTPhS4kf5ct8B9+2wi55OinbVD5pDKVAXhYlTw
uHWzkSA2JezZBabUUHjP/lfLDQ8VcxlIvAEz1BH2LKH2tvJgsKVsLFtOf6RxmDxN
F63XrTWJMj9QDQK3hFYjeQL6OvwxAKtdzP6uw96p68Wwz7BdRm1rrpvi0HBFrOPg
5piNKFH/LAhqESBPz6sDOJmI78OTMICyq37RPGcFV1h5gIWapuFQxrNykrN2Ufub
TjKus4K2E+ObnlPQPeoZs96yqOnZKzNi4OjNPZrMFB/aL2dIsCpXs3SbfkKj9wl0
n5WaNJ2l8qmtzGAmSLUtcVBqIs3E1zEr0TWlMO1xiDbGYXXCCb3i/nMbJXJwHEwq
veoMYrdG6PCi9fQtsZIHVSwECF5+7Cs5gkdwnQSZH1zDBm0RaKeAby7MGHW9kkHZ
37AvLzcMS//+NuBST1o6eblimAZiCNrFKLwQta/tjaBGWNtWLZ/Mit92tC/Fjn/2
u7ApHPfKZuJ6/OsC7HTtxnMjGCC3a6+areRWZFNZetFWjT5cvyGukKB03SBUagwI
5BzAJGD691/feT5B1I5XNmkb8nD2/Z2V0wCIpdVQUvkjAqG+zyTKJ8z/r6cjsKc+
DZdnE2pIa8CFK9hIlUhY8tAKVBGRVecAeAMHGiciXNNG/GZd5YLx9+26VFev8jx4
2v/bXORFTThrW4tj5Yeua9NVL5eJm378HI0GO51Kh15T0kvJ7eYJbosLIgJy7HJT
FHhK8O26evEN/lhao+yTdVarakqX30h48batBh4w6nPJYI8B+7Bk0P89tB5Qpvjd
GxHwuzbpV//nyTJS6iqWTfHktQFGcrmxyYHbRmeAA4kLNRAelfl1eR5L9WIqwRcF
GbMeSi4CJZ/9J6HPAyIqgfDeDQrTb+ePAv6amXWcYSoWYGJ9AjdgnM5QpGPIiqNC
Ba8cF1Ya4T0X93r1asHVBkmJwm3d9CQGJzCWsDLCOOdnWA+nB2N3vNilKzMM1IOg
4/fIhoJwLNjZT1K8s+ucWrJc/D4dnnBgSRoQZNLWpjBnKJZsrKuCvAa2CHkpJ9SA
LPkMF7/hNrNKPI5n+e9OYwbve2e4wS4dcSUbNz2B8wKXdRtwzPuptTCPpeWSJWtT
AbJ2eQrzeIriD9lzfh5rk32KHuBtziTq1SnEO14YYGZRyeeAe1Fn959R4N0zBZri
g0vkejiM7nVB5jACtg5LC0pt4fjKcfsmBlNsz/yNsjGj9PlDZKyNFqqnjyZORNqp
fq+18/q1l31xsPTU3BgCJNE8eT0nFeKxOWQSY77w2fVYoXEhzc57ECiCzCFVvhCW
Ul39suNOjoKAqt/vUcEpy/PSJ//Fzj5V/Npte5BGA4hefm+8Dvm/ru4NVJRth78j
dV76us43bgaQijXRmQ7lLEyOIzcdOBX/+pm1IWCK6+U/vnkcWTBpzCMvYTCV4A+S
X50P/mdoEnKJoa69Pzt86T/g6gcSjSOQ/Zjef/8Mp5l3u0Ms7u1vcMYSiiTytY6D
xOE8d2b4PYUqIerva81/Fn+fvUVbNvBOd6cNBjm/PhGjtKohnkHFYqP0+uJjZnfx
iAXFg6P+YLReCXfoCR/PlWD4ty8SZEZm0MDhwN43XM+YqTJMFhPm4PC1xQO1e7t/
mveDNJMxukWV7U4yyhPsOC8Aw5NKnd0d7FAN684GtxAdYF59yN9Tq1l5+UmP7rD4
t2YQv8w3ytWsANsIoJxdewi95MmkMe2EQ7FGRtyUJuMlNTnPaoWlGdhEz+x1/QAw
etRkWlXdMa6A47q9NGJUs4qoOdar0l5M/L7tShNnffPw9I86TkNhS8C5CKP2Z6rm
NJG8wS+IwNh3Qx1wdmUpaVFp1yCxCtsBB5NQfNuZNO6zW04RNZzIVYgWbDqpB9v6
5mbHUoBncj7NYftI23ZAdOQauqj72Lz2afulXIdvr2KFIddRbTgtM262DK0/FBSm
ryZK95GwIFcahndA/i5G88Y/6e/MY/v7cnOwziUSWHAgfXeTyiWN6O3rDosAAy8l
OHilvjOfUYkITp9FY9E6I6luFNrnkdjJbyfG7sTgmdqN9p9Lp/FwiU0QT12/Jjz7
4SR+F0lC0o3lLJcfGO8ODOzjebNwppOtzpXmYYbsu2bglvfKRifDcmU1FVTCVV3X
gQiig9vZ7rtkUmEcPg1bczbcIPPRxniZ3w6FkzT1H2Q5q8kBcpbD3yWlct7C00pt
bkJBbnABO8o0wz1ZqVgy6NWDxYWOyzxQ/WLpbp/9ujNEfo3q/g2ZeNzXQv+1BIER
c/aQnKhVs0FQO2UCjxMHAr8cJhb9tA2xn5hrd0Dwq0B0Wdme3e9zRmDW6Dt7yGYf
YWG6xR45/KnkcmCyXAPOhtlpt6YaOU5BJqWMtqwjswb7OfAsi/n2rOqTr68vnVFJ
d8otnn8tEivDHYWFWJ1i00JS3Bt9qx2Ks/sAzqEAtNTkTt89AnxaYm6AIvDf6/kT
N9mB2btGcUy2QavEqYR/X2giXhd1jo73SxogmNMl6kJsa/o2ZD+3bEUTH9QtZ2tq
hvYtEbKptrXIF8QAM8hxch3CX+xbQ/WVKG/Gkemmr9hpIm2Nb0xos5sWUDIQlSKn
tHfQvtNCDeFcEVUf1LKNSSUHc9nUWId4mWDdC3gaU7isBppwShDTGMBTOSxo1lQ8
yxPO9yrzVtYD2uru0TOfbFv8JdXb3bR+dvFxOGtknyOQQ9Cj70ELEiDFmEjUweQz
JwE2G7HvUxSab4BmrS0WZCWVrkWwa4iJLkW0sqDBbk5SxjUosfN9D5MSYl6Pf8TW
jAerI5U/dPpNWNfF+TRyUM8LUywNjCCnH0LvtZMnTx+N3Asj269rlvQwrImElPwb
veSdUgclOxj8Zle9ULQSSdcj7IjH6gJwIvgWTgqdUFAIjRwD4QE9CNffQMCqa/3b
0v7KxjykvzuEhjD2H5AinTC4qDsR394t2JqkTlNtoo8=
`pragma protect end_protected
