// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iPz9Y8ARKmvQ/sSEXUDeial1M/hWa/hu1ThRDZdxetHQ071DiN32FQgkwhpfMDuO
GWbjxu9NNJTDTjawqnOMekVcwICsEKLPZr+boV1pGBfpnl7jgINEzgtfvoRT2nps
XOsjQAtoNlIKAWML9G0qSy+2adVsuMl4BaEDBB5SVCk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20976)
Uh0MGGw3meF1D+5XRFenJWsLmpoC0ms2gBvzwY2gkP/z/vcUKEBuAZc7ovD5PPOt
vsVwW1F0l8TjFAgqDwlEhI3jVfQq6y1VWxWbCjxT1j1i73XAZNrMt4PQT8Fmz9St
/Ij6xiEgPJjaGSRowdU6QudmN7vd0XStBFpzfWuljz3EN73SgFiyu+nZ+/B8azeo
gkcHT3lJTFs5uVk+b/VUrv0pRYi7Dpr4yaGLODLJyI4yBhnQLX5K1UJBOGLW6VV5
EGqMYL94dC4amx1dEO8eL499SmsQ0gN+jUtXzOhNGbeiz3MliQsvJweFdDWrg2My
kuKbPubzPrmptXCgEc/jyGGfIQfOw/t+2TCswfK4Tnmg4lCVER79A/nqA8YrZV2w
QtcZLLiSeNwUaQRJZSZzLeEngdZlp36hhiYdR1lbBEuuctMjd+/WEyI9vkLDkR4N
KzKYeCrkBVFi+hFQSLiJaMg0hrB11mU3oWVbf5zq5lmOZuf+Jc4cb2TtRpYl6r9n
R12qeVM3e5ULfvSm+nOeBipiZizgum33HxMBPWsXj8UquXdhZ7G2A2mRGfCsiu+A
wMDjEqhIdUQ03J4KQVjbIwrMaegC1inNkkfJY5fX7UoC+xydK5qVWHPHlkeC5X3L
oR0fOTTx8BljWYKWeDioYXnH5q9DI7gTcYovRXAvWJQbpU2z+VlplUEilwWuz2Pn
obwTnqpXiBEd50IDVJ+h0bVtBCkpEnR9op7FdRUy2fccXFKbEfIx4OC1SyFcupfr
6vl1njXV67CyEsQbJVoeyAc8q82CFKaTstgFE2P2g/tx6Yt6FxIXjTY63Cvj/+E8
1r6LzvepJ+jVZQes76v6FzuxN2AtKn2Jjn28644QTHb9kRDjLkC7qvSGS2ZBiuno
Yj45j/+m6sxDW/V8CtF5qO3jxuN48Ugw6JhPlmneUex0NeLOHbtaJvmQYn30pWZ6
HZ8qgqOikQas8nvtidoaFdV8LQJ5hx1DrjhByrfrDOEVMHMgUseGnZuH8KsQMkgi
kPkNlDjjJM/oG0EHuAifqT/0QZE6gngeaNlziczD54ryv22crQ3xAWhrZvxxwvzH
5cMZqIP5s6yfIAGEzWC8WXmiVD2oKdbFsRSl0eztERYrcckhNO3SlcPn7AEVNDE0
OpZhWg/ksTEh7tajEmaiiZGKpcyK3Qq/oa6LqSuN1ke3v+BkCMtHCZNZPvsVPGn1
cIhT0zqgv6czMuSPRKUrWKeknVBaNlxPzxQUCzFfW4ZQ1V3Xojd7xn7UknpSRjkv
xgQVKhVsq33fQZNugSw01Ln6/X5Z7TPA6tSsfkBm02liIoDNdI56LHpN6tOowCDh
vnYplA2c9amJZUUedTw4uE9Urs5faNmUDaRfd057m5is+DJVOhklOrx4CkDduzNF
DsqiHAP1m5XWEE117CUnEvbuEECVv+Ayd3r96OiV87yvCRia4f7LFH5hCaymYuEV
cVXgi2d/LKn64dA6G7GIhwvE0/gE48O0/UtMnZEqeJS3AYCIvEG9T3koCCm/CJmc
ML97Tzr/rvjSxXlkioMfpMkGOanMqZz7yMVWZD7TnKeIh2QpU+K0eHrm/YKm3VpQ
hJ57d9wDhKH5Y7IK8VOlKz70RcuNSQGDY8RlKkbnpgOe/xA6i+UmHFwyBW+fe7KJ
D0yxG+Co0Jr6O3C9QmM9ip8OIVsfRJ6wCo+Bpk4f84XmHly7cYARGObADmhDHsqT
KEzw4IOhziiZQy9OOPJ6mgQTicGbAiNkJlKjeL+78TsY6FbskkJtihzaQKwApUwr
V+ZdJSmuFrZMleQBsYULD045d44T70H5Kd7khQdcSFZOHLod28J4VSz2fXtWVixJ
0TVfBbTdJJlMJRi5ENimUXHfPdWxyo3Gcm6qWYhQmi2igKRDPIvLg3hRJWT43hmn
DF371vRCw3CLzuLXRaJkpaFVW8kKT0e7MIPg0VP/Qmi4WY0CHr/D9PZ3B6KjInRZ
jTSTorycroEmsJ3cq0WWrtTeRUQ3VaG91Ve5M3P/RGfwK4naDXfGn1wjMyRCzWon
MaFSvhhbyB2+bR4F8pTvW+SPkYGGX5rsimp+8zEye9kqXJuxpBfv+7yJoKukmuxZ
0+gZDXpCxhpF8fRw9ckoSq8Cq3qlNKcwO0yZ++Ja3+LXiGyCOvFCmZ1x07A0vl8y
qcpUBzuxRKiV1Yl1qXBb9gade99+V5zZD4os5moTqhps+BldGULZO5xVz2K60VEP
NQtl1NlmEz1oX9JFe1a63doB5ep+mdUGuDy2dnNqrbBJAHmuC1ojU7tWNLVPus7Y
VIHoFTJ+F2geaWWSbUk+Y629leDFYU8bfmFrUm5X45VJpApWsRGsllXAOU3iFd6q
nyJr8fVz36CE1KjwTuy9zFX3SD7b78SfuHzngasmsoY7OYmfLQ1hAfXGBTp0pc0r
hX+VcAgsDnTdiRHuBvmlNXGejPD4NdiwWR3MWtItjmM6xzIq9i7QPxlxSIySnP6z
UW3wuBqpGjcjgu8zL3siaGsO/BUC6DNtR00e6kzf+PxeRKDOJkT3pFnv4w9shlRv
8g46HlkUUiodzOWJBsW4tUT2gTxiFF7JXv65xlj6Dp/iKe/NUspLn0iziuH5tT2k
SeoCWh4t9mahm0svVqYgXa0d6z+DnpuPM56GmeXLyPvVmRZVX+4D+4fkVHmyyoVc
aEPKRLjtlOYVvfjz13qo6HwZzrh2RqD2aht0n4vqQK37ImHNEtSwRySQPX1BTMGo
4Jy6AB3aNJcXQMw4XXW0zTiKJftCB+FLGSmFWxfdfoYIlH6AhB5Smmj56O9o/3pk
15LqOwrL7vXbHqNCmktrVVpT1UjMPq6bYkwMN5nv/aQ72IWzMPq/XZU74ii10ZBY
6F9CBxEIleRdEmZ+/9rG5GiFqGspPyIDyThsq3n1c5x8kcZp+VJlGjAt3dppGqbc
VZR6CsstZ9Jm9FLKpIV00wksOPL6uHeZ8BlwZLImFq2o24babLUV/bBzJHlrIL25
wcJXbKn/DsGwD39Y+CMmlCYBDiUkFaYxnMLP9m8RWsygqYGXTbXAz/NCsijwsBLs
acI4JcZyUKa3dKYLrrxfhefUSBxV8uU4gvgHsZcV8SpJNqwTY/C7OJJF0NHvhMB7
KivAItZQQXJUO9cT1PB9gX+g/Eojzp1xc0Puslv8G2Bk9C93pggEcZ3TZBSTXGfP
Oo+pLBFwb04ztECKJhw4McJsbzswhG8BHklYtibfH0OpMPL+SpCp59grUwSJ+nj/
BQ4LW5WbWTDYB780yUYMg3KyLdVLIDy504DcH+gDO+CilevnkG3njDLxQwv203wm
OSitUSnrF0cc1woJ3X0V8KWH6LptvdB2TZHsP7++DKWmE5OC2hZmqay22r3Go3rO
hiQDe7lY7h5axiO02vtQFWGaGEoobnw1BW7Cbas5Bc0VeEefIE5blL9Ox9MwUMA1
9aVtAwds1lzFNova3VKMTZvDak24gr8VuAsxn4cCmSyTWezXa5l35q4pPqb5dJPY
bHeiObosQt6S21LImsLLXenuN1ccFdw2O/E4vKN9No8J75DFisYAK9TszO/ZRp2R
DLIgDK38unuhd6ECzU+wv5xgEzDmJgkzjx8ENSGAUMeoC/YrW1+AiCEgQhFrm+ld
+6e8MllwsKp6vjnZV4SK2k1kgD0YE5E/fHuyqRPEN1onE927nkQFAb9fFla3pWt/
xhLxqNMuQ1jf0kIUwP0qoBq14hg/Lo8gDxu4epRGdQJCD5fOPnOfeOKzhDlchoOu
2zuwClQv7aDTrwsexjxk/Lqlb7Au42m+p0E9adHNWPLrvw1Mb5DDc+/cLWFX19Fx
8neM75ZRDdcGvICj9+FLRQsM87rpWoNKN824R0PQyaCM7oKMqplOzCnajQK6znOS
A1E6w2DYnlhzufX/NabJ3fBRS+Nu3ptVwvDLnPBO3/QFOASf6bmbCiugBC1Lh8Yb
jYoe+DnhKadi0tzZyFqCFH7lHkYYtQPJI4DVTIUzXjJH5D+JxrbltkP8cBRfeS+2
iexSRC5Chqd/qeCsJXQ0jAxDHtoenRa6eXqJKtVUnWyhAxPC42p0Igdf3KACTXDw
89d5KcTSLV1udeWwdjFkGPQuG7jWLETjP7n5VmIE9RKy3+Y9xK1QN5COgpAc69gD
Nd4vgvxTlH9kbT1LCpkbyOFz3zyQsvGlgb6NqrCeHM2pdfBOFSkadxEkHZF6cJDn
vT3LMu4CMZu5A1HGDFmbqCfu4z3It+ueHDjmPxPXDLzXaE5THoXtAzigGReqHvlr
/4PRCahOXJlyq9GniJUNqw9BEPfOjLzbd3j+FYrlXHND4j2Gh/hvp1DIRZXmmfxA
Fz89zwMOAkSPk3eGCQH4zMKNwJanLz0Ch3jNRnUFkA6HT2TY2UuzL0k8IilipZiv
64nvpksTjIVrbQjVA+75L13Ha1zuglD734DnExBkNtLK3zkF6/D2FHWaokjZeIio
uNh5WS5rKR/imbkzUlJP6/pERiB3QJw+KjxfAMdd1hpS4Ey8G+UBsA0kRvFWLcwf
iQIrxotkjVTZiDZ7bo50vlemInvTSgT6XlcqUeNLoVR3TgQ0vV+8MZRI1gwXYBfn
o+zrdP6bXrvneAlRrrODq8HNQqmNhYHpFkbDdHLANOnlvgYSTKoKDcfV8XULdKxl
0thk+XVLrGsUFIfqYcEXFMvgSnjwt06CZIOkpptJP6BflrV0sLXylB35kPT3HmCZ
Sy7JKhTKgrv+AE+lTql9NkNsvMSbAEKcY5JnhcAMyq+fBotL1rlhASAUnVwmvw+Z
LMzMSWszh8RaM6nrf1tF1rLj3R8wOoAgjXeFPYuwOfv3oXJymsQ6l+nk2alK/kwG
xfmtc6w8G2NaODTCwoy2vzNBI5v7hJcoWauxTI8qii+hrCVgu/QNZsm3E/62PZTS
SJq198FX2D6QebFVJ/SRSdcI+y537yhjdMmDIb1DaZNo32A/7dPPQGBKNkbPVowg
0UDzXBvyUyOaM6PB0Zm6oGccjchHznrw1cnQNT3gAFOV4H2a6dzNcix4r4qZiRFi
G7dpL7R5wmZON9jOFEBIfY22Wxs2d2swvyqSIaC/ZvPW61Esz3EW+E7BS7v+XdvH
Cd43dKkj5SXMQlikW3EkYq30exWS0Z+vnP5rHM3j9f8Q4c1db/3meNNWDnYaspab
WGhIv9E9fnemqa3EmRkNxjpdgcLSIN5qWydF/giiAQRwiDLjKsGUwtgVatLYEaKM
MdCozvWlxJuF0UX5QZKD6V+e0yjPk/os4i4qmLd3zYSagnGkVH4nJ26x2VGyoWRX
l9vThV6W5kNwYXj0jsk4tKQrx5Hz35dALxSU0sadZPnJ9mUhKy2UTE6vuCQ3OljY
Ri+X9z7+awWq2zXZbSymW7fDUHbKuyfIB1ky4Hf9siCSZZRM1xy22JmIVUGecdh9
JyPKZinRYbNpOXjAXMHMzP6kXzeUQanyC+qgHjvrcVGHQuBezDtWBPIObQ2EHyMN
AOadsFOSFzWEKxvO/B2sxVeSMm/PKGhry3ZacimFVFnjRwuRwEQ1sgtX6tYTQJTM
bZ08CWrU5aWiZGNFy7k3QDWfSbGk2USz6c/buxBsRkB4PEiM3SZ8oxJ1slnU5JR+
QCSR71+yzyOenjskcXDafEQtsNMLrZFPSUdjmAkffUbLmHlezuPh4qcwoX5I+Yoc
a+QdEwkwhYFBWCUsOKLOKY29UJLHixlq71G0kdhaPdNZEQ+6pKPM7V6vh8DXYDD8
sygAc8UlJR1Ca394j51zSbPUK69THkcNx+DffljJxy4rUHCypgutxWk22SV4yqyx
Rgw9lOh0ett234we+ItPYgtw1nND6WkbIBQJVj1/uYcr7dGJ3499JX3UjFCzZ6wJ
1/p2y6PNw4CngRWItn2N196BKIDy1ONKUp9opfPjSEWevvPVNN+qysn4YwrHCL1g
XhBS8bEBJB4nF2Mxye359X3WUvPr2I4NglTVvHN39+Tsh5TqUtxTcDcPKqNusOPh
cu3wabwscXLHtJxH20d4DDNOxOVirRX2fXsSId/DS699zs7j8aFP0CyuVYihCX/J
ryW1kv/ZfWGRsPpSp7gGzINW7Z6ok9vnB5EeTG8kuPAv7uGGlrokxXnhgsuGZVUB
yyCG1I58EP+kjo0KjbMWc3XCIjmYO7zuVSKs+QMTDFkRUlgHcDkycvZbL1Vria5D
07BGCdmsSZR96t/fgbDp4fUVG65cHhz3j63X4o6B9AgYHHtY7gBgvllEOISdidrE
mcz/KSAl5inDPqbw8/5oyIJuO0yKLD4ZQK/33DKq4xtCqH1gImYpgyKaL7d6XVej
Y3ATUuGCbLa5a1dJf12G/dm09WpU2RNfko0yCFWGOirvPjD47HY99aqiqA8sXMZM
suhkyHQIDKpbVu988LQYKjaUstpB/5ZNBHF5cwK4LsIqHacOjwJWGwXiuDyoh49B
NS3AlGIbxdSU4aK5E8Dei0TCW/aUzMkjtkgtzZ9ttsQ6T9pGWfKIMHAFsq2e5GMq
LyS1glNtPzllsuVc7wRP4hk6VyuVTERUl+Pya+0OxgMFp2zg2JHvVVovp1hSF1br
emC+4/SsYsuoZpD3jsiJ6QEKEWmtqm3n3Pg23cxvfHtdJf7qy2XrToQzZXxi5q8D
qVEbV4FjbHf43GEP6kE8r8wnhx85VTo0Rjiyoqw+3mwJVKd5Vt3NZfMj4EtDt7b8
WpeQpWVF9wy6TdC/5SMtkFza3c6GV5iJdudfb9+E2G5zYRNOiT2KKkifXNz45z+W
WnHq6nL36Y5lYph7RjSqXUXhl8SZimemXFpjAvHkZAUcU/+D+IUWYQPrLeq6WfNH
A92TXYhd+8Suob35Em0zk8vfCaF1dKV2gsyPxKmxgJM4yOTJtVOx7W5/MLrcL9e4
p3msq+99IotKA3g9BPFZMOjrZIwjwpfWs5AKD8ilDvEks/4iopAtN2mR6Uqx9/6U
4v2VhXAtGRN27bXGKJUPNz5es7grRttyHWmIxDipvP9LO675+6sRCuVd8807+Z+X
pAWDpTjMk6dLXZwO6znHFER418VXY4l6uVghzab/n8vOD8mpL2/Kl2XMVXmZkveD
lEOLDiUCIiReuehk5lo/MWuWkk72M32mlum9juLw461VoHgYivDD035pv2oc1qKV
qXs92gXra/4ge4YJbPelS3/ceR3cCb+2CsMrEhie6sGGwWpaUnUfwtrz3L3mejvZ
JvWz5Up4iU/j9vXApzGP/o1TAOnzGzSnpdB6vwajSjIzooGqTmb2Fpn4MaO+9Oj7
c1HZLUiVZHN/Q/i22EswWGNLAhIo0WVrnaoKZtO/SKVTI9tnw+Bb+GmIsBevnoOe
eqOEwP0ojVJD+HxA3zYGyjAJFlaUx3oxnd3sWJSfNI15gVe22EIkn9pNtHS0o1qj
DivO1TUNw5uN1duufSe6IGsk5bwN/wdHyWR1s9Y7eWNom+nJlQpcfn2i2pPoE1hu
a5oqDpTQn8WNySwEHjOtcnbKz6abyG7Hjd7F1i2cUjnThqYKnzfNzlf67qICG8LZ
po/xXUiPEo6r6gyalP/9rOfBGJR8Y3KHcpEfNxmOCRs/HibW2bdTlBGkasyqTRbt
UxdjOFhtOLfg3uDkiMIulwNtMGkHxc2MbElgtk3TUwGoTznJXc/yCznJ8txtbUID
FnAzeHmyIKX06fbsuuB1aYdmGsaDbq1ooo8COda7Wu531I7FBvY/WoIoxvclX2i8
5hAcVY/GFfx/oFNi5hPQ1O/OUlQrMcUk1UqOT5EOlnruh3YCbqa57+C5xWG269QI
LOZf+9UpbGgzD1W93zm9auGDX8454O2UKP1Fs+f+yxZ5xiZ5k8XDtZ6MNQRXScwP
mFM5w7fPE/rj430H6ZcwSS+bUAiL+DgI9rvbN8UU8sUGbfxjsxjei9zyp1YWKHWY
EgHqn1mbIYVgB/paFtVWDg/xY1m3WA2YVbbiNQdO1xDjSnZ+pYDAl2+ljDjjqozu
C3npQmkWpDCFZ8NFnyAfeyJHWgMDceZzxAnk4ZAHNxLyne5ec8hlyClqAFcist1r
nZah4NJGZmjk0GCvNKQLg7TuVrOxkwzpHRCDfU8/h5Oaf9eQ05rQPQBDc0GhGca5
P5PZ1bhFYHX+y5FQsyg9fS+H3qrvH6KHOoomnJe5Lcm4R4IydAD61VgZlt8JpGNf
KgXuldDBOQoHtFCulFCbGVIH8VxO18p/at+QHg+Uey85FYoAYNV0WLtBJ7aVzEo+
jDrxgX/AProUlbD/ZqobZB7+aI3+FjyH6VcQcv9ugcDk0ySfyY8au34Re91vIaD6
F5VNs7NoQOWXzc7N+9KTQ7UrASD1v6rLv7gWZmzY39MlKIJL2qXjXfAxBG10nzsK
XjBsApljlGxaXRn9/m0yaE0kFgpgV9b/cqqUeCPWn/EN0AK0VMqIkk+34br53FAc
AR2P1Aki77yKyfT2s3M1G4zbIJ7XU/F/YVNJbV4b8YU2hUUKIFt5imtHBCBDPipG
WXBgY6dEG7DytXaW35IynAxXXlQjCISRra6MgGMo3eqrnx6J4G4ow9m6AV3tLTN9
/muw/Lu2dxZMYNvNJa+Up+aSxgy+VqTq5O/JRvGm6GoMn4ew3yGUyQvnkJ9BZ18o
ITMug6HSWSjWMGg1ALKoSG+8htNByYMB3lIAMLHSUXIbMvTv8BDjSWJ8V/PPWFGO
lAm6YfNyUCEZ5tBDvGu/ntDiUh6QiSVfqUggZc/N/Ya4JJH8j5QCW8WbXbaarsv2
Eqz2l/N7p9bykECy+td95wDvse3JRbikw/rIwmXjauLuzuQW/18KCDZfiwy2oqZB
4m/ysG4h1njmcfq4Qu6WwVgnKI4noEISt5ullwCiHHUyz5geCgp5m9C0/TsPkB/I
LiDTmdU+tcTNmscdY6yOLhkkCbM4MpBEhKWwpS/7PLP+4XxSshV6s12xlf+LT9DF
9v/IaQqvDm7Jrbd/WMAyCwqI2s2Gcgjx+2EEHEU9IAbrEi2Gdml/0O4eylALXV9U
7UT69Li9Ui4jCFMOn+xJnMLom5xcSVBgt4+k0rvnxJbgrftKUNBOHz+4wAj5rglA
25dq/5hHSJqr6d+nDVDscuJBhU9VzEwGwBGcLbIUObrRui3sp9oQZEyZRNE+oHCB
FypSciNu1yrSpLUnYuNcQEKj7vWewLmegEfJvqLmKSmfcIqgg5dTkFdgCYzs60oT
Pwuc0y+tVD5uwZpP3Ypo2vAREJ6bmrJu18sdJwWP6PuIZxtC7xqeLNjVuFW7DF4m
hhxz4s3jsKmdb2yCGV7iUV4GoRd1fjhlqrNMeBgeV1KwOfWypRv1zjnExK1sLQ3O
/Shf/Q4hy4uBV9P8JlfL4InaYBjZcGNYV25HA6F2ks5s4HobONsftXcbHeSYte4E
6OC5rCtbu1wzD+WYKqTF7+Y1Qzk/nFHmX8vI8PpLpjzf9apf8qMSYLZA5UvnE4RC
VGbDcGqoCeuU8E0fxIrdbILrHyFeUPuGZYArHieazQp9vIKVygcD1YaPrLaNxXee
FEhOIIzGj5ma/t/1lUQIKPqM6ZfZHu+53ETHQvwCcGR8akj0DElCRh/rutcbHfBY
AJ1f1Tf5XNsYOHnMXEa8efLLLjuW5H+6a9mrktcsEu7y6BBs/+JmATokkf8gK+OP
LeTBpTSZxKrqopVIbNxCTlHQ+PY41WUTh0pkMr/iezYmcg7NHE7414u1DiBZFldp
iXrFB0hiDq4AZm2aOlGPWlxJxKPl9EVcBkea8X0/cXZG58sJqks2+HpnorkcOGhC
swavSDLxlXV6AH6WuaCgwEAZV3r/j40S68k8/59SGdD21SXYt82uLyDGeWCqVYKG
JaUywczspcQ6xyxoLsvA5+XDaghiPmiSQejMLh7qOi+6WTfT7cK8QjsCdvcEthOh
Ior/unxJ2NmjNarkLXsvnmJq8By1PyRb0lfKUnA8jJtDasRaEAyczQaC9Cz2RhMy
tUaOS3ScqM8bIplPJ5/asrKuzjSfkXLh/imeGT/bKVmYcmhI5LPSHRrFlKfkB4z0
okWhPcUoEZqEYiziMdKSRT5uk4+Mf3RYkW5ta9fgkvQ/jqHzBthD1AiVUtFQiOc9
hzfY2/hREWdf+rezSMWAVBbqs2Qh013EuRL5OoN8Q5m76VNwzz6yAGHx/jWkDu7s
0kXGbA4/UDQaRcm++izzaUFf3atpOCbSMFKiGfiNI1yzmfAre49d5jEVTYfSvkvo
Zl4RiTlR3KJle9bw3OC5T6e5/ZhMakDRy7wyIPtocrtUeJhpPj6aPzzO7I/33qMP
1xbjHeA7AreX22OT+r1YP4xWz8Vnxl+x+9//cn2P28wnWLWg9qXvlyS7phbEA/fq
vbH4AzcDBzoUFOSJOZGWIcIW+pm8JWLypnR6mCW+OvWkYM48TkG1KazlJh+VOl3W
dO+UzaB671uU+HLxNHoJiSE9aAwYJxQmErfHd5RorLeaE/HkEBcz427FmR0y8lMi
np+wEA374LZxFkicYNOYfXOiG7XtyTISCWH1TyitldslbyPvnf/OCheT5xL5gC8t
VElgj9v9KOOYZn/zTReTgMbRtT7VvPSoKBmbMlBE0TDIW8t7BQGB+fPyQeBoT526
XSnNpKn9o2V2yknz/Pe9nriHuqkieK6mPVPud4ol98zQnap4TNm/c5XK2Gcbp3nQ
jRO9pg4gXCBRBsHGO4CZ4YI3kGVDBlQMbwAw3+Z9985388C79MHL6pGjHjlUzTQE
rCf2VttSqUsxAmYraPguzrfNb/q8RSkSwij6fxonYjj/2J66Lb29NrE4Afie/Yfk
RXO/DcYm1yArlM+PzmhU1mjvOeKZeaZfgRmzaQ7DfMi7sYxaN55MIVwNGEcUJU/a
jv8Q+qkzVjuR1KtuhvVfSF349CWTiijmdle72mhSF0Sg4PMAuDeGRpQQbw/nSQgF
c1hW6OfiiVUSzEzuky0qUf4h8pQhOrxr9pn/C00vjtREIGqL4wFUkNzj5SLxpG6R
IMzmsBRK7sNCxrCW5SyiC/hRMzxMQMmQWzb4XfYXlmjU59Da9xoAktlUDG3I+899
POmrrnfCW63KlNWRqWw6UsPiYE+FjDb1z1CO6GL2NH8lwYKt+aMsbCgKN4oDwJaK
VuDBUUj3CMci2FkBJryliZ5t25/1+BhnFd1OcDqZcitYgd3zmAcSs3YzkCH6+TSq
eqHqZv0FUZP5qFNOaWI0YT4Jt8qOLrkwhxLPZ/IUfIpalLy9+Z3zq3KJd6BBSa0L
Ve/JlT3cyUhan6KqXAFXcXozeDeUODTECSrwsOrPWZ9pz6Qbmq6oBqGtsscOw6AQ
e3BECgG6C5WSTKmFVZ9qo4xu+WBADzgqMEZ/tW7RtQ5B2Vou2U08gWWtgePhPuhD
EZysOI4PQMybUjmnLylUUOnfg+E5ROHL/XAvxDLtRMIcx+53vxBsCodQSt+c9gBh
dhoX6RW9YJ7xxaahx0hNRzeEdP1G2vvkwoltW2MrFoC1p4LEsPo0O+l49K+1EjAh
b+E37gvE0b0U8TdVLYXgUHnqk2/4W5Rn471HtMJND+vQgY2pcBPVDlrJVhbHGmY/
XmC5USipDHJtRWWz8Y3CfafUK7+dUGvU2VFKRo4Zaw5qpi1qfJSlp0vjfEkOGP+R
20bYNN15jgB1IzRs6YcZMhlmkRIoPiTEcTimLImcrMEPorwuLx0ROVUrGarvRu2x
yrvassmEWVYH11sD8CsrM6Y2cU/B4p5Adfpu814ggxaCbsBkrkDGMm+Wytk7VaRe
UentvBKEuqs8qtRQzSI2Yef5XFKE+HqL326/4LPVOOANMFWQibih7xmN5lXeKEgg
N9ZsGUzHxnKlGT4OmoktQ3GUEsBLKVpGLS2m0Z/VmpzWBnS52KpU+6vNBOVtTGJa
kd08WqtNeZNt013CJczGGHCec8sQvgk+05A7FIb6HBmQ2wdSMFjXsXgevX330GCE
Zc/jkdS4V6tI2rbjy/pAt409KmS1sDM6/Bfv71g7fWeMoWsKyuItmOO56r0O9ZJJ
UxfV0sOxIp/PL3ANc6m10+aSxIDqoL6EsnG/yR5xKhaI1AaBZaoz5Cek5A8sD2Cf
ChgWLdYIZUDou2VW0AhHgniTuFFhVThxGJFzMnIt40btRtf+byCeLgRu2YcpxeKk
fRzovn0oxml/OHWNb3TXcy4W52Y5NAsiQ6aaMRlx7tNV36w5jF0CvObKrp15ZEyG
HKcgkkwWPGnJdjN/fF+yFUU+YCc8uWW8g9Bng3GKLlRoDZsiCyVkooESE9G5bdzU
67bsB0+QQzH9tFX5Sby686C40wL4Oio6fvVfOs5HDY8ovgCJePfMohHIb8JRtX7Q
v7XgVayZPIUBg8aqvqc61brx7geqYACzphM7tfHWbwPV8rEiGlm0hnXI+vf0k1eC
DuuDFz5fHDmaljTMyj4LhNx6r1i+5I9aOtKE+ytqfVAOn+g+zhS5IhR85iCmAkwO
5kopw/fNUGj9qMHpSpb5PmxBgaDl3o9gjfxhlB9sUUP0Y2VGvMsAGL99EwQzoLoc
3Y8VN4LaSVfRwbh5aPfSmrEkh9WYxCLoI9M8jKo+Qzs7n0k0fenESOtAI4MIXbDW
2JhdcWuXZfSHSwHeaDVkN2qEdLed8K1fFInouPnEW8DtFfP1O8TlUXnJfEzs7cOh
a+qX1L4447ZIeD3KX2uxXUZW8b2b+yzWZx45uip8CmwVBvXdtFmJJiPrtshpluDk
SV8qGbfEVSn8OlXatayVO6ccAfUoqpM871AxmShU89H3FQffTo9C7are8cVrNEbk
GYf/QzHGynBI2rVp1YuTyWKGRLDJQ+M0QLH63CKa3QehIHwoPO5evcXZYEcWAo5e
1guCwxfreBOQ6iTCKHaWUE2Y3/U5DhxfcZttrN46HfzuHNgcZD82yNVIG4NIxjK+
6DJF0yIKLffTZ4hcUJLSCkOhlTpYYj+NFx0NoBHCgyw0i670yrAabuwBQSnPpMf5
HuqKnHUgJRSkvYDT3yjyKPWDqyjh6A4EdNF7uLBA0T8+Xtdt0AgA2xKfTqjGBv+2
t1TeHOfslCgqgi41zI9iYacppf4Ka3FdAm4clsnCFMo66Z46WkYFIjo36VxcN5N5
1wqBEiriIMNdYkO2hEn0TQ8WFq+H5oP3SJcyC8AYFnK90dyGjyR7QW0FqBL0PLLN
OSa9oRpUzjX/fZN2VXAB2wqq+N6LlhS5KFvek9lrmYUVAuu8zEHjaCVVNUKdJhIe
dGm/0L0qe9QFWpbWqx2uTyPZLOT8fgP0rLX0Jrse5wjCJn6QwSUsCa7Na0kB/l95
oa/BNTyspmqtRypNUQF95IyLAdy59ux7TmPNAIwAF9ODx7crZ2nHzYnL85gEnc8H
nlLBzK+AdIqkEpto+OmrfiqmT85kK5ol8yhvaDsb2zZps26noRQ03hATu1ymd8KM
fDQfFgVSmuglwrBVhoUSMM842eLSddgwrUIoY6gPv5qHguh4+MrG9eDSrA9H5BAR
lDtTXJYG/DMYM6MYRfa4icDV8ck3QpGNhDIiMCxg184h9EoL26Noua9PQy5ldL2o
4n0qa13jZX1iBJLThUowDRSeSTTef1bAmT6est1bjKXTB19rf0QYNlCjOYbBX91f
qrXyG/BH9vXlePdAWlOv2LXpS2d66Q+h9tnGxJccnJI5iuwV2CSBugF/slPGOzO/
siAxSfeI8f/C7xVWwWinl2G2jGst92pmtynUxF3P7E3vaDTpEht7mHGWOD2Yl4Js
azAtHBN422eRJDZcfkru0Rzu09XqGQfew7oOHHPM9n2Qxpi+jXk0VkaCCt+a64LD
MrKojI9VKSKuekIGmWvIqSTHAb/fui9yD791WC4f/cHhuYBTXWFNC2uTEGq/h7Dp
e8Lzk8LKw6LIFdqE6zeAWZBBUVM9TMVUy5JZLh2/TbKWc6QUvOOyyO4hva1lc/34
KjFNYPtYkNLt9StOMfj3JGk4F9vQf3jeH3MGd+hOL4ejWHmTjJQjCXQqSlc9Vq6/
b8dviiJ3pY34VXyqHn1j6am48mP4AnzmYwNeumslfT7Zr/ayfyjAyXo2ZVLx1Axo
Kq9W6bXx+3p8IrTohyHPYKRxJGZXCi9YK4VA5UGioH8j9dEcZNmnPMmCiyXbR2I0
na2fbni5xcc5vSBpmRLhDzkYK+ycExjbnE8rfzf4qzH+nwTuVUvk4kWXfpOPjxwv
Qv+y0zV3GTqObtnOMCIFv7u1BZGPCUeRwE4MVVz8+CmKVJHBoTJTG4JvkjWzjxJ4
sVhmVnsW+cAjbSd/Qn16UxqmjLVGdQWy2mSP3Z3gTglawGekrO/5fGz+Z/kAGkHX
RXbrXg0Ht+jzk6Rj17f28YHptsC1fZvKEC7ekFjgWUm3gWAxUaV90uGA2HaVfAGa
1kyapuILb88fUjiXCVnZKQQ2yMBvliL9jwFR5S1RZAl8vFQsuBRz9zUunUIEIMBw
44nmXAHfHyG1fdAmlhI0x5SRZdR8Fo0sVBXgUwRfoH76l7WTv5lKOF7MrWjUh+sf
zyKoFTFQCkUV8DN83DKJ+aAFKZmN9dLvOh4XmjqT+ohXWw2iJ2RMzS3OTlDIdJHZ
r+qeAl9wzI4lgZ6ZsvCkvOhB5HMhQo+TKlXowdAEoYFUkFVFCNbdU4GZSTBe/lzU
Vl674hhgJWNR/V/yh8Dlj4ptINg4PrQvMQK9Div2TNUinjZM5TU8lCaN714MEAWE
NlBbBJ9qaUyzhykJX/14vY6XU2VO9fHieNGC/Q7Ym7UzmKZaR6SYoHAz7ZiqAz3N
2RlWN8njAYsQNxjCt3OqoxAbD1zZt4H1sa8ykGQM1B4XLRHp+EF/uYVqIFyJEIeu
339jADKQYOms6uKhkhMTT3UrOVh+qIJzK6yF1RJzIUw3WX/oeQUtCyLV+enwQ4bi
UlrPAsn5wjrP4lm5LLcvsv0MosFdnkUpSNUCvEN4Doqn5XMcJQlgohS8vnVZGyo/
RWO0aR3HDiMmTLdFtpzVWo3aULI4BECmyAl+wbdxgD7lm9eMpn+pme9r03qfO8Ww
B6BbEuYu4wZsvSy+Cc0Dvn7vTsR9ZYLBTxvCUOyRQTK+vEkTXUiyR9duM5zZP5hA
MXAYsZ/6abijEkVw35vqIeaUqrmWIDyX6OH2MXoHwxRT1973K3MiBlalngBmdwvU
7ORcCwd6stTFXojvoA5wuJLUEZ5vw68lYWzp5XvZZAhpVbQIFAtXR1quvoP+3nh6
iVRZptDvXraQkeldYUyyqw+7N7SB676FP+Z0acHOMdBa4OWGfD324MtUmyO+9v/k
Nx+dunlhAuaRciiTxEhmIFvDMCZ/4dCmGmFs2IFEHjfAJ+0qRz8ez6FE5HdaJHSk
qmaIU6738SvmmYGS8YMrMb5TDTAP+EXLde0mpqirdCyy2ZXTPJkPqHzTq3jrHUmP
0FV3uX5JKH5/N2OS1SgaLGttjJKKPmGUcQcWZRe/yJy4xysodAIQEyFbyrsG1Urb
JX1jLa/JwnIpmwyIyP0Fota0FR0PTvrFjanDQQ2USjdPMeWX0GF+T9JOVcXP3t0a
nP8wTqHg4NuPjsndJamDWn/zwzSAwNSeWRkXtWFqQk8HqVxHK3xO7NrJjPISWw8x
TdP7gCYHno5Ac5nd1rlv/OtAcytNyS4oufY3LAfekWJZhIK5GvZh0Pt/vCakXabg
GUKvBvcDMzIutaFqjjF8s+vRCizkm25KXcqm+I5OTZPQegnHxCnBgxYM153sSIar
hEa2QMagjzmHs+N11A6UpEKBGAzYnQ3N0Uxp8ERPzbOGLDWecE8Ywi527lFrkia4
BNkfucrfDNSnOLOXy5RtR/5EIrt+ybf9BdTKPKyazvcdfSviNcPK15sjLbsj6HKR
rZo8/tKUSlC4trjm3GDKIId5iSCreGRSh9hjyjod8Z+yq/UYnFjoYpBYu3daoYUj
02d1QvKldKiR12c7MpuB4ElL+qry4GTTc2LzfNF8n9tTvCBkEv7FFuOyQkdwMgKG
HUrFN/0AnsxP5JirzK2fTRWTPWRxvgoNMhqiC69uC/bwRKdpqJVOUPwSMlIYnJsY
VYwVEtS1bv2qL8jb06Zelw0F2lVJY6ChdFrFrpmw2bT4n42RLfvuLX+T53yejID2
1sud+Xr/Rv3amRTE/zR+2gNC59XYbTdnEL2i3SOvWqwZN0wRbV20f5hdjsVkR4Ws
dyBRKf6Vxjv4AFBcgW9+pf2cEE6FslDy/UNE0etSHj9KBtJUWTFOmwDSUiPtqcCP
eDOuaWkg46CxB3QXBuyjC4tdEQM7fzaay7NutevjCtydmTyMdqpUXSIe4cVsp8JK
SQ176kiBA1k4UW+wTLOFE/OvvYtEVnYi1F2ojZkR/66GnnW+E6/uMgZzLLvrteDo
lnAtH2NkenfC7cD+KrOjHyPi3plhQMB3CKDDncY9J4QyDFx4mrNGrxC6ae1gOdwt
/aTBA2gTTSRAYqfbvdOMcvKA7YToLQWVcjxdg1KMyD/ucPWTqA0Fq0y81KFnCJ+k
nmv0FWjq07U4YuhHbw0Gasa58/1GAbSEt+/trfBWVXQ6YZobjuz79AflIQip6rSE
hVi+t/aPiW+RDD3TDNats2/csD3a3AqHwjr0lCP0ermQX89HYNuGvuRwq833p8+w
fbPRLbeCcor3eY0dSb0XmdDxoCqzdBuBfG06RAgvSAqUYsC7arBxGRZ4toDeg6LD
Iv8zwc2UyRCn0I/tgYMA2l+I3XvZI3gKXpvxe+d+LdgSh3gnrQ9oYZ4STHKPaOl7
uYpc9sMf8cZ2s0AScskksmAIkfCkBIzkRqTCRYsh1sjzPya75Bhc51TZJ1gly9sv
OI1MwK31Zde1GsQ9Sq1v1ssR19ApAgDdWzqETmt3G5JIfEiP09d6zo3uTtd6aQeP
wYUvwrtZ/WnOZgFQ8MNEUuVmHKL5nwGVPh+dbtDvQPLKO1T/aDs5781aHep4GrQh
3Hg7hnRNbMVO4nMEGvPOYWAIBmO087BbAzWrJzzDJtgp+td9vTE0C/0e66IsRSsA
R9tsyDFxMIFmugG5/MThT1KxAhKIAYEdktNY8gFj1sHik8BE7YvWyJoq250juXZS
lfev1Rz2L+69YB6kVqJfTK9RZsyOcps52mHdik1i+T7ld+Ahqx4t4RyBQH+Bm9t9
Vpc4BaR5IybWRixdsMttgztCsW87rMvHS0LdnSkeNQUelD/wq2d80El/lNHQLJQu
E3o9754r3ju1xg8uVMfg/AaB48L0F7ljvpecQDzyyJDHdvkjcvOevdo4ij/HqDst
pXSDqgUZayVzUrXtnLG6kwdCvGrYspllexCwrzPRMCleS5WrwR7XF6tVPGW4suvl
6TWVBgH5X2Geq2MHbhr9lBxYE4p3yx3VRxA5nHbk8XnatAO8ZUfcM2eE7e4tkeFI
raCV8i/KvDnGDUijU7DkE5pEZKPh5vDWK1ieC89ERHLJSir84olsCj7czlfc/YyX
qATCscDy/KUGJzaGTlGEiFIUSMq11wPMxgHpXoh2rrsEcelK9W0GQBbc1+2cRVyU
tjX9PDXHJD7PO2m4IZBWtE4oi+ixLc+d116aYqEu75nFsLBFVKyYB5o1QAKqgEGa
qpRWCnVxQV/9JPLNGJiGFtHQNvrFT67egPY3/UJW1UHJjJp9rNA8d31vqNFN3x0w
ifW9FsSeX7ounkjMMGttpo20KUSJrPrq61ct6XLLt1EnCI+oGJ47rxmeCwEGygTt
lwjftHH/Yogz3poswE/4h1WhCAUaDFNpbFq6i3W8UixPJtShOZio/pt2KCZY5gR0
HZH85+GJaB9lZYcEuCAVKOcC+YAZ1HiIkFVZmHQUBYQFqMEQDpMUgIjJh0dD/yaT
sF/lTkrxb5O5Mo4lfpbYTGvipPsGyaL5rtwIHg/PdSmlSQd88B5rQfHy/RASWssE
yxtwyQ9uuR4qcnnrv77SExKmaPTlWJNIbLQruI0krRJvVWhO6jq09ooQpzINyXRG
nKdliC/RupbRwhsyOsB72tnucudnAPIwPiSPQIrKLOdwrCcokkGHX5/u47ivym12
046/GzfBJSLRGaAgq+s5SbNP5t+xOqztRLuyzbp0BHoHpboouWo+1kordga/wpQG
9jMn/kN7CKlnnz8CjGaVy5B5zd6qYON0qpZw3fddJyTmzrMi1c8UewKRkBCERDf+
w16xso5udBeFWi8Pg1tP4WwG4L0MpnZEd+XQCb7FfQbOQqc2VREXIha3KCDyQyZN
5lhDtivNlcEaM5bsnGisNoNuHNeq9yDGYAafnbeI4Ux2TokutEjPWx9BM/1bkqFc
cJekSxNgVZZ1d38ML2KEsCaZ9LkSpIE2vTweqvNdW96ydCtRsMatJV6omIHR5Uyq
Ll9QGkom1lP75/aBFYxh7468/gSmFTYbgOWprBosyOvswQGN1DwC00gCVx9ywxyb
+i4N3pKwVFx6oIMp7djHR1tynMXSgMki2Q4MN85PrDEsqYwhP8svNs75DzjEWS/f
UXbhugQCYHnBUFXnCSte9I3zucKQYOECKYWgJJjwGjkUbxghJR5p0DArn0ke0qhf
YqdkwhnkNK7buk9+RDPAVokX7SWK/GEaAfBs4Y9JVa4tNED7iL6EbcRxFL3PDicI
fZnaH9k3T8O2m2k9UghDDc7qCypfzzyPkkFyzz32Ed6ME4e7IMm+qRPWHvAx4wKm
n6IkxtAsuu/Z24Z14IDNHfUIybPecg5fkgIQF+gt5ahEAY9WackSzNhZzFQO6I38
JOmzzJvJSX5lWuLWL5mwcxTPQvtVsqy0vhcbvc+YtpwVScNciLpiqkdO1IhlEhAF
fUEfogrXBX8Y8j2bOc1bGEpOvUaq8QQq3vxxH/N+K7PnF+gLtouWpUuupSpQZv0J
4rPxxEB8nVcNeLq1BzxeSGdSk0Q5YUJadTBmgcxxo8w7RflTHMR3RHYfWwUXI6l4
rFFLPp3/rJhCLecuKu/SvbKnnRp0nJOgYHSj9am5VcyXNzps5RRj3LP98lZ/i5Ka
ukk/QkKm6W9mB6CJ25xqoAwp7jZjttI6ehLVMnCqeEtdEL0qA+krp9tcDn/UrBxm
LUXeHYVh9+WC5l7GufW187tiuJFxRVyZ2SUcuxReM0QZSVtlmtMQdJFekvngnFcQ
ZqbDBdCXge1rhRzFY27nnofyLaWtRboNYbgU1T1sWsbdBCj3O6oLmbByLtXmNXjj
a53g9HmxzhBpcy9KV0G3HM4/T/hj10IAdf1W6zNaw1Go4bJBDQofug221qXUhSfW
8THUWTdvMDPZki+sq6mSy1gr7aHDVBEUzG+vJ7sx3A7l+g8cMZTrBpnnySkDWtHO
Al3D4FYSKa4DYNsdD1oCzvbsQEIX/1J7HbBXBnjxkuJ4hYW2ORxwzDgHGkM6Jk+1
tdDfJeiSZ3xLXgpY9zhHS9P5EkRgWiNCaCNXeRlJs6VOAet9YxcrWnxGxtHTB2U1
lB+VCYsKPC0ZRJUMr35d+70vnkg+2bqUzti8JPFG9TrafYrMcUpyeXXZYJIZjGoP
7eGSKMXN5A/dvIn1ltxCjdW7F+8+Yvof+pNvy7WTpdaaEhzebryc4jzywie/4kgm
qb95HGmF2YiF4SbAkKjkClVkIaJT9+mUnJH6ZLeXY0gV0P8WyFQTmbbSYHDdKwD1
2zorrJEoex8rEg8wBaqZrVwkIuO49zy/4oEalbkK/hWCw75r9ajH1k3NvME+Kl20
uacR+AmusfdXsPsu+nN9WEq5Qfu8OCGNEQacSqSao5HGv5GCt8oZDLjMglJmPk4q
WfQj9/fXKXEzpodhRfIIPVwbIXL9RvDBVFMyOVjkEDo2csNkK6TyMgpvhRx/ZUVq
7/tGQt0GRi7qQDojWRYQuozDRPfL4bTYKa+rJPB9chrjr4l2tjEZf+6TrTayyOn1
Cy9uWnEeRruZP2CV2UYyFbzS9nah4lH4sr40tptHaeOvs+D7wYB418sGL4d2jIBf
XFYH255M7bLK6ibdUKZYiTinBVE1YQCdmz+XJKt/kuFf9xZv6r7e8cqhs0pM3vpP
yqaHyHmVNiIDclTsruZSn3MRp3mhJbe0wSWtjmVr11+E5RDjdkKxSKWoL3uVn3ON
YoTwb66nn3Hn2gw7TLTiniWzWnLf9QYbZT/iJh1w58O1UuPR58YWcUuutJIR3lnu
mj9IM1Ofdiq6Y/Zbw9cIIdJZI5+U3Zxht1uymgmUZlcvn/7wZ5DUIFKVUKNAyt0Z
BMVKvfL1FqaW4pe7uI/ICVaPXoqzr/WbEmz6FrO0DkYm2e68GmHI6QfSfmmnTFvV
gZz+5O0iqMOM7J1Z+CG+So1R5Fjz82r6rbhLs22UxZ3+xWvDKjKeZcq2RvH9TEtZ
qKnYdgdccv6bpR9TVJ08ui8fmc4V0XIk9Sh+UgoEbhGAniIpocw+8yrr2QWe2pmT
C3XdpDzH6jOpkWVqxwCpLYtXTpAN/BQ4Qzp5lrh9FLVmCjPiW1HlJAqKMMfHYA3/
hNe5DMjWQY+kJxSFUuW984vv27bMmbakDbyEwOmRnARbFtyk1UzC0W4r2TsyJaDJ
Eatb4tXFnzGk2BsW+AyQLtLH+ckhMwLyqzgP2J+q8Fs/f2IVK/c0DvrNwxVCMRAw
sS54YhnNuOct0m/Q1CYCTgOpfzP/ti3A85olV/ob8KrNSjoB5DzDLzfZUCRqhxuX
pI0TYdQpiUoyQIyvVaD+UGesm6H5hJZnoJspV/ngfux+/5Z+f4VkQyRa9GbGo/Du
WTVIHIrdAE9DK2ngKa1kkGKPuyz66lwj9X4tQXRXiVsto9kSR+P97cSnPKiiAa2/
PtLHZmcSlAYievoMxswAvXRTxO2YpDQfGojHL4HSmLoQ1IT+nYujJlVKn4zNXR72
ooJz2ec8/MVfHQW7j97JY+I/Ar7EH4G2QBdX0PyqKs0NnZ0v/rnb4O5AnN/u7eM6
KKueQ/nxV3tZbKpLHbXW3jB391i4SI+h0LPUzqh1YvLtPr24Opvda3D4OnAqqLYW
dxy7U5pj8IR1Bc89eIK+5Jmuz2V3jdfXpCXx0WUoXuqlfpWci3Cnn4XLBigXZ9+o
lgxV8g/t0KQ1jpEOXOa0IM/Q8+7w6mHlQ0Og2C6dOFmXBu5KUtiZPJixQUQ/VmPz
swMYSl/t6WvPEJw8iw0ezfy+8W4/r0Ppurqn+WxiEkZFwmoC1ovJd0Ch2KmdrjJw
vP1WFMhkts65xOeqbqZDJdpajvcHuAhHkP96YFCcylATM+A94dM3GLPgbraZm7Xv
D+Ga0iduZbLBqZvnUTNMn/26rAHQbb9y1MEs0lGT2Vcai77Jk1jQRxKhX+JReHwR
uuMxHy+sF3eeF1r5GH5oNxvPE54U9J0h9JjBvebaE9lzjXAn2FD9jxZj5ZfgbmQj
i/8c/ozg7adDrcjV8WkonYJD4+OZ5vUV75PQgTxl1d7eG3upa1nfQ5B/Ihy5t68F
J9CMC43Gq9DNdFRBYRT14PD5lXTuRt6JDoYWuKuYdUlLnzG4uoJOq4k0gpcjIPL4
WUAZLvDSmmbZbuWL4ZMl+zb03B//34NZ8Ih46nJGMqdPGeckGdtRiI9qkk9S0QaQ
yaM8h9Hzb0J9h8xllbNram3B17lnljRwPa0IUJn1QfbwoAxwL2ufI9e0zcCAHhY3
f3YQyhmfTnvVU0lIBUvZR+hqifpC11EjgwBKVCyziQve+uODt7vbY6XKLC/GfCxE
+YQWZj+Rqs5KL3TGLcaLIWffdqy3D1QeEGu71NN6HAXHdje2u3NAMWJYjkFNfEuv
ZTEzDunAlsNZIUIBwzw5kjugQsiPMUB27402T7LmP5ZOgw4807DWzd9i5q9Kv4m/
R6Iz4Q2qfVOEnW1w9j5+j1rppGfg0OqeIAqkap5QUfg5sIhcczg7TdTbhJ04RMO2
Dt/x7b3hTiOmxnndBnlcl21yFVtoKiMXeRSsQDVYLs7bUUtbFM01JuAcKc3r1Osx
SQK+POyArUwDYZBJlkRDQZbl8X4+7Ar0sUsw5tnK7GQGmrhpQpVCtBlh218xL2mB
VCYS6XwDJFWmoMSq5lrSo2TamamxVLA8J9YnbleE5qRtDiDZywSHkb3x7DgoPdTR
16ZtnkNk+AzjF0DbNAuUCLw0k6a6/vJ2HMJDs2AVvuwi0NiTrKJ/PcnDUBvbZlUB
B3PYzERrE5qUoa5A+jeyGu8T773+ZRr1/svNsUOiePj3lY4tOf44Ewyqh4XYLq4T
MWxge0eXaaA96S87P06xkmVjweAODOqS4sIg03S95whgDTAafEeMT1R5uA7LflG3
C0+2h2ZLcmkVuVIxpinP8Z4Fel1LDAmZIEHWJqBpjug0k+u4BEB6zBEAIh9UyCgv
ARAMhk4RsTrg1zaD3KRAfvYy0dy4kfkkoQY0VV92OzP4ulmA4nr3XomoL8u3zPB6
MGht75gv8h3TvDVR6+LjNCXD83qBA6ySTTKd4CUJ3MPHHbCugHj7ggf66alrXWjf
EgdLEdI+vNsJpEVSBF/9yBvkR8mKZyyMirnJswSfnZmsh7ZhvqbAWuXQ1Q/6XhGd
eGotES2tFHzNYImEKNVmHNDorjLmZ4ThDwzW+qS0LxwFN1JjQMTu2CDSeZlxLuQj
Dam49HEUImu4MfYVgL2fma5OKRnOkNSsiFjINFz4cZ6MyArnIBc1usnLsw+lFcpt
/Umw3XwKwYkrfTCFYCgp2UW3Tw4SkyD3DaImGcFO4pH+5tgcCrWnyh7plJwOQAhQ
s+YGpygMJxqT4BNz7YciLQOtQcrvVRAA4uj7c7p3zcwp6zjnLCddDppFk77JLSwO
E33Dg1wkpsYYJQMX+FBKrXqt82wwrzBLOtKUgdr1NZDYFnN1uHPff8ar1Zd22XjF
hwgjkNtkniSb1Nb5K8j8WsEcPQMJ346AuCgmUM0++op1tWzC9gR/TaYDPJ1cyaVJ
D774uLJflBWKGGvOzMGOmXRvIq2zJ2s8gqla46mSxDJC7NLc3VgkO681M7HaKrFD
QVGXhiuMxMnGg8H4rGAa6wJCfEayigDlyOAAt5P1HUMlwSYFMQCWo/wLKA769OXR
DeSPnJkeTLkqV43BjBLUOfDKsbmileDIN7MxnnIeaLFWmMI/T8OTccBJvWy/TiMa
YY596SAvKLO8X2wIGSjAyXPbS+dF/3Rrg7DNlHDWsGRXJziDazTrdzc4FX8cZZLV
p/GthuVMc0F+W/x6ZW6GnD9dPRxuHHaynSaIUgch3Mc1kpn5PvtlBaYrZxHD33zo
LGzrt8arFa2GhGPU1uiqHUfxDhXE7Sbw23bohhJcaGtAXf36LyNjyDKrG6ms6Kyp
hEWM/mS9x/3pm2NQ6tY5B10XJtvinJwpeyPr2xzBNnA4Koh9Uv+u/dWp4TN41y8C
x6icfvYulsDsN7/8j8lcCduVZRRTFk7X5Kj12CtGxXzTxvHWjW3pf6Fnr+wicjVl
FhMgDY69syzOdZJmiCar+/jTMM23jT0Ia6cMW5IPuLuqNK3oDLXfTjBznvRbTy4+
sLrFblhxRtNWs9L4TvEcmSwdYjB+L6bGff9QT7xf6Y4v4gC7yWhKFUcGY4/ySbby
1hB1OkVOtkiUFK0uETcgbVEBhxEBQ8vKanly5iydS46SuXpt9cZsRX1FQhc3T2Yz
/AHLwX7UfN2NzO8sDnqMODgqXw48WGFSxbDlqRdx6DZ0gMveVlod1/tjG9Mw3bcE
bJqhF3cQGONfSAjvYrSRvoZPcoEzV1Yc3xynjaxapEZk3IYj5cod3Dfx6lGsGtaP
ychW9JbK88m4aID1+mVBHACX9TvGa2C4sTcQefCgCDXgX/9JJ/6QQ6HcumKra4f/
GLxhaFpW166IdogD0qAdsdjt68VNOcug+bFAxclEqsarMcZnSLY9iUhJfmUzAJ8q
4TutP1cJ82ha9czzjd2CGk/JdzSpi970Q2Ztstym94BZn2vRgXE2uYbjpkf9RnBn
lNxOgyavhN1IyHzDi4O5y+3hCCCr8tO5SRxreEgNC5N2K0ynxaVfW3VS3EgGTx6M
PlgfAD2MXiC5Itvs3nTh0t5NDEQ2eiB+RO42XAV7Po9x3RhuDfDwJGX+Ok91nGzk
L4bNP6pjABdW0PbNLvF5I3+PB9nst5K8xfzk2LigllttA5XBFNrg7sAYEuzWOZiQ
B6Nn2ySJ8dcvk+ZVIVXziuIZmpU1+PuqDMdSRfSeEBw30u/IUoUtctUumXczMstR
XnIk/+U0EgsugSCFfysz50xJZdF5x4CF3sj1kBeyIqIEwB2Zw6MZSyoGVZgJSeTz
wXPHt49IR4p6YVMYJCm/haEyrn6S5KCYhYfSQ2xarHGHBL2F+XgECw6p8v1hvxte
m6Yd81hMgYkM8cdKdixnq58EQHp0/hkVEtHkfXupFvtvM03KNEHPSrD2WmePJbQn
WXftLD5xrgeJcPxi9S3u1HlK658QF/dABJZvfr2ZJD0oSyifCc4p7AFz7TItPRis
/dZ1b4A6Nf+lVceu77rXMcsxhjSh88J/FeQ2VXd5t+GF9txuR4IqsEUD4h5KFIDw
Xht2axij5ja2NSyPy1iXQ1uQ46rrz1FzyhhXcoBELksqH1dno1K1AYNxAgAyPWkD
JiSeVnvdcN1AL/94EYUL6H0kLlM+Gz4i8bEo6XoI0ARMs6aBQn5+tZxKVT22hWRe
PgxTlVNp82mzih/UvoavnYNXs/ImaGBz+4yd/1VAGbiwLA3SlrbWPB6NsD6f+ciz
j2Fe+kAr/P9bB1Je6t5X3JRQ/kj6QLjNPnJrrxi/tSdCkQlV9WUXjToZcbkrIezq
vyT9rVGgReRCV8n7EWV5cl7zHiXdpWO24ZgslgVgVe+651GLcsxUWO9H+NH8cXFS
Vy3ogHVU60J8TzXwrRnGFM1FnQf0mpyYFwCOKbb4t4h21C01o5A7wTejxBvD6V3k
68nzM81UUkqV62h4YChHvhx3JParB3mctEf2/T7AeLGxbCB5PzCZp/jw8tbSnAhE
2F/VizsYEd7VS+7Q4NO8xfNLt1ACdK8lhKZlZagwrJ1+vT24V+Vf4IGFrcKHliG9
7UOYLD4n8jgQCR4RJmUr816gGdk4Cceqf8tR9VqBusS4VqDoYwnTPNJS+oxK5wwN
hBILkWetYUDNvZa8pWUtwEETY3n2L663pvrjOOD88DWWi19YJHRhEqR2/mAdnELU
UTcwbzB+xiM1WlwTePVTh8G4wjYkGSauYiaToTuJpmLt9qb23tYN6RhkociqueCf
i+CJL+S7KKkmed8p+eS6cxlrfPFIDmFOQOCNcX5UJGQm9cuGhhX6cCicOzN7a0zA
xvrkZlpZZ1gnGf4XOTX21QH+wvt9+1n/sWBNdftK7RoKePQ4M0SBZAOAllzc4Gfd
R+cf+YJ6pMjO061WT6vbiC3Zb6sqQRLRx80W4Ol98e71AJZTz+3IK/6S9Iry9jmx
bdfH5wZMKgjeBCIimsP1qS60OsJvmZRI96w4Jm4X0eNyLQwR8SgKjjKaYJyCxuUT
c8sijEYVbU0UcdLdRT740f1YOSe4J7mqxKO6TB35Ch2O4hwGY6+aODlztcQaFl/X
d25rTX4VBY1P6b6OPIWNJ0bWiv/lSkNDWJvqOLCOVkCmqROC0uuzXVCmxtncCHhY
emViT3jOxa7PL1UujGIemjmsbFyBrB1Hs66bszhKA+mN3f6ZHaM0jfL6wwqHM1TO
SpD5Yj0gx619IB+C6x/2qZZ2i74K2ciHwsuNpwP8ITctXS/MgkxUj89AbT6xBN46
GNOeLt0wdSwzv8ivhmVhs5g0bS3rfAQFuVlhp8ZbPEFqvYfRxCNj1ifDw+FbwtnW
JzvWH9ddcvYcc2xOgB93tI65EQO9Gnc1E2wXgaYG/QGthweqAx7Z4RfeVtHoi4gg
caAn+GHgn89FRPe+AaHCalCw7ysY0CBUFIjun9hKWG4kd+ZMh7wOJBH9aeHDEE7v
MCMNN6Ne7v4P0TEkJI18ugqHVm3uVDORGWPMJUUs3npE392Dvk4zIiP5yBfxUlk6
TW3mYPozeGF4fqWdjJdSHZaDOGDy0JH8KC/8q50l52zCxB7JKJkJN0/VL6kHmRZo
KCFQshQDRHoycudaHbhD3LUBOcBFReZ0nES/LQxOtC36RNLtPruYe0zfjLAmvrDX
zerwmVysmbYuCj2FkRd9GY6hOxQVk7xDuv41yfSJA1f2zRAfc0WYOE0W4Z2MpBeM
ruwFKqPTmNSAoflQDSbKA+460x31nNddFNhAOq2t31uzreP4c3wcGSsL9EXhVRoD
+Kn50FIlVKcdlbofdOXPE2E/fxbuGGaOPOCbz/3hRPfh966V8kRh5Ldt866ZnPzT
i/iV+5g7HiwnY4J/1cEGxEQN8C1CC2rUePf6sz2Y4xyBt5AHjECleukmKIkxL+ew
CfJsFPkNx7xKgDC7FTm7oPeQqKd+B0Ypsb/WW7ebxtYZfkL45Qwfb/Md6yWl6Gyj
4B2/MUgJK7BJOOfhEFKgHyJfXMZTaG/jWm16SQ8I8swtgO9suYQnk1m51qKKkJ1k
nvxk6CcTKaoAkPBh+Qm7C1vAts+i4IV+Z/iTaC3IoEN+GZp5ZfDFbYL0uOmn+WgJ
CJXdAFbh9eSPlV1E20DR+itNvIyQN167dR/cF256AY3eTd2juG8fUBFuJPodh5BM
GRQt/cEgYqB17I4le8ZqUyBnQX1GJc96xyaGjKwTdZrFgpQamhTLUt96diIa3zmy
myb7vbBybWiASSAXd+p4NpYIPrT5NEnIYc2IWwBanWBMIRfXJ9nDsVs6qD5B8yOA
xqkF037wfiloYXy5D0bolTz81KewzQOiu47Bm549REfQ8bn1qa9Ie/Hbr+wpE6tX
YPHOhSpOxf1rzKmok0YG0/4Kp5VbkQzEE+kc8rjSA2PDNqX0Ubv6/BehY+0Y62kY
JYIj5LG1r6SuyjHCJih90keVuj2R5J5o3MoAcFIlJxZU351rzQAZXoCRfX2NghZZ
QZTmx3zStbkfKHHI5p4B8w+GvkzaqlS+HX5MTWodIB5jDUVgatWW0xDUytB3Of7U
UhnG7I10E17yWMYOMENvLt7/8LM2XXoy1HAwOidQ55ePPUqv32qivFI26171kdK3
QDObvvLY3QeoXxW28UwcUQK2j3l3JY1LDorGG0ZIIHJ0wmuS8Qm0qZw+Ei5fC5uC
5JkjJfF9jc7dvUweM0xDBhcAPquGgxqmpipozxCzhpr4lQ+L53kJUyXCUY+UJYk6
LnO0OdLCt+yM4XaiTH6+PD/I7TGXMg4ifXM/154V+trAYxd6kLbzHBx/igkuxR/R
BgHqjJoNq/yB1BCNp4w9M+O9xqa/FWxuQ5GL9mQUroB3mcb0n19yntME3mWH4OkR
Axk2L8qoDdeCj6p8SXq943wO/tK4CrOZCBA3j8wun9vADRhl0nFVGRl5ARRusXxl
lRGSCXWzzxRsxdIQYDHgJBz+hZ9/Kl9dvcGdXSbS0138uAHzbfzusQgfjNmp8RJh
/YidYIeCVVmwHelfQk6bTzEqTOtMebVEW5wDKbJeULNzHdUPRFP5LLmrcxH/e4Sf
oTDX5DKuNFXaVSXl4Enxjep9DBB1s7l11qYOv+ARayCl/7Ew0Wnp7z6eresTJ3Mf
GB9Dz80BoveeO/abjOC1lkLBNSwlnGhpErs8CLsBCFwdUBzzlLcWQBa/fjwk2QQv
nD4jvtinLNSI8Xspn05ck4KsQNoCz9LoY/uI2qY4hA81ELYk3yFpkULAT+mOL88H
EKyDDJN+f5gLL7186AbbzGHR37Ef/WeeOzPT+QhFGu7e8SpBAPVilhlY1bHPal2n
Y9w/WJPl3wuRlYiHAv4E7LO9Ju0FDsL9i5wz8h5EkiiYxEDqAvoGuUE6Aj1DJZ5a
RKUz9lK6qbVLc/ZSYyQYGa9rp0kjPB7sPpdkWHgVQYYdUTC2LM5dv0YLl2jhPpRF
7QVgDsTs0fM6nTyM7NRmEHgATQ+SU3+0zgX4URyWVf9UftduS9lnplBbmLNlhPbs
`pragma protect end_protected
