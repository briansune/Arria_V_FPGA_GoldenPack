��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t�ꎜD7���(6)oܹ�hQ���@d�79�T�8HntUt��ٛ-��@\Q����9��]Rn�����ä�:�"O�l�=�)��]�)�����;�cV9��]-�&R�4Yl⸩;p������1;�-3(�O�u�eg�i�~]9WiA�	�{��������Y�_uW]�*&�V��6R� �e��ٓ�f\�-�VS�[�=��|�U���ך�Y��;עȖhh]�����R�g϶��y)k�/{Ak�ba.q1����6�4�:�5��;O�Q�nӂp��L䣅�$ݗFC�G��S!�)<��v��rj�n�v��&,[Uj?�����[����Lq�}�Ϧ%q��л���I�gr���5#�<�iw�A��De�|��_r��7��G�T#���e�Y��OX�?��&�n�N<>q�a��V)��x�r0��΀A�핢���W�n�a��XX4�Sq��nB}�ߑѾǴW�� �����=ח��[�':��5���f;��n���ofd�J��D��r�^�h��Gs��&�/v1K����:6c�������� V�#n�<cHLQ��͏���q}�4�"y�O)�'�� ��{�x��l�Ev��H�'8���нp��r^�&�w�چ/G��y*ʻx�S�7<N������C�E�����oAM�뙼���ąp	(:�>��2�glo�`?-�)B�D�YV��|��ז��)bv����oS�u���ܐ!MJ���ϡw������&@6�F���`�E��K������,�Z�/ ��A\�q����k�1�nz�2d��]����E"�������"_3eܲ�\ET{��hׯ[����׽9K�����Ѳ��)n�O���%���FŖ�\ 7��N�Ǽ��C�)xn��|��2$�k{ɋ���෪��_��c���IY���x��$�$�E��˥7����=Z�k{�S�\��6�^�(�b�e�OVۦs��}){e&����SBKL��y��!�9�X�����k�[~}����\��}55t~�Q�G|����2}�(�q�hC��Fb����[�Z#[f3�d�V�zn񞙼h�/b���%�I��ya���D&�,&��z�C��|c�lP���o�{���U��+'�L�����ug��jh<�E���穩�N�.jm�ܳ��ʧ~��/]j�����R����B���������;7�z�YZ3Vg��4�����V&��I�pT]�h�|�k�p�������k�4��v��) Ya�9r
^�wt'��yٕ.��~ �:=���ʚ�x���/z��ˬ�E�x ;ˬd���jm#U-@��67�0!B��~@���s��9J�R`Oޔ&�P�,3I#�e���k2RP�|�A��Ie����I���������2Z��la��4<���S���Au�I�t�Q���8�jO��fyk�.~���C��Up�͎�R4HJ�7@�/��w�@�A}x,�RG@�3�ݬ?QfA;��D5�kz��,ᱳn�vtϔ�:�~�N^9Z �z�-�ׯ��f�#��������(z����$q�$��:Bq�VN�����Y�v85�F6��X��T���D�GU߽�v
��0��9�$W��[1$?��+��T3j�eO7���EѮ�������2J�;d�|h�Z�"�r3 �a%��ڠ^&�2W�:�g�߷߾�P5��P}�q3��¨��}\�a���(\�̬g�Y����d��
ʿW��ը�u��:�=~�<�J�'rd3�/�BbH����@1K�<!]��hqG�L2��ڹ8xX�Ф��&���� i��I�M5*O�9;v�����7{z�5�X�F�#��P�P@��#÷2��Ɣ� �l{u���n���K���6>��aM���FU�P�M_���!2r�k���,�S)t�iY�╫O�d�8/0}�0�'rX'o"�%2�^ ��O�����L.�VK]���:�B��Ԇt���͕�5v��Ɵ�r���G��?y\7@J�-t��k6�q��մ�7=[ҺAٍ�@�� �:���K�c�?p�ѤH��@��|CLxԋ?���~%�c�O)��5���^�$5���	s�{��m��M6E�,Y9v����wI�1Xu,��0�s��j�_��+�p��f�����"#q�)*=OtO	�s�P��-����6;f�'��~��龂HF��+ۍ��VX׿U(��x�o2�������`[V|�l�u������ڬA'�)��ٻA��mf$�Q��!��lk�`�4�&���S?C�6�}�N�OH~)�����D���_I~�+EW/�W�sf��Pog֯Tw��Yh��|7.D��뻑U4{�F)�p���qv"i�a�'Ը�[�v.ϴ�	��}M	͖�v�*����%�Cf�5��Z<W�ڥb�['�J��T�/�p�c��"�
�.@�[��C��-�42A��(F�����,~ݮ{[\�e,H���DM��a�$	��0�����c��I\#����+L�$�j����S�եZ]��#���e6%�o�5�P�*6�D�0��!�eM|������<6:�$J�ӕ�&΍��#���%�4���ʱ�6���ʹ��U�?֎��#*�ZM�IO�vu\X&�{m�KS���OW[ĵ+�^9��R&��N�T�tie�<)]�����c�_�/�D�յƲr�
	"���C�s�A9���T�1�h�C6�t���^~�����t���M��I^0�Di`��\\3���0��R�&�,��t��%\W�=� �-�r�a�jȸJ�
�L
����$��h*���fO�������`��4��]A��r��ap��e��qàR!�'�����|��w[1~�-6��]�(��Ii&�X=36��DU�&ILv:ו�0��4����!>�1Z6n@4�h�|�͇(V�.Lha�B�V��#�{�y
�Ȏ�;&�E���q\?�Q�������)�au�!*���kA�=Z?���_��x�wĢ���7����0�;���;]�l�����w����1����ű�H�����
����������*��y�9ԏ >���[�w�OEn>��ޑ�[!�9�cz�T_�Cϼ��;��)�C�̩패�OBFA��c��w��$���nL �6��B�dh�.��醮�~w߉�*q"��CsԄ�5  |��U�F=����1V�<��uI5"�i���<�Hf���i��̓ϔJ�e�`��ʏ���̽��MS3��/n�.́UjK���]���p$���� �PG�#b�݋��3�X����(�9���Y�{�>z��_�v֠�=0�;���i�K*_�F�l���Sk#���w�#n+hi�:ɪI�~���ڱ�)]v�1��~�_�]�%sUAxP��)]����*��}����*�%��3M ܃J�IֲL��-�}(ci�����l$AE,�sۆ���:�+��MEeL
s!�jo:�|ޢ���-��:8�x�x��P�,Q4_D�!��Q�����rv%[� �u3J4��a���(���#y�0� �}�.J��v��΀��H�m%7���zo�[�0�vW�7�n:���eն}�x�I����ۻxV=����GDu: �T 2j1͚~qQ����yr�%zB��|�"�w׉�^a��Џ