��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)���vG4��NB*v�^%��_�rG�v�2�H!�W��m�e��
H#�w�e|s�>?Џ���w@!��1�?��"Yʖj��ug�je!8z7�/��r̚��0{�4�%�C@�"2_��`�AL"�հ�fY;�R����ɏ~q�Ї�i���tqs`Z�abB�v�*�Il��a�A-�K�.�����Yި�[��q�֨W�a����1f^��$z�ٳ��@($
�^� �i���2�͚󘪷U��y=C;�	ZQ�{�_���S�6��L��aPW�a�����u�iG��g�.����>�C+q��KX���"q��;������;Uj�+D��L�'F��
��i�8\�b�L��[s�KN��T��<�(�+9�8>5�����>�I�8m�|�	���TSe$�=����r|���ֹL��y�e����� c��a��ve��`���$�;9��V��j}v���P�M��Kz��h��4dK�s6b�>�����Pt�Z��Z���7l0L�/F�?��a������x'��v@.-gx��d��{�t�~�M�3�%w��Qr+N�X�d@�hZ��<�$c��ڇ�5����䖢��C��)��d�zkmp8{^�D�cR/���Ƹ����4��E��梯p���m��( �r���2�J��i�tjfn�?��ih*%�� �,�����y��c|����d�r	�Xv4��})<�Nz����&���my��J��?4A���G� q�*���&��G�<ӣ!r���ڛ$��8�Ű8ї���1�e�V�Y��Wɀ
��X��*�х��Pӑ�Z��hW����|��"�%՛`�8֭��ZYo4���&�%B�X�EUOt��LB�Nﱒ|����	��ѝ�y�׳�t��h1أ=��qP�������7��6�xKo?ޭw�Fh#�\�]"�i5/�k�j�ћ{5�� �bHD�N���c�v��P1��Y)���\�8�	��!��IcmPf�8��� {՛�k�e/ӟ�ƛ�Ьs+S�X.�$�/3�7WWDӨ�1+��B�F1y��&�kPy���c���"��	c���J����H���8<�6��������Y�4ФMvk�j)�F�x�;o�]��� p�A��:�<����1�5Y7no���:���Qp�Yd�P�
ڌD0�DV/�Ͻ��y��=\�qw��7�x��T�(�QCM7IV1�d�{��6�cRˮ���ߨ�|��HjN���e%�5�����JWRR��K��q-1�>w5)g����pw;��ݹ*�uD������l�>��x*��Ff���&P�E� b�:;�c�m�}\|H�>hؾ$q{�[�id�g�D�) �'��l�,!�=��Xs�|�e)>�p�6��0��~i��hW�1���2�+w1�3�:��& ����8�P�;$�~������5�#�o0�$��1V���x��7A���W~%{��[C;f5b\��b������	1c,��[O4�'T�;�Z�5��H"��6}�Ȥ�2�������zn+�J�M�����zp���G vsQ�o?-0:�|�xP	2r�L����={O�6�W�6���Ռ"i0z��*J��nbG6(��˖��ߴ���D����2<<��|Tu�����g�a��Č?�_��pp�z`�eH��Jy����C̵X&�ԍ�j��a_��$��.��}%X�J�>D 6Gͬj���ی�Y�,7�-E�9���?�#�"����=� $���*�5��w��J��l��L����iX]IK�߃��]�n���*ݻ���%��Z���r�pN�		��Fg_u��H|De`�>I{�{	��y,�3�ы�p?���I��4sU�^��ܠ�x�;��v p6�����j��� u�A+����[�;��K8�r�m}7���ly���+&P>L�6��t��!�PCK��m�ŨD��P<�+0u�B�֛���,�C\���ΥA`i��_�Qؘ�O�������n2�,� �W�C)��\y �N��
�d���t��P�&�fz�Dk���4�����'�|�	���������R�����;)��ɯS��Z1�H ��c���،��:&��R�����3/��ϒ�:F�{��x�`�����XP��d���M�!r8G@ঙؼ,��8C����FO��3�q��5�MƿY���α��dEz���Y��>�Iy1��m*mw��iE�z����v��*F��i)�����>KЌ�*���dyy� Jjh#�23�Q�#��W�����b���e���τS���@�XG���YL3i�2T��}ﺌ:�ER�%Ud���*U`��Ѽ��(��<�:	C.�~E����ۮ�R6�׿m�ch+��(�� :��v��7_���Cx�h�9���m�4��*�Q�z,�[y�\�Ss�۽B��j��D��A�����Ơp|3&7��"#�q��)^�N�"��]-aːUa5��R}�NDF��_��3�����=�ťv�V-�$�q)&??A�����ܔ�)��\m��R�A��n�r�)+e�M���@b���ߑ��|��S��e0A�ɐ��_��fld96P��w�ʏ˂�ʴYШP�h.�)��O�w��!k�vYe�r�'M *5�A>�S;��6a����Q�»����î�t#Z��AAO �VP/W����4l�����Nų��>�N�����x&�#�;&RV��N �0ۓ���FP��A�@�8HG�����/y�,�q �ו�@���D�U�CN����8�"�`�����\?�h1�#9�!�;;�56��;O�a4�%s�w�
_�S7i"���,%}�6w�QG\��M�Y�`�)P �k�?��BoO��R�y�w7>}|w�Q�R3GE��$�e�H�L���AK���!����~̠�`��g���%gs���#�Zj����`?�瑟��g4NPH��Tz�@�ㄕ{[Y��OQ=ɉ�q�H�Sp|f��S��h�*R)��W�1�a.<_�6�B�^m"h�&t�=�����G����
r~D��>���t� "2���MO��o�n$���mn���)�~�Z�;m/���6�9��c��TbH�:�I�:�����R���0��W�:>��}mŴ�����ӕ��Ȍ���_	��n.t�H���N�{!c>n#�"'.eϏ�=�[�by� b1S��,w��}�?�9��r�%R��� ��ӿ�"�qHf�ˣ�xOA���^��"���/�Jt3���X��T�_[c3+�H�����
���w��	���J7�Ҧ�}��G�u1q��?4n�hy�g~��nuİK�?$�	s�=��q\�n��1�ЁȌ�L='!���D���q���m�(~ ���U����Tr		�����Fw1U�ǰ�~߼x09�}`4�W\.�y����j�4�߿�N.O-#���A*)xڋ8��F���ӄ���Nu�%:�n-N�9���tr*?�����pWJS�T�`�J>�nX�<̡n9f�%��:p���T� ��o�D�p(���c���!��2J�ȋ��dV�$���[|�I ������	� a�
K���TO&�"�	X�����`"]s�4�p�U�y"�Q�{JV>���}��Iv:�f��i�0�Zt��#l~�F;o�a�x�%��� �+�&�'!A�I�Z���g�$�'�[�kW%�i�!�)�dr�����=�of�3�S�[{�Q��Ur����Z�n+��4���T�`�Z��yդ�{/��n�k�U�}���C���b�?/"c^��=������إ��:��Z��JLmӑO}���_���lt@-���QdaA�B,B��K\�|��DB(N =Og�ߦle�ɺ�\f`2�b�OU�I]2Wbn��|z����R�T>��Jp�V����L��鈨r�k��V�PTv�f���¤^C�GE{�����C��Y���?�u���m�M�|�$<��.^q�r1~��1-x9���׿Jv��(�I�7��`V�eqSYo}��������lP�t��m��[�ƍ��'��kq�j�Ox���h���������5�<f2��5��h|���+�D�mbxZ6)VB@[�Y���������6fWM�Xd��a���rl����-�?Ե�TO5���|o�XA�����=z�4a6�K�W��AIK�}RgL��d�o��ݲR�`��z�x�w�Jm�S�棸~e�Հv%w��*ࣕ��d>�m,�$���%��1J1�W��<L�;.g1��x��\��í!���I^_�ؕ^��j�n��_n��jX��:�ߑ��E�/8�:L�Bc\�Qň���M��̦�Xdw:<���	h{y�T��� w��ծ+
�(�&��vU�Ԉ6�DW�)8*q�6=b;_�]M��a���w�x�4�Z[`-�x�G����3\���oƦ�p��Xf����m��,�U{�G�揤:T�T)! ��"=1�K]Џ�H�LCډ�##����L޹��]��֚GYA��6��+���5ڢgҒ�Q֖�ֶ�M��chE�Dn��x�@?ƣ�S[B��iL�^̬����3�E	g����JHi��Őd�:�:n˿Jǟ���'2�sh���4�NV]�D�ˎ� 3���Ќ���ܳF��I�N���m(���h1�^�)�5&p�O2b��z���[T��7�r?屩u����"��/��"HԦxX�_��6� �Q0s����G�ۀ�Q�ag��]�0��v��1sjQ0�d����M$�;n��RFQ{�P}�"��)ĳ���<L]+�0�o�R�~��TdΖz�-l9=��0Kw�w�[	IM�;#��KG�nr��nRf�.�%\�����L���Y�{
�'���f��o����Y->rD�z�I@l3pD�J���Th{(A�cc�
BlWS�:�� ַoB ��<�_�I���/Ʃ�h@��c[T{��m�RV\ħ�H�����u9+�^`b*ἒer��?���39C���e|�k� ���3��P��||#������i��"�}�0=)Ѽ���(��;ҿ�pX�~K:�aDǴ�v�d#Ӆa}$4�
�M(�X�$��)��fu�����p5�������֟���(��f�U l8&�}h���S{�9����vE�3Z2x�ﾈA���+V���O>zxr��� ;_��@I�:á�d�����_��Y����w�3��%����t�!��ך�+�ʙ*��BS��
��IE�J�vIg̽$����-_M7�Dț�{K[�'5���q��s�S�hN��,�Ï��3B�{���,܉�(g���rГ�j̑��p�0|B�T~�w���˥<{X{�)~y�9��"����j5�c%l���)��/�q���vji3@h��meH�&�
~��0yW��گ�҉b���C`���9A��Y�ru ��}�m�M��;=�����oAIk�P�JW���N��?�lc����u�Ӌ��Alx�Mj�)#F�n @H�����ސPC�	S\��G��"����n�V�$2�WD����>(���Ԕ�L��X���b�'g�+�Er�ʷt��%�Y��*i��
�"u,������#�/[#N���C�U����b���ȡ�3�q�U"�h�y:����`�V�ȝZ���.���I2�``�a[*W���|��R��m���^k+�?���Bِ�����UVA��fz�'~;�.�K��p!�V 5喎�f�ڀ�ěq�����⃻0���1>��EqE�4�Y�x��/��e��^�jK*3<;W�
���2
����⻪���k�P�)%h�X����BH3�T0ڮ�<J䱖��b�60^K���,�
qrS.��oLTg�o�</��8�h�^��5��V��p�PS^��#��u_�@�!��e�����������%���������q���r�\��O8(Qm,���o�Oe�0mт/�@�uY��C�o.��E?���:U/_3�_w����>f�$�7fJ�g�@qv�i&�{��>	���)�l��_�%��p�[2�C'�%�h:����A���B*@�C��p3x;tj|�5N&g��$��By��}k�Exȍ�q�U�\dl�_���\C�
J�*��
b��j�S�PCS�EXmS�c7��R�l���0X�MZM�T29�#�C��2��{3�X��^�(F��6+ٮ����uE�n�c�ǃ�@�,צ6 "�n�DmY�$��C=Ȧ �UB��Њ��h$&��k��#~�Ƭ�K���4��{�����/
�;��F�j�x�o*��0�,�>p
N���I0��<H�i|��9��f��M	�3Ȧq��� Ka��^h?�w��e'���t�cc۵T_�j��6 �h�mV���GHP�hy��m}f ���&�^�Z���S�
�Y�N�&,���������R�O]уJ/𵰛�ʽ�k"�浀D�������.�{��9�������~��Q����j��d~�-���qJ�G���n�����5'�f�[,<�ݑ%������"�\���7�����6��#��p�WJ�a�.}l���w���%�����#����17>�B�Ӑ��P� +�"��_9�����cܙP	+��T�>)��h����5ͯAb2eߍ���m�_�_�"P�z���
�^�n2~�f�݇O��+��<j+IU8�d��"�$r���l|+��u�|�o�⒟Y=۽��w~r.���� ���߂�&��!�d?RiyWs�x�kbKs�&��]����E;���D�o� ����H����^�4p�$(tlS�3�!���W�Y����)��&Q��+Tx!��)v|��k0h���S�.x�<�dU���,��v�[D3�l��?~"��є��P G	f�7�L�cn$��ؐ�Ϯ���fﴧ�#������m�L�{�e��zو_���S���N�v� ��ZR����g02'ʩ;`u�P�vϩI�{�YN���Y�8Ϣ��J�(^X��*)#�":� � �S�O}���S�AF�sݎ5@�h��&ސU���\�8�tЏ�����{�c%͂]��_��p?�7�ǳ�1��T"����NI�&��3��m>�
y4������p�[��ښ[��;�@�DÓ:��e�眗󔞐��aAl���%�Ы�N�eOO/w4�"���2A#���@s�������dj�i���z�<�G�T�@��wC���!�U������@��Z�L�U��?���n:;��w�S�c��ɜ���~�M�9�`L}-��g~�����G`���9L\�����*i��ϥ_}#'DG�^Y�l�y�p@x=dN5Y�4�/���,����:̐���xk{W��u��^���@��X.��Si�O�R?E�aȤx�d~���j_^?$:8C�p�eا1a��u/;�/���Ԥ���r7"�)ZҨ+�ȿ����#]�  0�(kۡ4M)j���oXU