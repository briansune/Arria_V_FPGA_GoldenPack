// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cgPXIQS+eaFQ1xhhhU4Niu/PfUbpSwz7l8H/LLuF/xPCioirOxHH9uS00nd0XIWKLnSjBGaza/Zd
4M6l4zvTS6LpvLE6tS6xObc34OeyMn1j3NFXug/pS9GhviyQxsSYELmWKYPs9O5+dpbQ54EnMSko
v4Pl9Wh+E21tQ+s5bp0FqWd6Og0rg7EiKdNa7CQIIpCMrYue64X0LRGRBMhG9GSfIpiIiuI7rrAn
scfGM1l5yAp45yRq3pTs8lv6lhJeB3NzWuGo00WJs0I0RB0Rjp4l9lhT/QUPguM/NL6LKSc++qjb
E9yQgZJFCARRKFZeyE90AWnXdBbGGhv4pRqegg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9584)
7H/QxC7E6BNIv55YDHW8ifvUG05UE/QHX3v3+GHOfiqhDGDt7h/xsIOTro7zhjc0vGXD5+z+o3Vr
cWROjbJChRICyjZMhUP+A7UitJ7ZvJKKGed0M4Ejn2aOYooTI6zOBvXF5hbxP7fgGjEIa5cP5I0u
t3za3DNr54eQGGKtFKFerFh0P/NchafA/pXQEwZXAMh32kFqjnJVrQlJWdyQxp7AGFDxrEExFjMS
f6O7v6kj1aiySoeHdLCGh9MiL9k/D1iXNVNisOlmE5SZ8GcnnpaZqbaHXgQz1Q9LgNO7Vxvz7KLq
DeI9V5nF7Y/ReGrSC6MmqcIVLIVnLQkR7baE4wplloGBnbUOiIBrN7oGu6T12MCRgplYXW/ME8xN
wOk4WPlD9sKrGhNvpVDRyvpKqN/pE5KxkRSTaW1EdIDHUaTityQGbdKg9R7mu1zRiAtYgGd/qkOG
wsSvnvHDYVSO+JzhT0S7gRQzn+gQfSKxMdjBsI/cH76QUrtKVhvfJwHY05oJ60gswu/HTI4YhaZM
Dx2PZtg5VEMmdeyqkDO05zUbO5VmO/kIeWM9/yZvN7I8nNMPJNFW5x2xKGKSQKKOxRX07x1M2cy2
Y+H+iQpi1Mq9yxskGXpNUGdw09LRMUmiZKzotWYn3IIwz8qT45JnE8wSvzm85bw3d7ysFjA/MVqE
z9ZyDmxDhHJoHzwnuwRbCAHaGhig2HC4ml5WBnsAR4MfE/IJGPC0qB+tAxXCdNWlk3EYBT/HDEcU
znI4lI1NFIWS91i5ryM0lQPipsfFdvJuUOWH8MsfDEHVieiyL0HdidwftiEnGkJzheo9waacuFfF
BCEohw8FpEUGz29jV7yE5O3yrnWLjDAai5hvxjei/JhluJJ3FBd42vCwn6UEFnHL/2MfOsuPWLNk
L+PjS+7gMJ4WMfUInqVNfN9cC9s9YLf1TiBid3Ta1oGh5e2FllCNlfZtXLLwNbcupqvFHPhtL5HH
NF7+W+NO+9Gygbsts8VPh2pHdSbyfbw3stP906SPTAYYfdE+NeStpGdGe1ExEXKO9oMP/OZXhGTf
Eubxq8eCLJy06PZZrE7g4z6yhVzkDMbRk1QF9qaH/RLv8vNGfrWfZTz3ceS1ZIprIqbcJNAIf+Io
ydGH2p4OLf7nitpDTIYPPi2AryyISeA09EPIs7MRXh2jfKJRMBrO+gBjhnJggnH7SXiVtnx00sL8
uDduTqHfAAVQxNc70NcDeS/VbxBc9x8SYyMC44gTWA3Rl12+W4ey6+t0Z8mYMwyKF4zm9jSdx6w5
m7P/zFMc+1hhdeYTNQ6oazkZX15wWHLF9ab+Mvd0e124VOv0ASr868h/oEVNhlm1aKozsa9GC3nw
uSo9asrLRDDZPIckT1c2iZtCTTAHoukXVUR3Zeim6x2dUmfQFsj3LgEgza9iP4kRUUeqPoqv4X8N
0yn0P9a0vmllnyjgBtQF3rfTx6lSxknLEWtqjS5ulvVmBmplP5Eyx9oAlfgdcmXtWVevcMoyJaeD
+7pRD9sfD5rNo8riNbSU8uU36Z0UnXzj0D7wRigcxK1OWNpABwWSvUHhSCmPy/z4iQcuF+ZrYMVb
5SCpzp+nhskOrCXUqK9V98rRuaVDBUfHUxIvHCaeAwjTbiEte7XC4OmrY8C8iHAIQE0BxRkHoOU0
eKr2TLhHt2irO5iGNRmqlkjkUCCoGfXHf5W0O+VKCcuetiLnD6ysB7cVgh5MCDYvkWZo4efJ+aYd
oeQOD1/Yu6PPZfVHNhjiL50Qhc1gNeoE1wi75N9+FbrzPMJhDU04C5uoPx2QzFw1yVxbsbcnbg5M
HRx6yIH6C0wMdzFFbKkx4246RU/nrKP0OzEtcgS5jgVWPG9Z/aJt4zuCTFkuoskb10m2RwJDMz6D
TrR2EB3l26tMQfsx+UF7PqX7VYKuEDXIjZQXKLfX1wk1HvGlK8NTC1ET1s7X8kJrbLpUAWJoC+sV
9TDTS0JRsSeAOE0wWd9srG2knX08Y3UsWj4z9HNVuHwTRqRtdROV/k1ktw45LXPKDyX1SvkVyZ+Z
jvBPdFpPu8UL7iSaCvDk8V52mfW3u8fqRvBl7NF3xNs//2rhKao/RAS/074HG1hFD4eC3rBEouXc
R2fUGWNtr9r6Q/O5lHoFJJdHIEbDmq1OwIITwuBgewpergzSjsk/ocF05sGByEhtWgWduz0brSFj
mzzUwTj0wgmV3FTutfbCNIw9RbdGKpilCW6CArjctxpDboJlYB2w4EUQsTAzfjrCDgtrjm2yFsre
wK+2ICvNvz1iHyZKmCFUuln1tGP4RwF0I5SaC6BRUttcjt03q2XXym1nzKg7eNw5AyTFpvKy3A8F
sEm/aJ/bXT2QFwcQIs+HUvHye7mCKcRP9TzHGyou/Al89rLwQ2En6LiPiyTkXlyzZroRw3G0sek5
7ocBRTEJYyp0dbCRBbWmfwNeVmhrPc9O5E+eokDz2XYsHWrXhysP3VnbjTTIMPOBPnOOaRHVTerL
r6Tsi69mpl+4wWhnQisZx5fLC0zVMOYKP1GG5qJzR4tZpa6NQNam0NAtCVY6KBS0hVET4ksAs7lp
WV2nsren7URQg8sjVqAKUGtg7y3JLIJGnAntbjUQd/meWroTecCA5pBjiN669ozewUEqSrub878v
YZpuXlU2dWvS06fjvhvHL3faqSDUU1BHAprE54ppfOP34dSV9HgdEdv0Hhj5OOIGqQ4GgBkkvT83
uhdL91l+FLdl2aDDQfSTbEx2vSDXfXNPuLJzVzQAANgNeG4yb/Bngjj1rklLRKoHkxk8eCiZH5wH
DUFCPKofG3Wnwz+Zd6BoAFBHHle3BdoXTLOS/+64RlSUF+e2BXHGbIv/FlB3jkET7ypZ+eyGxymk
ku1lC4LLI766DogT6cBgP/ohn7ahCrPuK7enEdQA2ycIByB/qkzWohMusNQ/dBlGBmNYcNAbbSSa
6467/AGK2qu6euvjFsuHE89aqRmLd52WcT2Hr3gB7xvUvisMFGYLlwb5ieNfcGcmeDEewoqyD0XJ
al3QVIw79JLUnjfA5ooxW75tdWsWPeCqYl8zSBYuahDHlivP3S+DoLmQJBai4DM2aXhOCuSO00L6
VtJlfUciuNIzVdjEeZdLkPp6AalHRukqBHBpYRL7thNCxIzxjIgxZYxa06DgtWKJa4qAIHaGLSjU
LuS0zyi9iBS08MdJhprVR0cxhgwE1E6gdlxt3pPOOrn4Qhv3JMSn2G2fZR5JXcJ9gqsW4CYwiUpi
L2Vf4FpgQmhtlBkpKY5eah9lIx4/ZGfTSXdkYb21TVAiMO8lPNk4roOk9w54cKR3OiElynvGVDFD
J4Oq4BXeWhDhqfN3yOM+SWSfRiR6VdSWGSXCEki/uqzOEHZWK5NgSNz2LyEyPJIz0E8BWFdigotR
8bTRb2W0SAOSyiRMIVOJGBXw37FEoekJAbhNzmN6XOht75dPFRH3E94FYC0VwXyKr7R+wtEy+7aB
OVpcJqYyiFT6x8uTe6NTqVODC/g3ykQ9DRR+5DqVs66ERxo4lt+55QoAQGPg+6eZBWs5dJuUcu0t
DgziZa1MxceeQ+bjD0SZOIsuHzzLbBmpDjBY3IsKzi58VHPSHDw7+smBMCLq4R1R9RJNYTFsx4SO
OMHSUHo28ceTkx2ThqlqESTj3wCqrpWxe5MUapwQpUqMA1/ilx0a4GMdOOvo1wdUy0dBWFcULhZU
66KfHehrgXN0D++Tp/sCA8VkgBdbzk5BbUtEIMGt9jVWNvVZToZfsTlCeDYtWOJ7mQQBubkemDt+
qhugLJywyO3lPbonUuZk5KW7X4VCpPI2lYTNQ/eml6YU4cX/Sifyd+GOiIYVzHnWEFp8m8/Tmvej
ev0JVRZi0ymUJYQ4A7cTMGHb7JjJxZTuUxkErzIMdcQVu+jJwA//I3idp6bTsGn5DwPQW0R4qXGz
PKLsj+I+r4Kkd2znl0FHyYrufGFTCjq/S17PeiLDkN3mDMMai99wJ2ZNCczzQKYLiaOJsRd8Vw36
WGYgZH9YiF/lOnbOiSIhmwv8wSdX4qXunWUv2FyyQpXE3v5rHSMwnw5mHAZfA1rnxdEz5qj7z4EZ
mCs+D7q7RrdzM+Q0Bs2Ml7PNqDVNIFl0a8hTSo0gMyMt9/aGj994YUnZ/UFezsaDkm0w4Amp5uR9
j1rgVTcvf6m5Kov+7pqf2DTntdMW9OuhPHyplvF1UmRt11b+Ejw2lSefkfyhRZ1LitqywEBOIhi1
OGZHhmX4/n6Oj3emyCvHAGkJm0oPkoyPMus61dlfsjuxDcfP2Nbf8OO4gfDmSi6EH60lmVtJP902
HDRWnb8SHSRmDB9KXNAQ/YH/XcrzO2ygCHiM8DHSb+i1/V31QJmNkvVdZsf9toQk1xKvJivEcp2M
nid7ltPABwfvMPRVzGoo/rVcOUVEZgvvn4zgVaYl4GwuT9qXVEF6MzB0trecG88myh7yrU5bk6OT
azBRhWVsveWBHJNModY6qfFJy5rUve95ktts0sZEGKlOtsnOxEComdJjnTgvJsSibA3/pEbMhBB4
TCFVee6qsmb0p1x1IQ1f+x91+35PI8didPYBzAyqRxwzokpjl9mye1lt47vL9FR00e+DdbjUEzoa
Aqh/Tn7ImIM8aQtlz3olb6RC8TWQH8VPo0FhN2cEMTLQU/WnS9FWaVoNSHZC55JcFAVs4YIoTtes
xNMJXT324h0yeiPDrgzOe3xBHSsYKW2LHL90ZQsr2v0wxPBQIySaVa5IurzRUm/CSf9zNGoXQQeS
tAwh/GO35sHgjBoO+IlAXG9J2oWNTc9h0M/Z4SqB5NcK1eVBL5kMOqlCulPtFhKDpRh3Y/O2yPak
FrKT+FCJ7sibcQTnf3kk8PSVIolKNWW4nr9pLHJrD0PMAumc3tl030AYQcQAoSiLYONzi9sGyhs4
E1HBplauns+hVEIpOcgWg4e3BhDBo6Jng6xd3PKKlj0U5s2gD3Mces2bIQUWdS+JOzldqQofIjiF
DyfRGZU4E7hnpKE+yJRSsRS6+OaP0vZmU+7HabPDuoce5H2cNzcq2zL7v+5GBPfDuN7i24e7ZEyQ
UOfZph0OPkfXarttTq4fptQmEem1/+MC3BqhQbziOvvo8sY8eQjVavgPUqC6ohzhbp77K4MSU0FT
bqqKQVJkEbTp0/AI452+GBoxQY8+n57DkRsGjCuSDc10YEHqxcjIzjnFfgA9BsrteZzHHr+9NnAW
CoF7Fgw1Fw7CCBVrrFb+Zh7U/QJaaaHdjBouxiVIa1VMPMj9vGyO1PCU8bYP27LmnIq971BmnJG6
vzNnYRzdyzuiauk734cm+GPNxFD5OLaCxdpx8m/hpORDHNqJQjAfRACEWq+eNNG0ABJOeCoXAFkB
RJCorqgJ2TAwV4kKo9blmFSrkzEQl3NvmKAEkC3jgPI9DfsttgcZG5VjMo4vTBC6KcbjzvPDoLiM
0yDixQa94eLSO6IZFt2DiutowlxFjh2879E6mDtfcJYfUbnKSpx0NQtcrUyLWo3idCYhH6PutrVa
9rChLvKQiML7IXqPdPNel753LBj8QhS8SDyxffQfLwvL0cPDYcMAYbL7etqp3WTDED20c5n9+Uex
SbCfcDhZT7vfBIYEiaToafuESVTpFDEc0o4yM/NtY2YG++1rl3m8dymZQ6yhMuItt/jE2ejtzZc1
qlE1xPLxAGSsFYr/ukbt8sKItnOxHjuUWdtsz5zMK7ugJlGcj+XZnxJGCmAbnSkHU3NnytnQKtjg
lhjfRqsybJPFpd2V2lWi6SD1P4PrMQ9BKjiFY5UaknsHhbZF9LMMpSRRZceKlYRFs/yl2NpTWwqu
Jmnfpv3ZNGQ8bbbXORr8uTe8JjUoMHfKN5BcHfHf9rN/+MKs8V66AXoVHsGjNgpc1qNYPvELJ2H+
hhyex/nRTMq/6SyPEWBSzpTRf2RwmPTLTLrhXuDxS5GgNx0FRSxIYB6fpbXsrg57jbN7ixHFusBH
deUFDRs+DBZKtrUgnqA/6dcoG0HIFFdKiyD8gCt0mIfDAOAbKmxtVhnWU3PWgLT44GCpbJCUxnHw
uMbZk/tpqsImLVwLFsIGe1slEz4noQowJ6n974VG3eoRKrLe0DR1UcgVs3AltQAKu7c0AXrIFeC9
G4YWGEOuf9d2q9oNRcVWhVCyD3jhCK5hIP1rDdNRlt4uz8i/AJqkk+SPeIg/Dplzdim8YJUbOKtT
MoD8u4RXLQOAAN1S4Ao6UrgrGtRbmQ5fQgx3teVRrGx/s7mWGRpD3jp1f8Rbs2rqecBDNbAQyJgT
4QSZZIPAmZhp9vzBfHaPe8wSqz1X6CQyr7ci464nygjrF+w0fcDhU2un1EdaLIFaXYHjQp84JUPK
/raGcsW7WQKrLr8dzcs1MsBvBZUeogNVMO+18ro7wnUFIMNDE4oKQqsTu7S2nGtxduSmZjcjgFkE
LU/kE/719itefz3xZt5Dk8PGx2t/+sHoCCLlpjklBWVL/2sP7qcbR52XWhIGADWPJJwtm1KgnSHs
9tPS5wd9SqVlOttGOSwaKt+G3uwEh3+eSLVTSz+ATbCn1fSm6vcEWf2LyNj6QdJbgqgokt7G7mhC
6VN+WYUIadcc28NBisGN9G+cxChXgV/WS+0h34hUKhciDuPgT/8SvZodZgVL3mbFkKlvPz8C5Uxc
GE1rluG3UqEKQeWJ4TMUmmXFdD5Ee6XiXrpbYEeP0mKVRlHeRW4Lm7q1krXw7H/giWvaZ1V7yRJe
RfX5Wd3wj9tS08x5eeJ2Yv5kkQVleOOaV+zxMW1VeEVfGUIr49johSXW6c35PxxuTgvGUwDhyOL1
24icJ3y3eSQBUD6vEUMOR6fZ3iczdrKJoXhE5VmrA8wcJxB930vTAECz4b3PSeGjiqsNQuKyq3VY
Z03I3YFxdqPgDl7WMPKZjNaZ6qJzs4uxRHG6VjuW/9yAV3/CruYLnPAGPn+XuDLo7jjxQC4UyYtL
BDeYHu2qT+83ogPAUtBeyVgT+Z4/sAbhuffdPqu/j+49krj6Zg2Ux/mMwHj9O1RyKp3QOdKj6z5n
hh9DglYXSuJTcdrNS8L/AgPrDYZj4feallHqFTQUs7upKiF4Cv1X4/Vjd/tlZOjezsSA4rfL8p7l
tOn8Lhbmeddi5Xq6AHIBQBeoQHWBqSkU4hAYmkTzX6uLmFF5acpOHd3SsIgnESUDGOx+w+HClvnD
4TnMeF0YhhVr91uwl6yIVzOmVyuR8UdyIDTc/m1X/mHelk+1OrcvwykhWlzm92A1rDowycGKGql0
E3ZMRo5Mstc3x6rdjRpPoiokXcUnfPWoV/Vp3shlEGpsk4DARcTeQ0eL8TPo0qW/9C4AtkOM55lL
gSRbeB2lH0MPuzdgVAqJmWp35PXmucrpJAhxx+xxclu7wyxPc73gZ3x934NBisVljuvRp4lNff09
RH8Je/KuflyOiFgzC0ONz/Vf4GxnILx+jHCiN2r1DURER3Nt1DD77WCt29uBA86k3pNK6UbUwdxW
Hb4o194tZJ/5apnEABirYsF7OEYlSp5i5XEmDksGmSbAmBXnTdrY4WWVJOkZEIDTyVCext0tqD7/
gYvHYrFLmtnJsEY81YmX4687nTZ5tnfA20nHutUTKU310Jw0fOYJzMDTdK2Db2w4oFfpKsIcTp2k
+WMsRz54WSJHaY3xYZC9RacqNMkOBl7HwHaIb7m4cU3FQ1KPRNMxvY+VS8zzIbaQ3XLihXes4ucD
pPvD7kgO/W3E56gucr0o9ejVbGifAIdYpWnr+r6jAdkh7ftcfEzpvXT3O+u7xvkvRQ33Kwi7tcn+
iyqfLhYWu5QCVUPlz+ZP+R/6qXCJ6T8hT8jpXWuqwHq8auO4n6GxQUurdX4xf5PCbNo0Ckr4XS0x
MZKBvYBzNy5Pphc2KNfbo8A6azc/jsQdjkUrH0Zk2P49CJXBcYA7LiBhbPfIHrmkoRS7Mz0KzZwA
UopUIyp5lUCbiW/NGVvaGaXrevBwYGYDSILYChxzZioUtTALdERug8NmEnEk+eY3KMvPpiSqkME7
3YhERk6F4xiwXwRdi1iVS1n8ep3vPGSnQaoKJwazRxtsmQcAKe86NuN9zJM3iH1jWe6bOfDTG5p1
8bbSFbPfCoOkfCLai4Z3j20Ni4qJWD2ks2ZetAwwEAMCeApLTKaM0530uG1nkDstpGsMs76Uzl02
ZkuXxdS0YCHZKi0XwMufbH8kSn0WhNXtTXO5+uJbWxghfzQI709P+M//BAdtnQwCBbRmbThCX/BP
6u1RAf2iagO4B5HUNJjnHgVBeoaEHvTcogIE5FiCAQvZrexbX6CiNW1eSnBzBvDAJf8252WazSQP
xfXcVeUpXWeW3dizjGwp1tlHl09M5iHZqYDO0ZjjSCppJgYMe8Gt77qGuDz3azsUxkqLsxas38Vm
I0LaEO3Ppq7HwDGSkkMm2QLjnplndD6657+1lqec8/m7c4bQThf0wjGxy3rArOXpppJGI5MyQAS0
/S2x4E45/8FHbtA1BoGnk+JVYfung0jwcwNkKmglPQW6V8GDXyhTdjDec0Y5mZWXeMf1ANqF1UXN
B6NucW/U+9lO4iIboJ6DDHUeEIIGcjY7XwbQdJ6oDW/cVJtYnB/zVQ87dn9/pKR89CrhKEPU+XCz
SrFJn8xf2P3B2AKHSmFdczlEK4Tbs5rvQjrWw/DG9ips6c2zkEIQBRjS3kMAmd99K3PLjT/qTy9/
FmRnK2gdLJxn1PZrhE8HDdmwvnXDO8NCFnRBVTw4v1CQWrKM4sTTSeVdZUqkJfKbialh4geQuT24
W2vyOjwKMweFG1x3FcQD8mbDtVoUL4VE1q/4lFskqdh0XFAPGL8sJdAKT6NOe4h3P8nwMBNfePBB
t65+HDQ68UWGZqdMzCWBk8Y1SSyDW7nj1IAZndBb6yR+wX0EX4v/SK89nIYZisu4jmvDBgZ2UoNy
1U+sb6+Z0X5NOY2QOa+F9X1nrDd8QQBI1BXFzvoH9HFcTpd/yPmOU/q6Z9Lvym4HOiEhc8pVENoN
62FPpTRZKtaceo/aKCMjW8eHZgguhjWpl869WHvobS1R4YXaVOlERc2O7b6Hy7OksRtThsjI1JNc
D86FECNAsk1tgFlczFfSRuMK493bWiKk5bIl1s8HrZVKywnfkMOLWXHzzOZ7HVm/4lga1DOg007n
YEU1tzgoG08Df3zYFNUzzMVSNMX00Vdh6IqfPnDqjCZazr9u4uPny3WZ+9OnwDg7So4qU+htCm+n
nB0TbKQE0X9y7AY5xkqZ33xO/TqMtcJ95AOgS68lVo5z2QCaMxOlvQoYCpMikgU7GpfYtlZT16iK
+kWdiL+4T+qd59PNQ7sr6mCtFW97z8KsbyNHESO9UfdF7svjKjINXKeowXC8w/wXyRgALxG/d6k9
spx09FjNrRKhtiaOeMGFWaBqowCZUN/IH5EQWb7aNw72MGRdQEdOAwBj/uGcYwJMjJ5vACvSgS+u
pLHShLurv6DPI7M2tIE/lm6+kK63ZwYvwex4MKG2c/I5hG2qltjhxfoM0riV8Fbp9YbBIEc6Xqyg
mJp5aEpo1PQti+vNfdc9cZfp/gTzWYWhhHIbfv/xSABs7ypcP8b99q8kdUtHD+UL6NGG+sN4TdRz
+0oXny6rpjO8JdejsqZK4jJMDIfzAFTuYgxufqJ5viG2BwvFT2aEb4D0rKGvjKEfvaQA0VVOagDM
+QCitkz7+tisqeBOL6+OjWO7Mk65y/VmrKdFbev3wefTiktgjtfBIbQs4umReIUdGEpsfFjVkRno
yG4z3yX/29oDU3Mu6HmU27E1aSoI7RpmiVZj0KoPYRUvP1IJSIwN6i/dzA7pM/VXKO97qH0ZYTYV
WewXyomiys6qWsZeNYOwqdZSLJWvSVMDXng8YKQ/XWtgWqOtqDdYOQv1bipGyHv8YsBtKWCAfH7Y
l00FTTaqZR/p1mrx2FtSkFXFYB2MOMNq4f7tM8hztCU+vDJ/7OOZezQvy3D3IEny0+XHB3GCIYWx
D+Mp+ZDT3URKDv/G3/GnLHRJwcESgwjw3048Ft38RR7NIpJL7n50EhSelZ0sLIZYVeLsQiS40a0i
RcRApYOCaBcEmzlUs16wex4GP83Gpbyjh6XNwsIbpnjuKPsPVl4tUF+iaic8dKgZgpBys4aP+bvG
i7IAmHEzh/xwSLzvyVct1ZLr9YsF7cvvtD9R+v6S9AQezAY+UDjcBvKz0//x6wr7jeeI/+jsff2p
8PpkHzIpUilmozomcPlmFyV1CphBZNtmCPkb6TJzx0YsGi9OOmySP5sX6GFMnRcoB9LqqXy2N4g6
kS2seSL8BCNHuKAMXFxieA+ge/0Xb/orYpMAF54ZUHvJQgB2Y591tgje8Cw290j7mzdtu1glpfsk
qDq86T1TXKVQb9EnSTP1WCeUMPzC7qS/orXRlxLURhWeBu1q0MsMMO522LnHGpw1e9jOigjsB219
PK/Kya/+mWe1xRKz/5e0HiR9dt6tub4GSfimbKiE90pkKsV7bBDg4Kvg/TNDyME5EPMy4BYcbw++
YLTZsHFKXq5w2O47PzJ90j3hA3Trvsm7kNJ82pg2bqfWyjCLqFultyn17prIsrC8Eg5LhWchnG2o
fb2AeXzGK6jtAOr4Bq5Crojl/YKFPLyUkKlXCsVkPTZfth9BwmxyUQ1Hs2XyX6MJKqE9Oa9Dvij2
LRIz9xyMAyvzQt8Agfto8lfhKBtbM73kvXkFx3vobJ9Fg/vWBoV0jxnTs5Ip29EwP1ID7ibmqpWP
s1WiWw8xXhvskdncrvr0lM23tvbDUjBu8rCNNc007zTwJLW6mIH7YlD//skfsqH+zMVwYWXFKcqV
sDjXyukTRwtdGV2Pzo5C8fq5yi8U1pQ8m9DvQBaEDgyfEbO0EMDvHnI2fKm2RW7dOvCh6Yz5i+MI
FW4NBF2wXEg/MEiVumxQr97SGaghpHTJS6/9s1bl5Qe5zGnPTyP1KEJWRur8aI+DOwxknOnxh8bn
7vP4Nn5LH1ACH+TeACksIAk4Vlfsx2koJn232fYzeiD8y19TIv4I4RxpFUQPLeQHOdoDOeC2d3Pk
/uqsYt5B+gECJVfJIqQTnJeEuiBACnhUSRY006GoH7FFou+RLaomprxMlifRQTaxU/8IQK+Yb57E
zAGaH6NZu6kumWcrjSwypmuye04gCsinR9tjtka9aWwCuWyXHqUNGH2AQlf0/nm8UIIVKOmNaIlr
Xxc5fdeHKWR4gbALOpA1N8ooYDoRPkvX+JRE1yinXmvomLlFIAEAi5hZvEt4reQ/E8lP7zUODaDg
Ti8s9YhbbqVlVjVrYni+n11jGtbPTFqiZXp4KYhdugjVxZJTaX9jFYtFlYFR1EVYRY+wvARJizB1
JeqsMizw2bp4RxUFdgs0p8c3XKwi/UcslzuE3/vuc8g7kzwHW+OcWZjBIqEq+aA45MH7n6sXpizg
FZLjEIMGQVTtpI+G68Hjb9ReBf83kN90ik+umYLgJysCgseQQhcJoM4k+jsp1blvt4hNCx5suYQP
eVROXx9BMprZZQ1jhZFUX2EOrIyIl6x5yh5Nj9Uw7gDT0EW0D+AB5SvXdX4p1QjwrBNya4COa4+P
g6kMyyB4ZsmSyqzjfoG4JgmUdrjrMvM0qMrRYHNrtKtUkOOWUqQp7Tto3jbgtNHlDlIi5ccT0wpp
jDuJ6BVWS68037nIfFc49Z59EyvkWyh9XoaJEOWQ6KezYm2absAR4OC7RcPaBDLg7yBcI4i4EhL8
fQTyJMUNo0QRuB6LOBCkDyW+7fcDWDEW136cb7/R/DqfgBfcgYUF9RIaUSZSVe7b0z6WbXSDt9ZD
O9+7TvXyrEMy6r+rhhE9h5xRqBrV4hHT9I2yFnvS1T73Q2YyqMvx0N6ZNdLI9cl4jkHDzUTs0TK8
8Sb/fHd5kRlU8zFvHvaTJBHnLXRYJ4AtucI0iXEmeIP722KCIJxXac/Y7Y93gHX9YwLX7c++efz/
Vw8qalScLp9VrjzTC2+z6sA2QvFefBHxSoNjt0DfmEGalQCd2ynudOwedA3UAEj2ak4ldrxZZfxY
g4gktcKmQv3oMhkV2N1aEbYUEoFKxtEEHojufThAPStRvxc82nUsePtZ8+Oj1ip1squHZG1FniI4
I+f9bRZKQ4QwRuHSN9zvgQifZuG58skioom+4cKTWpW8S8sE7VbboCS0Kdx5c0ZfITWAK0OLQlzX
yKbX3qPvdAxgDva3JOZzhrqJxReBAViHWA/NkRkLQWxBRYbUfwdypar/cTlSSLW3fuyrw1DEamk1
W5h6rDEFmvWjrf04l6jdXx0l2vVFdbP6tZUAXPT01I7XhOTqGRWY+jhh9PvyAYny+QNVvYi8o8NN
Ksq4DSRUYWBzrK23SdNwwwxSHOI6LmQ5o+yXCL+/xDBsxppcjNoTluFAKpn5eLM73TMniKMo0FWc
yurmzYCwzmx4vbUOrzOsnkVLJsvAY9qO15Yu4qnEf0yHa2blBHbxEguhFt3bMfiRUKt6Vxp4oDav
ZzKwW3rRRgIRdNie4e9JeSEQngMWaNR8q0VmOuCU/soSxBMbxgAjnHkbtiRMBjjzebVvki4oY0jR
6JRDHBwN0x49wSlP8PxxQ6VPcJmWqFEnhXgrWfbCPVnfyu883Cw26PunERvbSJ/itVtrOTtirQpU
tfzCXQQESCz/sTZXCeYFnA9ZfveZjo7NWES2RLaOOUIMwt2X4s9HksxSR8duVHFu8Z0ROiVCP8Tb
aJ7GwWT0tyM=
`pragma protect end_protected
