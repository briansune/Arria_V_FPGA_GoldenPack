// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:30 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B4eJK3MPMm2tpAOGpTZPgBWg+uqY7x+a0sWL7G153G0s1r2tKmjVL+LCBLVtjB6T
R/jliWFUc0py5sOCyOIc0fA8lc69i1rENplA/6WoeRGI6+lY+Kx7fmY/U9jwW0rV
djPEcK80myYz5tAFhvqG/qsfwNvk9V8KePMVVCxJqKI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5200)
aPUf0+pA6mtnuJ7mPVgTs8bOUO/Jk0JwzsK2Ap5d0NInf2OXaCOozu1rvaJN42TE
atrPGwAnhWNMSK/bPIOlnaQygcYflPVD3gzJtdHAFvH0hE0fvzoSjN+xyFcGLIbh
qM+6MQ2lu7N5Qtp+8cbuC7qbdDj7UNzxy48uTsbhTmVX0Ukc2G8L9I6GQSHNT8zd
5h64YniOeFpdZ3K1mDo+Z510/JEd/RvJT7A/xjx/yNveBxIYdzGJgNu0PAtkX60d
8Iuc9VFwmt0nAcpag+46mPBmnNqo6cgahPXBvQHSXVa8IooluZRGmMxeCGj0SQxF
jWepUegiUeb/Jm9ZPX1a7Ni45ibsu4mn0mB8vQCNMlBACLKJ0n06Sb71WO9G6Da2
EP6u2PcQPO3eKQ1iPVW6JfMJRb8cQ4MmI9MdgHgJzKzjxzspLVFldaLdTouHtbn1
VjfWTbENWM3bnr5hC/w9Fu/YYcyvJNmWbGHv70pseVfUH84i8ChuUHbDePzP70Jp
98X7rnupUQvPNkuiXEnVjxV8r/a8OwdjIhC/jbrJsR/C9FZB2MX06ozeg1HjEoW/
KBCrKkg8hflNlCmaWUlsjWQ2TWJC4Ux/2YeHVQoy4lg/Oh14/Fe/Gjw7AS/9MIH6
maEMnraFfXmRvrRe1CSiH+g+xFL2bA5GfuDM96VZ3cxViFNNaa5Zv/QCuBDmUVsE
V9IKa1nU9yhtxp8XTwY6UjZjkYW7SBKX4YW6YsdD2z3dQkXPDWbJEpk/NMEu2V1o
ds4mOZgcjrH6LrVvXPw8Eh9qelS+Sa0K+ZMSh6THgcTd141xFKpC6yOwXIyuMMov
znZfQ2qO3XW2SXY9n2lmQDl5W8GSqAqMQfvA8RcZlb41CvggMGmTtLK+80X1Z5e6
cJxi5l1qjwI0Pv9sVxOrZD5t1rqYrytY/Ns+gd1zG4Ns0YMw5p0KJGRxb1/P1psC
xQTL6r3AeXd7rZ7lhjjJxXIyneyubSNQeB40cJYQ/AXBll5oTu6GA6wA9Hy9ma4Z
kqtcma3PXgTGs2JdF2pgzf7x5fM27U87NxOgVNVM+KBtZUmaX8YUwK7tyIqxx+NB
k8iilKJ08L2M5DpwFMTXrRqZqwGnLfWMdhmsgiSRrTrbmwHtQk5gH/eeZyQMmNBi
D4fmkEkMJUIXOfyZv6xDTdcARC0W1/lM3uktazF6zUEMyAVG2pyG2eblUQMUssAg
+6wV3RZCWty6etMRFf50J99vNiKtV4y/TUpZgVHS0nzJhWFwrMgIezkQRtoXNCFL
z2YEYW/TBkDKXni4sjHg5TbZo5KWOO1rZytexGLiftCFzVduWXeL5JSm7lFPDi5j
ZK1YxNW5BJgKsFh4S4rDiAmBQ671UU75aLHlLaGDLWIG4IBmDHw/CeUEwvGzpQUx
5tDAi9436hF0eD4eJzRYeFdWZlUgm7xf4xgz2RMQtWotBjmJ76vVoOsAnIkncYvY
bWLRv2ewuvbE6NXJ7IIRMnQ1skGDhHwLvgPEv3ZnNJIbGoEY2QId29ZSahxzF6JT
1/ETeHVEx/xMhJVAJwFIerxzYZv6uHgEX2AUjMorsCOjnzGXoytX9i69y74oYCKc
SHRVIy5tObuowg8gNSPSaT3V+EPpey9ylBcWWkGR3f2Ca3MTiL4PaZphlAwg128E
0C0/eHvz1dkftlx0s8CNjre81TQ1WrZWmhQsSUAHcCHpfH4ICjVUTDNR94uqku9h
vWap1vTAOr7HXcCv4Aviwswvx6iY1U7viFuZ+IRpfwx+zRvVKx5B1z3s9vOqdDxC
jl5QmzzUvDe5lMyjYMOV7uDpnCWNzUDcJnFyiBq0K65NAf30JMHQlQRqrurR4+9P
UQp8FpuXZH8iulNHEg0v+AL976ao7Uf6z+likP6TapuJ3A3U0du7W+MCh2ktckh1
YYKq/HKHDLRTvkdpkm8z5yOGZitHAQXaUjhsqSojwT84kxAzpVzj9t58MaMkBslw
8om/i5oJVrXCBV2oUVbtubrVMWR4J2QzVyOWDc9rBmfGT6cNgwQLdq3MOs9FuYR4
BMm5WZKI9dxw6RcVm/VpT0dQS1ihxgeUjSGhgBSZUPaqTAttOtVj+oidvbVndk1R
UkHsXuQiBh2EDNAgsdviqgdN+hlsumkukorM9tw8dm5unNjW1GnDDp90dAXC3SK6
CGHNsa2VW70xXK4nv1VpQBW16mvohU6s6a/MfnIy0dElyAxRu6RkaFqyfg2thDRK
rNUo/NmpccuRisKItRKXFA6ARN+/vyObeHI+i8HH2Y3mXr1NY7n+fTtbtzmJS6PX
HeGzOSwfNhnPfATsmg/gekZyJr7k3t9Esq0G4sR3OudzezjgoFM7j9QyCdVW8chj
pNvMUk11Ht3EnstyjSj3htd2iT2L+nXmMYhee5QdbSKNnL3Xp140C8WsHWa+zGX4
M6tQLqWFrQ1bvZ+6xpNnFX/SgUrzBjK0scJAq1xOENj4/E0B/v8yslbRSvFes8Vb
T/mN0uYkYklc4lW1UUd1esbXmRDdokUYpqH6Gcsw5GVb5+9yDMzxvWVl8ZfDo1sd
QFt0wfkQKTXE4fZDWE0voW4IOgZGnzi/TFvyW4NLrLmg6YReYchsM5vb/uQwPMUb
wLRiNwnSLy2skbV1iCz1By3JPLYy1XwVDJNS8LJ+RuZPXSp4rK/ZBKNZQSuc6kKY
a5xLK/9NMkUKaG8czodkyDE0grOH9l+n8EFSSG+z71RS/Bz8OMwUIm9cawA22/fW
HjQ6oXZwW5d2wZe1saIl7pTTHUvLFAtF7Ekszm4W3F0iM10kot80crIt/Uf6TtHh
as5MyorzOZdXFLQXjID+QcVa43oBxWOPLgmMRC44a3D4uTcSyuEW5qCbIonFDR9m
H/DcOWNY3Gf723sw4eh+RPfBv8SugteyF9+OkPfisr/1KK/dKS0PpeDCB+mjWC9W
VaOfQCFsW5UwWmTN7CZs7tpks2JvvgjyyUF669r86oJ9PbL5W4/BZHAcZ+MYTFez
siFzPjUf2cMBayVHGvCAsMwmMFdGghXc/sROvFquFRSxWyG15RDigM40wbh1O/L8
oahmYFOlInTLNjOkfD/+J75wx/a5+6uBFWmtr7e6hxjvYT93P4PGu59FfMlZ++jq
LY1u0N5h7HPyBucter22lO7UBEpW6BV7wM7yHYAJDp7QljXJf/bdDPki2jAPIUlB
rIjetSbv7ncGgiFIXqR/SYrEw4jd3XrJbCEUW1N7ziae9l8cMaRV9pca1ag6xkAP
PAH+aK1T3WdQy5GF8mSb2Tsri8WAE26TXkuGpfCS3Cw6n1/zI+ZaG8paI5hR+XGK
1kkBtzLEGuhn+mNw26X2XgSRmoIKpYEckTLCvEQ2ksQmV5cKorKsJNslV3gMMB/H
0KtkNTVdRXvsi0w8mMFgfu8A0SBf2Php3vhb/ANmUdwx+pRLERBfHfXD1u/PSOPW
FncJG1PIQrxkxTCm+1Ska6rCQc471brXESRu7q3AkV7CF4GD0/l3FNPbeLNW+jU/
BuDUgIDx2GpY9t+NuCwJHHIPfY0H8PJ+Mu7oL6YMZ4m81vKm0zjhXBCIKJl1DOv+
HEaEhRerlATM2qyM3vAz0wFwcexzYqCY/saaC9YGpDBvyJk+pKE/OVsz6WXzq9d+
uUnpt5Cx+QuoE/bS4PLV/YmREjT705orpyf/sTkQsUXLVgr/lbTz8SkOQ54KjOA3
X2wdmryM7BAVwR5YOzb9h9HmKvUc5shwpIHsuqu3xBMWfyfl21Ogvw4aa86Z7JCa
A7S3cg996V/nFImVknSqiyPH0qLAURSpZfrS9b+nf6DHabn907MQF2YwkZXMHMtg
DDg6uZ/yDx/vOwb+shZO6CpMRxYzhzz6gSrlHEB1hUrhZwzPqh1pfZufRL0KCGd7
sgDFT6yfpquSwysCbdBu2DuY5GydkbCgrFELjMYSjChTlgiWDg7J9u2ew/h3Jrhp
1e+mENXJlFHnZcA9/S1ydWeLpkw5qBZ5kli/yRCkonyMC/oXCF38UwsONxZ21KI9
QAj4FQc8TGNSrasimpIyfFmBvaFe8EXtYUtgWSWS8aexpCphQR8agDuD5D1dtltK
/NfkQDUUcBC/sSbBRblqjpdbA++h7gkfKAs2AaxFyv6YsxNXwxflzROH8siMp5OZ
4GuxlI8J0cmukX7C7SEEUaM+3zXuTV23rLNq/OmfUDcG9Qf4XAHmfRZf5cvAPfNT
+HAIbk0wDUi4kGwtmPTBOEXbhP45vjXcJtxt8cIayU3AhOnWhFbcL5OtXPl2cOT7
SVsYdVxH8iMDCK8S7bGl6TaZUMHnURdGZV833Xgk2MWLSPLx/n4U8/4UFGQYLfEh
dTj/hqxjqk0hIGPy81yXSYZds4SIaqe+U7TR+hGNvypw3q+KAf9tM35k9pfN+sK5
SQN+oI4ZFXL/367T9B6f4c322DWKbYOzwXYRRjLEJ0OwUApFhvaSMELqUZwjr94/
wOGg/qFVct9YfpFF2EEzQtdbcf0u+5qfCj/8829kDMoeAtgvAh4qwoScuxdcycbp
lQ2MUJS+obj2n7/AKsJ7wu4x3AD/9qpuqjomOSVhFDRAPH66fyHcINYHQtV6Ea23
X79ING4433pleXPTUYUFhOqNwxYtEAZVpfIq2v621U4Yw8jXnksmckxewP8huUr+
a8TWTUlbflkdXy6ribXuiaECkH6iTNafP4ZIKHLLumHsMIPRuUhy5XD46C3QgLPg
kI0sZ7s1DP/HkyYq/G76p+CMG8p3VMi1x49Ho17lvHTibfuowJYWGafnb6G3/F6Q
m5n37qNaSmKDvd5lIFNJJ0m1GsdpO2P8sP1J/3FW30fY59TtTwNmw8aMSks2MyNq
CoeIqCd3q2E+3aE0qGz1jf7cBkZoFqyQ/qhghd/2ApZgTtAFs8nn3WMIr5KLDWk7
uXlCKJON594Al9emBF/hCh2nU/93MSLXQGpwRGvxFgSlDe9IKafCAmtIcMO90ORm
Tdjs6QthgvT46etfYrtd+5hVMPBiFZUVwsQu5vHIIa7L+IjtLQv03dCBWX9MaC8B
Q1HRR9wLvr3aBBasUGHAtthbzvHaTmAhTmKIxW267WxdDsq9aN2MaIHnQUVu6QI5
c9Thm0NBHrCjtozbNYIBHURsLu3Wnh43CRlx4k2y9haBdxBtE/tSzb4iwxMW0Pz+
9bgy896zmNFnKx3CrMuOmMFLFbwnqjFxtN10m1m4pA4zW71zvxKJcnkqzn2bhMIA
deY5ye3Fnz+m4xEF5Ln4PLRo8kOzq3D6FrS7TxagFg3Ed1851Xfxnj9kHkk3NUuy
JbRtDzcah/0baKgqTZ5wYRkF7XDpXG/rqProrNEpS567vFmOvdnYnnHDI+V21ItA
3VGrAT8tjGjcrdwdTPCG0kS+PXkFuz2NricBaGcAkmvHZZ7TKPJQ7uVt5M4tgdlG
hHskN75HpI8xxwI3lJR5ooV3IHKRO5PNbg7skriohEhNe44/EtaAEy99GeTRCp+7
dI7S4RX9Z/sUybk542pP84pl10iFvSkS4WK/BjdN5Stp5kDtT4xocLmrzWO9B7aY
OSYMjtvreM39LPsqm1W2uJdtSjMaO6Q/gG+BLAR5uBMd766ExREWLEemIoqHgyfc
oXd0ngodZ13Ijm6X50ojLyGY8qbylj+TwU8eZo0yMCWDyBgRgINYt0tNZenm49jE
pVcKDl71QCYKWEmHzJCLzQeU/6hfzh/hgu4yJ5xxzfcQm2ZOEOzqYfLlYag8eKkE
e8x08Ww2tqou3m8WrYaKpxRQTqZKGeGBE1TN5SuxeciDjwSEG9yunUnRVjjhXZOH
9v15Nq2cN/PXds2eN0hZxukwoprccd2TgijNNW456S4kBmgWM/B8RWwz4Wet3aNB
Y8lQSMg9Srt8tIiEIIVaRLimazYKPnXxwBIcrGS7QxNGxFKJX5OqW4On3MMZdmhs
oR6yLRNZCEh7CJ4hxvt60WukF1gAOWzPPkmHiih3Zq2do3JNetItmjaUZTKq5itX
MIrBCaQP5JJl6K28KoyZkubsV2R0/uSF7xWAvjiYMDH+Aa+z0pWU+qE9bHmwX37C
vezykmee8y3o13NyhjjrEI9Hjk+85PxV23I7sOLBOJu1CBrer9z1g+Uduq2/AJCZ
CEl/3G+HMedbWUl7hRV/oIMIGxi7ctvJ5z6LG78WASb2PczzByVU+BoxRR3lU0+x
wGPIQZoXxmk0TWiVzSkhjhjy3BtUjXKH3Qd3p5hFYLXOQi/7XfYwr9XjNpXKYoE/
UDfr35yjTwu+XEOVKJhtGkl+M3bFOsBSADB78IUilPZI36GWDve8lSxQIOwkvF76
GV9JMe6cQ3PXyCxztQyW6/+C+BbB0cwojVtxtzwJNy7st5G96cmyJj9OTCboKdJG
eN//JS7Ml/uja8V+6Si4qh8P7AyZu71p4Wm+1/V5xTGpmcsRRLxsK/vSKyoD9Yv1
8tx4DEOBLqrxlWKB+FIwI7KOVH2JTakpsOsruYfoilSJImdoysgVYYjG0JcmuCM/
1JVq6fUIrjxwj7BoC+Et+NCODMmnupIkvCpFkAmTS98GitfpyzGAH4W84aHIL80e
c8vVEVoVoG7lZCDz6pL3oG4KzuPrU4sL9/5TmmZKtwRml0Ksbs9WgCFjR64ICeAq
ew5Sasoj154PtMiU7YIW0lW0S0AieGBoBpRDy27prCdI5vXeyMaigYBuXjG85JAS
AZG5Msee0qAhj6cvdkP52b8e42zIxpD7g3uUCKu0FR6moI3ZS0dKqCIvGsHStxss
2hbwN/HWBwYwGVQY9IgiZ0Zl1YWoodUObO66I7GyqRYQ898+LqAYql6Lrvj7JCdC
rF9BIMCe37NVP/YGcmVx70GLWJPqw4ZP6Kzd+d2QLCy0ChY7eJUd7pVpxDXp/Lzl
qTanjepzxSTHIi+D5PH0mA==
`pragma protect end_protected
