// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:28 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gGeWXuJ6AJX+4hT87oyyTFX6mfGtSGuSEY4ZLCAm7EFPMM+xHoObr67Jg8UsGtbG
X+mhLZ8aheK7i+dBs3BglyNWfcOQO757Sr8YmPCEHSlrkIaHEq9/90Lsl/kmPXxe
765u/n5VfwOif/35uhroGtvWxjZcKRmbWvIfUcvV7ZU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
BPcebfmzGqYJStT10JWoLrU+q3/uk55bubs6gdCa6BQxArovDEw69/0a6t+MEHY8
WKBYcFVBtuIgBMkqwD8Dzg9ue6HtyA3fiQuci4msWEA4q8ywWwKjtgwo7HJ8Alkk
0vzf/Nb3YolUE5qo8fUjBwr9ynw5x/ZHVzz7IqILinIAtzcs7pVCoFxbSRhd98NC
7EUIlIGuGCuDM/UsEUW826UnjN/8QZJBvgUeeBqfxqu9gfC6g1fCaE7KBmrLaSRx
gCQG+VVZ1EBiumFqvQiU5PyigQEunkckT5tvVSc3zZnmeZ9Cu3XWup3J18zohMNH
YWCcEHGP2mp6ZEdQkvpOgiaSkZSSrKApA9JhMMjRDkGebiavFdvDSxFxOXrbkR0N
ecaUcH4qi0LWIReRCs7y6iQ2RwBq2cShLRFQF8mBbM+nJEI0S9wVY2Wysy/++IKH
k6iQ8y0i1KMxcYu1q6lgwS2M7h28hRHciEjxUulJWL5YrOLPQhHMgVe8BpvmZnsn
z1nvjY3xErGDocUtQjgmqWvXuosWl30vbJsiL1l179Mu4KHGtgEJYJ17UBeqhH1f
56TdO+8q36cI6NiLuF6Q1JgZ8RZcr5Z1hzfwZOG32t4JRZV6zCZQZQrP4FSZ7mf9
FNDohtido57O1Fla5d/H7rA4vkLnr2COcZxhT2AP3qnbt5wVoACyTZuTaJxpejkf
vyGfs+HKMQxv4B/zoMvsSuYxNpI+5/biDrGp8MIG4BG6iJnNWu/xsDrzTUoimB0G
zPaNsNOEHWc+mgcRiR9Io9LcczUYspMJfk7W5uS6OFfPolX9GJ/a8sK2EK+ba0O2
Z5zbK1gM1XnnWOdDJ4rttapYeUUuaxlBDkIOFiBKn09NQYk0uhLzNlkxZ/pxYfAb
8/OltQ1Zg/reWCbV8qU0GhCf9AmeDTDOil+5c8D4rYdCOVHzdkXWX6qEECltONnS
fFRGQzMAWyx/e28ASWioHx4ipmfPw2T4anGhXb3ezwQKGCLXFOricuMotkn5i5bk
JVXYpcBDCpVkr6Rd0XFLxlk5Tek5xRG395n7bmGeK7iZotwYghP633HIQXqPPBsI
ibkr7iary6eEb3mQcLnrBYTVzzMRxy/ZS2otgyn3CFMLh64v8a2i3LZ33d3eEMoC
3TDVutsVJzCNHQl//kYNEc9PxZBK6iogOdvzt271kLVuDRku1dPfNlPPhFWufBQJ
6FEIHIsph8nJREedrYaDyM4g+UnP6o8ZpoQ/mz8ZmzQ6hscEdT2pQ+02wI2G8r+v
TL8RZeNZLovCgAU9dUknloXg1xg2hURN+JqrGGC2mbE/zz6gX+yfssBRN7fIkjll
I1yYDFkGEQobEx/XF7r0ELlZFzZF/8XHZnCW5tIxEHFkZdGt7z4qW0rQk83z06Ef
f2EXmThK14lDM+ghpqIbWUYz0rbw/U3lsnvOsPYrlq6oq6mbPGEAXM6DdwHxVz2n
X0DM0Xq8J7I7klqEI4fiecGOZpvwHa33HbJoUwd5mLO40dx2yEh09LOE1AUQZ+wL
fIUreh/c+Aai7/IL45LA6wFzwrSwITcqD0Zs1m753k58GvFLLJwdUB2tYJO8wj9E
46xEe8K0NzIg4gjNULLDnLOu3mrNWoaemtu62SBaK+oLECtim5Sg7VN0zYfWZoBl
lMCZeGOHXEF/FZSb1aE5liS71Cn0FDpye6ml+vXWCPmqmSxhmuJUekGZn48SP0JA
Nk9B4o+pvaZ+/SkkvEQIdj2pzVk6HAYK0WM4EhsOhDIo+2QjumgD8TAK/Qv0KY6b
GIFEPXI9wtdrMnojoAl9J5JjtHxopevPYx1Bgkd9XKspIksA2A+nrY68pLeJ/dHz
PZJKpr95cIibR9iQLQEtHHLoxhxgsLtIgDbApG5OkDEJqABt2XegrDkn1/S2qnmz
i7X2vHst6PPS7aKf7zutGY2QG9TocC0n6nlr/WKbmsDzb7CvpDsAtinSnLrjSosc
Ii8Grr4ZG1Gotucz45m8PdWbmTOSlvPSmHChH5deSKvpj3IRppJ6pXoeXTUST072
5rGZanFO9qCxzBFFtRQ//xnnEO/HZrbpzAu8Q69LobVOgMgNDq0ni8co/Cg0acEk
Y23ZGdlwz3T9AjKrFSTyQc2atvB09+VCYt6y2C0ZspUAp5zQsqYwvw+X2UlTa+X5
kK3lIHIig44l3415wlWJNHXJmkT7DXumdr8td2Daszh3NkHTe9+UmwtN674PzxXA
T6jWudgRyz6urrVU3lzKS06wSYvA8XQoH3daEo/lbbsz9O/QzaR/xOrxolJiOZ3C
XQxrLmKkj/M69pHlbOC97En4J/uBFdCRB8AkYlHMWQk=
`pragma protect end_protected
