// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:36 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YUodXIKI3rd9UgYJQP15hlodoWp7CVpxqkB1hJDpOI4h/PZXk4NYOBmhScBD4FGZ
MVx0Dc9Dzup6J8Q54gOZL4DADhPuCkoDUK7++HFQgxvItB9/ApHd9jBAQR1nCHeO
iH2fH50cGsflDFte49n8Ld+oK55TD8zG8iIC/m3XagY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11472)
Trm/+eCaKLRZVTEtINgJbj8TFa+/GtFzLiL8rjswSWzrg58FLeHJkfRTzgvSsLYP
atWxxLQRwZu577NXGi9AqyOl+3Rv3q4Y9/Q1b+dyKKuJyCuwpoM2bnpvv1NTxpFN
GfKyyigLN0W1OsO8uLhbPFOtLa71o+y7lsU6e4X690L0893ZQnywhCYb5O7YrwWB
TKXj1BqK6aX9Dl2ELteXMcvfVlV9UP90eaYb/EwNEz+HSblzhNofmfGCNCFeeSC/
ZnF7yDMUZIdXUTdBr07/lBPnQfFmK5CBw4UW9chcmlNkNUHQRr5hD3zVliQMLXtp
Ev0Y/yy/j2jeEYp/bzrkuhC66XGFuP7eeNa4zdI5oUF767f2J4Ga3gE2JYPULWZg
6ljuLxrzq5HanwUYNFcHteLfCBT2XrydYkOLjsYy1XaqqFMrmER2Lop9Odold4FB
w1M1AbiCwo+oe2xyAW3311wXzl8IabmiQVYfOo1wVRZgTnXZko6sugss0w7jHmr1
LuHB46TL8n0h8MAebLTvsVlpgQWQ6TYW8mKTq1b3r+Pr1xJI9E1jXmUVouqr6m9M
N+72lCCGYxsIHmyps9EbC1NI0L/mq7eQRpdX2zXbMn5CXC4L6dL5PE2DRqPHLzFv
6zRqce3adlB4xLfrkOU5Ypnj9LiwCB9yXpSU7ecAltW51pCZsF1IN1GFkpRQRuu9
NyOqoelV1sRAm3Q9xywXijWeqp9vY66LvrHmrSSBeS6msjaju+BbWbtwJt3nDIEj
5n5wST4V2nnaM3w+/P+dzQFfTz/puRxYj36lDOUWlb4LC+OiLG3gXFrUEjZy2yA6
S42+ldEkdYiZCvAsa8hl4ZxlCKmS1LvzX5ttTUZCuq7jTHP+ELFNQkHIIn5YUtJU
8tq15KuWgarMNQ2uyfFbMyUQIj8yVXQmZwNWZyt4erkg4OvZk95H9gLy8ZNVeq5v
7exyguDdZj5JBNAnj+stZBK/+jSSv7LzTG5LnKH971GoqtLcn8OdEcWMa4hN+0DO
4YSJzJtpsmPh72zHW923btX7f2Ozm7OTcRqzjnvRRcen42XKGoRGgmDislgmboD/
MNmwbKgWuZ+ErWbRqQbyjG8ptlj+7XSfrR3XagAW69EDtaosxbRHBEuhNY8X9m82
AREl9kxtKvHmcEktQA0wfDEWdI/KNkEgTYLQx67A4GPUiE26KSTXkm/m/0oyLTqd
Y/IpgXU7vedbGSqwTBcJQbmvgh4+isvOBRSyRXn21EqCIldeI3RXsnP9X8wMssTH
pdsKTjhwZdF8px6C6IlZesZQRkc8oG/GBbIM95CrZPV+qmkQwl7oPlf20zLxFiAF
6A/TxIjBd8LKGciq0h0VQtlJTeoxmhQwsxsZlsbt1tTZ+qwFmIoK0sc/27sM4UEt
GCtd/pxBSh8/tfn0XhhTH06ia2+gAt2lvFa1SXtirqpggCYZ+bh4bSItZdFVpaa3
sL1riMRSjqd6yVDB0oPUTrmyrurKbGmkFAHoj5FaXbEzxjj/70GHmtjvA5YowuvR
IegJUYOwNO4G3Tbkby5k9BWtg4brDS97GfxCY/T1HkSzbHke+jMFIAict4Wbu3Zm
Y94jazKpuhmT/fSzD3PHGQtFSS7OBnfsfRhqU831CpQWMFCYAJmoPfdx44NbQ/WF
9BdV81ZPsNVIsXZlt7qKs/Oiyz6+JFXiVY8CA333ANBYNOCW/6osO/oAw+2RiKNg
vUzo5czFKbx1I0C2DgdQ50gkYwKPhns7frSQHyEFKORUHRRS4rOzq4LvBJNVxjBi
gZcvr5xJPUYgLib1fk43PJcCibB6Y2h75CAjNRsKFJ4xPzngvXlp+cqWh86dPXKQ
phYf7Fl+V9993SkwEmKbC/tn3znvSJlVCts6gLdRjg7JR9786RqxSUcDzZYot+tE
KEQ32HbT8eDGCBCXnTZ9IbFQhjHA8eXjM6ZPd5VM2i8bnsPrWW3lsV9rM1O/0cEe
4ikQ+vIvSkEykUjSG4vtrwpEXzD9E64bEP0rzSX31RWATh+kZkgaXDSoPKFocdyE
DqEmY7bhrVA0bDiLhrmwGeNp7XQAqu2AeEQHRfYBfYfsfNKeaDKvs1CSPnGPVSQn
eebN2N2t/NIVpsiOXeEiikgSv7rJyp99v7fICoDuWVzUnTUXlI4YY4ATEjVJwHI7
wOgo9+saVgm8WEAbGVPLuTsahnRk5CuAbMIJ/8McYW8u3C5Eal56Yhf6Sl76UT0A
gfjYV+7VyiKJ5aMAnofNpXzEUe/vPDINDFlLS1lQdUE1OaY6pOqdkpi56BHBAI6Q
GMCHMKBuUQa8+yb2e8WA5w3o593h379Z/LHrAOhVeuWfV0lviLbFRubuNWeRGqTu
N7i8OLEzK21pnEb+eNE/q50hW731JjNidsnPezlMBnACFH2Ap+TbTrrRGrmGiUF+
W4AyvXkZTg3wM0zFmAzI5nYF1ZQBQNrdhgSD9f1s4EALWMa0sNIB7cNHviVRHdrd
fzICTNmcsJh6NH+xOVHTtELB29rZjLzyxtHkk8k9XsrcsQzN2wD45sWsENeT9rpa
ORR6KVgIYkBCq80fZvJ8B9oS7wS9wDNKYD1z1j2sq4JKGN6aELA74opum4sqRXz/
QgD0kZdZZTXZIGzcBlli7VPI0OrGmmiW0x5JnxtGWrpthqLASTfR3AjZV0biSdJt
I6pVJ/l4FuUe+iUa6Le/oeAIsvOpR7gACCC0YVmOqhdWRFIpaNcQIHhQIiDV7LpH
EI33nZ0wgN+ViU8j34l+kaJmSsuR6PTv9qndfyn6tflUvjeWit1mB5MQ7DtMs1hH
F4SCQ9F+9B+mpdw4ghgJA6V3zHo2EzxA5lcGGIBnAhOs5XJ/d7dAsoBgnIPOkCg3
7S2kk25tcr6r9QtSnkvQAS+i47O/GytcAGzg8GrswwuQaoUvEVoayRwHTPmeosWr
IrK2VKjJEiT0Pg3qM3EqcVWdDmQgaycHQjQsphtVfQlhsA0XOKEuUIVVi5JMhME2
V2Ys4Zs4nUIWp6vLVJi1g4eYJb3Ou0eKXntIQrYudnxOTtqnfDbRpoYSkPRQ5drn
+FfdcGEoxAQ3TY0Y4ugOKfYOInY7oJzZB9nXWGHRxQvMM5roKx67C8BGolit+3N9
rlXg43EF2yVZnvIlgEXpczC3nZFZBk8IGn7qj/9vyfSYkPhjaBqnfIPw7XN2eNnO
dy9aAyvEi+7KlpUeahWHEhvlt0esFh7gW6Nx5BNaoJAmLQlLp3n2LnemkIdU0wYF
pmAUE04FkmCpJN0XzQ0XoA95HAgJCqMS7+zdwkQN0GYQaMooNapBnJeb+incdz42
LGLwlbPCcPkprqa5+jEtagfUTe/pNAYzHZ7x7NbSAUNC6ewmUccfJh3D1HrxS8Oj
xNHhZ6dwylmBC1houCnuFXxv8c9u8YpgkcXjIo094U0JOkdGsj0MzFi91pnOgHs0
45VTB3ANPiEdmVDL7/V0MJhQTBklPMsueM7eblmZzXLt9c1J2horYdPYuqtjtIyE
t9NqKPGcpjbGSITtj37qXWMu6zHMrseLwLLczebgIoilUhvJSf+NLXhJ4MEwrr4B
H9XNyA/VmsKuJVJaoqkFSLn07eOfD/2W/ucsTpv2zujr5V2CoaWzMfPvQz1JQRhJ
1R4nW4Os3rjTUaXdX1+puqUtD6tVT/BFbyjc2sP5Aut58F5URO49j04yVD21Rumt
wM84x7uP3r3XBQ/cKSFclqp2iyt+kosQ170CsAkXO5SEJoMNEzIP4RhSl7zgDV+k
CKDRfIBtQHbzHFuOVZMPZe+3H2MsZncL5VoedkzhvBdIGKnyCz/fwWSdyAA9gwwc
a1As9Xdsd5FaaSjLKL2Y+IUV1dn3XphzGQZ0IGKcYEDQuncMxEDSviU285Qkf0kS
nOM8wEboAtLd46PHEbtSZMUM79/f2E463yoZ4DrqLVE38z5vjdpOOpDZkjtl8vwz
4bUB5O1Ii7UM7so6R0kvBlymQ/UTaTRfMvhmhqogVTruQAHjwddMQ9hrLCetEyGl
iEeixxMMxTAE/+pcesY4RJ500PRwrHuHLT1jZMvXA6Y9Z2+yC+nczqfd8tbOHiZF
xaq3uZzDLoEi6T/POl94CDbkdLVrv3QerURtIZtiuKp/nKgTJIUFHpkTKFYOwcll
7mU+Ze+3MrNHyZg2SWdhTI9fuCklmLw/WR7vrh1Qyz+iEkLtA6OYImEmid6hYmnN
ZbOgFbpl72IkhGCiHHbsXPaBKn4vDvCBxehd/uejf9hLJEwceRFshEoX0fr/cayX
YZHat5w5Ey7EE50/H/S7jRn2d3OuhjBWU603cSyuYDz5CGhLR2J3hGYMVUCh0heP
laNJZLF1QKIH5cqDeV3RKdaIotmhel8CWivKgnXz5gNZBSopvP6c+QSfEq0VvXcd
SsdgoAPGwBbgyBPxRlZRPpcHBQTNCXycCng7gGqaHopMLeiPPT4cqZ6EY2tuMht1
I5USzg3wdjAL6KElPi0La+rm39gvy/K+MoVzPjoROg1GUwxEl8wnIsbDsHKK01RO
KlF1mCD177QfgRa/Y0mpDHBwrlMxxaXZd3Pse8/63ry06gKDQyztYpRTpfPa3+y2
GCrwsLm9rQ2c1y4w82zYuW3mpGRJCulo8FYIXjGayGrkA7XL8u+fJMDV4yJSvd1I
wo9ZbuwVRnT1quc1UR4/CikbQd5jT8R+VKJSg4qHE+N/mU85oVQ+NovPpsq8Tdu2
vEWm25yKxpREyigfdZBlL+5fUcpQeQn0FOR+yymvSyLjuTUmIfP00djyYm3DodQl
6kDc54EecYN3eaivdubyGY00KYum9UBiNU5LoHpO5ytrHIvpN9mp1L0/x71URKS9
4Fi4H0JnDuhw3hk8OkreSHkQp62aijTFPLpFPGSl6J7Ketxq5K+Nnql95tPl3bxY
W4bq2QscOaetljjClYE4Dz12txChtMQvM328YL1tUsVW10+yAHBGi1+b02R3IbC5
V0O11RnJwuDx4FF8awtwC/AmYAE+qrRSNe4BYIMPSjN+lcxO9NjevMMPLmga4+zC
fqE+ix30uxpr/cqZ0bgi9xhJiCWE1J52kQ+DZz1GIx+icajRALD+tlznjuE2zzW6
EgnA5jAmoFzbro/pU6yrOccdvj8PSwLzsUpbSgMGKgWRxNcNj829ds9IfKEzdrR6
edRxw6EgS3f5Z4W6AqTTesFinoiqKaI+f6DHrftp4f1dHgEmYk6G4Ah0nSAtS9MP
RdVWldLfA34BwbZqihJDpxK5QrKlv8v8NY2CuT8xfuFtXT8S+9GtRKvKkb+tJKlz
cOsbuk2ofoKISqrjGZfMK8fvCJQ7LicIv1J4KTJFM3OJZRCSKTcWLHGnWHNlBpoA
5AKfUNdCUPRSnnpdjZOzU0UDuRP32/HG7O44vengZYT8l61FrjoPe6CscSgpOser
OwdRrGLXIpRkC37yv0lF02e2OZ0GNFp1WoZHdbTK2cQB5hQI5X9KNDPX08bXgiPW
L4HCYMzS+Ukl3kykz1dynG+ar97sw2rdJ7ofvKpf6MFAicq/2HSJukqHrfzu7kxx
uHwO4uptqszqKv4bx4ckArxObbv5/NyEzwmU1CM9a1seyhUMeQnq+DgcLvfIf2fT
Yn9+LidYJ2DM5kVdvWDOZZ7Tr/2+xROEev3+188cOsA9iav9ovHN1vYLz0WqR5VT
Tn7FlJMBGn2S+10zBq5h+zJ8eRbLkMjIKShNKhoNC1QAWN4ZF9nktD4ewCd3rRz7
o3N6Y5d3ZuC3q19Hlu0EA+axJtzxEqjnuYRW7gBZVWeZC85vkZgH/I9IkFteLxg+
Lk52ZK6r1DGEJbUmqIDJ6AigrQ+yP4qnGZinqOgGWQVWaz+C30ZoGmm9eXDuEAbh
Cxx+O7+dww/WXCoczCtRQyrii0TgKOUVjBhtqWI3WqhaXGhc9QLcQG9dKiVv+tnL
M0NzerKJfXdOfAhrdkcHwAFoQczupFhs7kTrW0G3Wt/zaBd8HVc9GvuDK4yd6Ekp
4w2w9PhvIJi/QU/h4WoO7I2jZYzhirA6GeiOcmUoz3Ae8/lpXU5hDZR2fAUn17Qh
3JuhbGHj3M37KrwEvYM9KSI17xmhV2vrKYuh2DA5C/hyhUIzOZJiSSY4My4espRD
misEBvgwewn00Twbe9P/1fnBfrrzzvnp40AicXdJuGHkXs++m5CaDGlRaZU6+jRj
b7NpjnHRJHjlcVo5ZRhzNk8spP0L4Kam0MR5yvCPx6e97JFX26RwUDcx8lspUg6Q
It3qAPOL3iJKJ41k141IvLZXLoiPUNkqldtThysA3j0P/xX+avj3LbOtGqX2aWR6
mpi3706Apdoy4pxOYAfWHsNAtlQ80ek/chXDRSlqJjThLfoBrPEnKdanfYgFMw2G
37xur4s14JqleVwZnIC+mcqFMOUIO256X6Dztyf1FAvw6O8aFuuMZU/b3Z+mwTxz
Lhbgq7/K+Aih2eavdQAAWBsOKvokeJl99Rd9xF599Ld8IyTOy93gFophW3WPa/Td
7dfcahAd+OCLZMJzbtFXS2vyzN/M+Z/ntVgX0jilGR/ANpwkgHn+LRPNNqAzmI/S
D74c2E3vyMyCHfOcSI4sLzToXUjGkY5HgrUADW+zy4s2AvKWEcSOOvWD4j95YyLQ
wE+nWw59V/lKDN/P/Pi3TApiShbszKV21Tji+QYcChbQORGW5p2VLViOdCHPlnVw
VVJmve/kjrCFnidMQWY/UtRiHGZ07KAE/cUzvwoPTRCQGRixHKvsf24eDiWry7GU
f/gs5vGEIAboaOiWpplXnwedRxanSsC49N1NQ6f9RiAFBPoUYZKapd2yfyzSWk5N
C3W2d4Yc5oAEgdih7YSRnBGG8mGmfAQ9NvLZsCCAtywhMcQk/A+uu8ClTAmGy4Ja
vVM/ihGeE3MTbXp5yRrB+VIjUX06ECTvjuo/wqeLq+fkj+LsG55yc1V5Ls4+DCae
WBWyB7pNeP1IrDmnMUiRAMMgGfSMiTESsJjqGVYGrWCxzUJbp7mmcTIg3aSq3KZG
DyOhG1llBkSgVLoaH6VFNxJzom4/mcx/k1tIiCZExlSsavS1wsrMYyHUtCPZ+4dW
MyBU8giaYWERkc0XYw0Fhb96vTmpGGnhkBIHycLLkVhzlKklk2Nsd4X9W0nomIKh
reFn/fF2TS4vi/RCCg10NPg1jps3TMhLhXmPFRVhA/KW4bcJhVJWzJLlsgI13RFv
bza3CPRvSKmtpoev2cmrtis4LgSerAAjGP1JRPB+Ltv/Ht3dpvpe4sffDnTOiZdj
NZXgYUY93gg/aAy+IGZTN4JwQ7ghurjN0umN5OoyLbsnJT3vstErtzN2zxg32tB4
o63eOcWrEEnfWVPLqRAkj3ac1LQqQYAoBXEDjc3ScubMjZwKIVXQdOAcFfbMATrv
UZ5FhPSrycfJbB8JW05AsbS3JPfolnuIOmDgl1Nd3uNGWLi9/iWAFfJxC4HxkLhm
8krwMp6QFVcFzRPjqZnNfMz7oZ05d+dwDbEiT/EGb1DDqD5AdmdApiiPKhvlrgJs
+pCkIVY1TMHEhepXIQuRxQaYEkb3gUxb6MAU+eLL0n73ntRsK/PHNtlTecCgMarG
VQLW6I/4DLdrhmArL+58wPQilCz+ks0GmhDkgWv9hIuNCr0jjNDKwoLlK/9y9bfQ
JAmsJ3pS6Xivf1dT7kRodzhHH9ORiNAAFIhZ0g4WbvadmTRBQ/lVWEboCl2hDdDm
SWNqlmHopRDvOL551Tavu393WnR0QLGiz0FIyt5fjhyeU/caK7Q+7eUTqwp6BAh8
qwAbZtIneqgPS/7dYI7bYFAZxMyGmn6+xSTc9L1H5GWvWoMlwdbcr55Iquy2yank
HGmSZBUmJe3KNUuT8ptaji45DJ0m3Qq1aLaXkUV55U298te0D3pT8sS8IbYyE2bs
85qcf/c/TFt80+0QTc/jOvccJwD6tUglWb7GecEE+o2vlLFrQasOGNQruuhByFvY
sJJL1aXvGZaohSS1//nmTxv+37c9ReblOaq71/pRVJ7ChrCcHyBL44NjcbcYQQc0
QZmSTDoI0OKgba/kVFY8b2VM+q7SMCknlkLR0VUd+Pb2VnVrOgnT4NR970b0fhOv
oTf4rImonpxoiopntpGVhH1iHvI9EtD9EFb4yHTjR0uh1HTt+PRplBl7HdYu2Ed7
MnXo0RTATd/dfSwnBh1Wot4wO0PtlUqBsRr7INgciUPirX10TCIqtpffzMabtOiw
RIYJPUIdbGFCo3CgSGglZJKkuLbh618iERslMJBA0Qj90OLWE7LCnHfBKSSc2Uwe
c6pgSs0Gej1EtTg6HrGhhqlEGwczVqMk6q0l7jNIbfAUT5/QtKkoMwQPa48DXsm6
i0Wsf1XhnWCAr/MLLhCK4VzPlEKSKGmdTyVOnWu3R7yMHz3vppAhI7SLCfoC2TqD
XkuPtztDaclXngssMidgLJI49tgRhLT3ZwUpGdux2DhuhY8SI0sOGcdP31CfiApL
+AjbxJSJb9LUIv3/01ChBfZ60LrTYEd+qjmyoRdDCtKYUfDuh1S0KaffdTjaqrxL
WJ2khguG0p2R0F+KRUpMhAz6/NxLMNr20uyb6y1ccJUEUc6Oe1hGcb9ed1clou1I
rz4uH16l8wedF39HdYNvTBFFi1ekE5y/OfEnOCguCgcxHgF+YvDlxW0RWNWIg6k9
EpD1B6bBpf1ud1u9sa2VxfoNg6o/ISGg6yXFVH+letGopa/OsKLsjfmERcve8WhQ
GhGdZ9plofJWaQPeS0BpFk4WZ2+ji4XLvYPkke3gP/00KxJumy2xPDd7eqvGz8OU
mIH+R+1da+9xq0RiPbfD5/03rUkazXq98WQV7t/Kwfvs25AJFdYpDEE3LXp7QvLk
dtSh7LNlEpZAlPBDzkmXmWNTkRLaIBFlmOf55VwhVRFy6UYiKCvtvKgeeXEpWZiA
dJHaR9rHVB1xrnvjZUtpHW84bWYQKKaP7bWK7saWWnwIamfq5Zxa9e7diUgXFK9x
zAyQpxAaZYcYBcd/kHhtwomXYRIUEC2/pevCvYX/Ad0esZjYVWFWcpXd6poGJRm/
SnhNOSiY+LAxV1grO+jGjQJSfcJJeAf8HRxDQZG8D5MeXEvHzvY+3IhpoWawdq/U
KhzwEyP9+cOyCmBeDVNfgwlLr/aPY9J4CiMPZ4eWHE1+iN15I5cKzk++GdS5B7kl
kinMAeqM1BcIz2zTBOLocjHwzr2HIBPpVmgVGAeWzKNiTwVPSjhV1+5CSJ5drBZg
F2/Rh30VUNqEQaxEKQrAwrsYwd6xuGdTwWUGHjTHJGO7no16NCjWizbbprQ6zTdS
D8AMuAoVZtfsDYeue2qVAkt8gTmHvGykOjeZDTEd3DixWMONzKXRtCQ9DpeLoazI
8OOby1I1IXx3+ajqgPRppyNqGquR1gEypQXk43COD8yPukVi0FOTwWW/xJZeVxMu
hIxS3DgtzpDsTPsx8UPgjrrRF+9t72ZzN0gVnOAlF0QSvGMqwU8FrGdFNcSof4Q2
+DZz8uO6pYSJEc4IQ2/gmJuMezYT2eYHvMgVmmr8tn0oULLkQ/lQO7L741cVAxgO
CB2fQQr1scPZGX1NApBuIjCGhsinueSZEbi1R7I2rGDkDIx0mD5bvoPbTn/vZvHk
E2ZBEr86bZKLS0UynIlblDbuk6oxyqzG95zQIYpAqvFb78dcl2l2Zvya1svbGtTF
0/ZJoj/EGQJkWc7rY04C+a/0QcKsIomt4LDJds8MbnmAlS79TExj++vBydwTG6Pq
uMxoiAzJa05y+oPA8ZTs111NtzVvlMEjHuio92U45qCo0sinsYKsf40qI9dYdn/F
gVLDojiVK37e2jFNvLOk0XQwJXvVTbmvC3N2pLSN9IzkcX0t1v0Gw2L4ml6NXLvM
WTQSUFF8Sv9P2qNotbR89Kk/vukPlnsz5jTUwle1KXmAtR7rq7X0BKN1t6V6mZ6p
hIiIdQF2JPGoZI/3EJSMPp6v7wKB4xGjaCL0/yRo5fhvqvNI8U2icJP8H8SOK+4g
2mi3PikZoF6RdUBQRX/i7+RwTXgF+3ACE2Mp507lb858xXcdX41NRrdNDd66/jTr
WS2d9yhsYabCafifue2zXcPeMT5ZiwVi68pNH8gJ/X9u0s6AhpTdmWYGYKvlz6RI
G+yKiOauVR3HrPTZAWtga7GPnfprlTpd44Q8p/ixbyfXSPiZV2Lo0pNF6HMGGqBA
GSIlHaLesBrWJjIQts8tlBlKwbdyUfdkSEN5/zWnrKGa79/tLwllSqSRTkXelrA+
HzN4TZlALulBqDT4vN/jgkYcCet5RIe1BITLK9i4OR2eNCvbF1vKoe4iv8FhSUYO
V4Dvu79mBDPbw0hS6n/LmjgzRHyOnW7cVQRVefVEoocbGvhrkUtK169ns5yxzt90
Dslwy6ISJOLwWHrAJMI46Z3lXrwiwAhjCAa6WKkP2d6MTQzvIPM+minJuUr8Uucy
2a28XH1NqAmTkwU2wJgabXsKEJfSP5/cGU/Pdnos+sDyHGzepAmJ58RnCXG7FS2B
1rSGWXdVHuMFLnRheuDzn8KcAfqU81NUnbL2OE+AF2yWKz441I5Ca4+Te/wjznB9
sJdvNfFoHg12OVuT1Zi9/uANrX+XnF05VxkC978XBJ0uX8Lfz4rZnqxaOw3mhqtB
2CKWM2Q1iocvQIqeOzuhG4jCrQxenINkSDEdKrm6aELOZFMjjoTE9bQaP3cUPcvc
xe9jaLCz+2dx6Ejnl3iPXs5cLFEhIvjNwUkONHn0nX/dnx67sRjmditooWa+OONZ
Hi8aGhBuUvxR8K9FY/wGjS+ObP++g0I/8WXzSVsJjonqRGOc9RLW+1OUFshXkde/
G0KfKGjvk9mRXNMjhepdPCfNJIhdEYqx1rQCWfhc51n+So87o2h1Gf7fmNoUfU40
bHkk3FKSUlz4UpyROKf0CZXcWWHw7h4tP0SkdJAzF8LavQN3AAv/VgTCnabAsXK5
mdbssCRY5m+7e6521Jx8ZEH9kyEYukbgXnJ5/qrKG2RXiyWvc8hwKBzMSG6K67V2
ZCo/eTrvS3oWFtXMsiuSMfxc4WhjKyfeDUr2aq+NhXxDseXNqae0FbyKxEmF9WVp
If1W1+lP/9a30OaNovt+4MWskZV9CSoeB9LmwV6ogCfOeSNQumFJRbvVKJpx7MQL
C6oFrleTcIlcwT0OmunHn2au+5pInYH2l7w8oV9CzknK6XxKcG8+e/jHTamkvf/2
To7xUsEeX9DmtrJq+ogetd+UcIFsVHRSh8AUTM02e3C+Siueps+pff/0gFPcU1R3
0QM8vMPN/fXMMuFAVPBOvWL9mWHHPPF0YpzkQj4W1PuCeY9Rj5F+RXL0U7IqYm0f
kjiksN5vVBQyppNSpB7pF2mE3X4pqRoaJYeLKTe0JVR1aGIKq5dtJNBOxJrfRiUM
LsILFjEEcIwklCdO+DnsPY1OHsKT5X/8sfxBg0etEp8yk4C7gJbG5VOY2xSECNFM
doRyFBHuaQDTMtewIEnKgpge1gxuaduxsQLb9w+JafryoEkWl2Hck5U16/KL3vNf
x+kTGSJGRo+kl4eYmIYsI1kYPBAPLlOn5iiJ8IBL0WsAoQIOPhVVMBA/TiCbixlu
Po5JWYXhsEVAeuce2Kpf/QUtxFZHBHEHT0vBT/Mk1rPvkYo4p6RyS688Qa/8IRLf
UTZqEYoqQBu97aO3kCcWC5sC4vFSEjzbq3M26i56Vsryve8Az3cB/e/ZOFeW34m6
usYt8Kbga4le4huNhcXRppkZ2Gqq8+9re9Qjxv7sjGMn4o8mmnCgJRj//5PqFRs6
imXLAJ/L5r7hWrrC3RzweoheCPCredd75I3+6XR0x8d1tFkX9BtsY5fMLgPnzoRE
/WAJd3Wiln0hICZw757ZIjqpL63WHNPhZKcokrpK+DTutAaN0z5oMzkaQzWgj7G6
ekKYl4XBCe9Txjpl03Y8kpWrswZOKRmvvwSgh8vYnaUyPgZp+lqnUXKce4gArgWL
8UxWjoHM8yNjBNn5zTjZDGheKWqxv8mvYjQ2ejnnKqSiHKQ2R4TW5/XbgHm7yoPt
828GoeU6ONVO6rdAq5a5M9moKjCkirmfcQbr0CcOSiKGx+8XCj5VxM4l/+Rm0XSw
tgqCN6WxIdy485FghWnnIzl60emuqol/gNptNS1kPCh7KMDZWCXpvxSoas0mzHPI
SHsohDLiPjQEkI82RJjH/Q7zJpqRw8c+eNXZRbFff2vJWEzCJyflOvtlSAiIUrZ3
wMK2r4/wibHh6Zd4rqHfvskmAJcXUMUmGQ3lXzof9XKXA3yraiVxWDuYZRowcnj1
5yYtbLaWJ/qJJuinaTrZItQDfQLslf+9v6UbSaZtu9Dio0770XM2zBieLp324uVg
56JBJX7OHsU0KCfUEfh693WX1x4IoWcJEZ7pzcoAxiNu75kS0cnq2Pn1cxrDyc+Q
wj8lexC+d2Ts9eMwGRQtYGKr7Mikyofozg/sRlCv7poELjvuqbDaseqpyiMcQhYO
yyDj8yxVtIMohRrfbOqmcHFF16LTDmMwnbLElIX01r8xjPc3twO8lBOVb/dyRh1H
Jdo3YZi3oqMWeItlnhViWuUu+sRLXeIRZhgrq/npnaLx/JGVF6ViFm1EQ6Ffc2G4
jP31YfZzAFvCkU4kZSAo2vCBO5y65p6waHGcA38fEV8BgdOHG1XvXXqLHqTdNP3M
tgKAPCic6DsliLusKh+Y940xZJtnSJBgrXKWgBupDZ6TUBj79hS0RTYgKWWfBmEO
sMLgtKbk9YdBJsTi0iNUBHo7fPEOv6zszpIhP4hefE4PkBolOW/ksqEeucb2f5wi
bkCvcvh+D3jNEQjNHexpyCOa1jboP8PaB2EMJAwPbbmSCszKep54SnqMqS1N7Kdi
1uYcGbzFE/O3zDN6rqn3fwW4uwuuhf1n/BxwE5ErV8q4bA2EsM+IhOTxniNRHoQm
/uQfOXYQuM02bmjR1KgstXZDkS/F4dy42XWq32CuPRTHxtnD92USdZXhd0+fj+ZN
Wcdr8JYXLto2ZZgXY56eXCo0wCgHhIMmNCJG0PEStGKoev+UJltc+BFWECjRERad
4b66t4vEQ7sOhCGe0Wh7EseONofZkiDfHjuZ+q2atGSXfhLi0KuufCLtmGEeahzh
ylRKGp2Gq5M+tUt1LV8ISFm1NjnhmQFUhFrgt8cPDtj6YJ9HAGITfOBAWmiYUxX9
WJ/LiJy6mee1KtGNMXRBdDxHXi5fs+RU+XTNTU5nSojJyBj1PphZXHcbdTyqSTBb
KSazGRpnDDlhT1bLCfZQt7ojPWKOrV/eLh5oz1eEbYjw+W9teAq8ULehf86utYtH
VgQgjMn+Jr0mW2Xq1k5TlZEo1cIKb2F0Atw0cMCb2E5D1o0Y4YlezdU1F9TGU/pf
Rh2zWvlHjsEmABUWo9Rcgqp233FWQAoH1F4bj7YhhgtlsR//um5JCQsm5uLFEYN0
yE/aUm6O3s1yiCpreSKqJ0imGpllGHhZzX8wknrGqFf6pjAPqYfLE/OcSk2/c2ur
cFQ5kDva4tgAOf3Uqh7mtMQcyLWY6Or9daY/xkzvwBJl1lvomiUoHqXYVjCv4Bts
cQBJ++bPdmiD7Z5Rwh8ToRQCMi7lKRe255QsFa7zXbPLFgM92phtojE0ux2iKaMA
/v9Xdi6vgwxE9MetPNACJPzQ5frLYc94hvftZNm+sQhEQ5QkeeTHjDdZ7mcb5mP7
cw//MgE069kB60k23XOKOQmlbgIijTKSoLGnpAD5MOUTj4uyw8uNv+tMq/DaevSk
bEVEeRm1hKeQOpctoGG5oESRQgLxoBpHJ5AUGnqcl0CiByFRWbJza0bPZn8AOYN3
KsgHFLw55WsvtPdi47oyW4so7Aym24rOZW2sy5LHA7T4Zxy18CllZdaxOWavG/bc
jdrwgtFClyQulUAEwla37z7FidIEwMlW1QROuXLXj1IWhDEHjjOie3uK5rpUIIm3
ovTwVcb6cuirdN76/+tG5kdUNYhkKBgYynpTkdeunrfIMvTqgQVR8xRaUNiYN193
n+jcesnWSkixoSpCb9CG8jltNHVUgd3cmCZrrXVZJJntwVe+3OR+7mxbQfT92NOD
nnct3/X2pThFuW4ulVcEOc85n+pVozKk324oKWLdv0hJy6DpfLLnpmy80ZQu0mbo
lt7q6YatZ8UAHrIjNrQYQGjvahp0msVWCBQ7gRDHertR7ZJb9w8Qsc0QLaEO+Xln
hrx255SSiHl0F9I6kopd5ZGZbYXVjL/PqJikZ1DEgNOQFaU04oL7UDkxBv/Y7UcC
k1Kru5FoBlEYkZzTyS76xRQ74uh6lOij5ceEXRkYbzD3+urYBTehep8eKRlR4B19
eS4YoG/Qth0Y93Q8ocpb/G69aJ2G75eAc8hEhw3REmYFaiiQD5tmIG0Uh9OP2E0o
OpUGXVfGmvYewYxqr8flZh36gpvEl+iKTZh2r+sb9mpBsxYM0RAMqFx2xvCRYFF3
RAIRBiS2eR8FAFIIqW7WpTKJHFT+PjmgisvrCLgOqplWguP9pbXiKWEFFQik80nq
krTnnzwHGZSvulfv4nF0dlY8uGRGQHqMAMQMHwoi6WlA+/zXgljCznX1ywr/B/h/
D8BaTU2DS1324byVwzfR9ck4vETG6ATar7HVnowAleDGTO1/TKLaNvpSksyElXCn
fvimYy6vpsNX+Tpj6bMWbTwUup/BAbu6o6E6pcxGe/jRZyxRE/byObSgW4nIv5br
eaZG0pOUomSqgixXeBrNxkEKDTz3O5BNUQ02SbV2zUFRqnTIltPFTgMsiwFsMnS0
uu/hi/4UOL2ZeBbBf72/M0BJlk+6RtEIy8qpHXKLc8bVXHwAJz1Evzr+7i2auQSF
FGk1TAlKM5Eehjth2MZ5hNlGq6vNPeWQU3kflhNYaV4tstPXIzTKDY9/5+4h7tj7
VGs26SoUrDzmvHNYjrnnonjCMjIaD+ekusmG+wh0GcG7bQZsA29PnfNcYfaOredd
Row6kaLZS+gq8blzzv7346/CUbV8d4iu0CUldu6VHPmxW1ZhLBZO6Jt22jSGhQoK
HR23aheHtmRmOFHZ44kVmS+wJNi6BMXaUSnCy6nfml5DeWIdP/gcZ4XgyIK4PnnE
yS2u7Yfcb7HGzuIxdQNCwdo5Pmu63kU07dXZpPzq6IY0X9J+dVmYcVjW7tA7v4ZK
d+slieQSjHGZI9jQOx+RQf4gOQyP/yPzeP244myfvF5Uj76SShRleWL4gdhojgX1
`pragma protect end_protected
