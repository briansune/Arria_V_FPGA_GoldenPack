// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:28:06 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RTrJkVL+bhPAQPRzGIHWIzI8RV5yb35YA3rHJaxoqV1jPxaqJ2A3TBWjLOtkezJi
Y99346wmmeHr7GYkzmGcNcb7g1A+Qi+YpcfzC4Q1qXQt2idg/jlSYnonlGghEJr/
TNsSPHfcxRrX2BfGB4Pw01tbbsdFneWQJED4MACODkU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4416)
kmuDh+0LDHR8CMIdKzVSGQK+hM+0bVXsyEz6Sjl/swUT+D7eIcJocwmPQQO9OEu2
neqaOkGeDlkY7OIbZeYuLUKnSmvRvWziwtWE4CRQLORDL90yiz8101pENqrKSNpG
HqgBrx8vf2J5tT7fuFbPzVGyavxcfy0+1TkG7toVPd1mAeZ0brC+bqFezWQp9Uk/
706H4jLRadtghtDJVAzJnS1oxCkxtoaZ790QLXoDiIaLGsn+J4v2lrGgxB/3f2P4
6EWRdLf21OPmUMPOBN2h8g0+04MUig606Mf22Qc5NpEMXlyy5+v2vmyPSp6axE5T
uytcH+d7AHSDIP11EbChXTYZH9D5EVXRSnjb842sVzGM1E9Uuvb4XB+aBxSnLiWH
vjENFdIh5ip6CDrk3tN4EaXzCf2Pi1vDJ5t2nfcMyTzvCmm293xbLbpDBx0/C3+R
TlTDoiMAy/pE8CJ+bGagAq1L3Jiw0DvmBBQ40M5fSFiYN95oRI9q7+RBwt2ICQ2r
6rzKvYNDdnB7vU8gwmkRw8Ln6WnLQVQ8yT7cURW7eoEAbFAl8QU9o3NMPa3yEkpG
MGtAvwP2SzqLJiiSqnllvulOJYNBPUPfmBvZwNqOQPhsQpaJilYjGo9elgi3QUkt
QLbXmg79p8HTFmKVQTV5M5OsMEuSIPIsECoXd/k4OYIuRn9X/+kKYjW8wmaCYS4f
F/Cfi8FjSSUIC4u83wPrkI8x8bbzweHOoL3z0c3602j5KyOsKd/4YiSRkppbQOWx
DSUPzrq5eZj2O0R8ve1HxZXNbmGBTS7V7e1wm0gaWXLQ52L+5qSzQXH5H/K2iEbY
w7zbmMNBnKMO06ltFhOF3QWpkI50wWSYDFB7AZZ0hHjmLbun18luchG5fYZx/FKS
JGcQegX0Baa2Tea9Pj/JN/+piDSltS2BRukTlriDyXBmPndVyChMH+sm5n+5t2dp
rGEa/WTfu9sBupPzgGogzvVlc1ccLqR5K2N873wql+oNxd+KfsXANE6ee23LDHEw
SkeWLaDm6VvkhthHWM2OauZ5oT8BEADojxwaVzYVKH83UnRNQYqxkExJCdEA9p/8
MktN5pMnoV2LnxYpkI8h8B/E50+bXDG+HqMgEf3q2OgMWcd7k2EEgMXlQhblRR0Z
yw/9ya7sFmVavgN7a80n9LZo2u0rPKFzHbLDtdJS37CWvSFaRHYlERl8LuCZzWZ2
F7Ck5OXl+jFlSgEyx3V0XHu3xAaBFXvmId2Tnx0Oa6JoGtV8RHISiHjh0WCVU1XP
L0ZDjDqYYJsg7I4Gk8k2BltdVQ5D/eTaqf0vrKPGzUCM1zOjQgd8sYGAfhKfnawH
OB7AXeoGNBu7t0YArC7LI9Py+Dl9C///71P4C6NqSuN91BId2ki7uMbjQYShcVu1
rcspAGFXu1YqBvYYMHqG2rYdhlrV90t77NUIGaT/JW6DAlwwEnK/Z5RVL0j1/78K
79PAX3Xb9n1ujv4tgj7z2Bg/wVYDR8Sarka8bkIJ9EFEIwRkLEG2U+n2wvbw3qu5
iab+lZ0R6/T4tXgXsGheFdREzhWR+2UpInDW0gQxa0SUKnUaEXWn+wRGmOujAXFb
Cz9sNu9MMn/il5x2xqBfFom3ybg2QAYHoFHBrLKHPdnMNEPHWq1EXpuwOo+m8M8G
iQs+gODM6Est0Wo+dOEKj3SaWyRCbzbSCmQZKbWoAaG8NjibN3qNDJY9r80OG9rL
savKKYZd2dKMLnLT/b4aY7tuRuAlIr+hHov7efHCm9aSDGume5z6bRJ2UXagBM34
rufCyIQburpw4+TkcS8823CosWEx0PxKCLdLj1MQhGwASD/ll1c/ccitVk2FTjsD
smR2EuysfCEGcxGTAwS+inmbMb3UlFqyym4gG/M0SAGwjb1/dfV/SGHV5NC2Z1hG
ieQzwelYRrWUVN5UnXVJP9escBTWe/NvpC29HwhdrTAHuu9XDViT9n1yHRadWA0d
Y7EcUJvu2vT6IHkyWlC5wyQOio6470lsSHjoeAenHkpF6qvnMMCJNxqHvCQDMKEi
59pO/I/2pT2PHXu4sNkGB08HmNX6Xmrc8H8jSvevT1LLk8IRorX7Ep0yp4K38SoU
QJB2aD6CQhWMoruPNWsmwzzONhOCCwhdX9rrp7p4XKGhEwVksn/nF1M5ADJcqQ2d
e0tLZ+Ww5ERojmcSwhaMlogZTH6CG9mcBZYt2Qq6s4yRG8eDDWH1aCWfGQdGO373
oTG6PysoAqdbeX070je1wWaoGao3EbM1whJ+8VMXpBAyeXXxNtq1pJqqHKSkGAoc
WpchRIVOBMLwsglyPxhNRqRpw3p9OniqRqEJeBRXmcVPEm4aq4bwCav3V7ZRkPdr
BY6DPikie21q/n9lN2lenM62+FxWKyB6r7zIAnn3/xWgHKtctY0hVqTegmotrSCY
lTDYzFnMHLeG4QssgHI3wLaQF02BcA75kCI7iABfZwNh0WQdDd/j+u1FjZFhsdXR
PWCqFntkzXiYZBOENXfnU2bd5jK0Mk/g3lEijUoLuLrUqq41UtIzzD8LySkfG88+
HFunvBS0ZTFcj/d+bTjjyUJ4zfTdT87VqExFhR2IHz8q2LBmwbYe2EgB3XWdaBww
nqVCRvl+R7vVLtBtbH60IJMVlJ7RqMY6x2iUTmMxOxc4BS8FHD3pQWcGrzj0EwJQ
YJ+E92PYpMx4xClZLrdkdjsfHHcDI9NWB7lyzJebTModZMxNTektE875hWkQ3zW1
lkqAxdCZPNy5+1Ioo+Vy7aGKOiLdaAQ/hBfHI5UTJ4JTKjL0ymlMhV+fFlOHoiwh
O8U16E0nQdrT58Cgzi7XdNMsMj0G7jA1IdgBpSKrYyhPcpgYsp8rnrfjMA0omUGm
oDxRhlN+s5IdXoFU1Gue9M1F7oFlx4F4Keii+gTjB1U+KnKFRxdzMrHG9H/uHW5i
4LQuWeyeswMltHh17zbWxv6xWP6bEIKXYw7YjwY5cttg8fpy5RU0C+eoJWohzj98
yvCaWa2n1lhh6YXAa6p6CUrromN/S7feKZnlPeDsKgoNoTMXhj2lm9+qq0WmKoxX
3YAAVqvzDeoIL1hzJleK5qIh6LfD6PC7ZVZSCdBLIDng4uubsRuZJA5NVcMaNned
DSp/G1pi3ir+tGHhEW+z7Qz32K7kFuluGjdFpJJqMHIkYwxJgLSG/zW9y0TZHrNh
1+hyodP9hEINynPYwa/yqf6+BX7x4J51bkEadfYHQyVpGz8YYZiEA1aUkJ/anBLu
ckkEV5JVWvfJYWMuGCcs7fIJbjfQH/E3EvZOhE7CouimMJB2FkBkCDlqRt3selRD
O4LzmPftpb1FOE+p1E6Jf2rvbwsAv1NnL8vTL4z2/+E5tOlVkf2moJk/dY9Mc/Ck
90pHhLqCLCg3pgPzkA7NOT6kAiqdiImEJwpyGKsdq5hgfoNMZficE2ZdO8HhlvrO
INkDoFpCUbcqoaYtjudBkKqhzpMaxMYnbevHY4Khc3Zk45ic4jlCmrSrBFot2s87
zc6PH6cZPqqw8Ykcmb5n+fIzObUtAuM+3RwN35eCw/AlolHX6D05WgKOwzBv2r90
FTI/BxQToY0QX6/zSbvhZubuBUzKtNDBC8PrBry7SyfAvWTw4vWRKdyaUKjf1Wy7
Yg02sq0vf513nMBH+6d6xq5zBhbYImeIu+M0QQiOFEoroZ6og9Yya3r7RL+17Fhz
JJdPfxQ4VJjAOcGixvw+ZFPM1tnE/WN8uQpd8LN+wP+w25cyvqumwmSU74pEoq6t
FGwdlATnLHyTKlLXQCwAX3nRjphyMQ21BmRbJQK3Biq+H373WU1y5y6Fj74Njm+i
yoOJ60lbByVgZlULDPLaABAgmrNOXIux64YyYoKS/uR9gJUHXPLlDsfwpQY6NSV1
W8LJ01t0IOTYPhdfKnfr/U9abKXMgZ39howiQHgstnnjeheEeBKCspxh9L7n1tL9
d8N7BzygcxnSxZ9fffNmVHDWBRiiXR35ohPISNwXgesH7hPuGzwpZmkTY5TWnJhF
J3f1pzBh5VECi/fvdooXKRrjJle4PP4PI+14T1SwTdO4aD6K+vsARG3ex8ZMH14Q
wApvU/AdakUba7eHgUbqogysKNcbRBcrtgC2te5VjgkqGXGb6Q21/1MRZpHQ54yR
3F6ulcNZhVL5drfn5ZhJWR2H/fTS1ljdIAJSMm+septNN/PLAfshCcvQJDLDM6sk
avsJ4E/K592KVNqsaLuAUrgDMN1Tm6ID0AwmKLiYPtq4WAcIfCBTP3KJLztRxnhL
h/uXme46sPi6W1Wyzevg/0Jzr1i5MXHdU/C0ti371rEhpoE1GNHAYETFnLS7HqJ3
v+0AXqG6NVaaK1OS4SbdHvuLOS2Fjhq2F47ni8ZeEDO3AuVC/tjU84O3Kfc74Rfy
X1OB10XhoNaavFven98RV3Mqi8e2FMm6kSmQYg+I02x9QNTfMwym5BdvRvu+41aU
wMITkwgzPrgF0SvLA0xUcs0ZoafeghCb+XQ35C/JVcEpBW5r7kmcZq+z6ioFm/t6
lWtBZfXYx2Z0KgLQ/mogrOPfkRh01Mkq4g+UEjbeOJMGcavmFU6dkQn5ip8IU/Qy
SXN/3C9dCMyPh5TJN4/K+pYF8yA/Evbs/ogQHyw2LbifKELHWGnfQDCTKPRqbqV9
GjWUS5jcxWCXuxEUPkzXdLh7MzEL6ShDdJLyIIs5MryE+Sy4PNEtfLmWXNfeuo/V
gm9akhsh8f+SYg4i3ewfYLBb1RN5EX6KoJaMk4HVj5cBfksEpP62MVlerfGX85RL
PdUiSmMdmv420N1d9Ulm6je994Z3bH4GmTFSusmhpl7VisqNS6HKxT0sIH4e1xrr
QohMSQgHeYLztMkzTc9oomvbjn8eNXbxB7hM9IGvbRdQaEoB/NHw+lC2yP2CPhCr
ClHePC3J19irmmSDkO3/Bqw6k+unCUw0xjTADs32SWM0NVI+chyXpsHg5xObaO8w
IgqhglVFRRE3VjnBvyynMe6XVGRB8Ob3NrSUzfyeG08PLXlHbO5n63fu8g1FlCwv
n+/WKuZ6LynYyYxhkwlZgxqG0KKR3svBnuOPPudTjRi49ojK5ENzLZiyN0oZUbj5
TO4kA63Qg3PMfkUpKeGUh9lFbKfGhP61FB4dB26uKySIPz0+jlmuzMVN3M/WDJ0O
K1VL80d9R8BKMJrY8yz2sTCnquUzC0ndKbmrcFEYFj+C5mMqD2TW+5swsmnX/as6
UkTk9/G/++b+39AazBJqR8qMxSE/kZjt3jWRLVacvYM/7tOXnLua24nHOlPaqkfm
05TiOVscpKs0QcTTrGBq4m+9Ui3oekbDkavD03PL9xAVQvFQGAOjkmGP78IrkfB0
INsd4+7cEPtKnx9kcxa6cOAJOBQzI6aYukgqL6Fc8w4GsfxSmBZnzyjtE4mx5zWK
vUll/AoQeWJTBgkE9A6tDwmOdLreGnkuQVUexizJg1uxSf9fHTrYy5njTSKeCSPs
RsGTtB2wxLgmCA2Fnj4TincClKSGpBDJNEWzbIUCHo9hwlW7tXDAhXPdK33Ys+q+
lOVnRU6gnHyIO4qtxat26EjwtB63T3vIqqf9HYY5AIVSVX1csJ7fCbzzbSckiKcj
MQeyx2qdXixUjQFSj0S7bRONjqJhcH3ev9txwqRTBBpzudGsiq4NMmhHxYHWGeNI
9K5hVgp5Z1VoO0O6spAAY3wtXaUxMmGZRk5o8v7hMnA4ImlcLtMUNJZkk6rvFHVE
09TahEZx16i+dVtcHMHUzRVDDOBhOUIukH8VMRhcVX7ch0/cYhf+jhB0EPsaSRaQ
UkuVmHIpcERuh5Qm9CLr5EpCcUZF7gdx1PYODFzVXsuuXYtKCv9jozNRKeTVlVs0
`pragma protect end_protected
