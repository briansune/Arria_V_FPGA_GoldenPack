// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:28 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CYRHArzhkJ8TSnlfbwo1eE64rpZCI9KY7RbwYfKACJ7VNATaqb98WnH+4On9qlD0
ybmLFf0aA1m8JAj+Rh1yMDg3B3ECmjbc9JnGYmYn32XhqHVVb+g9R15jdZOm+PLQ
Amub0YuwVgBXZht3mDTiumq40annake8KpEjEVffbQ4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10256)
DAp4cyWBI0DoXja0J83cDwTS6tp7OhpxSyigqeKBCcxMADK0Gi7AdK4EKss7pFcY
CZy9f06bQgG2OknQEmJyr11fev5UOqvjdl8U/HmP1sQR/sNa+qfcf+Cx0k1Y/AKu
ATXvGYlX8EkeWNjBaNx/doQ/66Ri3HV2BqyAK21+cSWyCyUIlxkCeDFQZ+PIHzJh
1aqjLDpBoMt+6F59Nr61hC3OSqXBbEd/4WRiW5W88+WHchMBapiSgWvQZk91soo3
uTWuurnpAMB9aH6vLBdv5i+X9Ka66Xnl3YTWkbZ8fn5xM+uoeT2IZT+X4v2Y2TRx
/MOwTzaVp2hly10ocCVst17lRSwTXP03vttJJlOkYNbVyDEudN2Q3f3HCoUUZVMI
5wD4jUxq+ER6YdtVnuSE0bjAmrMsBQUAZWEFYNDu58bt7XP5xEaEr8Un1XPeWpml
i2XGhrpu6GhGfwSUVA/oCTj4C12N90RXbp1LrQK5oOMZwQrx6pqMCWfCiNAniQVm
jDO707Ji7M9WGRDJwp24dpxyugWeef3qck+3pVaI6GVlYslsdCIdUt5Vzk2HZp9m
ZlgA/nLWsP3wrkMpsoblrVDcWLV9Bm+FVJOPzXPT7gQSdDLpfCaRjntNIiwILUx+
B/zPvn4l/WbGyYhd1Oz3hJRllw4BPgQJbD3qohXhuGMRDUVM+FUqzALx6C3EER3v
5HtikEUJeAb68ZPLBy0GClh97GJcLca18tsD9rvHFICgzuHFBcQcZ3gp69GcnzUH
rAFodC3gFAQUNgZW3ufKw2I1LkrGa4WEooHkK3ycf8sUv83MwCLDTr0lNoaM8r7k
I1mqizzjMCq0zOz8+ACumcgARA8YvXDP+E0ShIlELeCwQsAx5o16UpyBfYGpCczl
4fWH3OTbsHLhvkbdNgyPzKWgnRAljJmFU65bphafGV1k/ByziOiyEKRgwm0N9rfw
Wd8RGM3Gc20x7RoSWZkdgo9NpKFdVbNYSZv+KtavYajFOfEvAGWh9nTcSSWwG65G
wBMRqXOx3WKoMveBz7F61w46dtDwUDscdZGI5fw0Cz/qvXcihdbo50waTjHoDR/Q
E5haTyxVe4mI4Ipa0ZFRYilE2d5ZI8c59mDgfLCqkS6mF7GrWOIPASr5z9Wwpnfc
lK+7zpOV4i36e+llEug1W61purhlsYM0K2Oiop+aYCS87cudT4C7Mex1eXh9g+C3
KOU8BducYW7zdKpuzqJQ8n1VadWU9Uw667eKH8zPp4iLTryXlPO5TNIQ8AXnXjMr
xdSP7EC/QNjWWnnSHidoOI3m1XxTA/GmNtHZqJnA5uybm5BFXRiO8xNsS+hyYguS
nkFqkutT6RO5gMeQiaPP7Ffjm58WTRLFvndgVgSPSTcNvLDCEKuR7pfDkusvJyJV
op7PZQ1SK+QYl1gQXdljDUR2a7cYv3X097371zQwmW03gRRgcjMsiq8O93ZJ66b1
BiimuYki1/MvsbHOLSnpzhC+TVnsnEV6pn0SGJorf4Sy7/QhQl3MLVZ5UqUQGfJD
+IyXCFksc+Ldm4wUsywCfgUh5mYjyuum+iknga+2IdLw9a+YKVtDGQ/O96C6uIYx
jiTcjxkUuAX9srJo4T9N55s8KXE1nfQvMYwE3pYmDFdr+08Hd3MlsDXDzksvwTKh
mUZgwdwPSvrXYzndF7jRMb4nDGM8G1Czso99FyE0iGSdcOQ8RvHHL6CdweRjD3PM
XlE2f5wlp1CMfFGoXnPbnJBXxcUQlttQIyKaG5pROx7i/Cl1eH8qqDQUcvD0O18i
5G/0X4bYaaV6m38IhKC70oY3E8yG76Ke2kOJlEPH+ToqEV+tp5SbHQ+lBIUAq/LJ
mb6xWB9QsAk8xYdbSvU4/gh5j7NJeonpns0c5V6QtrbeQCbetxky0zlavlOmtoCw
MxGxc7JUCjaigGq47Z3D4PFtae/xGitgvlo2qs56vVrsHeJYlBcfXQ58cd30Zs5Q
ol6WbGl49k+UNl3vjnGhEAaawyDuHYIm8jNd/1KohZXq/v7nwRJPJHCLbjx/+417
3l8k5LXmkmzY2SRpw4JslXDWU8/zXlOteDCFaogut0ipiE2DLl4st7OhlB+ymw4y
PqI0GkV7CKZzL/H8fku7gdvqK6c9RndR19BCfo8Ydu8VGcHibO69OxUL0JF00xtZ
rQbS3Wi+PZZ02YHk4pQ4MmoO1zD1wlmNtruWPpl5DGEBXwLZB8xhSiw9OEfakWBX
uFiEbQ/v7xeh8tRTJAkPE7THlR/2MFiFgWERRByziGht8YX2H4H9nqTjooICerED
2rtM7HRWd1wcY1xtSkTq47VyYgprOqnQmY1gnHE035Le36OX+Rhnng9ClCapaWic
JTkh3ZfRjXowIu6ofJ8iSSTi380uGbXVA1ko9TCgmvCEO79QKTM7zEjrgdk1s3n1
tZzbY/D5xGvbbUnOrjBkkjh8vIuH23HQflwPi0pwUp0voH5x8m6pWPDI/n+/APz7
cM1Tqu6sXrw0T2Qf1K8ZiL1TIGVuCRtLRHyhHe1GFbagqOHzFdjKizFiN5aKPrNv
LGleqoZPo9x3n6JXnSfeCmz4NYDiNTr7Eyt2x1ypZcLeq2frBMmPH7atkkTVFPol
KHmk8a42JjBkOc3iS89BgKFsCgh5mzO8jsNKUbu+R3I4TYdH8Lspc8nbMVHTaeZh
PaPCmHnYIRvVH49eihWDZStmlJjwWfpb6XNnQnk0j7poQFsmR62WzKSKy4yx+09O
gHefBUtRpEqD1TdZmwm2Xz4WfXVpTY3/amIbTNR+Hgk9UbQmvbV+DDzskYxQVhbk
kpsJgupguE3B7NpKBoOB/koRUES1mc4lvufhzKNk7zw+Krrm7u/zR/BaUn8Z4Aoq
qparCBeoajxMVkX4ZsiUWM9+1VaxYhVT+X4OKYPKJDoOvO0cK21nN4ujK+lPm0eG
vyJhBSksesAheYLy07VZAY+mgKMAvAj6eEDc/a4jCQa1IDr4FajxayAqUAnrU67V
uTmzlqFTIeUTBxcBVeAfU/RJMGnHmZia28nArSFExwJ/2/jOm4+visj26fqJK+A6
mtKFJ0jFxdyehtQtkkJqOZLhUUikdqxZ0DR1vJUC5rbC/97gWjqpecKZLsF9J+GS
3Ha62IG9GQFF7J3MPuzDHR4wpPb11kAnCItd6tn3NFaNcEUoRuL+3Qq8hFGdY5tp
Nbn1AbOF9JO+MHJ63XFPXa0CfqA7Mld/YyQ1Jy4vpbe1HzPqgYbP/IEbCveZm3JZ
7UTXobwxn+Pai35teAXQMJy4Fb9WULcjbAnseQs7q0YliKeI/f2oTsfvXGC/RHO2
L5io2yMcBOBdmk87DQ+72XqEFuZxd2HiB6+oBkezuNi9SCmX8fj8u4eKxH5sQTaL
gZ5bqaYiuShRqwTdnsTdVEa+4R7VcToyeEyD7mUj/55qvR1T8/EdDJ+l595swm91
k1wewzrAJ4XuPMqmOAso6EfAqVAyfCIH0/Cf2IyFEtIwthoAsGdDkADo8FyVUpsL
89S7IO/XsH7GNLqjTJJXEi7Cws0awGsmKoW0mBstz5zFFYH1s41eCsR6FPsnpyHn
BN4ZnYalQw0zNqL/P1WB3OrBv0WC/KhLM+IpNSGE0PfHyYVVMzCevhsiasrE5Jww
c3aEt7BXWLoIysnmxj3QNGV9KDcBBJ/G5Z9ZqbeQqzpJp1KZuQmT+CSWfIfzljl4
AQBvZVhjLFOf491SdAntqB8FL3QDlSotf/I4Cw7a1HSfnyIW3/HAMvgKT4BBftox
cA/Mqjj1kC37NYFGUomfr5d1G4M3teBZfTerPL9oXLhH+BjDdQPiS0o2VAjnn3W9
Inr1g3ZZVg7qSzwFXw7uWoGnfiMsAkROytviV8ReyeJeo6+DVTJ0m6zEceQxcPIk
T3lws2Lyz4dMO2g6HkelMJXTIS28Ms79iNK6hndvnnP5UpquRy0JDBBJlmeKpIW5
ev1R1dEQjB4eKC4W1baqtuN4+c338ncx4xvJd2oercECdMH1vCusOhQZRXOvFfcE
4D0lD7aevTxe5jVUVREevC6gkWdc6mdVimTz/r2K2818A0RJ2lUtf8z2W8YNeVxl
AB/sTx1s4eukyYPD76J+B4WPW9cPnNSFmuC51yHR/v33iXdQT3e+7jXuVOJwvYw7
iQCJO2I3Fh5x6xpqEUNuyETW3uv5jZlgNPDc+cKvpIGDkfSOHdf8VsrjEZXGzfEB
mm5B5XxMLyZArdVDGX4Rw0F68/E5mtNxOXH7E6ENNmdx9ybxzjQRlm+Ng3nwtk4P
y3Bohh6MqnPh+1bMoWMf1wS865ZIa8VaZODidLIX69xfbpoDkbOpfabcqDagwL0w
lUR9APVAz5CpNA8sGK5+DmDW3amenXl2W8CacBJLhEWJnm8bbSSgCOIdgG50wrwW
KQcQ5MEcaANisP9odOF3REpJwbmwqxtGN25v5sJfil2Kw/Z5xdf1DlA6+SbVW5Hx
OBfsRkJuevc8MtUXu9X+xeAR8h4Z8vQ8N4tu45L1IJ9OyMsHSUWB/I98AOsfoMHa
1flujYaI9ZrS9EVPbt1F426kGtcJQUX0QTXoRrtG1zXRvvAs1t6qS1lzpsFFZ526
mjcXUIHo5vJiAhE181du7IEYqkBeq04cZu4USozwCh07VlqQqm+Vbr/rIEzjhmIk
Ef7GqtYdweTp67YIYImdSQOyTCJutBaIYLMov7N2FqB+2zpP6NSYYbY0ORyXPStk
7CTiUTP/jXB8tuyNoho3G24eQWo6BiHxyWv9one3cFfzi/mrz1fA93N6W/d6I8xQ
k8lfeFwkFF0Bb2V250dTVsrJgTbJTFrZeCNBLVUIzChCPMfs8KT1C8FE8dkypvX+
CRzCvMcULlh5mTv1DpD1j8z4cygVe0g/hbbe/y/f6VsnQRCcsPzn6SUJXsvU82MA
x3/6TkDYX8lBCwYvrBxyhcf81G3XIvIfZ+QRshzq9yOPmI9wdhDKXrhWMUsrxOcq
vlm2BX6Q+mKTJCxj6GWdm8w7KIu6xPRY7elEFyjqVstM1BLUG58oxiBXjq9X/ekf
0J5zETulXyehbPIR4ihqj52kIXoEtE0FkrtVhvFS/7Nh/jWqGEHENH3qrKmPOR2c
YCs9lKLWGMBxtCztPsufaFqwDkKa9IJjjarrhOtCdWKTgG65OtigB1lpvkw8KoKH
aHGL2nCNfWHtPtPlqhbi2mrZZR95hj2EdruGPNXQLtFJubDk7aCIPayMuk0sai7/
3TD69Dd6XThtjraVGbrZyLybM4GAviF0+uJWx9r//O/wqQQHSBJjK5ySlCichQbs
pr1v9BgXT1mp3onJ5zFoO4p/CJMuw99U+omu0TD7XYKpzZlZUkARInF3YxpIkyVn
7lco8rE2iaysjUHg3SVxhOdkE6YW9Fz/NrlxdGgZDmnOPOwrIslVwqXhIiJA50ke
Doc86bWpOREiYK8T12knS3nV/eDicL4FrxJtXIMf0N5cPHPrQslfRlZ5lTLjJa3H
opQz5F49QACSbPk/aHVSUE63RQsaGZ2b/Q/dKGiUDCdyDNrMLp8L/3f6uHi1iDV4
Ol8jqrfapv3azoUJ3OhpkEJ+7XjekjyCIP08sIX6lZtz5brdbVygpJppWpByG+6F
HDkhM33gMTGP8SRRe19zvhZDwUSgkAJYOVLOKZiRm5kLmalXJSr5nC62Ljo9rTHp
TZuHRUOhscaE4Wn5mHGPuLu/qVL89FFxY0fDyNi93ISbKVJqDQf+ohYUpYootXPx
mrFv7PupzVHrBweDQdTL8yWibG0OGkXrVnmMNbidK1+VrCmFxwyTxttiNpJLP1NW
VsW/+AnpO6uCXBTk46WDJ2jtEvgJFcd9+P7/tkxoIoSjkygx/SqUiMyQehW1dsXM
bb9VeiZbwJ9gffFD6wQ15jz/CWc5EbYQP2EixD/B77JLRBOgrn8C7P+1U5RpAyfb
IopVUTWXaw6irn1SLBJwgeEqT4iNYJpeN2Q9kctNApNpSFMpJ6KVLtnNOuq2xcB4
BYI8YSe2eME+zMU1e7FwwT7L5DeP0vQD1taPiL+pHiKepVlw9ZXOCTuYXr9GKtev
8LVeKJ5UE4zGQCe5mdxqqcmnVKIH5gdRlOo/FWqKo+FhU8FY4bMQmE6yeEdBG0XS
CEDTojOz7o0ViOdhbq7Jw3GHjPrmkj+KjRncxc+D9o+7rq/Hy+RAnjOO9SRJEKpk
5R4N8Nq5TjiYbeYCqt3sUXDS/7ft+lEJiyZuVssNxu7ghN3luxGe99zDSFUL2jdn
rpuozVmk/7fPpUf6T9l0RRw+Hj4H/NT0wknb7fFyTd8pll8DIAf2zRXBa58wOAh1
EUUzxdSj/bF9uHAiyO6qRDjr0AaIOX4m4nvOD2rj0B//XiA6sQUVhlfg68dwLnp2
WKvNPOujoqpNYbJwRVPmNjp401QSPoBhy7FOPwXKEArfbUsmH48XS10Xuf6/6FpP
TLbBCn/rFWMnnV+YTN7SYSWg4a6g34DelvB40plPjEEBEsaGnie/xWeXXifqYQgl
u73pFeHL1DIV2/NZOtkcUTN6YZ9LrvZbNUr6WtQqm11xxpJRL382Kr4EBY2WlV/J
bjULd7dJIVcP3dAGjM3Q/GAAn/bPfE1R+seB39O8/c1Kx99ufrHhZaAAqOez3oyR
i2O7tWeuDkfrm8BAjf1dMBVmdsKOlYVuDYMww8ubnAhq7pds6rZSpYePu2dB4+O0
7eOtaj8qWtmK8Xlb6vUNfvQWWCwRWXhbAz46M7HUxZdw3IqKzCDfHhud4mm2rvOR
nQPI43Nk+a2FcKpLh4wRXMqq5HLu5tykA+pXLvkKT4YIXFmZchehBSw355ee359G
T8R6bSJ99iwMml6M5lGlHrXQ0EfnFlhSKyPl0Vkm43xiXk0/puh0k1u5lSPxb4O/
XUn0TfxNQC+geMZzmo7B5rb/E0b3c73HEaa8cakX8PsEZex357VB6wQiN1edfeQq
rym9oeN8kc41FStJIwspOvM+fV/t/WY0JUZkK2MQB3//2E9hU0BUQD29em9VhY/J
1EMf7CFxZu2hWv86hG0BsdzVrFUL/4bz2nQ4+e+uoVP13mKDS+IUHr1a9JEih3jM
vqo5f0LsCMAopEL3XRzDIhgUecpM38NGSAmWtxK5LcXP/tAxq61FbsLotkyVKxNx
GSUZEiZZ+eCSE2iMrwbaunwX/vFwPWfIqHEhnN3pba8M+D7rwIcKSxeVvMjVz98y
eObF6/IB5mUzzz1t9HZPc+la8/Ql0nK4Cer1p/w/UXnsbuxKAEfg93JOq1qwU8kJ
iAzfXpt8zAo384zh1+MRgKV36q1gVVjoDCHGoj/iLKoZuIPHgGDh1aYs3k74PguN
UjAapaBsb8Qn2J51xc0AeExmyqImfeVU0gNdPWZDq/hXtVue/q8Mz4nhYun03O3F
/wrow4jtVSdUsiMKINkOHVDQUhlD5YGKs1nU82cXuEckry7kdKk5guFOoQ5whH4l
T3mmLH8BR3TrUVXj2M4+swEWNQ6M8HnT3sXcPETzXPr8DMs/U3VPTjHb46Qkzf3Q
WMryGhL20kqQaaFpIWOJ64R9wBEzO2lfxaFdfYDUacbMgGWl81ziP/LUHl2Pn/zV
9SZuE2S3qKbujE3M2RGFmhYL1xt+X2OPjYW1mqJ2+GSX1cchwzWs8pKXtO1aR11z
E7TJ4IYHT0zY484wXzmY/LfluNYtPI7HttR2Ukv6kMr/1HGom445DWcAFDSdVnOJ
eWVlgXLMR4W9pIMG+4kVXSik2akJLBUC1g+7TdqSDqQo8SVSIv6i5bnnkvRMBft3
kaIrXRE80GFWO0x9uIw8Iaem50VU7x6pooJ0Ki+8eWtIoCkcAN/xouwM8haaw+XD
HTMI/Y2m9VTLsPdu0IlVZZPB8Glk5yBRJDevucL12TX/vh5l7qRMvJ8+YAJy4ahO
GUTskxdqSDtsUWFCtp4hQOh6y/dN5CVE2d3pcAM2N+kJEjRttZALC0GSUJ2mu6zQ
u31OqL5N5JcNt/2pikP5NMPAJlhkTGG3HCHWtds9YMVRWXxfl7K9aIco9DBZzHjS
zqFfAamvSCl6S/C28cBH2s3Wu5ydQoHrOIz9LX7yk+oAxJm5+gypHpijUmJ2btH0
A18Q7fDqdnZDcw4TX+iuJ+6RMdiiyR8sIfB/IIOmpblhO/krxb/P3zlLv/9vJ1oQ
ybCgJqITKvmwWCFDDn1dTmqoaQLd0c7bjnDEnu+KsCZLF3hNKknoa45wTRr5t28C
rivGUehBsSynhEPmeO81DFhs/DRCB55FsCaps9jQ34AiM+s0I2s3jMWdoHr7RIG3
BOQLNlXGjXYjTrLiAjiR+QRLCX1emgZup3nk+oeLIkht0chhQOCTzJCaXwZ8i6KR
CY3CAnnjwpejosD0ICWM+0V5V/xNI41LDXb2CNZphvb1G6AUTebG7rLiFEGz1Mf/
FKfTnrx8kocS6BLkTdOrujcU814MVPOsp60O5oatEI3GABjq7NQ8kvs17rbpNS9u
+UOsljpuRf9XmhBnTXCWuxsLAQtQcJYMu17xNt+VFDAEZPqdGGoH0Ph/eNaxGmQX
zVPgaOu/PySxVDnxO9m4cO0tWh0GAEZcZF8pmM4T4mYPF8YvsD+ZkcArkpW2KLrz
OFHQZvXfCWw69h2EQqVWigHa4m23q1UflItvcy7Ssb6879D//gsH20J9irgkCTuH
9MK3fFupQKJ36w4NREk1Dly5/ST2gxfllKpArRcGEs87AsL34JDxgOWKzgqZ8pIe
RWmUJPnBf5syPXUeDRy+jY6Cl0juR0/4723CH5/t0JZeM0lWWJHIFnSWudMERrks
P5YjDk2B8V5VdMEXy0wmKEfh3/lURdOSG/PLUtyCN/l429YJG30Awk/SCbvlYpgc
Lo8l2CzqR7v/LTpacExKegKbkYR8YdqvQnnnaoxSXGBbkpzcsg0FN6y1YUxCYnNc
b7CIK9/N9yXSiHKDjxHqobf/O8LV3vxUNKGRMYS2aXyxPLXkQJFlsI8YP/hURAc4
4o6vtaSmRKNnByRFS4w5LMZa1CyfbIX+ODu1kKgmU0v8q9RC3yga50JG2h0feB5K
BR5kRYCMP3EnzpJeRjBlP9c5071eX3nq4ZqgDMF8YfJ4wDDbFIdWyv2d95dKiSNm
0tSPLdGEAIRjyE7R236vTjRjNhTw+A8BeBukdapk/1BTE6/Mpizi/q0oNBQ4RGSS
/jl7gK0Q96+d60UM+ojDpMmygLL3QHXDlktZsQyks1xLZhR872lhYB+OtdHl9/Kx
fhBgzBoFTtaaFK9+LbpzKJWMOgO0YU0doqWuY6px0ekXwLkAgiWJVyZyRA/F9Glh
nxAlHuusSQ84fwDI+wl0BKu0kVLjsW4GyZrQErCOHQcXYRU9SvV8satJ1wpmZuEd
CUqHHB9hWTqC6uraBljRsATqa+XFp8uYRQUBk9eeXJRUIlkS27TLjULfte/4obnr
UL7We7Lp4mbiMnNIY3h01N9pGH0SpmfSceVx9ZJltbAnGPqZ8Pq56HPY67ADTxhZ
VXDrXKtNZkIMBJjNJjzkHU0lfBsP6pcA/IQFZrUha0boOZRPpac9vwAnUyF4CsEt
5t9MjKtpzfDi4PMVtrk4T2XBfSlZxrBJ+y8CUUpKqDxjnRfl90/wvt3EcgyH5F55
kIIj7qz25Uqq14jbFKxhWr+WO9tbmymXnA6xbekF1SRA96kI/k2gngMqqJzfIXku
w0a3w8+gbxSjT0nAmUkVDmKU3YelSV8EEW0I9yQFMrkm8QAs9KPSFnF4FnYywuW7
ssJWn2AKkMvEnHeIF4jNp02Gq4hvTTFfI+nzmkw+wm7uonp0T/2riqwnBZUXK+aO
w42FXXboPTZ7FpVS1vc5gztxC4zd6J8XO/if64/zW72j72mQA66JLZiEiM6Pm+Ah
kILXyF+30hG3/E+tUEgrHCtff288+PlyPZs7UBArAf8o30fq6meEPJoZCeJ4zebm
Gd2inhqB+rNpcpcypIuYCYlQtWlIkYt5u5UhR2jywOM2+Wn5lOuSGHsLK3oRT+vQ
h6gDp7Gq+p36wpwJEE4YNiYW862jP9FvUEqHPDfnZL7+kCMWHB+4AigaszUkjF8T
NMeWdFLhCcAcfvcHM5vnrvg9TEdGz6OPfkrxKNf0uw79YUnAgUp51Qugq6RkXBsg
cyOL6fTg1ExX2ws0luKkob9ahJOKgO8nJDalLh/M5J1HNkZSKyaFXQVstpS36FVC
LcNFqZwrr0AMRLmK8Ft23lpyJs3KgTmXRJyLAUWg6fRsH68i4XL2DYYpglLtUBPl
y0KBb9irMj8iZcFMvGIhKbinnTLACxoW6nLz+Ta1Hz9kb282rdzMbhLjiHO2dTMs
KTdNYX8vsNEpPZ/wtNLI0sVKxX4f8TIBp4pKGtQTQ1TRSqkjjbxszT/+MiS629Az
+YTiz853I4AujuKwsurqmykjpuQN6+nxl9Z7hUAsnHC5R91ACjHb0lJmwnPjlgic
FTMXoDVtubaubseNqpz2YDSw5L/+gF7nN7GP931+U4GSQtZsQa4+MK5uw1Nc7LRw
Z7IMFkOi3icLF+kkfFhklMAGi2P4W/rU6Jcpz47P6fhhvh0+17ZgCmOQfrEbUXT/
lUSCbnBQRN4WxP5yupXjcNyEyJ0Hy++H/eIWVaRwkU91XivlaJaXx2+58bsb9qKs
GJJkocn1Y/75U3twXOXfj/NoH+HLMBfeY0tVo/GK4G/c6rXGBsYaOmlG03v/veY1
X45f7caur2I0B314hBtsQ4XJwayyoSIpKgq96S65TM+z0tPo71qApYE1+Sb+JPvZ
Okp7xOQS7w2W/swV2tiRF8ax0pAM22eZXmxs31kASD7yt8o7UAQp8DKYOAx/hHfY
YgQ7ORkJmBAlf0RckuK8qxxsVch5x4pokMoAbVTQkhw+LPxWMuxIYDPB+o6hS51P
CqFlRpJfkhCMg5HsuNXqxg3Rj9EY5iIg1NjhgrhzmvzCTvsKr1VwifsZiGnzHsrG
nEndXmzz41i/fhMpW/GDzpcUjQSV40hWuUs0FsZvEVUkv9o+unb7UKt4aGn8f9Zv
XoIz3oHOyHD6ZCspFwHrrlCzTF2UQLU/O091m33IPtJ51oixLWBxCj2N0CK92t/P
URzN63W+mvP0zQtvtHzCWjCrQ4uyC8eeIYCaV/nUmJG3aFu4Af7cFTDBRXkdxJzT
x6/4zpL0PHHJ1ZqGrtMz24sJl0uapnR77CFrpUeL49RTvCDVidPdQBV6mFD1YXRo
j5a6C88tzLxB3JDGDZ9LChNt51wct3KzndFA4/1H1uno0M+f+54Xr/74eG6rpQRc
XcK9J3ndE2ZPJRqQJ8t30ht6wXDeB/z+VETDTGMtrZoDpv5rsbEQpI1fVYD3ZdQR
UbDBx4joAnsjPcroZmBhOE4W2GLbPkSPm+SEX8jFTdntVllfUbYkDbenWeZQl9AQ
xxUJWLfkBc2ztX6AIf7XXmpx+0vtJi8odmYOk/YXHsrekjjo7Mr3o37TQSwWFqF+
aaI2TpQbq4TuomNM3rO0ItwoCsmLMjlbdxgiDorpnqCIdZXf1+OCyudxSAe5/Zzr
KPQYTzove/yWGjv9tg9+8NOfe2/+3rS9jWwQI8KH8HaB+3wL0XXgyp3HVjtEyAPE
0gDNaPeOo56QxDAYjihlRAEJqELlYGTgNkX39Ac2BajY+R+oUJZt7Ez8S5ApoJtp
7O5nErHIeCNYB7osTHxvtigMHgM9p0EFhIeKTYnevGBOcYbTyp/K7hqKTcUuVPWi
uOWJ3vt+xjj1M+k4AKsYQhwRMcDUKjUnHUzxb0t58oPDlHvoN/BDaH5F3CppDS7O
rhWHpm/b38yArNYUiJGLmFAJbU3BpuMFN+ZVSS4lzP3YrOOdg/05FlQLIHoZWZpq
ZkmRL3LuyFqeA/abdV0DsYu9iUlKGtBJjntnZAs7abmKfPGYwlb3Xsiq3jvu/HQv
IqhaalneYYRoudDFxVNuNFNXnO+Hkynd1heLtND9oMvtjKpJzBJSyNO8SOQxtO9e
wMrIP2GdNr/wyHqFY9FsCChs6aSjwPO+tMUDPRst1CT06vIa5pZIFMgQeBcEiFMe
q762pVbwyLsX5xBDHmQfX+G/f480gMiC0vhVy74Zq9vRKATwJduWweYhbvKd2vZk
x12pfUa0vJVGkdD8OiwfGKKCKwkYznlLclxjIrRltZC/tpCyFEq9u/4FjWXWxuba
R8/wfiw/qp3FK4dvQc8OuI+4uIv6tlwfmkkGo3HwyN51/LDpAm1Fv9oGcunBHxWD
kOp0ebCy9MXUtulwEyzxVc3R9qqLN0kqZabfKob9flJLxEQk3L2AKxrwZtqOSOaZ
j0iMELFwLhLk5CG7JDxpJx1cOjm2k2xXm/C8lnw0CgI/LIOBT7CFWD6hteDrMxdd
5kDFv+jKhfbb7YMqBTZ3ZEM9hku7iDacblUxlm3ceWbfwuQzpSf4iuTY1X0rm2rH
i03+AB6gmlvLfLn69IrZtuoHBbdxzDhI6OqD606+XEjYF9sZc93zBqgH9I1gEvPr
PUt/6uItaSroE2vCoWsz7RmAfdnVVc9OddTIIXTUu4PvS2tywnjYoMrf6MfxuTwV
J+1JljRwHM/Vn2aj5fizqqZEW4hT0Bsja371tl7ffRelxG60DmTAEEWt696NVvfn
I2sABlqIDKroIL1FuXsWlEJzg5vBNDdVfsxqsgb5gLGklDkqk6QUk1Qom2poxem2
DhvfY5XI1I2TWR3A+65Wx/EUkYRVEGtmK+9PBiZ2sDgfJiIv1WiXk5klWsQ1W1Zw
0e+Gzjcx6Lc6yvnASuMqClPOef0xLFr5l1Z9BRS3LKJxAu+TKsAF/jIQ88jUQkxB
/9sj+uwvUKEXRmGHOwn1F1wa024Alzc60OaKFR2YSR8BQYSuOn873WcrdkJkzEDa
pO3ZO0pZv3TPlfZANACbBAKTKg3e5SQ8Dp+gL+3dacIWMtxv1eEDMxZhPCYLh/NZ
PpV9eACKvzaH0gDf1VU9o9NsfVspsN/hRM1/PNDcJagd4fGmcaOTTU2g9XStHpsf
3xBd1aaRKAT6987xYKALVqWZ0LcYmdeQB/tDrNFwrO3uaqASnF/a8O9mSYj5VBon
5YqFpGkBCykGIdHN2pT/usEW8cK8/WKfiLaweZslpeaAKULDVWMQFz3SlurJDcn5
eewC+SJMsGCmEjMzZJM4LjUAnQreEOtNAMVsVew5XZg7sX8+8uEet+7H6y4B3178
HsDtbz9938sKNl1aJTENJ/ZvKnGzTHXfezP82PPxxq+rCCgmLZrZrYjneb/aWmWK
W2izHnN7we48fFLTXHZoS2QFBzZerElCS6ScGbn9LRRHqxRqOrHDWMNv/XcQwU5l
Gar5ASTwqEEdJqZGnlVZ33hxY1ZciFLrk+3sovelnaajKYXI0QyRv0Sts9vwfHxS
MQBVPI+rVj+03smTclC0CnH1QQJNJZuQ4HDvbwgQ3+GEivted4ikS8FykIUawlZt
OaSiziVOiuihRDYqquo0XloV43jfQlJCHYhfe5QhH2Ncn1Shl4U8hJD3yAIURcDA
3nlzKc4bA3f8bRK3F9ttHwgrGYn8jb1doJSFNN498dkqnyMrm4pRfnNJhCVvGEpo
DjjFFajE0pZO+8Y3U5et49FHlUjYMvoll1IfFwCJoUA=
`pragma protect end_protected
