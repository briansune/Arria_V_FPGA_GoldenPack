// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:19 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DWWfvr3Q0dTDdmFVmmrGSa11o/WEv6CGP2NBVrIXGXBWETBYBR7Mmhc7CJRTXDJh
bhJxlzpcGnTB4jjt6Aq2A6Vz4m0xbMc9FWt8mr9xX+ZaqnuFlYcQ3Z8AKxd1yWYQ
OpP/47K1A07D02q0B/if06rb+yJwHWgOX/SrgwGYMk8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46192)
2h/6UH0wVj01J7xXx2aWuxMjuw0Y0W7N6ncDUX8Yo42LD0qSEv0yPS3PylLgBf2G
qNpTr+SBZxR1hlNzW+zO/5iR3t0//SjicqPmg4qnGIJHaV2Bl6jvkbCmggZSMQSV
Y8Y7ySKSGe2CrLLX2w2AhOgckw+HNPzovliBfnkRSn5y4c/eag0vg8LUi3E1e8tt
YzCd2tPCW7+Yet1iGXfF6mqboQNP0ICmmKfX5hZG5d2lUCCoTgI4U2jzsQsvdnag
I0tdUN4Ejmun3lO22I4/UdCiNqIXQPbbL1+ujQF0Qc4U1cpt6zgENPzEv6yCwiAZ
iuPgV5tWFq4yYOBnuGGCnqDuWYpKFwnFrr2mKTtk7mWehj66HVO9e14HBvBsHcjx
XU4QDApxFhdFqKTqZVoDDu/nbias0yU765Qmj+vtikVIReA8omtq3jyiGx62W/0T
DI7rf5bTtiaj/x2Gzngs2IKUuVhBkiGMe7iOcL3jGpnMsg/c0CQLXulgwGbuSoIN
zbyVJjfVLa8nGdebDgOS05PzlkflvgCXR2DDsxCFYXAnbDxTfzn64sKLIVb3bxfW
VpPk4TEr0+EBJcsAo/zhcwQyCjcI8g9y4/DvWn7qeTLp4GFSLoSDxoIDtsefI2p4
NkJVq7kLqam67oGVnWPhjRVogV6vd3pjN5sUidG1o8mgIODzWp/EH3YwGG3GXQoL
ZtLUrK2Oc3AP5NOx4IAI4ze/2VrhpgQyJoRsrEAwSgZ7mJL3Fssbm9wi0wD6ELEh
tKM28Cg8i8vg+P+PbbAGTwgcz4Hd5XkrS3GknIqKqFSUZv3MzvFK/f/byXf3Fceu
K3pvuc7P+ETWohm2BPk/dwcKz+DyXEgt91kj4x6jv/cFBvFBc+kDE/KBUX9+U2Qx
7sq54KLPeGl5YEpA/fH/7r/uJRjsX1EtiXlNSEOxkfnzPLIyna96qKlwTGi6t32W
rBrUkM+gbChBK84OP4adLn+yFuvk0wsyVuLBb9YmCouXZoXTa3rzdyR0bJbfHUxb
MPH0YJHYQ9fI8k7p0/YmYuqZ743++0jpt2L0RskgOPAwJimYff2hUqAsBrY3ZXD4
Lgt9iVuSY7tfLUKOcjhloaCB01mGGkag2tvz8E+2dYXtvioTeKD+6oZFHXOqGXTA
kZzPmH2vq0DHmRQ62cAe36DHye+UJBHqwXuAAin38pxtlpNa17dM7SyVysIzY/gS
7gqPUA7mFjw2/CcIuOSD7fOJSWp6IVRcTf36pebsckuVtAL1cfWBA45EXADOaCPD
k4fNfMeUMNr8TudIygDc3AHofajJ5gEJuqJA9DhDRixQ9F3z5PvPGg2zcDSk5aFN
k4hmIOpNnhCZe4BQq+KC6DvWF+ywA+vJ5JiWBrSLrkbPs7RPezzahqB1kFxCJBya
3xO2dNK21AphR9MGDTsckwp3dBqZxR8rGMkIRfiApf51WWtl0JLXCm84wR9euT23
HQtWBOXIwFVCEXKto76WL14aNiegaK8FnB+0jSWt3uHa6eoAEtxDWTxUQ4KUoImD
l2Pw17QZshBAMBOFyv84yq68WHov0mcmc1jjhaGqkYR8cvGY4zqKoY9qJQN8uoMO
tjgkxDbV5LhIkcd8VZ5Vf2GLPuNIHOF2lU6bCEkCl0teOa7Zvk6QVPkU4dj7X1CE
ZVesQAJhwLiaXCmkaRWZ0YrMLphA4mDIagqbUD9bOOuT1GoaiRaRo2OkEflT88tp
PheAkpSaXHPgmssiOdbqwKDctz89kGNZR73neiAHDxOIcvN3SXbrgzBmyWf62y6F
qfGvxIWoIJc0ZCQZ6rgATWfDOrCI/JLJlA1a3gR6b2+I5poUd+BwALOnX08nVigU
vLQwQuoLEs6P093eiQ4Lpux/wHoK+Hy+KIQFnJmGjLyvXfG11MWd0ubH2U+cE1R+
XYuasSA64vnZgoeOFI+jcSQF8ZCt59qyEzWK1GX4SNWvUpIC0I5mv4vPRufhA5TK
h0W4aGFqxT2ZERr2K1bm0pG7w7zyY5kvpTZIRMVdhKaAga/aboiTV/9+Vu2tnSoV
rIce81m+KN6wEXvco7opzopKu+jygS1N95JI5LcrWRK1qHrfGIA5jCUrI5Gn469o
778vYECRuXiE8y62OdWLfBX3xOO+BcKC1sJsSyxvl3W1pyr673CtDG4iJC2iasfy
X7MpLfu+4m8vbG5pLQ/aJbqzjHoGjRXqcf+ExdlnH8fqFB1QYGWMLTrUH7OhLRCS
vDlvA+EswrS4EpQffVWqKWVx/Zptlcq0WD4n22Lk94dDRN32ex6quV2s3NjKQD8W
oVVTjRdPL26BgIe9Q+tV7My2s5ow+YR4XR+JDNqAoKKRKrl3HwY4dae19lW92LDt
SDlhpQgHs/jMl2oGjEPGK3GPRmZr7wgZmRCksA2mkFBbrPi67Kz5AwecOt3FNzE7
BNidQmrgSVOCDEc03FHREOTtDxzWPKV+ORRBuzNO+XcFhEf97y26j0ajVK+nohH8
S+8X+5Ya9Z2Mjfrpc7mZiWWk8UxBWNtDM2ji7bJuDgEm4dJTdUdHP/noBNQnaO9A
pNxYE6E9ZVejqj028I9eNxArnDQiIMBT1zRLLJoi5dK7Frcj0jyh7icZpwiasDEI
ypXBd0iWDCkwBL2vdMthvSrBt9IxaW4oNqe/Uq1a7/KkroKQ7IYZgu1LoJCvflMi
9uOklatY3p9m851pwVxuidbx3/fBBe97zk0AKngOEwDYwTjiGBPXeys3lIs3KE+i
0xlNhESZeZTs8/n3P4bt74mw8Z264532lqszAcYCpR3pFWWawtmzPv29SalHE+ie
p+5G/y89IxNbNIfQenMVFoonTsapfGm2MUXyvblfyC0cjWg0jU3yQyRmmmYPCglH
fzkxxm3qWauCN1xAD8qo72i5GmG9Vw+GWAPR8cZcswqCQ+5aGTBbukeKbcbUfxI7
5O3IUBt1iitAKgX/7jkFjShCSx/sS2pnptHvPuvad2fkwcVznLgYmPq2Eyf1AqZA
j4npIfiPJY4MXVY2DMQv8Y1zZur3aeXLN5Ge9DLG5mLZQdaUC/+EmGoRbOQRkPVm
L4CLU9gswAbFsS67LtFCHVrkViEOg99919iDMhv7LTZgyXgoYb7oZE6W7//9IXyn
FZdODKhtlycmcSPH/rSSVv4CEC7EZguqPH0VkNLp5C5QCE3227Z/mo7u+zr85U2g
3eVDKwiLwKgvjyCBN19VW9vQ4FpambawU4bMr6nWKhfJDUEziUFLvwCrTk7lL6s/
M2jVSDNyFON1O9lMgxDu8IzcR+2C8tcK/V+1BM4BCcJzPt44iCGD2jnW8WNchGZj
5HUNTII0UHq2J70ZLm5ZpyTXvVYhgcenNNdhin/2lZre+M0K4BVIQpJZtfKl9xsk
uFUK0Q98BGGT7f+DoQlI9lZgfv1/lAq8aAaMj8NZjB/SHGtX+B0G4ZIXgQgyT59r
GmG1oBbkASPb20ufEVDDvn1uydQhWh4m/ayDz4iHJKf33sSfN5m/vhFJYLnkB/Vm
hX6LStZIcBD81MEEcwb/L7GwSp5JZUTTdFnNkUc//7UAwRgix8I9eMROcOJp6Ubk
kxYtPuCL+xTd6PHV/D8kjp/m3nXt3RTETFwyvphNeGwQ+lqWtLQQ3DXD0XdDcP3S
Q1SXQSCCWQ7anYrl5hdpRN/8hOexhaLu2wSVsVnZ3lIUgNwlCHcl+2dSDjoAeere
XTD6erfAMUpZX9dq5Vein0cinv3b6QckSrFFFvfpXsJKHlS6irn9WwCyIElZS8U2
Ndz8vH+XHuCk3vfC2UDkE1obPX+w23bYtOgjD5eCB990j48kDp9Za613QOF8bfgP
jTi9pKCXQVnXOoptD7nn6cLx5r4sdAm2CBippRK1Ee6rasMMu2poiLOUGHX5MYRC
d2CVRpSz8aJmb2tcL7hsakVRJSOpbicPyTKurarhS5LLrdnqEJKTvI5xYzSxTRXJ
XDV+yK14U3Wwi9nvwQCgonZzo3I/MXHRjQNpWp9WQcf2TaNm4nUMmrKLxYvXKDDo
kLfFEjtM2CeihFjLGdi3AfVxYebBH3MMrP/yt0adKQZoWjklprDaiDSYIYaY8DN3
Y1CC+5Snexw9QVF41soSKUOjlJgih1quTFNMMB+inFOIzEY5AzPEiqKLYQSTwnzc
Z0usIpddFFg6UL1/16NV68F4svrLi8wIO4D9W2W5sFitzPCUOoYVrk6QoOm2idSr
kEJnnFpS/iMUbyxY9/rvRpRiWz2llT/NfBzOl/YE0TJBATiHLrUw6LQD9gczi1xL
Vmio2DGv5+WoI5QL3Ca9JGGSsNb9EWEdUVOybpbdDexBE2AHsnliB2NH5mVFpLf9
S7DdT53uWs4N6CNFlyDY9JCKf3om27PpZeU+Av0VHsui9CUV2R7Eh0T8HhDYwUQJ
rvZRf5r3OsZlhhzwXcaz4nOUmW97sKZ/1R8AsOHA+4Jnl8VjY3b94rbIKtZh6Hlu
jEr1sptp9+cxWXyCBfFqOQR70M9DWU0gDO5IQgU81W9orWt188zlwi3IU480pMLZ
sbVIjYysuN5aPWJ/31ztjtoInWOLsEMtDEblYEaHDjNJnL9CmhEvqgbFlZ2lfTFc
CQj98RsUa4AQT+LAAT0OIM9jM2SHtFM2M0LKvrj8eOjbS+93mBHVyJ0Np8jHBHuI
cWXYJ4k7D3MwrT1Ah538vXgxhGAe1fH0K2EWGGlzVQwXQwiRhbT6rNdqBGe6XFl1
QSDO0rDkr6O3Q4/HRhLXq5eUuYz+pIkRZKRfeun2QNqb1MDtO9i4ZSfSyZOUCZsF
wmBIlTMmLrvOEY713nfXK9axRGCu3t6HEQLfKLupRMnLgVwZLKCjwKak8AvX2hgk
aOEG5+aw6ogtBzBbO4DN/uwvtL21bR6eG5wJ3qUSdKsivj/y10Wx8MJTW4UsAJsc
6WHN/sbBu/0KPT7GEG+4u8GDEJY+g0SXBZdMdBW7pr0QdZJUd58U+OV+NmTq9TNI
5eR5KObs0C0JPSCA2rSOjmwUzX+PUYRwog4V3gOUvzHj6f9mMJZp/23VMHA0tDld
nuM7UCgntlYXiHuazYofq/TZ6b8j0A5N7kbYaE6UZHg8k6msleOug3AF9SxR4Nmr
4fTAmCqb9werhpk/JVxF2dD4JrDEdMRe8N1BS1fMMsISA+Bpe8sNc2eSjTkw9tKp
CkrcCaZJy2wLD0p+UXvNkia08XeBllOdMa2BkPjesESNo9IdkD6LrsJYHICGOh4d
Rw/h0RKVFBEoiQwtDgCoPIY+NB0Byun9WObYBwYN3MkSSONR0GKcKO74/ykKn446
InfOWDtZDH0CjBdFhM/hyL68qQVzJbbp9KpUE/ubqnT392fLZi71JRGX8azefvSg
NoYdF4nx1E7a4dB4pGas+kkAiRlp1C0AUtCf0HJa53r/ayKFyCig005ccMXMfChU
va3U+ImrSZml/l1P+t/d/IIivkUIndvKT+2YkC+RbysI44+0t4vlarfH7nq/6q4o
ojZMhjsXoBV84rRJRYPErh4MOotV0HPoK3JdzF7+c7Os9gB0YyPls2FS0LHHEIAf
gaqGV1Db8VtFKoALJ0Le27xmZ9Ajg5v2vm6o3UunF41V3oZwWOQsztNfX3SYlvq1
jKIwMX6Z6WjyakwS2W8aqxWWT2wRq1OEDMoRax+MRd6ZpDRmsZoFMCdp8C9z7EHa
hZyMkf3kmflYX2jEqm29NrPzfOFCvtmIF6PRuIRc0+BXlAuzV3d6jBdFZr6GNxP9
LjC28F7Hg2mumHPHq6cOPbiT0zt/1jdJQkbvI7p2CPb34OFUczsZw0mapQjq1cYl
HQrBR+9i6IH/nfuzr50qgSNM0/+BFkWdI9wOIJzr9/HiAFwmxCTocp2/UAyrN26q
PsXdEhN10Hd1E6OSqh+l0r423LFXIW0lPX+e956BP10pOzwv6kP+V0kV5xAHDULH
pm2Sdw+SIHQoGJDYPXavRw6sO/KKRx+c0QrmZwNHtQFKkpCf2AFMsny+W6xaXjBi
CZSCYE1fLMFpkGBKA1UHBhDmr5gtcyurdbXfTaDN5s17Om833XpGH7qGYeFlJsXp
0yWmhY/uEQxp+6NVk2prnME4qwNDhnbwByYWKUDM5VbqtUmeU7lZod/kVHTJpMnd
bOH7iZIWg1n8wWmxWExIYS05J8Kpd0VykPvtwbvl1IozbSBH+fPXyyPKOQ+QWNB0
QMF0/Y1Au13s+QZunMQ5eEDASpVmwbWq3oJKdKJ3rzkbBFOuQTrsJIUV8Yk5zOw+
lnz749wHlkKWhhH7uDx6hOjH/cb8E4IR0yV/ong4vF704/ASgLktvmhdfXQIq2oy
8tKsscw5JpXwjB1/rfjC55Di+rgX/nDDBYzDKpldBCM7OqT2CfIQhJyB5jVqJmeJ
90LwYGXZGFsyBtBm9ssi43gxM2IVv/A3cV1PF6BXPR6elex8Orh3PCHz9429GAB6
7I+eMZRwOa7QZ+zTzFaJEZHBxzMd0n/wqndzlV2SX3fYA8AqXLk6LRH68PdfJBca
goxktY9G0uBHdc6zfilGeaOIH0teOz25mlPYckzsLRdpCv0FR3l+u7oq4MpS9Y58
PH8AdrF4shLjf1lH8yGZGE4EBLd69hXIH7kHUD+k/98C0dYMfgOED8kJgHAnwlCq
A/oeFXv+gzczjhQ6EIwPrb6zRDbdz5fk8pA0OfWE36KcDvNN8IB6v+cPMplFMPv3
FC4apr65F2t63sTGEROAjqHGLVx6CT0M8swR7rE8xYpcFhXbiCG+9jjuY1R6qG/J
rBt1mzW4MfTqOsXRCi9adUmSrtKjdXWBiUejNwxzeDm7RJTBy9BJcHpane0MNZxG
07/Wv2nEDDXttW1G7A0w9nPWLvwpnPkJApSepRWzpj1hThQkSMuJQKIifs1KeJn7
Qf2Q8x002jjvmnpr6AvFBeuGpZgQhFCnGwi+ABnjUs8jShoweuTAZ8aEYB7VZgv3
29kTS9ruAVxNp5eP1RwR+0QbN3sAooo5dVOdcAP8uvPY13ZnOozmIUOgVixTETNY
Mz3pQ0wBSb4PMY25+6KNdx2B1cIWIPgJp67SVwrN75M1x4IHJx6e25i/r82iy2gu
0emsRAkjTxxBP/ZEabQb8I9AWQp7MOVeYf+aiffH27mSWU9n0hLbJxWtvOofBZKa
+NJGgf9yLOMlqQiGQEjoq2K1AP7uMl2iJspoBHbZJH53Uz2iETzZnXe1ueTK0UlH
6S5PX6haf1/jJcn1v/NnUMGm1ZeULw9m8fT4omnaOXUh30RFpGIfKPipSexOQfnt
OqrvR3X9s3OyDg/tkqChaj3UpxkZOljOpJ+eB5WS5wLfFtuD2kOua4jYqJ2+7Ds5
sh3LOiJ4AIViZYmW2Kpj6WqR0wJ4FaXtNFf+bz37Mg/qW9YSyTGzqzDNQyI8kjVJ
k9Y3ocmaSFIv1ykl5KYIw/oWNvE35Yic0H1CLf/LLqNbpU5LIIpGx/KO0EOvrU8y
XPr6fFO6Fo0l3Lz7ZdQLInp2AXjJwo54rhH5xcTb7xFf/ve3DJaSIZWPRSBvuL/m
lsdaETwKSLgmadT/lwqGyUNq1THRFyCiZw6GXPDNd1MLbCO6oKjg0pMHqu1wnzJm
TSWC0ywFEVlVDspCgSxPwPpzS6rmRCnXv/TFedevqZvBZF2Vku3QuPEUB5NvWBlp
ltnvoJrQFzxdsP6E7clJNi5yKuLRXi+XHqZmJHMJbPUntsnI8oYj4hHyKffhBlIa
XcPv2KXgT38irszwzTwaLt4pMn62j1mQ68fZqulHeXAATX/q4uyHY18ojrDoDzvx
NC4RIFobsRRb5+ckumIyAoXkQKRfsZoaI5/Z/iEM5EJqVekqw+dz9yhrDT4nPp95
vhA8Q4hfsS5Jv6Z/MRXC6WvT121Iee5haqOWdwW7+1yPZXhAVLbBLfiJBGn0tYC4
Q3KWx0IhMC4lXugbevzBRZXs4gTfLIW4bMHv2Yj/UdTopbddZFgHPAbwQ974Bfzt
EeUL6yNvUbfUb36ifIhOJsn4nzFjvgIwkPCpkx8ameJH5uQaqxS11YX+7ptxrAyb
7EGfgJi2KjxZo7mk8/Xn0dhgj1D2GSN9UbGKCu7iqx8YaQhL3Cq1rjmmK8fNP5de
58TAJVeUJFiwsKMHbqwfCa+ela692DB0Ao5R2ZKSUbICBePPr/wx4OXDxTT61zcP
On95oL6oZvMA75NaLZCWVcFHWjfyC6tJeSh05Gt+J5wW3EQegnEh3+yq1C16effB
8lP0t1XiDJ0RVvkMK7b5kCH+9owOtOcJHjNYGsML33XDJfkVKiFZA34i05xkj5Tn
rExPa0fZsjXzSJlzQuxcelVVBQ6udfeeSpBp8YCrvbvwDX3wjjnKHrHNszktu/uJ
OjBKXBbIf9t3U1wWc/BjKgRMvZdSlYXqutOFKncQSAvrMkO/kXj3DZYZYZD8NiHp
zx8hI7MsNfkJY50OA82rfEpUeSNaSmxjXAIMRZXQm3hSXGXwwYrYqv1cInXLEW7Q
03/rMUqp8p1k8eyr92AeeH0vz3owBqEJfeLN/Irsm0Liw5k2bqzQMarCVO0UjPgs
0cHb82gEkP+nseXJJoswVDJ85g3NcVA+qoHhFzJoKzugagzNU7c9qGZIOY4RwEu9
pcqS9zZuZd/BWeq7P+EPlRQOPtu8v9kLrJQ36VX9U7D1HnhCJNlAh0CcQ78RbZQt
C5UgOv50aLjZDqxx7pKWoiPTpSYc2yHCprKEyKbiJdL/CUOTxAANYxf0v67fSOZf
qMAY7BRhF0bK0NwZzXf5UxZyQavhAKqQJ74un/lPE+TsPo2tvSHWKo+nG62Wyrxa
bN1zIbX12/M+ZBSkMO43mfxW8LfUmKEacyVPbA4Lu+Fvhtyn1Sj79JxRdAVhuMiY
DF8Al3ny95QcXeU8/9r0pAyUNdArowwNmp2O4PfP5jAMopR/6f5/15b9Cj8aBZyS
sUA7Ej2ZUnYvs8eNt/eEDZzxBANCelCGOKXrLoB3Xtj+AAHys+BRGYLo/lnFy7+0
PB6hjhTU+qnfNP9Iwr//CwTU5YOxCGkwP8U2EpaqFGcbrajyK0cw7nrLMzHTKMDu
X8aToEU646Tw7yelUx2AsVPHWwRqsT2AYVIKTEI0ON0Fuuskq1XFQghiEYSbE/xt
rRmsXP5XkDXqPWK1OdvlOb8csR4/vDc/UKdD/mRHmjioJJU3Eym5KVXgvzCRfOvL
6sIXQMwpREjHoWCMNy7NMRk6TZ0FhHMDLHYyDXXCBF5cYF4qWEZ1quvegc4dGxZe
k8I8PWih1NDrw32ZVWH81g+UhDrus98PbkLqERUU1uigklPZolcbS0h2+6V7EvL8
EO/jnl01YwTPZrauxso4OebgWauu2S+iCghJV50CPYpd/q4Pu6ij8UNPNm1pW1Q4
kfz5rs6iGc9a2X3AAzouE/ljkT2+eGdFTa6EO5XNHthFJ059dUWFsG5zJVdHlz5Z
uFItr6dKVjijBojRBoot3g2JWGtYpw4wl+rv3kCEkJlp7NJKh+WXCVDxFVUjp1Je
nBFlejPsMXyFecu2/En8/UuZmnWjPQs9BTA5OFbdKf+3cU/djWYyBzy7uZD6qaOx
o5V9+ZvnMaAFmmizDbQATSVM+Xq6h4uHiH0P2VN6Ok8reEQ06wJX7G8TDM6wRisG
0tqDznQlcE4JKQybQvzwp5EPBNxUu9+TCqJ6flXmR6q3ijVeag6HNUbK2PWpfjuI
93n9OM5duvjaW1Zo7Ih5SADc6w5wRw3V5BdR0LL1CEtb+nJeeCl8gwKwctZzcExG
QEakhkV9PFYbC/NRgt708vmLfvwTRm+PwgefLphkyjNGRdAo9Yytjr0JKV1SlvyO
Rot0wVyf1CyNtwBVs8EEsWcgb7KdQRqFv+6/rFznYnt+DCb5RW1osvF7PR+FvREh
WTnU/gziyIVOBPB9OyXxjvb5Su2x51UkamiOh3fZdIczNqiDju0EI8SMK+RzHc5S
WNcTcJcJHUqmr22fY1PpC4X7auS5d4VxvIkFqdv+3VvbwAsWqIYXaKMtxYrZWw0I
b0zr0X4DAjgHM3fORO1+JiRRtD73ws+qIytDey/+k8kWeQ0tcKkwqZ3MvC0ze3iZ
icexlX2ctjICL9LJpd6S8TUi0oC/3poVDic8umv36BpFwBNiUhDtec31rdlheXGX
JyAJRToqQF7G+4oQmnKpPIMeM/khfHGA8AkqC1yMsYIE4CgH3lYMXJgE2Lb62i3O
9h2aRXMppRJ08tNeYRkvbhIDRRVfod6kVLBtnJE0I4gg0Wu/4r8YEaFtgVXOuSIq
uxASTD8nQAgaIaDP5/veTelHhTuZrs2tE67c+ZeJybcMe1RWtRxZaY4wsDq9sy5l
1jAJtRy5z4hEuhBBNGo+GYx2zP6Tr8kBifQ6iSJsCZ6HzI4wj5di0g+/Emlttu+t
CGUlzldf0PWf67nDQ4pE4o6R9JrFWnpV5EX4WMo8N+NAmY4ruQLl8pKpR1yvP6d2
A2u6I5pDpSwjRflklJxSpGQrDM9u4zp+a85GFA19shQj25cjNBQmWSoIppTJJzWo
2c2HDuSQauswJ34B5ErxH4F/ND+OEFdEvsC8qRXGDDnD7JevMMop7ZVUKvoRMEem
HVdX1EsQUylZwfpqsY4Gwe1V/64yUd5a+sCVHWjVfl9xWADxt6wG/wm9c4rkvpEH
3LyH9VHxzUfoAhd719DrLybLSSjA/1wz6TLxRaxgv5EZhHI6KN07IkakOzGhOBvK
esWnSKf8dcvzxjvlkoUAdpKZ4Je74Oi/U89au68morow8OKT9oApnHlrNM59bKPB
mFii1ZMAy3WnA/udp+nLA+x0ApTq1XUZERZvekRTWXyCEJeiDXK4oZNIt+KhbaWD
nL2EKI2RX+giWDhNGy9OlF52mkbwCacvPiEBqT3OtqySFwK9oQMhxxXgJ9oCEZdB
eLbfhGXHeI2B+M2eVGTLfFp+YsZtskxHkIlkto1eTVWKwhKLh11ZzxwayHUL6KrH
MmIg44bY9aCzhKY/ruLb75OPf4d1DnVdgedL/2jLJERLgZ2jQaGP4EWaKe6qJ8ln
Miqp83ne02wksUaJEV4BVC2g635hZ1f/1odgjOYPvGbwZwRhppc/7FmVDvpw8Pxu
/qA7Z24r0m11oyepB4A/TrrFImGxlXcPo0IwUO+ihKoTP2I8ADIChAkzVRl3irbY
NdKATHjl/KmJgePf6IjaGy9uPpYX60AcWwLWKN3hur/kUIF2RZ9Xl+r/v3qJrd7b
jfZKqG/5eBb1fMiE9VWxyg9MYRaV/Qr4KgPqRkjti+9BiWhNX0ks7xwElzslSvkC
3Wg8YpXtIWL/fHZFgXtIcyU6pnWXEzQmoe0P0sc+BzUNMYO5Zx2KRr8wKv+IvbnU
+p09GRCHukb2fo88r8L5wnBRj40j2F8wXsqzxDSxVHhBXOlndCfm2H/BYGmSllRf
9UF4M0Plwi1ca6cXnS0wxAxfX2WkjjUu1oGxehhdeeMjS+hqspZk0kROuWub8RL/
hIv3I84NPyUhA6ynTlTFj+Fez0JV0WvyskEwCP/HjNLR3mtCa+N2NxAyKaUSYJqC
0eB//3/zeSeW4RuVKWbfXVnsWvloaVVAY0KVv9H82sh1FwFpvtxbjXEMxLyTaeer
NbtrlOabhEA2HIJUPhmOOlq/iVtmulH/c7R4bQJIdNkwGt+TJqVyFtsXqRtRCcX0
bPj6+euwsJmhMJNZDQBDEkXfIvKvT1dj39+Hu3JJY0gAaf8yNHnMftJf0YGFN7bT
y85AZR5B0rMk0wFHWmbd+1kSTjWWsjaSTktGYAnTExzaiHuwZ3R2n/whMX+Tvp3v
2PVTB++vx5oq1r3nvQ6j8tPLmTnlQ1GiEt4tWP8m686Cr577v7veXH+Y/yNhkbig
CUEw7vlXOULXdiqJ/68kn6uK8kN4m6oY85ViTZZJHMugn0iKqRGZ5NyEckw0/u3h
DfzBjFRfnx9WgsSkoSxTUiDdW6cGRf+29K1sushyQzr2EtmtlhTQ3PmkWypToOnC
0IM9l23g61A0MwMakfCVGIOXK7RIHpVSXK6QMIWRZ42+i/lIJDPFGyDhowYUqPMa
s+ibb1YgI4C6L8zUuXSyJoqLBO8jJB0sdOYhEeFIsir4SycBFhF9fKvwJU/Exu9s
NaZc8KJbKIgaLv+fY8VxlWxENXlkF3LgLL23dVzETHEdl3u/0ZcMSawc96In1WHw
TugPJjdHWf1IHCTzdFT7+rMPEgZ/5VUG3d1KawI/sZfAiUDlKwM90aigh1tqL/Ol
sq0Z5B7ssfVuVJXYs7AsrL3qYGXdajY3MOu+LUelI0G5jzTnHFYZnql/Xmuk0SRn
SoAdJ1nK+VstnX+yvqU6l82ieO4MZSOARSqa5auIXgCuATsHefXwRPCHPjCOzRQT
ic9ojajUxLxeQVehmsQFMB9ciNN4//cl0xrO1LBjS5AnCizPKLTvhRKt06J2T7lP
K4PR3iodwNdmANfQqnVPSeBSEgmdmW7VGCvj0cwSKceYSq0oI7T+mt/uwMBV7fGW
CyqtgMoc0I1Bc51/j/fi+M+EyiVc2k36g1eVPq/Ri9YYD+y/dYdRzJYeAU8GOEF8
RjFCSVd5ogxliADSfKTsHrhE40Gh9QK/3TFGK1/qzqDV8Q1mfnZvjULQvCMCZgSJ
xfDJzuc0ztvBZe2fb1wgxSsAqFImYyUCK6s+/h1rFkYSDjBXwyIv1OF0JaR4fUsL
BQU6gd12qUQGamRZVkAH5TJe4nF8W0j8PugG8GHIHKJLvQYyE/g1pKdRHW1Y/7FP
o5DL7iJUtlcTnus4AczWZIUX4koHs0YXQuoDJWvAMv7wJNjf0qtN1oKeCc8kNNRf
EaRDagPNvY8cS5303mEkJbPlL+nNAHONRiZAaEegja9bWpp+dBT/UZBBu4tOHxNH
zYx10OT9ceRDrfa8VZA2xICr7z5s3oqmzbYmTosYYadB2gL5SfozJYXKd1AY2ntF
2cPmip6Ib2iAL69itcC7U7gEDDH6xHiPIVNqjYPaZ+bmzTPw0Oqq2XaFH7c63wLl
Af5XQsKFtSifzA4biAAkUxqtSIR7ROaje7NeS9Z9wm91Igqe87NPVMWiwT9rv5nE
zunDJWT0iUvZ5g58SaDsYSDpfCcKiFMmPExRYMNkK/kz7363RcqZ9h9xuldisUKc
PUi72fAlaURXOO0H89s2o9t05EP2miAXjQJjps6mHJVRL4Qua7pOxE3mmD9s7cPR
Za77+rKVu97gUEL602GXQuA0csT0GbcmCHkPQKtZcADAAga64r4bwrBk64OCyTzm
QKzZwr4jYvmur7CGt8fLVzTEedNCjzH4qe1y1LpD3hCKouRWx2RIJUrDG5bgRHyV
c/NcymqpuJkJO5XkFhFctlDpMVdiC1CHoV9cPvLX4Udc7wtnQ1IewXYonDfKTG5c
+U4LU/d1Y7aMahs1y3AmCNUW89qHl55242gpLno/HN/A48cicvcDmp/yTKO195Mp
EGr51LOc2w9O6BnIHOXfriQ1Ko5ty1Ph1kpVIDgIQYE65VeCOcAp+QLnEOhiLA7S
RneP1mp4ILmQwanWcqfgL9YtZKW4NR3DwblixjxfQE79x0vUIraWpR4+I+JOzUCO
2awWbtA9sIbh7v7bfQxAewQiaGo6OOABF6c3ygCfYje1UwN3R88Knrx867txoVcW
N7iiVswq8mQrzrviJqs5a29c+BhMq9MyMOVhhBd6I4cu7msPg2pnaVtPn2zyGOXO
DRW8wa1weIIyV9RYR60EuK6N1zMjCQdcelhPqNCJgIucYzwQtBGyATZfS3iHkY0i
MdGYxJmtrEKSY8pkAWQ5PRUFLSCalTCkIETfMFWZo7e/+7Oq8u1EpIf4Qtr+xhe2
gOjHSySFmpgQ7XaY+aISdP12+Lr3MQTlcscXlmioDnpbP+P7kA23UeYfc7N4uX9+
zpfa4WvrfUKTk0KqomPXeavZHgAJDCARBihGRFyBqQkPUWgoZeZb5VUJRWH09VfZ
mhdZjcRs0NIUq1gccH8Iac7wcjUwCXQ4nMvHxpT1O+GzBjx7P+tLcaWrP6tdka7n
D6QGpIRzSo3HBg0y/XPcs15oM8bqhx3d9xk4LcLKSpagoGzV6vaS1Lcz0cbLzazQ
cDPX8SG89EPq1pN/FuV/KUODchpT/TUmKvxDYAUHj6CPaKUlznUIMPpEi3DH8dCz
O6cmaHLCTOrSOTD3BSep64RlrxTBIenh9xOkeOwhC4m65A0q3exDgwv8xkwsV+Ib
j0W1MTF17005KIwRSPdQhU9y6fNrNQ1Pk/pence7u5q9cp92uk/C44B9iwqcp+tG
hp9errwbBACuB5lpHgFHdOBQnoFPyvkUSUbNaGsl26qjwXX4DLUYo1DPi7/7vkeI
jwrSjGMecuCjjrrxZOBwYcBqGspezM+gJvK4YpUYOpM7A0wBtx3qVReTcNlCc8nu
5D8kDeovumJ5b1clu1SfVrBeFgF6ddIG8xcE+xWjHF/QexpUcGWqb/0kDVo083NO
wRdP3lAiYbYiS3ypONP7QbwjNe/fTEijT5YHhuWTa7stCJyWR82kEiPDoCiE+rO0
7iAGlJW3FtjsyKEj6x/BJ83HyoSoS3O44XTU8T+7e+ufBg22kS86lPK3JWNaJVUq
wqCBIW5KT+OZSdgXKFjacZXQ+pCOhFS2LIWEna3k8bcwxn04p/6hQGM4MuAGv3j2
/G7wizwz84VR75HrhKAK+QBYrUTMy1uq1PAeZFzQyw9vffznowiShPaaDgIeJCVj
XVWPz2/5s1JaaugwBcMuPalG61T5VlzuAgcC7XspcVtyPL1wqPq9SSnkZNNp48eg
JpVUdWfS3xNlKlMnesYVUIYrEBaGO5k67JJVJ/tHABMpGmXbkIVCKjfkp/RihgmT
hG9eUzW60o3BQwllSY5wEl9wceuVBRXHjavLOT9ewjtlUQRItuP4uhWio7qvL4n7
oBvPpA1HL4WJzKDxUG/ahVPpYEWkCUVsTFk1wefzN0CaXZwRdZH65knUbrxlQD65
twO0oBtrVuiurDHqUCbQHYgTQKYBjHInUrh2DrB0JODki9P0RusdaDqSxDO3HcQy
DBAs4atJ0wqufpKKNF0579xqBzwvPfPRb8Bv2O2kT341FokDzQO13rl0e5VX08gu
NkcH74ZkPqtRAd9jgvS6ZU5aMJHewmXoJwBWYzJPD5YzoTqrFJl2NZhHSBEVfFZq
3vn1bmz8GMb9hTvEgKmViCGNr9X7ty/c/JVz586rrWD7V56Mmhk+mVIWBy8Z3Z2a
SQQOc9pwYM8K/WyLJt+GCBFL6jTekz74uLHzSVgyUq67j6qCLwMJO6RQ5ff3hIjF
y9GbUG4x75JJASZkfrkTSD1srOwZASaGQE4XxONTqfnpNA2GHpZmWbWXIFLHkRts
ldU3+v3dJMzDo0EpMShT1Pq7NoSHzyIXJIxGzwT3dA+YvbGs6+VBFfcZN3jTvY5a
lB8FzJAyK/KD5bewYR6uOxyCwzQFhoRJF2xBjBCHHVNYDPID0I4WpRFhrQr1DFNz
/u8ANjsGvQZigjfXB/AGBY7+7opSXPnn4KCmodwtdtWOateOtYRPTjOB90ow8jJL
E36nItucXR/zQBH39HUc0mE1DlCpyS7b82fZS/vDoLDEGI3M0mlB8BhDKUwGhN6c
G2UmGiMDoVgS9tHoZZyxHo/QWAJL/5eel/eMO37bHeBiORq4i/VdK2+z/d+hga8F
xNV3yNPg7oZWsVZ7G3eL5RNYbKM2hoJCxQrvzyvIaUlCoLm1R5MnYsWIKi0s/ick
gMwKVO4PKF7hIlzUgTQ/GY7TLbiBnVh4Jt2OIX7cFqd1Ynbsj26ycutuGMkX6K+V
xVfKwPEOx1z1LUjJu45oZCUTLxqikPI431x7Pz8WyxfNSYDPURCWOstfq2sOIvf2
5t48aL5mJZQhosQgRxFbz5TpjcNlGxaDDvAifIwkdCZUrrBKRf4yEMfkbV/S3U08
IaEhxVuvXVo+bsdx2u9Kfe57EYK75u2/tC2H0rVJsOi0ZEPN0g0lfIwO/0PdLki0
bgXz7WBQyktZxn2mR340B47HO+jPIHhzNF/pX0OJmHtjfkXmYNR7CCeeeONqrCCP
h1vOtFqTmW3ExaQFTiHNHW6+YX+Ha9YnCzwmxJ8R8h9CBLrHNVy85TojUF4vuuJ1
8OjuoK8opQFPGqM3ehvFJW5tTfOB2G7yAkfR4Bd0QcITUXQ/rDCwu9UEQISaxDRq
2CnLa0FHbbrl2dwbYQ6ymc+AjRV7Oo9PEX1G1p/p0GJZuXyRUUVdVmDhRZk+t8u6
L/gT600ERGSgirfwwROkRj5BBkRsYbVeHjNDg5Bh+ib5ttaXiCv06np2FIzEwhJO
/e0rGWV8EcXVXvLJw5ET8qDN0zMJ9zZ7F/6oJdfbn6bxf9cu3XIQbzce2120AZdb
hjEjmfpDyWE5mtkdS+VQL0NYkvxvKt994wGDCL28UnUSODkoBrgXT/40kA6PaXsX
oXCCs37xL6MTAbQbvr46BqzxYd9JOtAXlQTiijGWMlV7Au8Bxc388Id0GKUmqdtK
oWe+viit/KQ5b17t0Q8+3AxU9iwjQZVfsFsIyFNMMsVgrTg6WolLxreEcqBjaDNw
VlPoaWJm6yAYMja5kyXCyFQKDohJvJ5OnmtWACMveTeIw05hAgf+eZi3YlmGsEY5
Gh+eRkdXjGr0sOUKaz6Hjz6QjpeZ1UHAzww+8Wq5YOAh6rvlKCTUei9t/sgVPAdz
S/I3SpjlETmKZPfx4CA8OtFmmuoOC6rWCYA6Q/tCyyw0/f+orjflBZkmni/CJHtA
95bC+95iZxwKL9LEi+5QjzExaol3+FekO9k0/7+p+4Ic22JxUp6237Si1ssf9UKI
gV6Wd2LVftLoqwVolDXH8QDbGv3dfK9MyL/cIbhl/8/MjLcwV4IiK7EfNoflJmgW
Slv3M6QrFPU88pbwONFcXHts49RdOvhpe4eGfDF7r6YJp08B1N/OLEJm6LROInes
0enqLIwPlPyMkzXdpFXv0vpZKqgQ4SJQF4MKdLn/YTu1kFdFAF7nLiR/8boijyw/
Lw9eb7dcMrVfGhrNgyWhN5VuQY4NavzCbZRFvQQpg8tCbbuWnuLtvr2Iu5Ss3Gff
UdBEcTL3RUWOJzFa56in0N0/PG/NwShmk53o4EL+Bi0Lv3BE8/9WyDXmmbyJEoB2
7oXQCWA/nqEORNY+MFbhDMUnT50KZojIZ4nrmG2KoVAxd9j0d04QhGCc7XLmpDf5
8b1Y7i06V59pHVadS0seeaOs/qiV7UMk+HXtadS1v52L14waCUUldzJYh+pTrBzJ
vxDCxr3dDxr/4dCqxJO8rhqJqP64EOgdYxOGG+7W79vmlmxFhdSP8NbU2FDYM5tK
zouS5Q0lqBElPoJkFUUvFUMyLMsLATDiQG+/XOw91j2uo2HZgD+YlkKJ/EA1cjD7
3AshP4i89G1BqCUFd+O/cteZtgWZIMnwtEN641sAlTKMm82AElJxOWloEsBXKQgB
ZwlvlM2A6mZ4O8haWlShGbUW2X9efZ4//QpGJIwYWqPyQLGfBaslUxqcP6gGlApn
fW0p95MF0SfvCPOQl0wLB7u3gHI9d1ygsHTRGn2lnXZyqlD0wnS2QOqa/5Gjvadv
IJEyoJdo6YDOlV+VBDgpRAeBqPqWojqfzdBJasSqcQ4njvxUtuEKeqFbRjF3W29h
X5zkbOdfbsvFYtK3lxMS0TyaQ50d1IkqBRfO4PKeNTJ5vi0pMtSRQmRYj1N5WccP
AILddsho42amV1nn9znD9u+kJT2NJ4ksvQOUfwf51E/H6N6riBvg1aLGuE8b9nrF
KDxTVRNq6AzcLzlHHo07VaqFOA/zhhZR7M+tw3SHxaq0tVOodfWXTnYRp4OLgSJU
ksFuyZNTm2z8rJ9XPm1u5hhXEpWdIdqIAVMeMu4xA1/dFF0P8WB0UVUzvvbVP29A
4nmHh4WZuD2YoUcA/VmXgb+RIwkhOGE+SwJG8FYPjoapAZTZInLEU27j3Y1c7QK1
+jAt2tMqHMQTFavSUuifkfCZO05cTlDREr79Hna09jQpbuOUbR9q90zgEEDtvVgs
csvuBFV60Yl0rsvK8y+2pCW2L+KQM6dRRjU03saXyaZ0vR5Y2aWuDHcFeh1EjkDZ
UBFrzmBjKK2PXgs4JjT5vIYPPYf5NGIYsjyROWQMKPKECl+mywnE6vW1iIo1SsYd
zA8xDAFYVrKGpvGJOTfAgMBzTW7lmMZLddPoyVX2kPSQ2SURT8nf2FdXuxXBB9DA
prGn/cyBOuqHYCA68uvjEFcGLjk6y/obK60UiRiaBs4poJSsEOHifmSRrFmbYAJ6
IrDWAGqXRpB/ie0r1KLi/7MnG0QeqtzQDOODZd0tdzW/sbI1pVIbB3aQEPZdDYDS
TTN1XPeG+2OKLq2/fEBZpr36TffPSHCzuAgO9qLJ6asaN5nilHVtkq0R5HMnzVcy
kdX18TKXclukuGESIUFKLruLO+g8zi37GaQtnHHh2Z5wVx1vbBbcMMI8Je5J84dJ
+zV2QoDgaGRzjXv+DcOm3JuwsQDD+QIXN8Ppo3iZs07q0hSrFqZroElvG0MTIcMV
k8XDjkDJABkDfCXraphxK+bBnoCykn1RyAwTLuC0DYRiDrMHySu9cNOzw7EWccqI
l0+xgXGD8xgg6RUadOJ2xVOL2Jwcv3PJCtl2hcT21azpTnVEIB+6bQx1rNnKWCPw
kmqS8lzLi959eJFdkad5/qDCPoOf1ThljZaFMBjusozdILdYQjpe6hDuMJxMFRlr
QWEjS/6U77ZIigInlQuzXp4O6qZ26IgWseD2RW7npnPFA2Bz4YB5aV+7/C6n/yv/
FVXGVZ23wE5NlJCd0Y0T3qxC/jbvhBw+b1o00n0abRyWAjtwHAwxyu8jZSlRdS0g
FXGRWZ74EYipJOKP2yvQYjl4CvPRANup2Y1DntRC/kR/2snVeLRE0gsRoeVeYSTO
Xl8GkqCa04yhTPz5z5kzJvx+LI0xlat+Y0jSqlapgMiWTdITgXXt8l09MDZIs77X
hbwieW4i4AzqH4i/l2B6x7xyc2O9mn5xjjP+rN9nj2q7H5W7mb2EG9jgGP5RbLDk
enjkI+TtosmpOxdz0DfkUD4hBQC8Y9nRn2CsFbh0vOVhDUnIgtrcTY3+q8tzJqCP
5VyK8tuXu9q+YhDO5huQLanGjcCh8VWmD+K42obT1bdRk4y9uuIAC7j2s6xGPESM
DPN8xewh4+sqZpFlnkKt+8plNtM2siGrhrLoSEW53XBaVlosGcyNKKvOPPNayT0u
5fB0ABKJPeoaGK7LD2GHROof+jmpivgF+sv8RyTzHlhEzLB+FB502mrR9wTtxl2V
5lf9/Dqeu4zM3Y61dXObzMWQcugf6NnpfjGmYK1EdT8NUbQAkgc8z2PWwlO0T52z
QzsiUttlnyDM34flp6G0+31ohROdZTD3L02SM8q26cS6Zs/IVYVuF/T2nwRCsveR
KwqC+V9Wr3z14G9FNz90AhrmWw8NCdFMaWV7sb51LDpESITlBh95oP1p4UyTmzVl
wkahRgyOWdCsKEJUyY2qvaktkcuZ6W0hBpvt9ab/N/WH6vS8NuDdGakbkZPRB3Lw
lArrlwAZpZD/8yGchZViu+dvclLTDgMeaT83lamIlz3dz3XnNwvmz27CJiguISkS
Mvxw5NhxeCXs0yTNuERuBuuZFK4sKQNgvMtn9c4p7T2z2uKvhJFE4aTfFSqODIKF
MA06pXUsuOerSl347QSOczsK5+7/bMD1jGDGO+GQ732ONGHaRT1S5SwUEXonKZ7L
7UsUKKBuISN/sg8lPJcVSHFAhIvaAYT4jiWHNAuyaKst10+iAN/G11EyRBcz8L7D
lzXu7Zmw3CJARYwehUYPdtAeWC6DISW4bg7rxCeBNijnk1rdPh0v1RJxAEhs9GOA
c/rQRGntD4Kpxlp2YZe5sAtwQdyudHWYbhNm+zv9Gjti0PKdXMNvXLyg6ZKYS0Ig
D0CYoIkPpqwgR6jh7hx9mJMACwu7pXevH2CagXDZ/v2G6+zU0vNZhbnRUY3l5QNb
06UOBQ1GIrOybe5SJpGe5d0PmNpILDZMpxsuSvRA/kvux6b8tHxUWcP6LXbUlZ1k
En84DeWjLp6Rs2BIAPMFr6mLd25y5Rs1EkOWB+EjiI2mwUAfUCQl1TRRxqgnPaUx
/CkOA6MapcmSJ2JW6HwcojSNDxo1Yz8vJj3um9zZ9EjvH9XO0XvS8WINs0G6fiUW
Hcoyis76qAMOO78lJ1lezLo6NFSjFw2dZl5XYmPQXeYPpxnYiOKCHAfZNEbcpurz
WPBwX06j7U0joxbSGnr7Tb4C4U+Vs2hVV1xMCHvbsYee/7XFNCNwQIeRy7jrbji0
vELHQDc85Oaueu/pOKQc0iYyw0AAF15GR+2WGkLLckqwbDVAoBKfGVE80RUS8Qlr
w07b9AUWfaw2qh25F8g701p/zyNwh17zdken4OtpfzzAjQEqV6hm61gCfz3xaUsu
i7jRtv26L4l34cXrrfXliuCa4bM2HIvysiOVo5lJg36cPUmwDPYL2sjvtIiKjUZV
UIYNESK2AgolL8kGK1csGZfpb9RASZR2qN/BFvrxiBU2+6ctSsHroQJUHZL2tUUp
wE6Yp3kjmI721Y8/63S+XKvbC8LVH/+uPYXaKQLoqMgY3cL4cFSwQQ4ndbEDxRhK
utC9xl+dufaFnPWTfYt2Kznx8Xij0Fa0ufWUruNllr8OsdSXxeNq2D9j20FVticV
ciJtrAHXIC+6u8kqCpPN5gr9e1mhzt1WneOR1qPs2P9OiJtz8XRoKynPTDaktsSo
RdIof4AofN3M/VhwMiFP47OH2vqWZueNg9mG9TVi0C4wkn9keyIIVdoaGfs29mPC
xU5kb6bTF0io6QxRd+uN2v1ZGzI4oyy6UUTAoieBCJY/Llvs/UCo1yzwCdgG/Kmh
4hprl+eMaAKnbOxjCQBh9NDrbUfD2ffaHDPK5ymI90zsub1JOH0Sy7LhbcPDhEDg
PSeeNRE8lOZFjgYOP1G4TKbWEwHeYdTRG3O4BTyMyF9soI3KimIoCRtVecOXjTQP
HaSXA1Kwd3PUi9c6hpdXfE8S/3WWPQwVs4fcfecZ2eXrjx9k0WlgZOBp7kumDQtk
Og6DSBhshks48iJIyKtcKxjjraVNnVs/JkJLvjuAT7ne+2u5xHPA2mzTvqk1f+mE
gEOz7liifL/r39mQ3gjhfPNwUwHbANNHen0DkCJ6zM15EHbD6ljI0d+fOoTpP9/P
nQ/5cTxzCYxwV1mz0dLxcRyOSG8rAZnyP+nkD0tshUHsu78SeArY7scXIZftW24I
rYU0xdi+kOTGLVZnyGiY5hV8LPoThskKf2E4bP1mtLjoOd5FKQiB3poxuURndtt1
FfwCEQ7+wxWHuUHK2x1bxC0ASsnIutQsBayZjoTxP6Y3d53hz/OWAkb6zaRdS/nV
qa3Eu0AZ/NjD8mUl39b5RFoDEKw9LcjEbx/50mLv/qGqT7kYo/gALVGCCRqCE2D/
GQYYyc9devR98+ZhFUolhAQtrNu4WqkVMINXvvJrO4Ln58yl6xLkLIQD9FGFf5pw
nU5ct4O3ndILkxQliXfLpOAOGwD0aHpXU3cq2Hkb0DjI/04OJO4oLf9i4ATRzg3U
M3E4UFSGjv8kZED+vuBF609LeMx7vAGqitcBFJkvfn9uYt2O9LSK9SB8zAUtLg0t
1cVQEPpHJMkeueLr+RIt1U/fwCxRRns4VbhVeuDzN7d45D8QZyVhb9nmXWBXuwKT
jCdyASRmGjmjL7TSe7PISb8UN/+z0m7bw5b5xQ9Gw0xtb6//RDrX/lqMaI9SKsR/
Hslqa8AJkYzjpYv2QvEZelHN01MoGWbi4plxC3SYeIrQSnXXZsKwWJWYLAJm3pA+
3nR0+LasGhyTQ7eMQSgq0Nmqa4NDIUf6hhH9tvDuYmwsj2HtWNI7UP3Ide8o424r
EtMhQ2IhOENaYimfz9tJY0hPLmm2/I3BnQhpD9EDmDO7KXmUwpFS2EPpWQ9FGSKT
ljbEr/rvPQbRQooz0VR0+FdKTzkOZrgYgNFW+1q0D9XlVdku+K2AhXairqzBLZVA
kbpq1McelxsVkbJXjZfenmwmDx1crQ7nYvoTaVzEZavKAWTMOTijFLCuD4UiNG9e
UOhI+WWN+Zdfa9ftauFQN63I/LvgCogn/kPM8nb1R5lUyQL/zS08P6UUKstY60eq
x7nALfFJ45YBCRBt8v56PxY/DSosWtS44I5EXKNKd5bURj0qFyald6kdTuVjlr7L
f2UkatB0ANzHlcSlYC5U3cHE2hefSpLYJWZ6JPxyQBianIXgr4kLguAm64W5k84p
X98kZqEpBxp5TWkFAr/2J7g2IADRLcFgcRiThSrQFvu/L8pLvXwYz+/wGY7kL1yT
7eojXaDOx6TnXC1WW6aHABcGETnCBx/13sjnKxX02A3h22+1IkpLWMilFUigQR9V
KqCJcJOrLJVzIr+SSmIvYZrY2y7+RSVExK2o/DtRGK8MD1dkB/2n8gcPUJdmMhkZ
MTDGzDEXqABRJN6PuiftMUvqVjKo04+q/8+adgJx/fd+A0cn8tgsbX7MvkKTJ9pR
ix+8G0aArP3Aqh29LyF05NmzY60ayZfh0KPULRicBwBEys4yzApBhtp6l/Wgyvbc
QtZExbFfQ0xkZbgPkY32gNG2twwbNyBa8L+FAPU9qi/0OA+idHN6k+a1lOYAvFYa
QzsUnJcN5Z4tC33YTq1oVvuwXkq35ubhhUSMXPROZa+J8Th75uK1BhFtHnvB3UhF
H8LkbsPysRkyHOHiPUh601jdTD5Hm4FrD021jaP7DO8BYOcMSRVMwkzi3K74xdMK
KiOvyhaaV9ANDLHRsHNtnDsLZfmCFU+ZQYqhnf9mNdmMd4upeY7fYqdQUUI9wMky
M2+CedwiF9edCRATTBflnpR4l+3fbEJF6iZZ6i710NOnwtczwp52fwU7XkO8EAYw
LppKjjCfZ0S7Ztpmvbzryqx0esZ3e3x4H1Gah7o6XjOMVm9PJYL1zQ4gQSoABj+s
EBrZH+hWAUgHJVgFqlj8ZQaxpSY8wNFfPg50O9SIUgzY923qjmS/7DBzmIva5Ix1
S/462dPqjy1DSthUuslm2cXpL8PUMk1hEEOYpGHCSJNX7P7wcC2c4eOJXMoTZNvK
9IrR3yi2Xs8imPCEfDyaPaPeMpAtEwBb1+qpwRIW/PcBZ8k3Z6KHSo0IY1T8cTgw
KRprMKl2ctcnGYRDpW/oVwc0iy2paiEAB0gg4WDP5oDpEvtEmbX+5T3cNTPVGOAl
boSrV0TrUwtv4jnqnjh+X25wf6gMtFc+0vwhsoMBbOVwIjnlQcN1BGiNtizuF9UL
2/OOnS+mzOhd/edKYGG/VyfMvKTcvDPB5mrYgo3yOyk7BmFH4ETs+WYdcK9TxfLv
xSENn7Wnu8p9DpuUtDaXCEpt/h0jin1cWNP/v36nfGR5vKuu4IH2vRctwzBhXcdt
xzDXuivPBMyBQnIQG7y8M/EaicwiVK+lebAFogvHXcJi6a9MT65I/KHI3jIyg6q+
/wPa1YP6gghio+cQ+SorIsMn3B0Jx/6kkwA6l9Kw0uuoe8TRdOJPUUWpUTiFKtkw
dv+ub/uYeqSgKU0LD3ZLV4FxNfNcyl85sMy40k5MfvJ1BbzlOxQdoIazo650dBR+
xKtDAo0Sz4hXVaatFtLLwFzdQHqw3VqQ8FwZ29HN+lu9K6fBK9TLT8tYVq5HjHyF
c7zRGr9CTgMZxGAhfvW6/K2GpbLMNX+8hihdF00okojKubtpE/El7mRuj3DW0OcR
PPGzGgzF8J201YqnbNPaKIBe/LzXd1PxOTXc9rySeRThrfWYzx+bXjnTc65FAwag
S5gkuUdB6jcs0Jfzys48BXm0twzf7WQdfmaV4P5rjAYupFOYFXq5JNqgjd8FPW78
O9vf1WOtv40dikPHZvspuDqkCwAicuYy23Mrqur4RU9hkiWzLSXtcN77SpUAd803
p4Y6EubcEWFoBsNUS1Tu0v+mMjZgluqiPf413nnR9GGMbKEgk54crcQ6DyyI0J9w
EqHVNeBAKRnKQ+a0Z8KRcUm/8Tp62l+3gIhN4gt3wWfMS1zCp+g2ULrJJ0wzqDpb
zc0Ci2BBqRVnHHpPw5pL+oAK9exjWyqbTD2w1O/oW0FtgvLx8Vo/aoHQZLdXza8P
5UHoLD8QI2f82sT1xrTpKt8VJz2Rw4if/YUcRzK+4EnCFwEMka9hwBacJMihOCU/
rqP/tqYhqDrnUNDPA/0x32XLCk6DnlUwJIIOWukxOninNszxRYvR6kr9CiNybloq
nbYeD+fwVbi3ZO9qROC+2VKzcL4ZU8+gYVZW0xHLN4oQXBpW53pr/G5FSjUPlC75
tTMgI62e0BFPb7/327aV3WheKgThDpv2mniP2DouNZSAoTCNKQ3VxBsv5CJG8CwQ
nacsWgmV3kL7P2aEMQU5QodmoIa9uAfJgDUKIIxVJh0y/fKeWX19EedhBWw7Tb4v
/ECqPzw22TOBvRWcOQWFBQcCpK+MhnSYMU+FKHes8Kcg1t77agZMcgzP1bOGLdtH
6wTZpUKPsTGbnVV0qiQvtQvabZ8kCk3jSGVe25f7rSe2xg4puol+JlJT9t2IaAnG
/fmISFwAK3pnXKlJFyKd6mZ5UUBnmhJxP9pQgnqDIZVQI3X6lAnzhz/VL6eRyTVq
7iGCn5sQmtpvqK9xIC07Dsq1qg3p4Wp7TuQPfFpYG6ZuIsEV2h4zKT9f/veDFb04
gbV+SoLoegoDqeMjS3PzYvg3L7dw1mkzmWWrzEYleDiKBjTLtu8Sy6EHKJFc5CQ5
pueDnjie9XaAo8KX+wxFb8V9Mf/wcT9FM/UO0Pt90H4FggpT6jjo81GxHUQ0sQAG
JhvpI6dFsEnbq+PnG3dac73jgQMdQflCL1220JJTkFWyJglEuxjMtCpqXG0m/LXL
qbLD+5br+wAo1iC+TpgiC8p2fc97OD2b4I8vWSMUhn8CPutZfkZJTdFpD2dmdr+9
4pAmk9HgPPSo68y9urY+MdhqMPInPj+fF0HvoJOMVSmAIDO5K1KI/LArcqFTl1/J
eqyeYQH4Ys+cYL+ulDflHTqGFN+CLs6Rlcx3J3Z+nCrpKNvRxIDjYiGdhfwo/axa
tBZXOLjdm3hoPtyPsCTC84bHFa941JGia3xBesiQmy+hbWcmKC16S/+DbvY67qMU
M03+3HgOoRQjsKdEuB+w190VTX42hfNURyygIeUh8xOGHcbc1n6Ioq8T+FWyktFW
Ek0r1USs9nByxJEi7yetKSZz94jC8OCD9cliLn/8L/9cd+A196dyvBbRjXe7xVGn
79DSQ4PV1LXVr4V18z2Yx6hWAHHKJVH3xRF3yZ7GjXOP0EdgEbtI8fI5NX8DWgvV
lDFlcJv1bEh8tX5D2zG33v5UsHV3IdSo2oOhe+wpQqPetUEhrlv/Uq0Hw3sVLzdh
apz47yYx6FXaqYThOueYU1WTF3OCkOECJ4ttB+Ir4Pfe1w9Uqv6MJMhsBGYVD3ar
eCIbdNJbWNBfwSdkVpiKpZVvsTP3utRQKGwh3tgK8KbLGDjqSYLvmgnG0gryNuxj
dZCYFlX4AGFva2J9iRyyr8fWuqtGS298AHdpbwvKbAzoUwL4V2LyU7jHmPioc77g
/pko6aWQ4gkn7TcxnI9XWWBkJumqBkP4sNQR2dw/By1mPtFQxa3UAG2Hl522+eJF
6e2vklEclXiRefWakRq0MxEDLEc6T+Hd6dLeh4ltayEfaFrLQ6vJT0QztbG9ZSzt
kgkwitGzgOHiVDiEa6hTjODBm2YQ9ydVi5Ugrkgc7V+BKzq1KWVD7KW1tFUf5Fb0
HQgh0mlvT2zamKnWfPfGP9rXKXWeq/WgmchQhUhx5HDG3fs2UnazVC7CHerjL4Lz
yRCHTZcS4xMJDHehLTVI4kqLwSEDl7vFr44Y8IsaIxoFt7jBdPUpN4DMWjh/9q4P
ECq3k4uRnqhtzyH2HAwoypzCXI+VOMTwaJDsymbUNtzyKr1Y4gVHFhcvK6mXFP5q
qLuk42H/j2y/Ugkr70/r9gL/ZbVHaxL7bZ9cJa7s+dqtd6wc5A1VQlA9bFW6Y+sx
B8670KmfyqG7m59GSJc+C/yCJwMqTgQIdUdffY+GZZNRESM4Z/xVF8m3grJGs5Em
+H7Q8qS+DHX8UPI9ph6fBvaWMjUoD/kDLGsj9aJ99kzzgD5pC2sZYQ5rlQpbow+C
nP4ZLtsXtZ7237DKMHDlg1Xy+mBmDKhgaAN2q0pvGWfiqdQ41xQWFpNohS1PIeNm
E+dKW6bp3ZVkSJoB8BbbpZMC2L59DxM9eZJ01FXQsEkka6IORqfLiRpD+mcVMF6s
XmZdhCG3qq8vinq/HiEKC77HKJXUR1xUGhj3WK71v2znAtFtCLEwJQtiOMfX/c+K
OBE47HudCeghyawfB2ss570NHv9e+7yPb6IyOVsFwUF6x1wvHHD7gPCiiXfrlnWK
6KLef+NBfpFKrHmRouy7pNgqa1n5kDmJYPQVW0jxZkiOeBr5q9LtrhavF69KaZrM
0cSPtsTkIesJGVztSlc//XcsyufWsu1JNxGMQY4gm7yYT6eX0oTIUHlzmk/j1kh7
kKbpelJmWSbuMfSPj5d6cowialDtjb7C8LPUwaDvsr1IrRDGsFpupfeOhf/736ch
IfFzRJ8DISYnqGRCDohQtuDGDHia9tRbg4XRJB7d8H1iq8YIdpHVwL1Jrs8n9iBk
Ms3Cc1yc/M7PtVEDeP5wNGSqEVFMec5rRabN10MwPhXqMprQasxFwJZWtehU6I5Y
LF6K0Dd+NuWYgo+ZdDfYOZJis5gI8xF0MAamgAB3mL7Y23uSUWfTHg1wGAtXwvXs
SnRJDXbkTSW//+P+B31p+UtoHFqZyaxNIfI2rOKTkyMr1wRj/wRS8ijw2nJDObaP
wGP9ZLwJBc1hhNulccUroa6Z+aGa3M6/6zSObkIpG8QOC3YYIR4V34A8RIABVJ5d
hjsjWNs0QK5rnJapVI5kB1bBtrHQLJJiCTzgO3IE1MCRkhZWNeVqbL34lmFHuOFm
K/5rCwcy6RwkWQ+ZFS/Cu21aAoHM0IcGpD/QxeNbaCCkYFKmUDMOJklLUSRakWIE
MIPwp/iqP3wdnRrYbsbCDQMLarFCTcnUYFnMe/DfMnl6uvOWhloZ6oQYzHUynvha
Z4ZPLTlhtjQXc93SRnSfaiQ5l8yE6HtIsOoaKBQOFF1ca/NWFwpDzfdP0c33cwc/
Mp60wyXyzOExRDM9OdgFYQDlu40eIZwGPEboZJA+XqtifUFKnoBq9ENGbeC40hER
DsS1PskvXvd69NRYHQT5pA9F8W7sHyMOdho2G/aqysQBpt/r/e4jlAwdp0LIAHzx
WlisKdg5TWs3eDnLF5vaZD/5ToipEVxf3jTZ4K24dZX4BeAIbD/G+2ajekQNMXWI
ObLFL4KnxJFvBxHBTtFqZbdz52El7ArSRKrvx5lZBboJsnYtk+Hwadl5P+jWdUFl
9e8Eu5QbkJ6O0lH1Kp2xxd9j8gSyR2ay/feL698pu9B9djGRUIuHa7A1tBctuCoS
ikffUtgs49lZCJAYLgmvmKj8LKezTMa4m3nbOVTlxXnyoPiXPOi8VfttQO5Uph8m
2HS3+HQ6uoRH/XbxL3eCm8LZ/+sPUD3tZqQSvJ5Fezb2xk/2buLBe/u10f5nF6QZ
zB7UfZBPwJUOoJZfcXUYTPqGUA3npQ0phhMkP3sSbLDV8gjMPaGmHRMsC0cP5P75
I+1zzeKXIDGmUTBqF6Y52JQHoCDP97/61zoZpBtq6VWa2GVURsjCnc+KLJAl6bnO
lrs9OcwhnKHHVL99I6I3V4hDV9cpfPjRrzxyAqpjGJmOc10SMKIi7VvuUAiNhrsd
jo94UmwPPmdqX2cXdg+HLMCRQwx88k0ATaXGjxRCldh+n/Icz7JvXj7iK4rR4+X0
59oHvyL12+CxnMCzAgtwGJPUz9SCWF0udg0C3c+n23JDJbXOqlq8hOPqa0Q0oE72
GltqQ5CiQMKPTj1z2Angr7QZbbijWF3tJ2M7ch71yn1TWdM9ykJjp67axd6K1E6q
Fz4wJUwo5t0dZwBE4y0p1d3T0rqXtN395wcEWyD+TkRPXrlqA3sJ9iVsqYlg+MCR
8StIZ1491gto0yIJ34/yjvPw9L9MZmM0Kv9pGkBbPTFc17HUBIMIn6h0DbzqEzpl
ytn4w8RjPUu2Gi6nWdtSDavoGNogfzHKIDoqxOVCmw48nTn0i4R52/ybPWYKB7gv
yWciuIfILlso7etwGwKSpNAUuKaAMu6Otg4W+BanpQSgcGa+GJUvrMAAXBqaLc7M
hf4H2cYCCYAGx5FWnnGyjhfBPNldYwGnDofXULE25Sc64P6E4xdjIJH78fatGDZN
xmZJoQbBAkEsiNM/KoFFD6CcHMIbxztQnGrmaRI2qRWgQSZi3p9Z6TTHVc/LI+Gp
TU/dFdhmWqNJZePQLNPuMYhGZWi+8++1s6hVscSInbjT8RSqNqes7XBNoxcROi3s
Ottpx2UG0bCTOVTXwUBmQhHme4srtuLn9Yu5TE0QSxXzp+KEHprfm1SvsyT0ToMT
f8yI+mSqW7Tt9UGVjWvWuzsNnW+lcpzJopmYZfddA5Q+MVtx9930W3AtPxgaG5s4
YTYM2SJBtbg7+xT150Bh+t6pcSa9mhnfYkK68CqJ2R3scP3yiPyxhF5eKTtYFmS5
ZJGEddg6iVIfxrC1t1cyhjrpbAlcJWtLEBj5y6jFYt45qcXNDXNKTy4EcrGtPX2i
v/RDat+DmGfg1Lb1MWW73fhdOxkjAC89wm4vQQiTOML3k/w+Q46SHIrB/XVnbipj
wsqOcFeFaGVMHOb1UzmG+ph9p3nKfSMmpbQbQ+n0f8M+ynbr+pAzfdhui9JK8TWg
voFNL/vV9WUI6oOFLahq7LKjjF/635dhD3A6oS2lfvhfGwYslEiU8LyAeL72e92i
XD7Mj349XlTZWH5d+nM2nx1/FL0VZOWa2Hq61HemLF+PN0OawcOqfB1xMwV41hYj
Ya1e8z8tMa/nC/0uMODwNagT2ZstpbiGLQK9up93MkmlcutictzGjLfNT/StrPwE
ZmU5Ul3hfEaIKs+2/Jer5KlMJpmMN/GAMwJ+/caBjzE5y+0t7azS9SU3hl2CPwrI
gDnNQy3GPtiJ5zeC0CnWfUZwZ74UBXTGfgtEdREnvl/ifLf2m21jiyUHGcwCbTSJ
sbWOq+6W3UiawdOYFJzr9iRB4ol/yUYWq6QMmE5/WGWjhsxfthzrkrBFXZzF3GKT
Fl8BKJQYL49x6ZeZWiurrHl63Lz1iLKiWlD2vCH/XNk0VSAjGnkrwR3569qID0gQ
sHVRtCUmhlOeH/l//OsMuu+josmwbTEjFTY2X2lsFpbLa+iCc/7VOgLa5Qlk38X2
6AnpHY1M10Ub++3auR6Q9Azj2NQC0vLgzHkphk3Fp7+hQQjGHr9uitcBipBrnP7D
KNj41/W8brH+yPW6bgpiLIBkJZiaSzigi2luU9eEo4tn7YYTriHmr6pSXlQwrSEM
A8oXm4c1th8Iyex5HsewK19kbmK8XjG1HTuQ0z7tpigmfI0qEQRST5qHsmYJ07EA
C1GqtRdD1C+YA7V5AHtku0jujTtb6wuU+ILZQZ0e06IJNQWEyVt6d7oxx4Fb8bUA
kZ2QRtczEz2oElWNeo0Xh7W2oz2aEZXOQTCDOaRhZg1vTUZl2fw4MZc7o37DxFWB
8HtmdCrqH5KN+TEbGccwhw/cCPgA8SpPFvEJUYNrC9rSSCva2wB+6t7utcNKB5aq
NS/zZw7UgkjDxrCR0St3hgkxyInAGsxcjb8zdjnCqrVJ7zSw5ngch6ChwtDcF2M4
QJmpdAG5LI1taRkXwuU9IBZvOAroGWp1Mrng4hchkNqjG3qxWEx5LxnDoRf0KZ1N
Xcqh+0+DS84h7r6WIb8B8pILFt9x/2huZ9a6/de2P7X35+D7VpbCgV30UXs79oDy
VJ+mHRXI5t2uPtd5eJmIFeEUCx0WrlMVQyGC38J05cnln4DtuY+igx/x4EHuAgCA
21MGD3R85duqTXNcolD3R18br1Ve0B61nZ4Z1Xc3q733wkqlPHi0bgediOzZGC8a
CRhPioN7E/LgoqSO5xBCV8Uq+wJDvASeqzO6wpyxoWSpD4mNJ2+/ZtKJyjuVY7HB
1PBVkCUFs/DY0ir9nvwEsRm22WEdrphT6rzvnChbX32KLEzH9yWxSW939kGFda2u
vQDBQ1iRJYB/MkKv2neB3y1s/OJNBgkjI9LkSwZd+Du6z6o2uGq3yHtQg/PZJV4F
TowQJOGLDouJHNQaMZI1Mat9AXnXDce6Ns4ftJs/YNlWaOqYpOkHqHo2uS5t7l8X
Q50/6PPCLkaOH78ltW+x7bjIRccettr4wJfoe5KP8MmCsBVULPZ7kIiLVjPbLHFj
PBK1Xi3FkuoOhEwL7JzV3+v0pixwQsHYvOaVZUjmaMYj0kTZ4wcx1LvD/PmOWdQJ
C/OurJelxDLhcSAu3d6ermz6RBnBstrS2M0I9lDpYbHGAlsrVbGWUgDO4KoD8lJI
mkDJuw2B/B3rdT/MwcdNVUZwTTmZjFCicN7xFvKr6+nDhPgx03DZpOWq971PtOuP
WvnNU5joQ1LoiOIrs92IQnfPRJ+K2V3L61jY5t4OiWtDDnytiDJwuSeDW8gYf1Ji
8vyqabco9Yihh3dA4c/Il6V96iYunHNjCkbKiy+o51oB73NZ/eHqad7mDnmbLN5e
mUuck3Ue/xoLSEnqcsmrMkCLI2m1NmbHK4fXcAmkbPRQKBmQyf1Hg8i9hPp78JG+
bvDe0dot1mlJjFbsUfrnwynXYUgUggW5N78NctBAUbW8OQwngK44BuUchTcUEB0O
gU4TR58ruzlUQQo/dY+WXaEpfUF18gHn6tFLZmoL8dhKNl+sxp4Xkk0zd/PyRRWC
56ZNZua9E9LZ0PMQnr2AceHTOyyLKYuZnKkpwOVL6dJznzENWpVD7JR9j7Nrx9QM
MNLHfvUn7W9vQqXdPROK06dg9jvEnVZttNTJd7sqzA+r8PR5oBJMIrvSweYuWmMo
kGuBgnrTzkevUsy4S3d3OWuNuu+sU7Ej+FqH26o+gHetLanpha7oy6+ugSjN2CJ2
t7hihk2Ni/yengFRQtA0ZCVMCrQ0D6UkV26htcWrM1PjgnQJqcdRRuRRfdIOSgaT
OsAXOLFpX/bx2UZ3cZfhWtb1SaIUoON/8RwToVsNx9ATcbnB9IKmYgijvp6GGPeq
XHcrvHkHTrKOWvVHtR0/8NYwZgKaH1FXvAsNuIDgS/qP/CKxX0TRBYoaTxmrEogC
Ar6OYU1v4ftkwFofdN3Xpyd1IeXKmX6CgRJ4vsvoBQXwyu18yMSykrtlWuXhezxt
vdwxj5qvdCfVklBivhLhM46mb+9OYWj/BfTBp3O6n9JnsDqgyf9qUMAL8NGofuvH
wLC7+upvZYT/OeQOIVML/YxDFSauLmQd61r02ZKtokHvSIpRGqbnZOXb6+fBWZiK
fH9hiAqlv6AcQXm+dFfQw3zd3oFQ3hdamBNJU7IKb6AZEc0cDzJG9Ecxdw7wddWo
S9rHMmE4pMohRTI6DckRp9rU67HgDZ6X9izS1/o+mcM6GrbRGI1CPp9AY288Xn+x
TPXj0Ym/+GEcnJLT293N9mEKqRtkdjG09ZzdrSIb/oJ31b1Re8i5ko8OZgXL9n7E
njO0UnMqrb2OfPt4MNo+oX/tWWzBCq5jJ3n4/KD2GIaNaXsPcT+xrugnu2jpdK9H
qXg5/e56Bh/T/tMeEHgWTXknBMzKhoB5jxkZdawJPSzTeC312Ju05U7UZEbQnrH0
qZFrA938qcIIey+PI9POfO4yin3TVs8VDLvRvh4TVcYtcsDOL/pwwYDOOFDhkr+w
4od/LXdqVQommiTCxiZixz9nLcNFfSCDWeuc8bHe5XLnk9pWHfyO6b434fJT+YgF
CcaxRnzZEsMacuf+NkiyKkOp5MWjd6DJTxhwZWIAJc1VMFkgO+1l4shQ6ffDrRxy
z4MPfKBfoUcjB1vIizcI9B2ojQjT4Pf3yFZVMhpNzSu5so3MRAvD1a4r8ucinyxx
UAn89/eVMHWwicEc7qg5E5QZLVT6cU9dbTvj5N5cpFBCHlWMoLubNYJSQ5xm0/lv
unGI8ZPx4U+S3apJxDw1N84t44xqX7NhAPfpJ2fRy+sHD8VWQm94qNW5YHDSCjC6
WkluDcYulKWK0ChPwz6VHcwSA4bAQ178CiOt11sL2p+j7kkXXcDwli4OUHZkKV9y
xDruqr7tjxSO5t5HFOZ0cocTp31ZyMplfvM6HGKMzng8J8zxDNFfPLe78x+Bos7n
0GkFpO/FSiN07ZeBG6+1gdlh+whmvsrR+i61tAW7RI1T52DPUPtd9Eo/JkqFyiAY
OcN49dmTi21320Z++iq8OQRqeCIhODZXdq/KDAOSU3Hd0UxYJltcfKFt3insIQZP
xfKLwtQg9yb8WWNRummA4sqWCwVmxOvFCWTsxoLiB1KyduEVwK4cH63FgWD3oDhd
eHAYbg+SgxNoZrAbDLogmHG+CV1sLu67IxXCOIVuhrefX836+I4XWW3zs4i6OiU4
xyrcFCv2v1CwpEmyEHciKAGVMrHsLomO4Iyv+RnUIz+f18tXxf6lANpbygmymQ3i
u8PjN8URfy8XXsqdUZPcSF5sMzkChty5j0vTADjU47Tnu9P5bIgcfaclDTCsPhQ4
96e4fz94J0Xj4hG+xASPxsVJl8s8IK3po+A/f6vScgmotIqhyvRsibiI6gdsXSDQ
uj6BUbVgL/MyMVoWFZw9GoRTv9SpmgbiCpfQCR/DeYDoYopYACry4Y/3DLdRqt5p
Q33E7COPxAn73VAV8KXHQqgaeHnwQQOUYfI4nX2LyJOTxpAH4184nAErqx/w2eEP
76T9ifS+Xpxw7S1E2tkHOezrlZvaMWmPfwFSHpLZtcKA1NKN2A11JhpIjfnNrB/T
y+VqudckiNL3ZPf7QQDGy+sleeKlZ7TjR4q01j9+evILsdf/g15HYLN4zFQbfwuw
5xVng2aj9sWFOLLT9HrrPU+gwv6iaDMktPx+UuYFispgdTulzyIv3XUHRecaK13I
oQHQ9rli3DKjKRb3KwMuVWjb7InXA1XY3gI8xws+pkSXtziwtO6EWQX+4k8+Ksax
aGzpcgan0fcBopvzAYJOFT6r2jsEIROJ34Zfh5f3eh/r2DYpysUnwNKt32uzzHGA
y6pEUtCRSrjvLE9zS/sun+/KcUIBaCVkRrlFCM9XAPR7Cgb8ujF3HSn4KQt1JsVO
3AtSg4e9s15+KT6ej1C9bs0JHkD46MgNkAeAOAKDKGYmfYu0rY+fn95HeKRllD1F
YDBI4m1XkgONfI9PKvkuEQSLnuGiQkpSdWh7BNEDI5OEKyme9FEzSv1zlY1H4qDg
u1P6bI2nbq5hcplgKRMhh80qhdyKhuMtNxrny5BCLH5ZUSX4v3BRraQNzhNUfuo3
0RHgFIswmaOxpaH5m0O+vuecl+0rjL3gjSthmLO4ekrbgRIBbtiuKqobGyB414FM
+amoprTS3onTBIXo21WNDOzxxecMFK6zm3DVEcru+2FzUOG1akR33MxuU5skCR8P
CbWzakjSav16wOEfBsXgVoS5LAe7UpaWzDnB0YUIqLBBUetga1UnNK5+Rs1Zvv0m
jx1S3O5ar1l6zaH4EhkbKVo637R3BPY35XstHBhntYTfGaO9K3gV/C+SWfvLOAcI
NZy39XhHV6/YQIyxO/rI6FkhZeJrNYPA/+Ah4ay+P/XQcp0yQUSx3Nb5ikwIQm2Z
5AZmB+fjowalyfGmwu+dYrq74iANmZQ7Jw2o/i6t9B20hd4tXGMlYsH6VgBbeWw2
mOT54TI4KqzY1TMU3Sch6+taeEbA3mhAUWtENacJTfVQlj0kBvdgPyt2ncIUIUfG
MtM3pNJ9yeUSPPU2kk5ueF5cpLRN8Jc9BPPXLGQYqeGlaoXTWs3akg1Y4lGsyw1M
uMmqMTht026+Cm8pylEluWStuM+rVVIeBT/L6/cdHFMl84LqRV6RUTxOYiRW6awh
BtwKBYInMGzl5HLcrBu/hxQDGjAQcYbpOihdGxz1MGxZxu4oarnVN6LJO3b96gDl
GNC24JJPjA4p0OoiFNuH1/rRqXyJhYbDXquqg1siDxJIx7wjdo6JgokcNdMq3wTG
4cKo7Mo1t6qQcmtcz//aGYgzTW9l+s2r+PfLq7VphjMpiNTR2b/aKlAWRegs9HQw
oJpU3iNFLoi73qIm8+yR0NqzSjZDb72XTCSYjVKTUkdTQkdHOucHU1ZqVpg8VM2/
KfwQqtnO0qzvVk2iNyv31RURq4zAY+ESXWXiGMzxR5LE6qNZnf+HVM25AOov8W6j
bYck/NBIe8hJw7VPekk5+5UfCDvLwxpuJB9SHQUfL7ipd+Hy3mdNRfK6fZql0cbR
W0iDQ31dmUhp4bNUjxyGCylzwSNFLml6Cj64v2pjsX/w7x7/U8AE8NQ6WLtJOb3Z
BAKhMSFwyLv7otIgqsUyYGGLLPeBvdmqnjxR9qT72Mm3pvNpjEHRUPcJjUt1CqbC
w82fM3Cc8LrZ9JVd3F1I4gPF8eku8ARHegWsGESi38RuO1ajJo4LwQDDKBTYlBz+
H9XtFDHa5aTtTK9K4hYProDvi9ikPF3FxJpvykOuXf+QdVHnVwDVvd6HSHyb9EUn
rR2f2cWU7dkrh4vFZkpNHtfW2JZ7oZNT/OOhOM6ZrgHM8vusnvHkPJZJItB6UxWO
C6Ej66M9ntXzMyeQ+qH9A0RsxIN8NJDAiN4oVET8bIl7ybi+SXrgqy8sztUyoiTZ
iLDKi7xYisFgYilny7zKv/01tE2p/Nx8lCu30zoIGZldrw3ngkra6jKj1nbBwdYJ
Zl5IO5jc5FAGN1sQBGOmSCWtSQdOAs6vYVO+0mUz4oHIfJYE2ywVMnaSpOdZtov7
lGi6x38IMomMhADDPFzz10N6a+Qh9FXyyFYxKT43PQzaILOtSBLCb2ttT14XmD4l
j7ISB7R6qxG+3VOl7ZuWVd9EGX8rJg3Jp8YUN7llTqgy7tktJxi5oa5Xt1Lf9J3P
HrG+Bzs8te5EwYctJ44Swsv8ACXAZQE2nuyzFkNXKjNLOW4yvxhrAH6lDUYbKiCQ
wIFtwwn+t7Vid7R/qTKarEXg4izeyZ13F3sx+FEBotL+iMlArICzVqUxpLQgpukC
sLm7YKMDoqhhgwNdB8W1v7xgCkxoUvRAQZlkREbwgCHOfPG3GTE9/i12/rdxs/o3
b0KrRgw858HPPxdgPIgu7Vn0aj541867peLQVHEZJV/yFNthVQMOTsG5R46UebjB
ad1NbFrGNN8ZnFt6RzeVPEim4dJHiCMFJJLVTkJPGCqcys8G3G1y/+I7n2tYeLtj
S7qKPZ8/oFiqIso6cmaNKji7NFVALZwHOnR93s+di5KomB1iyZ673sPeGv28A/dh
+igeP8AJs8njvLvRgL23YsBcZkpbQszkKlk5ZOX1NXOlLopKU5ijQww0sEatChql
xTt3khBL4sDRZ7wQ+AiinJpWEb5wqQo83MjAIHtvCAOm996aQhMtWY95vvLpKTMB
2Mq6UhtPwDFtWu3dd3BkzfiEx6k1npqD9s8ua5B7m1mxF2z0DU+QMERGYL5917pF
BRQafb/4NWuQVCyb1lCh2QfZZ2CmAtyf/dSESCLg4i+k3/XsDTz+gq0dHX/g98Mi
oWN8Bkfo6K1peOXxE67jlVCGriJtgCx5lpwYOlhTybGrFFHDwGh4+jZ5p0CR4oVp
evN1HJdlmrWF6EuoDr/pux3tUTcUUfsijG+8K568YWN9kQwbQ6a+RdCbX4XaBDxd
55PZkS0132cS3h6NHiortlfzKS1W/k/yrhVaEcTHIIvjDm+0jUr/TO+QLU4GfgZH
su5zRvk6vy46gLbRIF6bVYdg+8Xdn3bg5Tzyi5tm5jWTuDNZT38UulDfBnAjRngN
+lR507E5cjrK89l0zFK1UmTHSwQhJDn/eCv4CI9eP0j0OqqX7+yNrTvS+OSUQZSv
J3m8lpZM2i8ggdySKTROTQx938mxAqgeAuJU1Ar5FSIRRNJBl0d41K+LJSdzh2PQ
qt+ChsgBQbd28jitM2X4FP4o1pxtPbF/EHa+6Hq4y2IVNvg5VrDMZhibwxw914yD
XEhNo18scOCIkzoEErciLvwKSAmDd6yIOLzHbFdyscRCno4BIi85+MPyhkPg21w8
fd6ZEF2gpaOKS0l+bE06cXk37aE9dgL20aPimSuKsIx6Ad9ENLAhoXWxelbOkUBE
CpKXianc20dcpPhOr8SXYy4owiaxvdE6wR2LL/HadVN/liVm9fQ/tw0reVCuicbA
h9RqH7kG2Z7UB4jq4RAD+hc41I/fbjqk3T6BIYQa3asKlWywCq4eUAOhxwFgqfaZ
nu6OYNq8ua1SHjGKUOsDBPlYC55uW0uuCz8M3qGQ+xCQH7SJAu72oH7j4KN6bjJX
egH7gfM+3+WG2jVk+uG7YFa+FWkBX0S32qhi1UoAOxU8kFF1ePULi8ilso7s6sZp
v3cWX8mIvU9BiUWFQFGZFUQLg47AxvdHUPEMpLrnmDrOzEITblnAn3uQYPwwGXtH
lmwSHe87+Le5fCe1962n8aLzxwP7C38vpr+sx4UtKl8HYpdEfLvyVfzB+RqSmmYN
R/zQ9+F6TbsfsPxYHtHuSq9LBdEornLuhlFoARbCKilMOZhOFELCL4RM9d2YTI5Z
cDb8NU375WrjXG0SB6UQ3l2zrflaWhz8C0hOpe2/QqtoeCg8MhT913hHDY7Qmi+W
tVius4cYj5bE6UJ2NkKZ0gY1iTikn8snJb5FcQeRN4xN+VhjNnMhTCXyKVv3T7u/
URrJ6Lv2fl1RrzGVeTClaa3v51ESW9apl5B4Oquz9J3PUkHshVGVZ2IStLHxsLmP
vPv90KRYOjS+kdVD0fPXKCJ43k/XaaQyNLXu+RUNxGYBj/xieZx4jHEeXomep2q7
Vvt3wnYOjHnGiE31eUUv7qi29nkMouVCfGXmW8+2WLkV3vFl6jzyyQj3pxDrWXdz
yi+B9Yc6qOKt/fPYqcza2rGgLeFx4+eQCGensIRSUODRxN+IwmvoFVdKeta4+w/3
i/7gp2w3c6hbACsef1+TN+djfiRsoStJM9mUdWtQBcVRKZWTtwrtYVdb/XEh53Jw
vsnyzl8TGoNC2H5YXLyNaHU2fKnC0bWAsU37kiQJ7NzJEACaAxjF0A8nYq56yJ3+
GCwzpb5HMh+/r2IaXyEbyRsb2pX+t9ePGJ2IE2sHJ6uj37cpAzLoLYshIzPYDkez
TIdU2mwGxpoQ9ZKAsv40dopL56sqw9+Wqh27QNYefTKRFVzjHaNA/zsZfvuN46BL
wn0uA6uiZ21AZChNwv30VZq3rbY6stKhmeqa1vEwI0KaLU2dPA4zrmUA2thdEUcj
50/jeBQBjZKvrVhslYqZQ8S0DUZaadAHwYOW4euVdU0ZH+hmTE1HM1kgto4fVCt5
a5fU9PG117YaiRpPmSUtNhGZRHPfoONuAPK1kIBlrRsUerztIeoCbtRWwqIG0nfc
N6crUDxy4sWHhIlx0UnT9lp0pIEfp5061onD2zefJmW1ysOyIPYQZf+KeGpgs6lT
y/wKOOyMMbyFtJ39SbF2AJT24JcWftj9bBou85juCGWjjKkOV7Qo4LPapanEFrJa
5n7BhZIKsCJ+Rf7msRvCTE1t6Lg77dr6cCVkSlpoa1rb9CTWw1mU3lPeq2ZywzYz
5IBHC4CQSp3yTd4KH3rO+HneuXrbe+RQgVlnX5+tJUUs1q+OMgp/NgfcsYrbkB2a
nx4rIBvoj0zw/t69OTFaytmWJjlQ2Kx1e2csrOJ/stodem0AItM6hE6i8Iir0yMm
CdTboMKMYhcRLOIulrP+TOqahyhEwerIyxuCyVfW9HeWOL1/WMceANR5nKi7hnr7
CCZLSDmxCjosTDNBrOrzoW2Lou0DHcezXI9X2uuSV+0N8hoDE0IugnxwXZ+b8xF3
3PBVCkLWWzXAZLDJn/IhEW0+FQBnQLjwMQDhGV1xEojGP1FeYl+Vh4OTyCAq3rYF
0lJT9MiL8TpHjMXdH8mnMBgC4WIgZ8t87Qx/F1xV9uuZHcO559iYfG3tGSPlt//X
VpZ813IuV4C1BX/T8KLXISxFhT9NPUhDXRTmlpm30RTz/l2+ykTVLzMn7PIiEJAM
qcFJsCUcxDdJFeA0W4EaJbAZfx5LnV/6pHSAk1Jk+MtmCCJixwvnS4flsToKSfCW
qyrsPp72A72vS+yJM5pfHfRyjpL9sGIE9D2781I9UbG7w9eAAkXJq5pX05f7zcRU
9Fmth3A+ZvYLgAsjcY/uGbzmeThit5fJ9p5E9mcpj+ughwje4Yz1HdedMetKnhOl
TG8ye6CQoxKaIdwvtCviBNb1vHfapHgt+neym3i0ihWDDKYOUf2qVPEjOEZuaSer
9dWLg+vI5smId3dvkI9tpVnOLylTpHCS93gzemZWG6MTsMCLvG2pEXKSPmT6zGEU
BOa1NjsjTOfrCkAXK5sF6bLdFUKfMl2mSyGiUSu2IOrzc+382pwn2Z7J/DD9CpjG
RYSyAW6H3z7U4//oRj+U8ZrbfpO0aTRI1jmVYL88Relx12enc/zTiK5mAdjrR2DD
VLD8QX4ymqATCilx2zuJXPCtuzNSsCPLbRWT1o0387nosVGD+mAg877U+SKoG0xR
ShlpHUjzxWWp/HwaH4Hd2REfv/uazSCeR7s4pDyAG77e7KGLUznagca4IwCYAcxA
S2ViIYOl4Uv8rPfajsf81Ew14dTO+lfGRNTjnkgSNScYRmw6hkYI7BBeb60MZBY3
Fwpzi3JukIrpT+pPimrUO+MUas6s4sMSVqtuZN2E86oPu5ecTGja/EPww5EOBGXg
Cy3we7QJ9RT6JAq1q2stPRyauHR0Ckumwz6dnia6Ag5H0FTZIHrBA4+XP3zqy+0T
5eFY7WaV6nEznJIx4NolFIwPvOwWO7K/xUBPGWW1q9L92XVqPBNQTkm8PfbdGZFm
41KcvyU8Ta0j4dmANELbuKeQlDl2ttu0ITYHBH/ySKDU9rM4WqeD0s3IW/1HvXoH
KsT4cAn4MDjx5GbUKHw6EWpD6T6h3SfqCWL+nVqXxermMPOhlqfLYQuX9mlqGW8i
et5VH92p6DIjhy1wJO1Fgrr8BfOXBkdFwV4i9IsdBLQj6hez0GFs1hTndkGH4YTm
09Nufylu5wiMZQJfYOQEkCwWMs62AV3UT1XWMdCO8Y1v4FEBoNASrnKpL8G24Dot
8RLqLAOIj7rP9UYwm+QO2XDf+mirtemTr7IpVH65sss9ykep6F++uzh225f5IByt
691+M95pOuyzpuMUww8/TJTwNshvN2pHW8qd6RTaR85UG8ySI7RBp6gl9R5nTvLj
G7gYopgO8IJRpqqQ7kRHVVIZOqgBKPYXaAWVBBSd+seGupLHgcUZazorpsqAha9d
No62EAL8j3V972aXq/qiD/gxs3c3yglooF4vHeAXKhxhbW5TFzuFjVE1m29kfLm2
QwgTTKWA3uxDKmqkEKZjOBgpQG3/rA+YBjWeweon9WRvDnOGwOGIzqEYClQsc3vU
WW8qXokilwsJdmKL0yjJhzgCSvQjPw0cfaDxSNl+5+jahAhQNrSePUHi+tFqreAN
uxgH6V6SGF+uyX3GlT9iokj2PPbOobaM6Gz4eXyDMi6Ogf+jE/r8vf5id0fZ85b3
uT5pz8+J6CD3EgqXs/7nmXr9aZk/JSn8FAN8AATKsVOO0v+XcRHarr5ds6z0V8OV
5gY739cwvXpqVijh80HB9Yo+dEfSRlztrtiewNfO5n7g//2B9oBLge+W4749RxiN
C6SV4NDpmFfCakCui928qyaH0jLOmdgtW2Swz3YrPEvSQXl+BfYFaVsKI2jyleIm
Jb0uyAYDsOG8pkXbi1t3PNflBfxBhTUzYboXBPkOZnf0L1E/1ZnBe1JjGJd3ZK5T
I/GX34PQ/IUVCDSdGF7JfaqlX6pRHAv9oNfUeokz3VOHUGCgeWpLMJL5kQUeECiq
fXp8fANIqSMNEBud0NJbQxHI9K5NQ4nCHWqV9YlJgK9f6mboR4uNXel+SR9Xurbd
XqoSaRMzpIhg7nYJ1a4Wrcu7xSA0u+TrL0Uu+WWhcMq7HXriB34Fox5Spzr7HWKh
UVF9AHiyNuqauS/y+JqmDYrpTbBXTrWHt0JWcM2XeJzxnQyk0lyTp/n78weDzb8c
OjjWqwd0ysp5iS+o/TzVpu/XWpYgrmu2+C7B8RMJs4yV/dRACvIEw65E4g/kYlcI
vMLNwjEKmXfnb/A15qaYqnLT6pGjEGVgdQ7jeB7W4EwYtlxTVf2nFRNalu7kOD96
n2XQuOzmYzqZoSBcANx/9eDX2gkmjVwip/dmcxfej1nT5NIsyszSJQn22QprXqod
IJ4jxNb4sJd0kkfMazBqRMzK+OiF2P/qm3D8//lTm9EsJ9+3AYdyM7lmQOfv4yJi
MjlB3PFSPGNQxU9+rDCw6iM+jvmZow8M7StVjADSgChaHojnAsdJMEIr20+NbbG0
fqL5Qg0K4nI43ZcAMIdNdnRt/dCygkr5mWdLdsTox/9XYMYyscy0LwwX/TLj4HD4
8269kb3Haoah5hukr7O8qVzx5RcBLr/cgHIz55MbGExVn7sI5E/AEAtTq5QsYUXS
hOttq0K3aXf9wariDLfwBRQJgcZAM7xuSMsN9Pz0/kNRoKUik1N80tSMmQzaWsnT
uO5hPV825PR+bEAQpbKQFiI9NmX5YjbXAs9E938QBr130ufnIFTjViP5gEpm/5wE
aKuOk8WU06gYq+rWkw7Us2BdJwXlYNAdmfML5lWnG6OZnxjtKh/MiNUn5BGnTxiD
WDTwgw6OiMRU8UmXDG8bPeti5HxuYgAXmPA5TkhfS5N2k8ToP/F6wDMqUSPFgs/q
GoR904CLBu+xvB4tQjsBuLFO7TcjZA8TiJBVDWL390LWDoBDit5vWl6qKESV/5On
XoJuYKFqXGGQ/9Tzj8SVK52E8S6eak4VUWuNKQjdHSW3jPqLAYSr9T+cK55jxTPB
wLe3QnhGf21VJq+OeSviaxjrKtxyX+G55OMoYnrbvYGfVyJ39GvfImv8DyYP996T
D0rHDiBu4xWxYkISurP9csjk+cApMAI2d0cbshr9/BtgvlqmFlNHyfPHch+9eiyV
gkCwFdFirflmlMhW5Ip4in3ameXIMf0+Ilv6dPYQAoh0T9KnZZfT44TMW7ZDqKy/
iq/bPDWiLL774LGxethDNsHD61r6RX+58QPoI1RG1p9z3KQ4OxEACqUTDkhsKRI8
AFIzcTuLdu297aZzt1cpp/2pTc1wPJoRgDPcpFCBv8fvmSqNPpBuElELtJ7HwBfj
pXVYiMPXy+JX8PFacvgVihdvRmyk6+9ld+WDyQP0Zibdz+9NROZhMXojCQOvdRgP
FjzxcVc+wuN3R23noWykUHbauJB/BGWdn/DD+qqqE3OVGoDEK4g0okcYYMfZQ4qT
rkFCJuaobUpWZnvMhVFFq7YPf0lpcMNZKptC/VfCKGO5ZaUQYpMSyUrqXDxdgAta
ok7Id1tWvlJQ98x/jZehs53OHbO0vhsV+fyhMI9jQ40scXvnv35GMxcNs40JUt7L
QwNt/CH7qjqfnowZwQ22/Ash/D5CqlisW0ZzWwTSUZTpNLdXbk1XP8t6g+x9o+Oa
YyaJR1FhXFHF8CjVkQh/F/moM3R8RMCOCvuOB02KqndGRgBdz7bq8rMCYHb9oHU5
hJ4SwW1udFPK+C9bPol2GIj4qRMmyXiISlhSAg0LJwf7fmwRMo0tNH9CVuscQLCT
8gaY2WWvmfDahWCvXS+v3iqj727DDPjkWvg4HG8h0OXCpYlXM/iYDsus1OPRBYBB
86CX8W5RTGR09V295Bsc7WMPKW5CqTVi13n8qj+uRQd3ddx+VPDwwJ8Zy+4b7Gis
GWFDSKJ+FxhE0aXaWMQat+eG1P9kb/Jv4MX37Iet/iLMRUM0WNpkjWh9VLhFtNMC
7YN6l1RX5RRioWY5YrksLy5WfP0hbF7jaLfHjCF0npDqKTODdXYXMpR9Kx02P3NA
XGE56IP1+UjOWFsmVGmwMmnK/EfNK2aD54rUhErxFbptEzVd4z5aXSQWzDT0LAtx
1W2Az2JPzbnIsaKAXmIHRXn+4C8I8UwIQd8hy7Ayc17/LoH1MFwCRV4GtM1BW6Rr
8wpQ2nbfmZ1xF+CrHppMgYvZHQKd8s5n2IkEQ20pZO28orsCQeyONHytD+K/HSdR
fqQfhlKgVIuzUDKlHU9eidFMcTo78GeuOLbMIXvvEhBIgAATDhgnjrQDJh+tWvMi
yRzlvDaBsNzNxLAypZsefWx4MO8ZwuzD2T4aJ25cJOd/JSJWlXfngKfYAMJAA+Xs
QB/Dpxq0GZcPs6ZBa8YuUeguvrI1EOPR3Vssjbd3RcYstnex8HuOFVGs6ZZ9lNGT
2iUUfejyFhKSjPNgqjO/UL78b/B4XHR4iUo7Iwsuyrshoek1JwshZsyw9vnCUjtm
xh3oRhK6D0RXAkWyWYFaopWZ7efmRabY68EdwXsz4jt/D7RVjwnQMy/g+HGRayTe
8IZ+hxUGlQEqD8xZ9N4AwJ7k8PlJM62KrmIion0HOSP9+/coJU+H5P11izQEvIIT
qCe0aHJAl8DmUYm1wLKijjuZW6OOCMIcfM2e0xFt4OdAzXjzxzgEmRaG2wh9oKmp
Q2WkMg8h2FSH47uZ7ey9IbxVYSO+8f81RLXfHqzEv8A7od1rDGz/N4+/RZVWNG/i
7KjyoX2ZCJa37GejYnnXrkOXu21tB6YzyDfTfQvnWao6m3aQujtYyydNgD9wxn7l
Yje9H8T/NFq5KeWFt3CSPhy3ffEzuNUrnKNEp/Bd6IZeAYVhdTVTyXAKkxwLBf2V
dRB0oDqA93QgUJ7qwOJqkEbx1nl77sGNyvmsMBxaE3Uio9yZmupRYT6wnlbkQLw8
Q+bHXT/Al0a7m+9p6VLjmeP3XO+/gogqmnbDrNgJczhmB3uvwHQCy3Jj3A1Ocwkz
mOsGIKGDGt0/ZL/YJ7P9m//45dn5lNI4XLWz3ap/AKDc9cpL1ReBj4Il59sB9xOJ
R9b255Vddl2W5KyN7hHGSZvq/0DJ2AVgfxGHkNMBezxW+8TSzjYdOR0+YfJi12Nb
vCHgObs9y/aWvGf6BMeVrne2cVZUBVO39A5ShPnicRi/X013LLhlQtci6lN21Ion
gcidHzaU+toG/qoU3kBPNoCzP1IpBlZeEFD8qe+/xeh6iLNIdKiQzztIL9hMwgf4
FT3FbQksbFQzjv4/LisMjLijQ+v4ayf88svpMeKj832O4Zcw8ciD2sRJeE/pkm71
Zpy+wXdhY61y3a4Egl/Qwf7uX4+03jbjS7rYhMOGmDQDv/BHcrDVNEzIRZ/wwoLu
1mD5b43J2QRe7lgTLWelkAi2d/NyHAXpxv/4I4UZ61mO27tZngHhY3rjZTNgGn4t
DftiEbeA2vd1K3gjHQtMSJ/fsLefBSrKqjp8vdM5UmdUEXA4GN0Jg7ogsJtnW5s5
NUAljdiw/P57S1kvIQD8jXwZv7ZWsOK6KBoCuIs1u5pMi0c7EsFHBpw4unOJLb35
GME1TLgoV34P9gTFZ0YeexN0KBWKUoTeds79239LGFjdXBwimcfKkxZr2z4gE83W
SeSeD1ewJh6Csb/PmY8LU2O/8huwdON58kEBQJSh5sRq8uxz8AKlJ1pDcz/We1uq
xqrKmWRG1OAz3ES/w1A3+3ES229leuK3BSaTiHDJlifrf1+GFRetjXrXxdWC5p09
+ssrUPmLKg4nZjOu0xKkykq9mZu3Gb2kWdmTBAiTpZ+LQA1ul5+PLSMltg+RDxKw
jNMJJdwhWj33y+7pvFdPnmIh1KFnujfQSyeiIptCWbQWsJ6HV60Cnnd8pvY+ikBM
OaLd0wEy+JQlpTtJ2rlzjuDYJLk0hVmHl+MLbR8HwJ7RQMAT9wxNJWN6c7yUmwhR
AiEzPT9zo7/50qFUYnh07gQG5IpMbsxDMHVAvPeks4f5yow1iqoYaaI+OVQCLzu2
SpqP5eGnwv2GBHHUHtD5HQGj6QBjmyE32gmuhpJdBau67BUnSClkFHiiSE4dwvXC
JvpjexY3V9WKQzd5i7/XYQEnP2QlM4R66i0sJNw0oxpHg29SdoTw4sJK5Gkhdf69
c8GjwHj9Coq11BUPtassQsAnX9Q93XSQzhPjo1K/H+ufw5MkOJvRL2LGQxP6LXaY
OGksIFvnwWo4aIFYUMfpDp+HTTA/42toUNMM29dc287vEZrXgZOEUmj+oP9GZ1B3
KQGBkjh035Dzi2i9hl9Hj+QqCgI9ldxUdCzgjjMPw4jN76zwMBtdoUphaul1bKMj
cesdN6eqA2DnelIdqQG+Ggm4OK5Q8dNJmgC0F39IGLCIgVHyFvbVfLwq4sAdSAzh
TAURcnO6bJvLbexZ7judUSmYTIL7ZJcvckEJwv1cnP0ceiu42SzyfvMVkqDE1lGg
jr5Kjr+LCvmyzaxxJRQyZ4Q9L4MxyKgfJPAoEwguZHYDJnPg0goHWDzZVaUUxAAs
3KUrVPwF2kKgIFQ56Y0T8yu8O1p4ukyVjmw60zunULIgI3CjHZEj808u84O7DgvQ
iQFL4UwPkvr5rnrWM3CeGAq5d7U+REOEl9XZ6J1dgqK2X0Rt9dqRi/yVhB5Vc/0L
vjhllNXsoV4N6UWfjISZJxng5nEr11rk8FEN+JpiqZQuQ3HfC73H+GPpiFFpN5Rd
UgLPOxisKl5Az3OTLx55FhmqBzDnpri4On6D7r4R2irU4XQoAgA1IRklcD6rqeJC
ZXddx14hWySgZptLxOCgO66mo63yP9ACAXUtv1rdMhvrCsQttw3iOzGtqMQiP0oU
CiwXe7LeiKoouhDXcVtT991PTeRllpd5LETpptdWLU4Ht5S9oiM03muEAgQeO+1W
V7uB3S48tOM3WF0FobwtWhkdi4MiR6MJ32eqe5HkRGWrBrEYM1WVp0Hl9IcKERHq
3lgncLeMVpMHhVmnOypoBCjYTvHcScjmGg+XHKzRYiroJU8nlil3SkZ+1rgw5GJt
KI8gbPy3ohjPaU4aCstvwqlvpqfthvrq9u/GoTYmVU2iBnO0jCaX0QN47pIR/0Ag
l9piIFv5uxVK2ZNJAIjLK9A3tsoRLjiiCAhvQnEeYS+eEDWn8N/O+lQ6cZ2gnX6M
nZlKuIGSKO1gg9Y7qvk8eHA7hOvUrh78/yahkm7PWGNnM1+GAnrKqTe5E8/mOZyG
JGiSv+XE24YsnlkKJSlpNhOl5fUciSPkc/tHE4+ZKY3BADqq4aiNipMdCzpdrAPV
uNmsrLRO3gzBnpX9hjKbF2IT3T4MwO33g3EMp7cjGRY/eH4v0RDXfpBJQB35wvag
qidkTg31ZRgoUV41enSnrXpdszViBDv8ARQmJENuAJEIcRYj9pa6O6UrFtjCA0pK
5da+LsZuRCmffKFr2tw1JMOHQNryL4vkmaysIrJ4GfUT5cmDSLvICw1MmzqsmA21
gcI3z7azBlAblDT/UxDswVo/j599OB+oRQcjOtx7ZPguCemv6nH21OJT9HhgfcBh
8DjtrJ/H3FlkYT/dWM+LAxIj7SIcBADGLBkZSBLhRUhRoR6ZV/4419tefxd3kgm3
HXe7vGquZp5GF3tl/jyDHTaVIXfKWTpLlBt4JJvCZQyvH1BdAMpz3vboYaFD+Xz3
mXfVfcjzgemJqQ7zxzzmiohWV6fR9IeNaMkJ+MlgpXSWSkSW0grJgdJIdZ5+/5I0
HJ5TvssOk5eGPC34bF9PMpaWChf/wRr9+mbBaArhts/DSCT0tNoTmqZMe7xBw35G
5M9ERk1g9QyBM0XvG9DHsp5Ttj9+rs2WxC1wuwq/uYzb5zge9+nZ7Tesuo6P4lJH
/beg+8L+pMJE/1OnPBr/kpOigI9XKBcEshDoLwA2kLVYmE01bcRqD9AWuSgAqut4
/zJ32jm5fEyaukUb/vI3rRPdwEEBoiDJhxS+gsuer9taH0cMKk5UkvKSSGJ1rA5i
8MxVVUAu+V3w6jnkQONT0tFUnC1+5V2/hxbWZboAphV2cFKmtmxCgK5z40V3VJy0
7xmoK7GH29+kMRRYWgxkqLg5YPfT0Vj6mskE/2w4+Am9mINrjrzQZBi2zFFLcy85
/+1WOiafDNMqDE6wPKqa56ZV00f+rPFQDiny2eO38wNBehCjCLfWPFthAnhh1/pn
C9PpU7gJ/xO0XIsvpUElM4Y5HuMPuP/dConH1MHkvZX9xz0TnYL69xqDtsUYRDfm
cnWNF75Gu12n0buZlCZWVns9cMb55XdKQrsXQ97bXDj2A8XiGew6dB5yJqoE0C/l
fTKRhWk7f5OoB6RkvvBYxSfzmZ7ReTXI9TKDVVFCbbbkK5MZTRuR4t8ZJtLbeGed
WbGGVgt6uGJ22uiFmeaOqZ5zkNvk2OajnwwMNPY6NtcdXy4ae9tbcHgJaWMEBMjA
tlEWEr2BJezod/jB8LDLEwEdjP7ZS4fcoONgyA4Ow/vI76fHyDOb9/1RElWrI6mg
HdmRRPYjOa2Z/fQbdZefI/pdNZMwDV4SO/IaDrDOnsdICce2rpmvWivytol9hKX8
hHY0I/3mbNzindLSSVNBUxBlnV0IW/VSVtwZRl5Ij96MXYTSDlT0u5i+rHwLVeah
W13FYV74E4lZLZrgucGQrqQQc8VQzC6JtIgk4o21ZCvmoUEl7HfWzl3yvjAtIzYv
1mJ8sZjbV/SP3RCRhOLJ4WYZKsEw9ngdS5+uXTjjpSsF8zqU0PkZBV+Scc1XfCip
N6bFyBub6LbLZQdZV97jFNCUCrWDK2HXtEp1wxdO1O68KKChBqzA3yynYHzGuiJ3
1NPKoREiOMfwr8EZZsnPMoG2nXs1pATwAD/ZSU5xDHajArfTmIoM7XFgM/d8u3Zo
4dCoZMsaXQZsV7QsqfmRmojBJplEneFcxU9T+KoGhzptvCC8nLhG0vWINTp0uoNj
tNDIkBDD+5PBNmKE227bX4zrTowV15LZC5WRngBa9oEZ+sC7ZJeXTGVO8NYXIsUN
pGhX/Kwrs3+MewCyWCK/AEA2SQbtFN3aMSdOz9SHzY2bsKMayXcI2k8uIDZaey/N
Yj6xOk5Hj06zSBDLdjrcr4r/uUONbZDgI28iabAvDgydCZCXzGg/JHNuX8TlfsCp
c9XGq8nt05EP3gJGysv5RLthVDLKVjdeWwURNPGEUpWwbcyaRF6muJioJlxB363q
x7wtt1aywkWC2bD6QUALOWpHk8i7v/c9YsPvbN4udUihsSiOCyxUo6eKes7E9mZd
LvvHjyW86FRYjS6Id2BV/mjR2xXa9bxmCNgQar6BsGSCroOS8ZTH6UQXjgqwShKA
3jA+hM81zgVfND9VgIUWS2pjWz039UH2PS1cpKoCSjWLjvBlUzzB9ANDSxTn6eT0
FHHNyWt02hf5dE+NRcyUubmcTvayK54dcNlu5jGrrS4yHcgrqwx8ho5VRdTelnzu
RIOBrdaW65jNn1hzNpPQW5UITlO2/8G2p7Ols5CFR9wPaax0ZbTkkptMJ+dmL26d
2sMEhEP5kfpnR90m+Abe6zsfld4HR2TRCRzpyPyxuDxpobFjKraO+w/c0ja/lu9N
CS8VqmT8LWL4LuGqO26iINbsLuhM8hgyU2N3SnH/vMAwvqrpNXCD/4svobCMTtCX
Vq033gHds9vALLq63cGbj9PFDc1G1Z1kgTWFLAIWzoY13ctSj7EPYExb/9f8EeWh
/NDJVwbydLQQzniGZzffz2xjOl9LgLyslJlVW7ucSAsHeXwwr9AbjFuEQDCNkfcu
NBupz6TTnxIn5nFROBHWNL79LIm7TOXt/KXaKL7cl75xLidy0xNebzSoSqM+BWcD
WIa7hNAAj9aeknU40jwJ6sw8bud7B1KgECiAo0V2KCAQTDN+4qWddiCynHuU0zYe
1NuOmhvwevnJy+1UehISXOjzIsZ83yoTEhULiYp5kUgJ1eEiQzpqyzLX8KihUi5s
/D/zSl0l3Ayky7UZ/DraNmgTIFDsQcjMNcqUDzJCsqtpduRZDvbHWPQe1w3+vbY3
/qQ88oVHOZ9lhhNLgctZ1o0077i0qmjNztKmiOEn05/xZx6lvXTj24fj5geHI2UV
p6QGSexWxhB2l96WoscVEWLsFaBpayfH2w1r87JtNaOKy2bENXwyXjA3yhyK6dkj
CdA2YoiJpotTuSTh85Y3KSCxK0UfWRp5M2VYNdsBVcdSyn0IqMjhmw84OJq/BYlw
HbY/KCRXOzDQnddtVkjpNLmnNgiYDOibkUMtK3e0UyfB4C+YjRWpPYHZ+k20rZ2z
GAE0N9tNpM2FDkP7nt9fmMZkb/rRbwQ9SloaO42Sldj+9xHlJRtW/XEJg12meu0a
/Wbb6yENxxvCHlxcpTGmK1BuKuJ7sHjHm33DV3kI71DazlIgx52nuXNVoHbjU0ZF
YjPCKPaFwp2IRBdQkWyAUESQChfD7h1WL1G5FLVfAqh+mjs34N//N1hvWbPbRv4j
CDVR/7u1h1ZMLssKw+wtqYCdZAwPAwq7bEhwtnU1KMDMDAfxwN6lxuSDTMm/peUz
WXtcbTwFnmzsk9H3IHKIZpsRXMkPsxQYh3g/VaKZqu5lh3M7qqUTxCCH0iB/m2U/
ckhkb4kzgOZB2Pqqe8X3Esiu9MSNf8pxY1PbGVPjSSDdMfvQZQydLGGlr0w4uoJ/
6iCUMWMRDG5cA4CSbOAYPeX8ymgyXWwNvA6H4slkIgfmBF2rKw5+7YXAoHMgobnv
/iOCD/l6xvlViJ+yN9fpI40htnyZxSRmZJ+E/T+5hjYVkkzO9/HM+ipdqbRmeOlq
BYt9ypoeHvCGhx2XNO8KeUai2nGl4+o0809L2crZoG1/ixKMCvgmsGZItK2Y+11A
uCV//AeYuHV8qKStzO2jAtMrrIB/NnXvdELQPJQddnuUbJMv8S5ccNwApFiyWc1I
MOVmN6wQy64MrkkcclJSmHLQoYXI+4deNStENH+BtYCO3kWntNdF4Qo+l96IsdlK
KDNRfmEvI6uKadgvTw+92GI+UUYMbfAt0tQ3iumYzdxIZZTUDqqm1lY+i7XKsdPK
B3ecXOVmvjE3pZaW5wQZHUTtIQIDH9oB7PN87BAEtm/1n3eOgcEVTUrnN7cevYUt
vpk9kOudObNqCRg5RVVL3jO7eGkUNmSpZYv9ewaQP8LxOLpUB1z5XDf29Sit7ia6
2ZpO8L6ufBkTrj3r7OWF64pzlwVd48tuCz96zllUkmFIjsuarPWz4atSVHRWe3Hi
zZLVLFSFMxFAOhT7ENYdsRntlKB2Op+6Al05/SwvaIg0ljdF3KHaNH2rvm7jZ8pl
/tCriekkiwJcTb0XtkpI8p4EkrfiIPFdQk2Y/olYBHzf7T3FWuG4trx9eqlOd96E
fxztS8C3sbomcotr70NoBLhjcpJ++8d7Pb365qbP3pYGUQXK08kJtrifyBevSOiy
sNoEjV2qMgc3NnnwVYLDJ2eVtVb0GjCfSsGDlTXhpL4s+DdjrXboy2MjjcbQjlVT
iZynPAqsOoDszEIMDVMfR5JJrsp1IexWaI9kUQdFG99W/YhdGd8Qv/9l5EMBTswc
+xKj166Bbzua/e60sn8oBG7RQ55xiqGNmibE/DFNoDrHlTJ52H6Unz0OXCBmzFR8
gw36Z7Tn+ajlUV0x+oFClvxVIDbzbJvlsY47HQeMAsrbkap9aqMItZVq5hGCJK9I
Nc5YGeGBnAkrTiWcB+5x8lfrm7UhVxxm6Rypm+ANTnDU0balkv7vkmSgwCbTRlhu
me3rOJ393d0Tb8iH5Z8HN/YiZafKksnsVFu7w7frn45ju1zqU5TKZWXuuiIrvqRJ
3CFIlzYmG6JMh2kP9Ki5IKSOIj7upBNZ4KoMX3ctNfVwoTnznfCVJmClgPA35NCp
BqBGslCnBWm4Q4+uHxdP8bzyDgoZvTwAbl4tsK/TklYTiNWsY41be1FCSQqz6p39
TzMaGCALsAoARa0UJ9sOXaCjQ4KKAvq7qL0N6xkqzVmO7fVKslipzKg4RvgBMhq2
sLB7wb2LzjeNMle5W8QZEzIaTTPdO3cLgerM6iIqYNSnZlYy91vsmWTtw/3N2uBw
mFvlRmOA1iFhWH5lHk51tjqwdKe6r08E9B8lfLzA0I3NFx8mmaxh1BwGLer5NHjT
/SYDLtqu+wPdEpEHLykOgQm/P4JEAw3wsvDtz/tGvknRvYiU5PbALif8e9H7fXpd
oucs7lJPSY3L2kOTIN8yUtuZUCFNgAe4hBiaGX5Bg1NDuDp5E6A79WztzhHhGKJj
z4IY2p6hvHqWBTrTD3xqGJ5SZEZQcxLu1Ku1vXcspzk+BIwgYVv4DwRqVdYat7Kr
9TvJgFhmiMs+MdRBD/THH0jOPhZsONcWl4chDpubOzPOzhMoGLuERNDkl/99pYyE
DlWLsrj7WfksnJRimg3xcLLOsw+6lrcgFLcUwil0hrraIc0tE9JDGrsSA9ao88K+
NoEt2zQPvR1Bf1hGNJn+KvXMCpE1Gpmmy4kWh49op8tJ9OlPOplaGuCVg/apXpsL
DjB5VrWgLdo+dDKcdvf0q4xBbSG1ZnQuUN3J6YufvEeohcUslhaiM5gCqLmqcOzj
07oPS+lDu29rPWZZj+qc+CEXv6ab6YH42xevhxS4lWtQYUFy32tVkvqqO+C8YST+
4zfB29i2t+kPEtDTH/e/vrmlZIqaYcg/LQ7JeXn1uqlkIWkA/20c+ncFOcVKKBph
nyOkUTc4vUuFje0BoAbMTeC23c9BZPtZx1Ptb6Vs7DWFS+MOYjXMXLrElTcabRcX
Nf/X2jvSiD/Z5bEo52bjk4aPxOnCwSSUT0Jel0Cm/pTRum7ox9OYimB8oCzSlS5T
bms8kzZ7ad0qAFyUYt7WEkw2nqYihErWBP7/f+b1cBBNxYysqJBfMYESjo+F+zjB
2xQReIEy7zXxkX7sMKLzL+k6G0CO6HprGPldSgHc0X4mPOxgynxAYZN8O18p02mx
k2v90MWiwgX4VT0dU/6zmAu4cFw5Xwi2Y+RdeLfI1nxvCW2GUTSIn62bXM6QK5LV
7fC4zXS3EBfHKrQQk3EHAatOlOOB4Dp0ugM0EJp9Tp/mTw2W89F/rOfHEEw+NFip
9vx6CrQWwHhgBYCiNWdFxSsAyMWecPMO+9cgiPDjQY8Li1lbY4lHQ9/6i4OUmKJZ
WKGLl7hQtFuy6NWaY76OO3YfvzQEDHjFhnXtumi3dWyAV42L+1llA33LxoAsq3bn
zmDUw7MOWom1eutF3CD+dzNVrmLofjSnONz0Vk907qfyKIHRAEiMMLBLrP94iqCa
hO52KCP6jwkWKi+52g+BkO5qwxUGoQloY8oNKo5XYO4hmro8qbURerCLSNRggZxB
0Iurx4nYnUf4cSdzpqOGT+y9iGMA13yk1ogmVYuq84I9YhhYWKmFHS3o4xmUreXa
aAs9fJ069VRiRmfLN4CMg9Ej0Q8l62y7XC6DkwAUaYRvoq7HZPWQ7RCTY2oeNZLX
G+XW9faOjLA8rk3xN02zqvLFxbhFr7XoB18cdrVCHJ01vA6gR1B0ktKU+OwhsPJF
VvAnpSZPEhnt0mnb0zoDiOGyRQfYk1HuQ46Qe+Xg/wXXKaTXQemSqRCFoBBsQojt
p9x9x01jt0Q544ZNJXm2deETmwfQZMFilczeUrKYRyYc0KnOqJzgm6s9u4FsdSuG
F5/3SMLC9SLeZ4F8gXoK9B9VoplIC5kgWRL8zOA1wWIChp16RRwZbpFaeRkT5EKj
hrTAIpO00PLQoZgEBcH/WmxHBMdY4wP/H9UU825hjW/6qGTJTCpGZjlMoUK15Nsb
AIrHcWltcFKhMFBeb4H4/6bmfdiy0v3SVHah+Mvm7LTqSllZg34zz5cbzPxZw/aj
tNF9rYyhRX8a9QzqIV54NN0etD4q/v7fQdqr2idnuX21Y3wmGAh5YKbm0RQfelct
DFLLXQBlLAcoWiQY1ZrZhf0RkZ0Gl+basg/bKlRkaCTJLzhBF4O3Em72DbBn4UkP
pEAUvboGlNBUSjQpWlbgAvbgY+JoBQbm8iBqpQojJBJJIE2Vbev0bh3YcT0Yzvtm
qjoJX/V8c82qUxbBt/nMkC9r8hweiZMpQlulKHH7Jlr5odXXfoaPbyEbWkUvYBrT
tcITUL6C466R2WPq586G5sOgR3HU3u1L05/ygmp9NZM47RDMT6gvJUEcjtFvrxGq
5L5hWLa4U1PWQ5qLLKbZ/KVc/kCy2uz3XEmg5hmwLqhX3B5UNIkrZ9l+EWqOff1O
pmHsK0ag3hcIfG7wQ+eVA3qpmRkCIk+Qx+VTIzQmj5MejP5RhCUzrZOEvYaiDpyD
+vUIfEZx4ukGXh4xRruoe8qQ3uuBXHmWe2C8slxV11y8gAyxoUEvZQOfflomIYvI
wJ6MpAoWk2pwoY22IOrDs1e5gUdELX7L2b9fYBqq437/mTer/wZB0gVhq760cIJb
3f2iyoGcnCSSWggKX3R0/qUWh68HtkuzM7qJNgrYEyzYWYOr1+dm/nsbXRorysAC
7xnL63EW9DMlwsS+ZVi9/LQdZqUnVNpe6NZl8bn0nvwUAv6j196cOMidF3Q6AB/A
YPHWrPrAPbLQyWLLUAePFmqcG+RAZiGnMRTCw1AzDRRtrpv8utrSQ/S4tA6bQFEQ
G9Lfvqx5GHS1UiPxge3lyMD0V8RkzX1VAlSNbNq5f5vZo/uRn2FmT2iuOsJyF3u3
24kH69o4FIRMVsjMPkhysQ2utgQPBoeX56gwCj/6FuBVGgeU6g3wgp/ukNguzx3S
9jL8Uz+IYr1SlaMaMoKive7x71x28AEdA+yXrxd549fMgZyvKrG4HoISyliVWzrC
flv4wz96ZG4fwRRcE6sxnIDwwEtY8iq1IQCVsZPtvUN89ovoFE0yjM6YiQlEKCa6
qYPor1VPOZFCklEp+f56ckAyUTYh+sMQa/gcl16wA+PrIXHzoQt2XuxrjaVDhen3
fjQr4vVEBjB1eD02dDZLy9otHc2QzMUjrKBzlZ4CDn3XOu1ARsQ+U8+Da+QACaUo
qIErQU1HnjWMHH0KL/R+4YZPbyaudwauHcQMo2f6EhQ11ni6RoIlEtpka2bg/ACa
CY1XqZELsOTJC38uPeQbYFscEdZO8bL0EzwRNlKKxIZnejoyhKQYGHELLptES6PX
0Yp+DOe9sQ8aO2qvMmgFWXWSQtp7LA1YohZDDwfx5tcHbd2l/GgrnQ4hWBCbQkqL
Q/FfV7D3DR6c7PrPnYz17mOZvRLAkCtODAza5n0CcfcL6N1uQxVvgUVgYKyK0f5z
eFwhxZ9afW0FHGWDguUmc600nOB19ZyZA7Da5DBhiJvZ4tPdqYclT4BXGS++zA0L
iJPQLz4OvSwXD+8/OImbFOXvPdHwpB89pIJeXz41luZ4PiowxeUPUO82//mHC4pO
HxaKuze6dpzXzn3n0BAJSvg+xmXjkIuP7FA6YsW/olH8Y54W/ET2OURWnQoGq6jd
lHdog3/FYXOmK01yRrm9p6nFPjsw0Tqg+Cfz84fBVXPaMb0vBZbQxwS5Y5ODCj5T
pKdHclFrxgRgHGq9S8H+aYIoqQ5t1zggVsacloom3hd1IXemDEn594zNqB44464B
zeS6J+PVzToTx2X7T/uZtavcY7rHQmwqEQEKVBql80Q/tm9wz2NOJnteRv+XtviT
iG50ZtAEJyhD1zvr7N5iX0L0IcchvQPmCG9HX9i8pQhd1oNuQzqBgeQs2dJaxFjh
samisNB6amHrpejpAasrgqBfU/xd+QAWMsphGLizHU9IqVhZqp5rUjA/iVz2zRAo
BGpWoBUXdtcjiULtGOXw2lFFfY4X4GsMoz2GQY0VsUVXnvWDmoqhG6sCg+yRCGLj
mRo9gKZTslcfMHCdcgMCYL8Rr8GxB2h9v614wMfQu+lTUPDtefRBkJ21DV4N6HL3
yfXeXQazXMXFXZ3J3p+/OK4ahocgjCo1r07ge03MGMQ9HjHuzFqwVMBNKhtNNlGR
OHiZklZIAJDpct9vFyB38ulmqkjVKampObLihKYVXPSZvaav2EpjVOhlaGsLn6U2
FDW5DFTjmUtZMMhQa79mAE1MWHKUBwXs342vWaHYQ02/EK7sj+95HTBuRmXkaER2
Zwm3I5mRXc0xF4R9arA+yguiZUd8qmAFBx845g1ICiit+Trf7wXi22A4sFu7OTYH
VZooetLE8bY3uUCY9HF1yc+w1k+naig+C4VHEDr5PmzGUsrztzzrX95C6ULCMV5S
YjBpHFVfjhxL60ALWHru8XU581Cyg1COKxdtKXQsUlgGROiHcV7/4DW9wclO08th
3Ym1K5OYIAB+gp6zvyfBVtYD+x6AQHCYGQqmwsosBcIOobvraHhzvZEaRArhBJub
kdq7E1MKQ5bF2yz1O1T9ykjgelEuaUfEw1xIU7/JfUDaCuL/BW5pk3S98cjVESI/
lW0czw9OsdRIfuNLMQd6aZcXJMEs9hW4ktHt/8fyGcrKf18tnlXiKFu0lELezaJ+
mt8Ykz4XH/dU4DsgfWrYfDe6irzASTcG2Tm7RqNrwXQ8wDDTyECpJlR5a7okAYFd
JHCIShscYCBkHY7dgwI3bhTjCAXggyTJCxIAz4HIMKtPpdSL7oFN401sLsgBdCVk
sWO7Pg3cfkmFAUWA3jCgXJC4IsH+TkCtn544eHImWw2mnjge7tgGkP2IgeuB2mUb
Y2NnyEe4SlPKH5iGSikCpVMRBqZ0lqUVDks+FXJJdIbnbjR96tsCfiVxEMUXmCnw
F/2Tu/EWET7ryP4NrucZRJXV0/mnjeDTwwRV6tlAtjqKP5jh4No7fJJ/Ub7EJIQY
Dfghp8IvIBRRWS3K2G5IqK7JbPZBygxwT8A7bxx4navn0NEJ4RE90RefW0vferZ0
JYvES/5gGzoUv+HurAXbJe8wRKFyAvkJCwa8NVzFFdo1TP4HDO7lLpRk1CtMJ7aR
RD+HTWru1X6TrksghpuETxx8FWm9jHfQdcWVrzSoJ4d4k5vL2q5+g3ysJcqPhO7G
w3Vd06e14afxDnUFaB66/HWCNV8aklxA+HVQKbweXWNxvIWWm/AJ68W9MBNUA4SP
JffOdDHfYIDqUXycJ75uNbw2BtZYTsthLRY/8hMoOaEfOhuRzaXfswbU1ZHYpEuv
B0rQ+1OkAHRgJsDo4U/26DjUFF0Ab3qRxuWIk1b7jpDGRGbsPizxb9X9qHODFjuW
TypbULaEKHfUFwPBHcImNEtSW+q8ZJh/1nNc9VddDe+E+Uk5DoK7W/yh19QC6ra3
5Do5ufOGgB4eU9cBkJEuyhHzAid5HaBJexD4eAeByGpjVTZS3LKRHTsSu5v8CQPs
JHWsCeeS1uvlmp8limkYGUT7ISb8P8B8f9zwL+XFgw5O8Zk8v52WBgHHXAvzzA/c
iPYPNI19hdhXSPDyIR01t9TmnROsR0ASAKnZ0foZ22ViqdQMICD4wR2JCMv7hpVw
sRbjBxsGcBDs+nvXXiu6d+JE0ZGXVGHNZeTetRIB/wn84Z5Di120LF7CHbesKbI9
gmzokb8MWqsqG8QFXTlb6p7g8yG1Ux1Rxi694VYowdeUhpT0nYy3yZad3EReX6t5
R4zRH7va3FN+ya2rXg2UWnhWGEk5tr7OCINK+/S0hbvrkOh2c5quHfh5UpWl1G2g
CHtHa/IZcGO7u73nzTLLKFpZXpqEjw45QCZukdlpMm+bQUkwvyfi0ojzYVEwgUWF
mCTVgu1kJtrt4oGn7O66++vuy4m1DjRRCz0nKIWKmFEJTW/SKwk07eh6rZX6LFhY
k2Nb8hTirv4ml2zYEtNvXeMJNRMAn+H5U3wo1NaJy8BIGqUMvpR2rbnYHN3j+eF8
+xYH1MydzWb/nLLCxpRzVTbG9S0hJuZ0gmuAL1p/txQbTE/jj50bK04YGrOn0z/B
B3aytjoL5WKIj4t49b3R/e5+Z27RtRIvqhos+KjnLT9xtlbti5foZYoBJnHjATC1
7a6zaiIW2Fu6A8zYjkxyls2NZJdfuQV63IaQKbgU5z+LwRy5nNFXZgvK0KpLT0kZ
4t9LFk54Py0yJYSaerokv8wH8aMT+/St2PKE3kzANlm2Fn2bpunJ1ADQaX7BgHke
X0zcpm8TWkrSwd7Eyakb/wz/J3Ay5mAhzgt4h3jz7ACg/FekL58xXKYR5PotLqq6
+YnvS2hG1Z1/PycOBuuCEliDlSoNUamqLS49cC2eFVxN+rvE51jP2v2AOJFUvqpM
lhMh3CBqy7sOAOtUrMwXJnbGmCi58DkAU0P7xTn0A6eAxHxtvFKSBvZ6W15xHlkY
uHP7+hvkrGL6NB0xF22HwYsqyKfZ9T6tYRwb1eu3Qvsnoe3SIovWQ3dtp5FhqDVG
dk+aZ6zOHNXjqr9zbk8mWvWnvKl7D4+nKv7e/dla9PLtCL9ZeRgo6/wkZPo2xUcg
NH0q5pkFwCedKDCSp/wg9IK+/jmi5xunHT2T8gI1vB05k+At5ktlxyBcKpTUbAcS
xfFiZieDdVkgxAvGhCnBSWJLqIZyHOO1FQlsKSn+4GPWlMCZ73/56CUsBzXaAcsn
7zyBgHTmDit1yEQj2FUVJQJ+5xLo4qiO47AHi+r/nVyaYoA4VDU7Vyhx10wG6y5h
qvJhNL8/4rXCcrriptLfuop9RLt0abZreDOj/L4RHe9WSHmZ2Luw7mNMyyi63MpS
q3EqgFFRv45YzI7I5mEDkScoYIRZID7kyc/k60al83lHkjHG4jjW+L/qStC6eWK3
ay2X74aM7wWTfGl+BhDNgVz5K+TIux6x7R+b/+VU4BFP2AMSSwTM+vokqnz02zS8
9j3UcVfBEfLOUbjIthukGl4GIREanEm3H+oOYvMbFz9fMseEriowurteM+4R9cKJ
c6+lO6/oZl6Dzi1/yPrmEQHPtwQxxUWXBmKdoqJ99SfT52OsPhKozQVioBXwcUP0
8LWKE+QShPnlTmCrNMsHtzJpmceKkZ8spJXAET94TidyJEQXy2JKvCjpDwb4CYZh
gCGZdcXqZ0U7RN4M8BcUCAom/vxqk8YWJnfRzbaV2ziWn4Y1bSrpZ2fePd0YFUM6
tp+geuO9UG67uKyyLJtXo7ipzUr8mK16LmXgarIfUUYH1dX53I5fSIO8blKY/sk3
nfqWGqYr1CefcweSxBaaJmgp2dpn9MWPcOJBUxVJvE0plFdblmeLvnMtxf/hU3zW
BdJmm4vURcEgpt1k3WwJj0eyi5+EwcurfBDqSU5dV3UYzeZb8q8qAOkmAwwR3x3P
P2WCDHCCMTPpwsZ9XjoKrhktMLoRH9sPNRrAtzK2vMNzGS7pBd9PupOmtqZt/6yU
H3YHlRn2SxxFVWHq98W2PVLPMKlgutcc/Fv4mptVVcV/ylUwPCRgRWSbnX+MKnci
pZ7PQq1Nr2FVH7CQoQj7di2pVBbyf6DH/VRgwqeQZUMEQ1x/zrN1r5wRdAQFi398
kszLVbx7vOUFfMtmvCuQwjipW1+QFNyTsmRwebTg4/Aw4ONDcWq1tA2T4D525SD/
0gQoNfZ4Dw+kVcqcXXjKAezluHWkJtAUR7xg9K3zpCjBPILq9LU9hTF/4hfKMLSG
Bbp9cJ525LteREZly2Az3inAADbeyD50y8hEWltI1qWS7sKn7GuUZ997ejsqDTL+
svrpfIBj27yR8wLxql2Dz+U4CCvJWQ3AJy+xm+/lGgIVora5x+UMSIcAzMreADEo
6r1F9N/ncc/oJi3glNt4geH3Zs+dE+WJ9CUpOTm6v/wfbcOBm6hJQQGZW9A2tSfp
KczbK/UF1WFJjEagGcTW5IK2b6DMA5i7DWRWm+rLl3EV4P9lvyMCJIEBf+uWbaTg
Bi/en64QYY9IDfXDXNJGwc2/W2nlORkWpp12pzYZ+Jno/o/J7+8WcLOq6WVAnvP3
yuk6lqTyifA9fStGjrhD/rSAWOXG9hpzzpyURCOipNiJjQL5/jIWM2x5f1lZO75i
vJgAdiqjPUd+Lap25WlCVEtQxr2kLRGj5gxHUznGPucbzJ012rqaGLkDH1WvhYkE
oX2Ufdi4VIL+WFM6gV5DEROdfrWoKIF0EzEhU5myyhvpQ6kX56RxgHqGkcslAIdR
cpr+TkayrK7nBP6I/w0D8yp0mjW0xA82kQeRDCkrn1MYqSR/7C0T1fdSZlOrnHpc
yonNoWDsvpfHulkl/NJCiWAGvjCr4ec++zDil9dyrHCETptB5LFeYKaZaxTzlpGh
oxtrQ4wzWTqLlB/lpYb9y5OQrFrppi/knpeRj+ZNIDyK0ZYwb0QfXbkyIAHpoh3i
FKbGXmqgV4z1NRoBOE7Jys9KVKPnprF4vT31b4njsJ7tLNaawGOwVJ/FtHn2W+hR
IYNnxL/1PDi50zBWM2tv1ZLyxnVUps+4v2C9vluflPkhiP+sLhl3AbwcsxCqxON4
UT0jX70z2Ahi44xgkgjS4nsNHGHu8FzD+bdcc6ckZOWydnH1oLa7aJ4zd22ByA7W
aHZccobzTwetDZeZSI/DjWDBsnw6hrCQoQjvI+5S1IfxP/Qa/aAp8uAcffAV82pv
P2liUTzmQVZg0eOUUCmpxA+xIHgH1l0Jr563NOoBUzHUAvljWCeOKfl51ZlYgObM
C2EPcBx/Yoyf4qcrI4v5yPJZQYnomEPfHJbRc33PYyWJe2QEKAbjGdCgvP7jnIXT
HsTqjWUpK0oan1cjmPSIRmpJBQz711LLTCsD2/vklbAzkOCRvTjLbDskx44G3ig0
U4LbivCacczM6t/cWH37PEnsADZA2TMwskLVGIzhLXTxJI1vbNlLQChSvI5s3dTM
X3GsZmHSSSfrbXWmxVKZaYoJEbXXrYyWRZHciub06ECbA0Uzp04rNrETpka18vhD
b0ogcKKk/JzQwVlzQOMENyCrY7wqZAy1gZ97gn5KZl4y6XAvJpnHfH61PSXt/0eA
SFBTSI4qxXlMdVDY84ASkNBZn6zl1V1K+w1Y4JFBM5uOrqhUqqsOgFtToeibfOXq
TxFiwjhs7eqMQbfWYjjL6UW0mQ6gl1l8at51ubUU6dDZgxY3Y7tMDQb1wEnTmn6y
BGN1M9j6BOMKUnuSX3bJ8iI3622SasTZUUcYIgD/+Ef0JDKu2MnPCucm2Jr7i5a6
KssqO7hhzZwWJRypB6Po2+pOdmPjxNbQal/NG1fy6Y/9IEhCEn+xIX4uO97Kr1h1
t48g6Db3fsfUC6vub28p0GcB0yNhEoOnhwhpPiv0oF8uA8ibGWIq28fp3PlX7L0R
xCOV7P/wfMLdgVSc1DieFT9IimYwAFMTJ/r/yslW95Saj4kL3LZFx6p17+yXC0L/
fQlDKZKUk+u+f+DGHg7xmPsZ0ps4C8iuCyodnOechLybIqxWlwAaALBNShPo+fWU
wtrQZOnYXteE8zF7hV6xjCZ2/mZFDcbBKewWjxBE1wRcqFSRXgCCyW0traIR7z2X
KcmuUwesZOg0BVIvhexpOdzULgYycqNvp4jioR8qf8HRrLci8rbcFQkPNs9C5/BG
mUBPxacR4k7S6TlgFMWten9LNzQ+Lr3Qmr/tBgCiYUgNA8tdqrgXKkoFptvBIqQg
nF6jAWG5NaCvnTqIx2IRsPWzms29hR0jGMWxHJlrWxVQd9TCi3EbdfX5M0lwtvhI
aKC9+f54tUf7grLlchMXvxayMEeunM0E5lIHsjFsvioBKu9HEeVgH+0+SpLJqCFV
Ss1gUm9MF+SymTrFQJKJbBcxi3uMZgGUsPWCTDQxadkyjvLGVgCPCe+Hu50tbL/8
h3wLhivxL9PTOcB+Qj4MZZ/rMfGojYTGWZxSJGTmNM+68TkwPwKtOMu1KaeUYJ2j
TJf1nTKWORwe/C1QN6RB4RujbDuHQ2k67YXki3P1UYtQAjcmV1Y7a8FUXNBi/vX4
hYaOXCe+PQpv3ZPenyRJD8myk2gFuybpNkNOmNUvzmQqtzrc7ThHWzUoYzMONp5S
Q8m0z5Cu0x97zDQJdie3qFAxaeU0vu5fZdnMVxvvCb3CvEr3MBcXfZc0dFCPZVDM
JBfX7BLAsqEj6TzWd9F999oDcNyQE1jv9bd6ptty9tcyOT/kfgRVQmgSEgrzQlr3
nEO+mIixdajqezjyd1Th4cBbxxBvlxNi6D6+av+KCMMBiK/j5mvun6NruPKU/cCd
Eck/z6/5oNZx5dKjEkNWgLzfoshhy4ivsitprbcWocf100TvkeyPIUuPCsoinCYi
+PtIZYm6ojb25xSkegdwKNQNBlN+ZSP8ArOX07dLiAderEBz7b7CmtZ/MrbN8bfo
ydO3J1y8T6aqKiLIQ+JVgnr60v5QusZVJKhMKUTE8ojSh+CV88wNgI9CI+SrEh9q
owYmCByTn9bis+wJR6zkwCNiDD9ZDhzUe1mime2d5F2j+T1hREXSkkKm938p5tqu
iITR4gAyXL7b5Pr3CGrP2FOL+drKTY2zWlLpzEZTFAQSkn9NTxvNyiDNkoYQtqh4
+YZf0bV0OsXGbAxGxCiZOC1k7yyEfVGAbYJvy/3LrZHh/5rm0SOrnDLuMo7vj+1w
ipZtCA4ZxM84cMwEPULTL4gtrhCdzCgjQfPb0cIJDdkSTEFXzHI5JVTa51ZrTlo+
B+5MH2DZ3zdXwvI4R1fE1XOyALDfX1Gm7omverSJokrp8sf3QO1Q/uyuO6HpEfVg
xSkcj8cL7SEkT2pfwPh73zaZ8yDPWgeMqNZIWTBYfmv9DnROKg+e/lMx63/K8Bk4
XAXN59qAUYVe02QvMY42FpXiQI3xZ72D3kAauWRrylPOstNRDN3vqftqL08e1WSm
/0ZP1KHmuB1IPVvYrG2dTCvPjSr30Nwm6E9dFhpl7hsAmIXAov96xz3g5UxL65Xx
2euxlOF5nkrA5SUm8IkobpwHl3c6+8Qu04+HZF6Fc3beKR0JMxQJ0mnuhe80WQyb
42ayigYB6egADKPsFojSE2crSbpSkwNe9fJULBS4EXcDvUmJZqYkjk74pu3LmbUy
qbeV6Q/ItTo8oH826DllYMCZXOi2CgU1KMPyUerB5IMumRdXJFirnlvEFuHczTnL
sT0abTAiOUbRJh6E8vtpzRcuSd+IcABFiynF2U7d0RdOiRPvdF7RQlEgt5j5YzTx
EIo2oY4fWW5Dp/FG4vZlZ7Zd2r1rr6pdD934ovCm4CtH9mAUQJPhcgu1ma58sv68
1VCZaxtEiYzWMpsg3nzFejJ/rdl7AHIeVuRXWOQKHqQG1rw3vyAjDMlFsUZMVxvY
byB2VYN0XlmjLStR2J8WRZrIEXUB/DP16uJNXBnZoPcMqrmBPuExSQGWfMijZCmS
TFXhZ40SzZgcjPKBpIxnW56p5cfg4hds9AW8Wr6ClGSgfq/BWwLipdqShFmt66UN
mFfde9Jz/XGRWiv8WS5q6g==
`pragma protect end_protected
