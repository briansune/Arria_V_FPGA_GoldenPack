// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bBapZex5GifsLdSup+sXCbamB29JT88OUgea64Bl8v+gwXZzF9m2QcAAwn0RGhKj
t368z3KrwZjhJZeaQ5btq/NrrAy4W3OoiT7GxyYJ8jqUpSWpIoIWwSVdSr9yuWlH
KOb4Iy/xa0FCna+CTujcVhlbDZSUrzgs6dE5KNzp3n8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22608)
QAIRNusV697o3535NWQIYqyP7KqjeU0uSAicL+BTE464cICrem6BGQoc5EBXjlAQ
hiPka+EXO/3QaxM/GOTtAVjUuXFjJAKjItjmblboCoshWSyWhrXFV5Q7543p9SU/
i85tFIN5kv6pwDBESkST6PXSjHdpcEay96jjF+B+Znb9KzwvGg0SiFDTShHbZrvG
+6zn6r8oedzm/46jG4djyytiOwjOELXlOjncrD0rTSEybo8ETigFM60nU4toVobt
Rtd/YJN+UH/b3mrXLWmzvysRUSOJ8FjMN/sOqxq2oj/g+rSnIIO6mbM4C2JlaBn5
LsI0OfPOZ6tNDia2W8b06E6cqRLd0EvSlwb4Iewa9oG5S7DwEgbkIc2qTVVg9TBf
+SXkSD0QK0mFSZMwHQ0SseD5YX7PXomwufHgcKQJuqGUXdiVF2Is2hX2uVslRuFM
cJQ2Gu4ie9KSuq2kKwM4YoZmdZcWVn5183QDUk1hxNsuFUuJPoAeu+Gs7XJ1zgtN
QfZo00WfeC0AntMnbZnVSMkL2YvT4UQQStkRWoTvPce1i4JAqAomC/MRYduqYe/g
PifgrmJnVBiDTLu5hFngDjw/hF3TT58w21FYkDKYxq+jLDCBRoL5dMEWEj7ze8Lw
J/K6KOdAYxCGbEyg9qeCu452sdGWwnDZ3inAxcmAjk2jN2Rqc40RfRydA5jy281G
SC5X5zmoEVzNJTgcAttXZFN9UP/ZQieI4VKYQ8YQ80TkA4uKDVXaKMZ8RSuiLyxA
/DaCBLIhqQGIYiyXF2w6MGRZOZMC6kHtQdYqzKgH5+KsEFmv6wO+twqERmpyxek1
bd7CMNms97U8+lE6FCH1xE81jI207JpIFR6oUiWzUj0DhnRsm0DRx7dZxEB0Wxmo
bx+ZTkM4QQZgQ6GrrFsudO9dQT4XJRNdV54OBBzRMb+WqXnjievH1GRPi+Ho0cYk
QDA5ybDY2U2NKvDvTNBErBdtlaCpYGVMHNQFCIWgPsZ/t7JXCS6rT2QvvY9oDrL7
z2JUcJkVOzht6yrxXqQwU0V7JKgme/ZqCL5abXM7uN78LPW08jUNYzBDC9eFpYXy
aoYWMW3/GsQVz2frkiWngTOjwnetCbZGHTyQBzzDM+P7/Akhdje6oXgmYV+aFy7b
q6qzMBDq4V+ndf9N1yndZDc29xUqKIwkg8V/3Vc8Qtmz5+xyveUwIwIApSSu+2MZ
GA2PjZhcTaFZvFFbphQxzXT4cmV8CjdJgcMjhvHoX4MsJidSpAc/aXpxkbRKk7Rx
x7k+ItJctt+WTagHsvITbHUJD7q8/X2MY1Bt6eFgSLVwKISRcWmGBWj+kqFIqeiV
hItxT0vT7iHs86g5zHtOmTatY0tGZdd/+Z2Sb3c+NIEjF0ecvLW7V6JIABDpEMD9
QO+9qiskUKZ5Lpfjyb/dF8sjfzk9qEZigMB8ALYBO7Anbhn6ygU24JsetLGz1/P9
+Ampg9Fa2LakmeDNbQVUtdYyFzLD95FHNGl5KDIkTWHGLN7uwviqzZeEQ3SQuqzL
0Bm+Yt839BhSQcMx8c1uvtCroV1RBBfFtBRneEtvx6zG+OWeQ1JpuNk+wQBExLV8
pf7IVwEhanY3lXhBMWI09O/nl0nXkQ4gOcfrAHNccsVyirt9aNs4AU/XydixMZjK
yZRqu1Vvk+3Tqoodv9n5N3W7xDvesXFMJTXJ/d2NtDtAAXxYAn9YuyqqMW/kOPm7
8P1tnAXOII6kOxAFCKRg1VHF49hejfanVuDE9KGDmQwUSv2QAu5bFaGgo7tdmtT9
oiX1AmVa/UcJLE6mlVjQMhPonuA1zj5mrV162mHOs/AZpohcakAYRVG0znmM2pAR
9xaTPiGRxSdtOcaqE7wIvX5h06tY/SSL1VVZN8f9djEOgYuZFD7z+FknnbWcHTJj
IjMX7rPsY1fMEuHyRHHHTUrwfL4m2StlVUA04iCe5IHuitpAYUyruOlIFTeeTtz1
8Z8y2zJgTfdHct7gqy8sfYvOtBNOlKpwvpTCc7zGKYMYP1alfeO62RGFeuenCTk0
74PNC0bgOqCoUww6/9k7po3O66/53DFdZtpC2TNl8vuctbedN+hgcOj2p2khI7tg
SvJMP9UIjUQNk14ZHMwqmDPLnbjZWbeYZ5Ib7bijFZyF4rpXhczfyUWeOlZA//va
+mmLlNqK19PjKqKiHTzGzFUpRRlHkAwTMUj31cU05uzaMFp7A4XC638PLGj1D3Oh
zq90x6TMMCRkF3kOUFLZ/gMiv1QWwCUUxhYbnVo/eiB2Bu6Y22dmXokXxR4Od1PH
DLENGIMnvjm8vcfqwhdkkT2LoNAiAllLEzyNL1XOjV1vtZPC6ACLZtG51JDPJ37W
fSC6TD+jrWmsXTEiiLSmIoD/1m0FjnZ71LkE/u9NrwjKMwokcCvaw9lgeXQGWJGN
Sh7840IrhDSoMEX+a0NUViy/wAbdH3r5b7slGsUDvdNhmmE6qNpor1C4n+ZQbQsh
rEpMUgmCqJBjSZBYxWfsjJh3jHKtL96uXMMM5amUXxHd65T6GuTqoPUrkqWVupzj
YbylmQ1Feq2w66ndVdQiZDCjgTZIbYSsUw2ZbQcsZBSU19rY4rRWMqcUOMTivxMA
40E/Qu7bVuTVPYQ8kGSXEbd71EPGv29Lm6KxHbbJsWaxYSjcF7FkqlJIuws7+JiI
/2ofdUMzytVnihYAR/c2BfYc6QRp38kpu7gseO5TclAMx67kCnKgwjVS3CBwX6/r
tUF6/r/RA4CXO5k7wC5YmuP1CuFNCLtz/FbENirdTy/e88jkMM0GoPxtNa47dYWN
tiwk2I5mi/fiYygqUXrLJztVLmJ+Jeoi/dMlM/VZvrThZ/sey9Cu9DLGPGQgoB7p
aUbe90Dxt8WARSqrTq/XeE8ShCXGUTN7DYWBPfdTnK75muZwDAVRRiVs9xyZzp5D
drSOzLcczM1adITnLLUFTJXQqElrXCncxp6iYc9chTQWRmqr/HMbankefNRYGwLg
eg/uWwsGm8iFrZmCJO9sqWoZq5W9lghdgpTFi4Phow0DRbrXHJwZT94wJSlWnzUc
VbU1qNybpISZiVBC7y4NEa7yqqyqE2SpPaN+56RHgALxXwGQWAVx5NurnoV2dYU5
BW8FOFoAdVGxx6DDXCK337FdpyBfyJvTUtWmVj5LgNSJooeKX1fnv8V+swZs6L23
gjGnEM2ihXSl3SOLC0RJCB0G+OKdy+JG1mFmJZAMyeLOkvhGOLb6yKCv17aGw/aA
RCPiwfDocvidBWNiTM2QELC36VZTZixy3Wl9xWEum4vnSajUm1XNQB5Ll/aiPo49
uFQ6/FZh7+yXiLqEgQ1pLAb7wPUvb5kS6bQ269Upo4JP9oaLpnPNNdiW0NW+sarY
NQT12QHGIyYn3XZMHqr7gZjTH7mPwnoLTpIWI9aAP55F+hiV054yrp2p4WHzbc+h
BH+n+b4OkxQlOp3p66S+qMPVDgMZeolb+sO6sCQz+rL7H/1kK5ITsriV8SDDx4r0
IT6+kb2e+nGjU1oSteS0W1z/3JdaEtqeRr+jd+E9rYky18mYqdjqIGlSiBpfdbNh
qUEdxZMty5oy/KUhJcL5WY5iIMOfVU9V5+H86EN73sBs+LGDkjbKskJzcJUhG0zi
8g48X3oLeivCB9zULjdWZaaxKTrGAZQMMssmWlpmSRCOwHblVcuLXWsN3cC+ikZ5
g777+hkFRmhgRHEXujCr2Imxzv4Fd7q0aJ5gSPvGAjIWiDJS3aAbbx1cKD9gHeV+
tZ1L2Kh1ybwrDVeR1l/9GIPG1rv4NZTnUEi/PLB4d8o+PpjLHeIWqA26qOf/zsr9
ye4SnU8AO5NYWRBAHEd3kp4BbfJh+ggotqFrZ/843Eat8lR6h2ziY3/St7Im6UZD
ckh8G324s+b/EVY+MEtJAz3DnZqRv5tb4sgj3OXS6h9RxmO0mqbx8AX3X+T26N43
u7XHE0S1CexTnM/IyXoWIkK92jYBM7MOSsQDVhidbykbJVCENBXZpo4EKLp/Av4l
fwxifrzHwBQvXR/ylM0EMEdy/veyaAXqHizF6l5JqAjceq2GxceAjrho+kuJckY9
1KY4Qg9Jjkuagk6NEoRylvFI/fLqNjMPOoKjwnKMj+KwER2ySawtFJyKdsI2W53+
WxUWrRiFKEBIuGY4OhdkQkz3cfRyXat+2mA/+pNqETuXPE16EnPwuXVksAfuqIIq
IsO2tPKq9XPJ4KushNU2czDwZMOeZMoaN16yYpjD7cTKP7YRyGJppgV584h5eJ/u
nSi4em34PuZN5DNGA3nWuPeW0O4C7rgQ4F935qaW7YbQh+/0Ii6DC5SmuGmUNLE5
h9yUBwoDeJbVZolNwUQVx4cO/nWZ4GFNEH89lne8qWHEK1Ex2N5BB3swFxWdm3sD
k2TDj15qREN5Xbs60VVrVtTsAXCWm8OZyUpcD6eHSLAQHH39+SDe8E+74HJe/pba
h3QPr3KAGQsAz1+puWh6e7Qf6C6Osr4FunRAAhpFY9BsB5btdMPQSjErWptdMAua
IM1e1dMyAPDiE+a9ECZLw4dosFESYrlrvrMCT0i4guKG9BUKZPKCkNWflZKX8gkn
Bg6wwod97OVDnE28m/nLhB4GEtodhfxJVxsQgk6lgmOphxQuWcAxDZM3Od86C0aG
mJnIGfu8Jq/Ic7InIvb9LsbNbuNPy2+FZr7VcWIiyNEeDTUJwkI+fmefT7/HecQ+
36cyTyEMWFsxVI79Z/14WGEO7k8hGIM1tz0/MHhA0044kO5PDoDkKypEdS3K4mnb
UhILB46i9wUyIA3tFGE/PAnulk8MrlQLi2WQmcnUYzwHSaTdr5qTEMQbNcZXXvz3
vStcOFprJKZlQcVPWrKGLwGjAKKfdsxcVbcF7kymDvTUNbVKX0eaMSyCrf1M/e9/
4AcFjXSyxE36Bc1k4GI90yRlDbaXr6ypUSMZfrVNZhUN68GYcGns5Tz57EU9Uj8P
UaFj3YCVbPW2xiavhC904gYOPxlTb36/s/brPXEDqtkP4kc/1uIXt3movzzSpDZs
Dq6U3LHntH77gXcfcd6iLgF1dTMiegsRpVQVxlhAeYz9l2Etdsqu007S2fFP5KkK
K4SrS4und0Dr5t/couV23LfK0wFZN9z4+LWbbbifZd8iHr22wMhQNIuqqFI6Y3Ju
6t0YRDOpFmSKOSGXenHX/Dqc8oHks0kcfcpQG9LzWyMvGy/3YRQjVBbLy55Uo73N
EmWPMJ55yqGZ6bWdyD72SYV/++o3AXmUoFis33EZBxY8moCECEuBKWUr5BcqmNog
gYLTfIZ9kmiE2s5VdZqI5CAiKx+OPUWPUqM8JzI9vfOQhjAKnO4+i7p18OIKLTdw
dPesbk0vShq2QUckJjYbFwPW1O6Llh2i22vOo9t+bXqEUwVrxAVvzCi0d/V+i57Y
llbRakgG2Oib8DfLKxWQYdl33JIy8m5lXDqAKg1Dib9wBu5E3Or8YaF0hLiqfLh/
ADJLcyCBCWEil60WMJ7axaTpTIVSqKcU7SmhHwVi9FS6KkQsoRdhV83SR1LeXS6a
y+4Fl+CVnNwiOGf1/2/qjv1UK0QawHe22CpROOeC7qX82wwJHZ3um2JErHX2ckd2
6MIxz1+q3ZY76I6l2GZL772RvpV5GFjdEItMzj6XsMgP9ZyFhZlBL6rdvkXx1gpW
80QFL6AqS0nK0TTN4nJX5dlhd/F4C/1AEx3sqqbyk+ZVwZULv8NtwGJ1Ds2vkTat
MbfLHwDKVjPsLip0DuOZ6HxfSBJqN08gsSLIOdQejZSyTfwvotBSinQaLIXHUS2S
RP+IHdJGXIBPxyeGq/uIvYgl11/ecHaJxy0qx6+I8kiKdAPpUwz6KFNlroK8/Qpx
6YwwBxN+vKIpeMHS0sBMEMcvM3pJSNmSw+/eQ3AKmg238Fpal0cJ9+HS/XpjGcNY
AtgLDDo+s0yFXnBjjFRJwQn3TQ2yC9/6yH7E5DpuJ7YtzjyiVJEjgj+/1Aabd4YE
T0zltZRlcgv0+Ud3bhUr3Ysw93Inh1NB0oBrAiA0jnq6yZLbKS75NVVdAe+zW7oI
wFSiEZ7PqkUqAnLUNJTazo1y7mUr5Djs02rIlhcjaI32FGZJRKR2bKQUVq3rj4kR
lRLjVjwrIPMpaWTCYnsjSOrk0UFIQqZswP4/BhJJwB/8mErXBFGaBsgrhu4u9/9v
npvak4eurXPGjmfvwXkjNMmzvCD787k8kZ94wFLyzwGXRIp0UGRkzQhsr7rlr2tF
ZtXuvoseYdXntoA01UCkIhhR8ESSvx+6+bvjIRlhwLLeBkszlFI1Svg1TY34cQ7i
J/g9LT+19B+YjWJgv5XrOsNXYlvNOoVwaBnuzxx/rT8a+0VM25G8J6ak5knBGC8r
APQES4qpnvg9yYNTOyFKT379YW8TyB+QyRh89b3WuMjnKFGEZRxS3HbyyhnvbZDn
Gc4bOJ/iuEH4b7MVsXmFq9noAEMoKTTPLt3BGgtf+YbHfMkx/GukyzmxY/kZ2+sY
VZ3mZkl2TmQi0pjYdJv5P5UPzMSZKJ9gugZ0r+f1n25+a/kKgnzn5QbkLGTPZmOr
clJYBy59gNKA7tsvjOaDI3VcHKJ0N1qo/4adqGm4OKJEWbMksgBUnWcLTVg76ft1
r4ZY63fMC2WOhtk6tU1OEyM6xXU0GPEIP2pIGMV9U9uebkacBICSOs8p/SR2oJOi
0P3b3n/VAd3tV7C0MQVc3PxrVkSVG9OBP/oWz0r0yZaam/zaKXO4PWP7SqJ8usDI
QHtXC8LY7tlvDudQtg7zxaJrsPXcgrgwMyfOUE0nRKpd1d6c5CctvgnYrYspzyuT
0stVcXQQAVZb5JNjwMCPPC02qR/lz6iDHpRypwPh7IF1LzoKCk7K4rt3rIVgCP60
39ksNnUnCSSsW7iq7yTSiP1BKHdlAujjU+qKZSqiJ8ekIX0EPXh4j7vdPpW1+sEq
8c1F9prpbCXuq17FdwMlQbcHfk9mc4Rzf0cX4sazhTFjQo5a8bY6A7PcefR0lNez
iTG91AexhthlEbXULiOj3ztEDSrXlG7OPn4l4LpBQ3/WUMg0PQ2bxTbCs+Rh27EL
6pU9KGFqLXDovsYBeac1rRz9csCx6frbAezHVBqT02IYjsnVZD9+VWDvwxUBqGd3
WLQC29fRA/wOeUbfEXH1KZc/00hxSknykylk+MhSV+Af3J7aDwstYqal5giwD7Lk
ceyqmkJpSumWAdHgGzW+RgM1jF8tK2bo8BhD/PlCXxmkljQAraZhTCbBzwNL9ob3
8i09B+DwEPxp8gSiMAQAuE9ctq+C8wjFYEB5DAFja+444f8YMeJYNcNK4fxq5Tow
midXsuv3T6FdF0PmRvrvcVP2Thg2jpHiuWfGJgOPhDrnNMDA2vw/HzHbBoEaPukM
o1YO34N6nalPRX91USgqk3TSN1iB/tHi/wNbGnZHRHBtVeIPhUd/GOlCueCiHO+4
H5zba1lYC8fMjMT9ozDvWIf6J2zdkOsJyi9FUZ/3a22iolqmBNgtHXIJO/K9PDO1
5gc44Pu0Xl98BY3EUYwXMknwNFLhuSRZe9D+fiwjZ6wRYL48JVQXcvdF8W321zGx
TUXE6XDUTr73HIrX6JRYxoAOPl6annR06+PVTDs+PEnvBw3a/1Kqv5FeIHJPQqyT
9Ausnil7LLbIFY1MFaQpFKjYSD+Am4uafJGixfy4sggcTCrQm49MikA14wjhOaO3
fw8G4jv5BF+GPQ592gEtMpYPYF4sMiGOuxaDZeKJkceFvlwPBMSC0VVpRnpWIxGo
/miX/pFR3TugLt2E20Cea16c8T5IWC4aIdvbODXtesPlbsKPRu4gnv1hkOKiIJs3
JNrMNVxfgqmYimC3GYwBedZnTFilJdIv5MsMltFqUfl8Cv8Iy5dh/IdNsroAmuof
3Qdtw5k81H1n0/1nuRFBlNxxfS7Mn2kVSpJG/6d+S5BKlOiun7iH6TySFlXbkNy1
rkUOqPxqNPw2RzYrdsbNvdSdYeWxrdnU3zoL2hcBqxnOfVacS+Xq4IREwzpZic5g
J7FnrQrxkKo2yHyL1fmJI39AF20ELBoWE7Aoq7HTTmV+ZK+lNeETkX6Knm1JdnhL
ZlXocS2COaNeQ9cCWmYYghjPSxHdtYtW5C/PjGQEowPRWe3xev3qCIKE7FypgT03
qvm3De/FfoyqgUNNUiKkeq28oDBkOhB+hDl9xShnraZZ0p4D7V0IokTG/EntWBgC
rr1anXwOM9Z/pfhgxBLcYRaHzC6BvKuVO/mClzEJQrVnxafIt51Z/jJTyOBbKIia
av4FV1vd0rZ8hubYR/uHvsmVUHKL6Dh9ANn/nkglZFnCVkXk31xb9FNdpAvE+8Mp
nkJjSYQGodb0o6xMLDuEWRWg4dGeMDprkDIt5JwV/u+mdzn3GmTU/jHH+a7iI9/4
JmnzFW8t3DDetj30QaLWU+XG95x+ZBlf0CmnKakse/oPcgvF4RMAaPFshR43XYMA
tzurBvK3R3kIniAMWT2JNbMRBqFInJ8V0/SOtULIEeBKXW3nIU8vS/wTIqu9y2af
YRi+heInT5rVYtgCCp+N09914y3So0eAPy6wD9vU+ImbGEacO20DqOJqibFxA8y2
E7itJQa/JFygZ7E8oI18hr02+itvIBhJasejXJt+o6qceNPi70eBSuVosviG2uuh
zXQtEn1VHmeOyIVyFeWNdx8Az1EkjBu83dBJfMq7cukXhJkFKzRHOiSSZDXEZSv4
gk47/bHUCp62pQRbYYthGUR6EkO2KrT8CHMghYEFZ3N+bSMwqm6et0kd3u6pHfZL
z5xGvVZKcDdQwq5r1OKzRy6ErRaBkHGFegHYe6oEyU4toYoQ7/Bm6l+uIhUmeh8b
UqaJ+liemqNrBadjIxcO/HBf9jQOVlMGLaV36XPZG8OG41ypzvvVTQkrYBp1NkGX
tZ0rFEDG3/PvR+00EbV9+LdukGiDmmrj0/+PmjXAUK6yQ4st3A4/jq9fs9IIjBee
v+b6M1LOoyLY1kCWwSxPr2P3xwDXQhQT4dVOngCZqxKIxN03zL0CJNbVExW14eiF
vqgF9uWdMZbgnaUAh9sLIbY1NeH3l5xxKqQaadEqfCdXD2WfR/7lhO3KULEtq5l1
+/fMPeD4TNAsWQCCB22rpKE5F5MHK4JWtpVEcZdUdQLPPS6JL1qU3FkNZlFDgMaG
lqpsI9atQ8S7jGOCTKkk5clS3CUdl9/AQ6uiPF1ghp6ZrMqYtyTIn5zTVvXjCweY
+dBqisbgKKx5s6YtLk1NlAuvvOaodnaAW98FvaLrJzcz+eOZqIz/hitGh1zcrYfI
EPYFvtgy2LU+19b8CNtP/7aatJHUQFyzhP9lhJAWt6WE9HbZ2RM0mKhInuAHuere
yfuEaEWtsbvOzA0nKG5QkJg4EVWsqo8mQIn1VL8zbgPURK4b5xrQsxyJgvSgGybk
BYdl1gst+IQk1S6FN+CNYZzwGJZH505Ttn0ouJKRv1pTkem875LUyiYiKSWL6qgm
l2FnsxMsMx5z7ssG3qUDMDFQvq19aS/qK6iBkOgQSC+MDrPTDQ24Khxo92suqGuT
GdaWLjKm10QF4rPWIeI/kOZbYics4Sz1poCYfgureegSm3JmIOOg/X5zHwCqJxqk
IkEdU57iRNVDpM6pVGmQEsAYNyz9BigPxOJ9X5qykdU9neciFV05xEv4dy7lYt+i
lPXuGajlpT2XpGhVZndeZoCQbKu5Muy31kaPWD5G6/u1vyWgaJhTCkB91blReFUT
twj/kNvHG1FaI03pFmmdBq1i58tG6kRee56yGA/NQCjjXz0hbFUpgtkw1Xwm94aQ
yjmcUP9XVhxCCN/3fwmqohQEGYjqdwCVzjRNoieCBs7z97ojsOJefKncx0cBol2x
jYMD4LBSSr+o2DNDgJaD09qXd+PDTwfn9PhZSLOET28qb/QTJR0nIJSnaULvT/VU
+8xrwHPgpJxtEjsrg4Ed3/obwWdqyBU/6VdFOCP+yUmLzZVYiGQ6IGuTeMyXop6e
acOrRGlsAvfTfeGctX2W7wB7AhGkfxAlVidxUBfiouLPmH/g/LkmOocTxav9FF8t
JPSCjO/W//ucstaFy6yaJkzo72dRfnjEQTDts/8vr6AqAYnDXdB+gAckIQcNJm6T
jzs7C6TKVmY8F0qDKuQaNuB0FppNjCCY3bdPYNdvSHzzw3h53tH0bCB4u4Bjrl0a
ddmBMBAlKNK2LFFk91vm2vFMptVNFyAnZPDJPX3gN8dQN+hzWMK84IRnYwoLUF3y
F5oXQM+wJjA+b/8J4PzZ7F+G91D8iZazmXTu89t9CMDZmicqdGwV/iH79Q2xAAF7
IwPlEK+7YfbPRw4nM+DVmFb3dIyNKXLJO5OlpiHZroUmVyntC4Ks3qoZ6sCQMfZ3
5LX+uK0shbexpIYzxtbO1EfJrtc0nuBJH8uknFnMbJw1vOC2JEsen1lk4sI0YLPM
VNDaQoyA2IN8tqJa3nJ5FTh9sYh1nvkHhWheZaqT039etXol2znr/h2ZChuvl35W
uWwbvNkjw89nC0GmyYXIZCUL+xsKb17f2pPha4Tw09TzYF3U/5fyBSJpe48gEVmt
Zi2M3UBgJYY+76dmk4z1I2520WNAd1DPozDF8mSW6bM0qrD0/AKDjrRGB+pBtXVQ
M2y6Jz5DJCvx355myqn/5v37QKPY/sdwko8RnemEtyvmCXzOW0cFmRCUjfhqWRcd
ttRcU3YQbVKRvdT2HdzIs2u4k0MzFmy7Ks1u66Qv+hvc7Y0Jah9appFTyxSURmO1
VrhWPAFysBIXbYiMhrAyEBtzBmcvj4hu3fVqyP8QS/KJOPWFSSigMHQh6lhT7Bx4
rlq//CukBSfHz7Ih6UvjDWTBCbCotSdMSNFXMT6ANhMbXOGJuAcIfPh8SdhQ+lA0
xwDcwp2M35967dSAa+PaGzj/WrIDzvuvx39+Ij691pulC935CLmHKsuVNj9Otz4v
0Lrke852PZIM3B5um4Vom+4UITN/vP2f5iy4YIVIM+CnVYwJBn6FEUsTJw8uG82w
oz2O0eHSKLG3RekN4tVIA5QIKhcXY6RFcNxu6XdfhJRpG0Dp3UCXZW1EgoLrYUd0
tpGlNw+rOP/ZdJTrRR5dUdoaImAkYQmhjnJCwqhTc0Nqj1svLaGYszJzGiaus042
zff6GCrFNYJJQgC9Rxuc3FsaH6tlwwzUSVDSqdV6Au5KsgaL5Fv6SUhoDPva5Y6A
iy5oayffcXE790yXxL5KFg7Rf6itUeXtKoaFDR+InpjpaAJ5nQd1K5/npTj9eBaj
jztxVyhixp9stsB8yVlt8U2pzPkcqKK4iXFZMzP/An6OFJ0cGWLYd21XLo9e5GhM
G687GVsSgqrNqI6TtJ++s+qsVau3uJbuMu8vJ3OJ2FFR5W4PhO8pd5j4Sh6Zl6Hz
BeoKeorjLtNDXAQDodcXXJ9pzQYLBpmNc9+0vSBF6HBYoZ8axkN1e9+IA4PZrtit
inOqf37NjH80kjEm6BC6IO6mezf/wgIKnjXhzmtqrp+LoABY35uF61DlOdKCRA3V
yRv6p9Pt4p6GtqAAxFvUMv+P8KDu7gZg3jkPFNODhFM6H2HxSJrZFxrx7Ys/ApdZ
hSbVZkgi39YJOlzI59MUM/liOMb5yOIC8XIdRuU6lzdPGNw6SjmjNAVIiEDk9qer
G1XMWja7XWpY2GZmNpBKAyRYEpwcg0u8l9lM1PTaqPQhIwllXt2qa38ux0fOp+Um
U4bKHXKCJGsKQt92u2CYkDS2O6QOrje0khOvQEV5QESpQEVLCJuCdOeLEkyIqXC1
zy9tc6eDOmr/pzQA8Gf5o2cm+1sTzD08LyoXWFNfW/E+1U30jgiGjSMDljR1AR5b
LytB9mqXiaRmS200IIhN5mBkcn9wxDkFE+r98f7cGiPIpLcqpyFUQrhKrpKIa0kq
bG+GsHTokfgol7TYvb0B5jLKkvfjTzockpQlUmLjAdhz8mvPfYilXDcvyc8PmF+i
KA+1OAZVwb3umv22QKgORGSgUR9jTWliU0CbeaWk6rSxAc4/N+N1mAuPbthZHpiR
ahY8ty5++Z8qnKhDQ5A8dACvnY3lYM43li386esmFhmKpW4aY+4VaKC50sO1wCaM
Z1V1Mgtfrtj0jZ4B6dFjQvyScj1YmCZe2C7aYMZ1ULxZkBCWSy0CPbsCyKBrQTkh
pzZxW65UQqN2Wgs20yDsZFXsMCHviMznw/zgfX6dGuCi6zCGDbAfeX79v3KbhORq
1WK6DoDSqi/0gQiSH1fesNKU1x/KSGvROJ4jViVbt0aj1QfDTncuG8WSAmk6ER9y
gHRxY7M3MqGPs1BOoZ0Og/KMrfPjg63WFf8FcibKjvd22nSFWqICaZob13/QhL5H
xjZYrFsjX6sP0u1fIm+lnUSXmMmh5CqojNInGZibpKQPATsTcjzxfcc2DeJPc9Hn
tF6Oe5jal4+lvLoluXYhDpn8aQjpO+Av/Jr2hX/VBIrigzxd9pOBZilpVINZW208
WRgFUtVjYjpTTBFEvaN0MRJDfPA78afxjaT72eOrdyo2m7atoOhii/6sPKwEGMRp
HqlSPECFkHR1zGkh+gsb30ff7/UV9YONSUQRaYVRvTGu6NyfYbLTL7DO5swTB3VR
OoNB2wDSVx1eKmI7wChYBmUGtNgV02fbc5cM/Dj7pR0iHvo0lVWDSlmus8ZPNN7g
5jVu3fy+zcD8xYm1e7kp4Pq7IjMULk3UUtcO2tO6dHmw9pTk3drel52/UTtO2EmZ
U1QTMRGvDAJfexv9H3eY9Jq5UUJuPqS5uD9h9HdIvH905dhO1MJsKeHT1NtuZfhi
H/3Gk7XRHRlvtV4zbhnrvT8iNBKgU9UJkFt8doo7j0lZBwXELqMQF/w9/57kbS9e
Xyh5IhboAwal0GvUnTMfGiZ8D6xzHnP62tDuz9Wfde4GbuKiXpRgKj73RNhjrOkA
jq+BsiTIvB/oHB8kAnbxokqTBomz3KIdlMstfiGzdx6Y/y3if0hZ8KWSE3o6b7lS
N7dOUeEFCuR9tBxhjBjl8Aolwwk4JSCnP1r5kYospCVatdccqQ5BS7TghCIx+1RO
4PfEiJyrXs8FTEJ5RkK8xHIChn/JxARnuQUVEN/esgMGuhW5e6DTZTCfsXdV3VUW
+lY+qHAGigP1jJdoWzYct29ReshD2aljv5oXpqhg3t3HF0LZBiSorJ7W05EqZVcG
J0/kSywgDHad5xS1YJW6DDnuV0mptNPSinZlyrpG9cqqidMmhUTXbTkWtd/AYsxx
ycKs/3e36cu38JOL6FEaGYdN5r+YZrX3VfrZAapBDH4ueyI1O+qHYRf8IWow09eh
cOqhWgTN/jGYEmctJU8fC6ciTF3eImcJkZIvVTxWediOmDI1WWW5N4uXQKQ4rHON
xbS6UgCPHRuvx9f5IvCsh5Q8guxflSfh2FVOxC+XL5uLQNaYOQNnp6/Sm1tlK6JX
m9rp75VQUIPbC2b6uZQib3mSOrJo46rV32VoLkvDxQg47+LQDVe9itZdN+l7C7Bh
0XZ2NrpkOzIruBRw3d+PU7oLv0qk/wSc3AV45CSuM8S4nGvsMnrFlZWB2w2JBtyG
fij2E2BvNdGN3IxMTOk8ciasiT4e3R+vFKDDM4ak5iDjZxDiOUgmr4Vb8OZYSbV5
pkHZoxHEAkSdOuCBBaRcGCQ0lp0voEMm85NoYKbUXSeJ+q/hAbNoYxiSqD/LlAel
42W7RlawI+y+kuC2OXCoEgmwkXn/gToOJKkz70lzzZpTiVm9S222gkmplwu0iVo9
6cUIoLj9hBAIPJV5Siccv2Fwwgx04ckioEDmjrMXxUsUi0T2r9bnoCeGA8cdoIYB
xWvQzsup9FLNm5zXzrWyDe60A82/hXRrbUNWR+GZC3MjtoRRRJwYP+zgMmVMYqAv
C3B4crEU/GkPZliFEbDeY3aVzGAJ8XjGRXsPejrhGfM0Q/rBKPdDddNG7kZ0G6YQ
nQKaWUqYz/eIeE0GUY+FdxbHCZOPWTPFq9ybC2cbiGUGXa7DGhI9KM6Sxp3l5L/c
69iwLNULpnG+LUaHghanVZibvTjQ3+tzCRbHPYjqLVzneGcLe3D4UV/12X+LWvZA
CWYQscRrNSSxGnERkK+i/utkeoHeZTPm5zqUk8YUDw/cHE5tnoDp1dGV3WPnJZGL
zCuuPK40bJqhUQWiFm53iLYp7LPkxy80tfBTQ4rzzHR9n3fWR1tWIzqPvm5rQEEg
VhmqUGR3J94LAQ6k+F01+GcJCz1mVOTwjir++haQf3LtvBeTtmw5DrRsfNWLUs3Q
ILarIIzfrWKKt4S3UBwVrwMXBi665umCi/X2ylxLRm3IDg0rIaeHqTWfXOHtirS3
qwB1pElnInaA6NalieV6j7ScoVrdL7YWfgG8EcCR1RNlRBBnRzNdcNcq2Zo6dox0
h9bwt8fxDspK28Wk9PpNeeCiCY/Oab0wrd23qZCViHOSFpybmA2eKIJHjkq05RHg
lHUqeCS/zOrQ6RELhr85YPIe3BY4xCCNxIrolR+NcMOzobeHWoSZGYIVTScg9sRi
Tty1s1eyvE9RESOgG/p+hu/QWcy1+4FRFeGxjEPmDOgtA+d6MbItxJiHlJqO8mqF
/U4OkvBe1frGI2qXyF9ZDORcHp5mG8YWKsPaVaRGxH3Lb9WuSciLZkAuWtTVHv1W
CUxu7o5JosPq/8Z5+Sx0A1vzGIsTAQAeiA4rz4Um+N6jXnpqL5/e/US3aCvD3gjn
hbPKwQkosTkuX3h/VrQpXqSlzND4nOiqYQC3PYFUtt4Pn+c/ohV6clM3IFshxgxo
hUhPG+Z/OClGlTzPPIXbSUtXRLfYIXoQD11R44tJqGcl0xCIf+YEGDRRxwQlhKtV
Lb502hWkAo3DLYvhs/VBHkrhb2fXkJ6b2NyItSSzqhIHj2MbyM/rJrJXkR4l0CdX
smdCRahYzjPt7WQpOvumup70mBjjErOG57xLdDx/8qfJn/w1bBRPWKG7ZEucCU7h
BDxRpkhTc4EVX0Kj7PvABwrfEKzWiZVp+11aoFFlZlucbYBSkOO6z6DCIoy1uH/Q
pcH0CegsewJ8b4OsEZhz53qiWKRScPPBwjcE0Qc+GPG8TOm8gtKQDHHvKWZWl9pb
/iT4K4EXO8/TLaRayih6Nf4V36iIHAeEg2d+n18l5Mbh5G83VgsvT2nihczu0emd
KOAR/beil22v1rRi6pJrTYZGC5B0HtLLLDrHR07EYJhF8cXk/p7Sh2gC1gCrLkEg
+w2viLhs53epvqTro9G9ylB24X17Ju0nfQGDJRCb8u/Oqd/lko+FAWlz2eyACy4V
Ans3oBwsMJEHhZ0td7n2Va/NtMPguiJohmJXIeLzcokWhalmr2HM6SAXUkDoIBiT
JcaNTi3rSc1ThP5di27uEkxurkC8RTY5GaGFK8nJXnOi6hvCHaQNLeXvJA/OIO/V
5QRbWu6elXcRo7Azyvpvk/F70RQGRjMUg0UpkGm4tGQH2roIPHtGElx5JAUtnWya
RFyaR6NGIALN4rOoBup7Xy6WdXGVRo4EmDFYCNebosfsG1kEnSFo+Uhv93IDI9ne
V84fvrAyndQhRjwyNvjrWEyMEurJpWYsUQqu4upttpjJ53LXipDW70i/u4HAa567
noq6RTSQpPy1zju/YKgMV3TmkTj/7T28PlR0x+8fFG4QLyuuOG9m6K3lGklKXw5K
+hxh2WrvhPL3MZH7ikMKWn57qhdAiUOUMnWLDECfYH8pubTerY04kXihKa1KiaG8
QXU/QeJBcWIO4T1ywMPHXHkZmUH5uTjbWZvxqapZk4FAQUJ18D0VYtyzYmFd9/qW
1hh+9NfiLdsRb0XRTm92XUdtGTLCDGoOLiJIYN1yroYOkhZW9bGxfp9a3grGdcJb
pvxvy5JS1FMOTHDEZn63UR14Fmp1zhF3KC1oJD9Hdyr1AEy5DYIO6TiDLjzBwl00
FSRqBJ+4rOBPahgnuw5iNoeXjNpDQSYOI2GCnC80m/ViWGZi7T830eVomvNpNyxz
1Bri8/IHg0Y2tmP4asyZMPXCkZUTrKZikLg2xAWFq8JiC5INaeTIQqXVRQrZr2U0
XvwqnUtzc+TYk6EFbjR8oVlP25Zt7xduigseYqLHEFGXhlD0sEB/XGERBn3ikqtP
ci9QwXfWB9UuZlvLVUzKipgC+/XeYNjpu6zQHtM+siuIBKKFd9nF3/dcJS38fBnE
ofhR0u+2xiZBOa+vb+7IzQqYRCf2jxOM3d8UVNIj9vgkmTPMUC+SYYDvpU10S3fH
qHWoUm/o7I3Hmr5IuJefcpxjVkfFHwUdW5AwWEqYbXjQ/CMbnhh6XqEqhNCRV30l
gmet2W1PXP6Xb0lEu1t9apElC+fs1C9MvZgbU334M3c9TW26/SWTYDv/Nhmuk0Xx
5wdmulU02JE8abUM+at+dSqN1UFigOKRiapgHBfOuYkZEXNst/DlCQtXHqocOBiD
PBR1i0S3+ca/wI3ggnolEomJdIHHz8s0QzkXExklnJDlxrKnR8DmhX3QqdHdvkjp
KKgSZKyeaycMLw/mY5/rZPpCru0ylwTYs6QZ1zuoAMFBBlva14vn3alLOresqWNP
CWrmHQifBr3sYw5eSEVZk+VjXCyKYNtoK8TFXWaDXmOs9hq/GySGnmIZ/wfurqxN
TTwXMqQlwX92aC3ZXiW2Ea9ol1wNtgG1fBOwlpFJAX/3Bm4iKWnkQj3ZVYP1bH0/
s0Ni7oLZaztRKW06QoSrvuAJXzEXYOc75HzJXR/fQE+yz7gFkQzC2WTO9j14sxnk
fZ9oRbWVOB1kk4JhDNPO1Hfgmj0x/JP685DMjd/0ii+ErMy51nBj6etzFfWBRvzc
pEEfS8jehcLUazf4BWus0ft2Pcs4DIv8tk7v9r+OZzgWKubqlZAurAMpBJydQipu
QWly7R/152HfRlsdQJHu8F8mUrTerAQetZbEd/d7/O77EtmoDWv5UqxIEQYuxg80
ICOEvsnDn2yjmUiTFuk6Mq9KCJAPh7DSKKqx18xbrno69YZ2+qc2FtrYmJWP686r
nHhGOUSqCGtxhCqLloLq0/G0qaZRHSkytakgXGGBiqdvdD162e7hIS3Uk6s/JUSO
O5poRb8z1ccuA1WZGQzC5ZrHNG/MtRedMczDQ/8WKTj7d32jtM0UoE/Sznyafg1a
UMcYYIdA+rcib5FczaylygOwsxy+zils547BDPfzZr9z+HyFP1/QnR+28X2XOQLC
kbVgs5RMrEnUmPiuinzG2M1vMu6/+ET9iIBWP6pW514575fx5DBJ4BVHdSm4XxC7
cicJP/7uW4sY2t54UKa5MIOv9eRdu/LXdn67WxU4RsrNRdHiWCqCmu1EYyHLzyK4
jbpUoSkH54Mw+IZoG3NG5NwjiuHQF1es/K4oUqS5GYu4fFl7ukEnCHDco8qkzuiR
DOFUGJ7PduLDkGL3qBhgJqizIHp4fvGUK2i3nX2x5GMeeD0GlRNmq7M/3XNbyFSq
XSvdw+/0ynfImrQgVUklD8oj1tQKEolxrAepKRpSP+zWC+0ONps0rmaMXsWlC/cv
SphsbjjSnhUGsJW8qH5CNQVDL9xjXleJUBvvz1iVE+Z8OgK7tA6SfWw6ePQembMn
PUWTjK6D/Ruj/ytMhD1v642R/UCgBVyR8x3rS3CViEZGuX5xWiu5xPhmuR33BDmB
2w7qf8gZ/5/0f0nHd9eYrH35Nl0n7iprafdLhfrQVwfmB/70MLMrbeApdtxgfHvw
TYtKPS/UkUrWuSu2BCj9jAdUMiLZAgiZ2cbM907r8fWuE1LJnkrmqErwHahkBBQe
rwOHa3jzXsKF4HFVUC5P15WKScppE6nh/T5Og1SFi5qP4Gn/3dtSsNudwJ8lx3wS
HxMcSVpgCwoxqQt/hJcYnWQN75wQmqN0udACyiV+XSQWC0z+y6xo6tL2C+ZoIZnG
7ebnvvP+3nH/yY0DNvPi8vjxWmukvA8/lCf2XMUEkzUpE5hQFY3xIM9n5SaD3/LH
ClsykH9k6YxZxgQubC39RNd97DfffQOMbHjWWgcYglPjutlQdxwGdigjPNNa/xCj
055kRDE8HleWrn/PiXtnQTMQzAtvhwE04IhzDys/I5gkHFGIlgfS70RgiFgTJ+cM
XRWB3n3+X7Qldr0pyiHNG6lwBODS5jB6zYaDwHUnAY5LzpcUbG93onTkqLiTDT6o
L+yzxquxh6DufuS1RpJrpByPcXMgq0R7UJykPpafoKa0ONMWxlUc+f0SrQqKr0IK
sQiYi+HFu8btTMEq8IXzZsM5bGIHN4HQaHUkysudeQ/yiWWzNjPFJSBF5yYbi4dk
AlpOXrYFMQVNyCnKuDB54vsGTOg/MqLW/CqICglPkNdYQmU09DD4LUmCeWtNnZmd
8LLcbyB4Vd1V19xVtmR7KAu0BmnRWehhAw9csfo4jZKFwLjhkG2vXkaBsVB3Zf6P
4o2u1C/buu7JMN1hyA3ye8tfFVLEccHR2YDTkqpOSG+f2EqwA0JU/exBcfByZEr8
mB3zLkoRCXbF9np2sCQEm8qvu6JucOqRg8sxDHAUkEROX8DuqpveQWWfW62jXjTx
DjbomrFEzvqgm6PSwcmEC/JSCqOsGoB43/Mb5qDLvQXRiQucGYl6OW4NAUi9ncZ5
7i/i/NLwUyTZOZkO93dosX+ok6LoOLlqdTmt/25s20YFGsBbVT/TeI0KBmezyq0z
zUj24c1FrPKV40gsKsWaGRABCfDgz0Ro6mgJs9TAAgm2Zg5/WbMaZtWCnfoiVRg2
DtathBw8WueDckXAn61FlDsteVnEG4c62IN9tnbwsZxTa0xzMFgxzUJf/X1XwDvs
ykoOuF5Ky5mscufeeWgSWwUiFqXBpDlC1A7MT45ZVLfc+dX3EboVqypZCrZvyq3M
ElhKAKIfVfP7yemEZBreHBlcc/ijhbp4+wrDK6BczPLnyIHLhAuCD2rSXmB6Dy6L
Wiw1Mh08EQzYrrodjmV7S2DLNuVSC8zlD/LwH5Xx7iD5ipI6uJlZgg+2XdHkkieA
TGDbVTgVEF/X/QpUOZcWk7zWu5j0B+yRUOZiI5k8wQ9TrPXFCsGQpnoLz+gIU6Sf
YyQq/um9tQGhhDflVU3U63gcw29+Wx/5V5p28+g/EtbiXWjYfuhhGNic6qrmHL01
ot1UWLs+v5bQrh4KDQSnKJKEYtXn36/5574WNtNinoDi1mLS3RusbecnE/3jmhPS
iqBvlLLCm887MNM1Y0DsnDmwDQIElv3V6/iGc3GiC8rhwchQ9wvyQiC9IFPPQvEp
Ol0O25vLeNl/DfN5Y/DGwEVVJWLXwB7Dz/IoX3pBjpsnZY0osVU/TADHnqIzXWCe
L52/NlwpHaXGu3+ceb9SGI1A59Rvl7uDq0yU6TiIgXg4z29RFCpbJ/pTiTVnpuy+
4c6qCCgY9oBBR/ywqvUod7nK/KoN2a6i744l910A0N0qkqy7VEKOyAecjIWLeERS
1J1hnYraQ6JaaPq/iOcGmie4maK+9aeLuL6/mTwzTetiV957FKu3Jcl8Qu+oqolD
kdczObsb3Q1m1R0KSSRkPs2nbJFddZVHrkIYiI+DGXpK7JPe81l0hnlbDn0kNGR/
BkH8QfB/7uAY/JKK853+bQ9PHx5tPJhltdqD3EzjQ/JFZJUkW3l4GLz7MhpCVjBy
1qI1Q39OOsIMfAE48val/6tm5wQsJvI6mWa0otgxkldYmFvTSwd5hg7rCsZGDio4
pMx/sJOyGPlwJ02qu7nFzNnXEClEtYlad12mquM+Zf3uWCay5SA2tBcNKqX2PpKE
8FvGeRBTlnSA1rIqe4EESpD4vC58fH48O0iNzT4vu5aV0a6eipaCi+bWxqYb8x7w
O4DfVElpy58HU1Qx1KzvEOOwDIPmljXv2ZetG2xRe2kQJEDm2Tb36aByxPTs5nPa
ERSnAwkBPBiJwE1iHPo5A6GyNTR2G4P9BxBE6LJPAM6CyeOtCrOSsq0PiNy2c1LD
iSqqJsAU/T/l5JlkAVe3v2wgHyWAxe8nDNTqjjW+Q363AnIOq+X/X+eCurWpRyES
nzAxZ7Wjko/b3icKkC9IhYUl6c9V2ypqLMFIIjbPMkKTJwjkIDbtSexoavRN1J9N
OHhVSaCiALsi8nJuc0m+wjhndpHCzWoAnGeNilkk31bnUE5NchMfdU9FRV7CmEP7
RdOFYRHcJB7pBZlVXOq++aQtgAJwK89jv00iK+L/hi5wQsfQSAALX6RViGc4wkVL
bBB/zUikvJaC+MG/Y3OJFZnqmKa31e6ufdHgciQCZ4bPtmCyvMDR35Ka7+1wbrqU
QQmYPgwtt1PYZMHtAbGgpu4SVflI8fIwKFdKMm3c/Anub76E5otf/57pjFpiUhsr
6o8RcxLKt10IgEsr+wLkH+Fkbhes3kJHggwSmQVvW3AqKpuBpmm1I+E+pWyQWo5m
3E3bZO5I6tIWuN2hXY9NesysiS0gcXQuQ28nMs32bTYOBNORQ04xDzocLYD0LkSq
B6XvE3XJ8xJUHcvCABxzrQn5Kj6AUgxXJRgEgKwCT+W77OTxngAFx9yyTiGR1NLC
m2l+PIrlT+V9/azbm9dgJLQjY0VVPw2PI4DGGxJVX+AqyT6iXejJnU2l0LH2PVJ5
NwsCgoDOMXlml1yyk5TZ/7ygWmeH5IMFkpf2OPtUe60T8msTG+HTZvt3m3ghic9a
F1PRcZlZ7Lg1HC0xl4x94S9azZgFaMSeAmD2fGwqymcNXEJ4NqWS5drsNHED0Iiz
DSpMvwG+690BHBgzr5oFvLbHai/a6kdC+PC5noLFvBBnO1JPZq7VI0+Rbt0tyJmr
A7y/UNMyDJ9qY8ljiE4RyeZ7y2dUyyYjJERWrLTKSosmr/ABqJCqd1Y056U5MwZH
Kt751+eFPwQXj2gU6mn6DLdwaniZ/OthOE2hBX8M34lePAK5XE35Rj8512svGCzl
SqCmTWhAaTxjaWOkwcYAfFlsIAo9ia8ew0a07UGNamx7vjCfJrp3RKjqfRndlK/W
wRh1FVgZHiw0JUMG5bmAfQYnintCa5mUFtD9nuHmBBpe/DdqV+Y2cpOMFrYwxrjC
5bzmeiF0/lD8CrBmSPVNNVyNb8JUZmdzGnqJ1x/V0Zwp344N+x0Gxj1ExHj4GIcG
b3hJ+FEEjysu8a5nbfv6xR1eHgbTMi3P0u5v+4qjAqzRN9wc4xnV/D2lwE1cZFMJ
eswH0myo/RJoIMGRLM1p/livkb/B447fDjze9ikpWTuRGpr/SEfIgnj3tuZYXBUp
IrRa7uhrt+hSFq34/hyD72VWAm5yEzN+a+EWWKpNv/R+25mLFIIPw3I8+QiNbKDU
n0G+4T5FO/hMyVcIHHjTvpqWm4I5Dm/VxOQJOA/fTxDlUdkR/rVv6iyHSRncMcD4
F7cFuZRo4Bxsi3MrJ9iRlRf1eEwZJIyqn+hlQfX7MuV25r4XJc+sGwZ4w7tQ2911
NvPROGsqcU0zWugVY0E/Qxc0YPR1O/PyJdtdLM6Nke0Otodo+Kk3ksKJBq4Vj7bW
XKMWp3dcMdBCnMHI9ReggOwnPa8Jw1m8CzL5SMqTpjH71R6/k22rueEP8sG6W3FK
j+sXeMULhQRtIBxGPFQ48l8Eh0Mh3OrZWx13j0v0/fWYmam5M7oUvh7tgHHxiuAq
v0bfbJcwSU6t7XE0uIgG0ohDSwo9cyX9b9zVW8f0PZPCvSxxex1IBmB9mpP58xz3
tRnj7CcfanCMLztBZdhEkhbN65j0jxtKfMo93abPsU1UIsxawr+7QSbnUmC0N+Hs
JuPO4Z7HAt5EFLcFlmPfiAM3immjoiFyB0de42qm+rc/VpFhTUu5R5j8qZ4+F9/o
UbPDax4L3YH6lSeZP+Qnwa2cfmzyqQHbk+WdCxmKCTjgg618HxZbQ6pE7fJRt2EE
nXjTJdhpDCgzuS4oS5YaBrBAvy1hMD+7JtjB7EuoQepMKVDESHBQw49ZWfXuRFHE
wIHSmtRoXx+uZsAacsxHfA9aMC7Sb2ohxVRxo9JedTVJL4oSrjlgal75SKqHS4v3
4DFfPj69vwLt/c+8uXIHan5oc0WU0iXKgHaF/LX5DOmbGgJ7KHIV5h1eBpCaKzic
udTGBLP/zO79d1pwkwzTaLa/mpaMx13k1tcFMX6zQOByp2Zp/yM4hP8PIcb4dTx4
EPW12/xWHVrijkCrdM+m7Z1wgaXzFCF4Urgnw6fj/2f1PmVbQm2oLv4H89NrOG4P
OIlyXbuRwpsAPoSOdmAAapZr3t4OFKSrCPtgXYgH7qp2IrHUPEfpXF48p79h7iDm
6UHlxQJRb2WJu9Z34hAwLL0CNQZsYPYw9nT2u620vC16zL+HdYkz8a/uavA4e156
qm/CTbruPK0fL/YjjPN9J3WuQPJW5YbjNfFXVPMsjPZ2waewGYK27R1vppV26z78
k6Kk95mivXLNaQn29x9cyE14v+7OZlrcuOcFcCBv84IFjWT5GwIfo5oQcTmYqd0j
jpBu++GBR8FI6HsCNzPubDmfk74wXS8dabHfpSBNt9Y1qor+5WP/L0/BYOo9KPEz
z8qAvIQOQAG7h8dC4kj8PfyZiGP9H/NcvDraROwQfttFQGlsjeLwZSn0G8VmTSlJ
3TYQxee/fGuZbBxA++1vE2Sgx1A4dLsQ1KibzdyC2wVTxgibykTl7Cr8x3HzAfVV
pbExqf2B/IXB4z8KO2ussM3G+cMjJX0drdOz4kUF/ZVuSOqY/adsdQ9OulyTQMTU
8qXDgJGacrtdLNC8WZsrfCJ0u5QIoFgu36Re0rK49E90pCPw7mT/uXrUrgY2xwCn
wiRtaZEtOZWExcFSIbZBVSN0O190MrN2hTLPiqfwZo4lfdDpj7ZLRrhTbi3wySvw
L5sQTGrGKyhoNoFr76S3lIU16KOrg3o25ZIrTf/KVsEThohvFNGC/hqzeo44XAm8
uWknb3Tz/egwRd+v5L+TWnstHPTs87pQ0n75Vf41fqbEv62RYWzH6/u2YKLNQAQd
Iksanej937cpZ8Z18VlTuLkyXuI9oSGyIldwnwb1EpKTCe4evxzSHRyF00ZIPko9
PFP0sEMsVXqdj83S6qC1cGGNiYLvOfTfXFNf+3yjWa9AkUKQf5cIkUW6V+M43a9X
qtEJImYD8MO5hBz1N/PNfG7bwwitZ4Y8Z43J3+BX3+fwFYaudyU3W3qr/bK5KS/S
pCAvD6lfpxwJhQqGHfGJEMKfUAVQ+oS7oA4v36TQUPZNisj12aq5xYDLPBmsA8N1
rEe0cw0HvQUJCNyBVQ/MVRQNCMXup0+WuOLj0tTIvMUmLc4fSeDK0mNZuzz8X2IF
0VFMFg9grOBenHcAjg60SR0ieGEs63rohvWHOzfClQqJvOXkNEYFaFzzp04bcfXP
S0V+f6SsiiOiRDKPLY36qf31OMmhtAj1tOmGGmNIuD/N0mWtpbsDdQIzvU1UmYGA
QpxJZhDi3ie89rUuJVQFTtCnyRStSMfWfI3beCz2pne2n5K2NvWB7J/k+38/k/QK
kj7zbJ4q3ab/+MJ9w4OJhiF3g69afFQRNkPXq0Lwz3xYCW+8HWSlauJGcqmbintK
VVFBtlCHToL2e38nRo0q129Uf7X3F8yB8Za5YYBKacLvyOyoXtXps5wm0/u8cFG2
XvAga/TtDnueFopj6yu6YgehSo9G+Z1PvrPjMKbo6ZlTaXb7uWXKnzN39QxAOvW2
FnY5mcyrZVWtimV5qpwirHMl8PGBscWiKnK/XSQ9Y3yEYMpqk+4XSHjAM4yyoC6E
ClzASqv4iWl9KkVwvSSsB8ucBa/pbnbYj3igGqEdJqIcgmoBEYQHof7+3Rk6NCxW
Wh830o+PjHZ7E7ypbiCKYkLgdea0jFV5H0fnKxrx25yOgfkIRvIx5gg9OVYXZ5hw
3OxtRKrY4gko7sIf6NYGkle1jTQiIa0a1rZHqZpW7fH/lal6kmO0VF3r+AXDKEC5
csAjJzKsC2/JoRjLqPWT6DR6FiyKRqE+mVFn0NB3wIHYGj7W4Wp+V9pKWXxgJumc
+x8edJvJ6+1AOsUP428ezeajZuQAklxykm2qsaFNKgTMPynmpIrA80XMYhgI8GEi
A98bkeYiXJ4vct8A1WOEtqj1YCjnwuOT3k1S2BL8D1CaIyzFgAIOo1/rIoq6V74d
kjJJZEgiomvvqhiWzxZlI7kyeMepB70TFjIH/YnjiFckhALpfAf/sWiDI6uBXvVz
JCYRhkrcqWTfM5qJZ5jrBOkZ5tCkeqTvYQvVz4H+4YAbbA1EaG6+bzgnV1WOroTy
b4+uKmHrR/+eqxs251Azeck1Mj0VqPXpSHbFKHYgah9yDRNDcNrNnwvhUJlO8/gn
ZRUtPASMHq9APDItitQJzCk553G0zNWREu3N2wMQdyZYmW3HMGTNWmUdnH9fpFJV
wPngxCjXEegLRpIMNk9IdXvb4IWI1vLEWbQIx+fl6GNXBntm5i1t/eALpgsU6cHU
3X/ViNSOQaqbY/Ri1P5eUnVaR3vmqUSfzUVq4yRqmmBsq75mivslzeC9UNxk+z8I
viLBrnR/gba7dlviP/vrOuvf5Af7MaBBuoHDRvAYiEalkDF0kubaMKzevqvP/EhB
cvn8wiUor6KBHDk20E+tsRteZg6PQ9fBa/voPOux+Un9Le8J4ptaD2LVqPkK4L1l
E4Zv7DAQPeB0FkV7iPQsIQUZHSUOeNIA1tW4MtpUoUKRHrjYc80hnO4sDlfUz12w
fY3HyB3Ezoiu5pe7YMwbgow1Xx8qFVeSshNQnUnHb862Pzep21hSGsl461FtZV6P
RFxBFIlDBLaDnGj6YfOfIjKvauRszGObCDDd84Qw+D1Cuzj4RgkIno4G/V893gRA
Q69yZJUenSfjqtOGvKXXQ90LEX1fLS3i1FyJPc6UD/rCkzUKA+vSIwNQJGC9OoPo
sKUHamCkjY3jWCXw2PnbHOfb2AR78Yhf8hr0dpFEH9YVdszuDOcnLYbJgijsmtoJ
OXGuwWEFrlgirVNKycTHIgk/HCHG0uhrWhXI3SlaOiYoZXm0QkZI6S1cbBss4X5l
4401iMl6+sPfGwZRD3lQGZ7Qw1OwqYWGdqKahM3noEMyWXRN97yuv83M0wtA1X9U
gxcaU5LdE7QYe9gapEXMZKY6qV2UZYpSc3Icunqto3fLZ9CoWFq98DHP7UQaX/EA
Yu76D2LD6HnwZ6/goUXONBuRxP9UxnhMb418xeJTzBW/jxwxSWBVW17/1ae26uvb
rQY5463yOu+un96F790MMoPS8WHyRjOBl1qfAVWile56rPN5j45ohj/1oeSDeTcX
TpOVzRj7P6k+2ELV1Wj94mQJWqd4/x/TpJ6wDvlVgfqvQyFdYLHRYrNn9gHFZr/N
xrUgSIDqEPUpgbducVWf2WzMfTkpiEek/j4NF5tDhgdY8VWsE8e+kBoZawMlQNVN
t8Hytl2TQSmFM0W+LiwbdrFBpiacYCzxKY4t8JhYT2Wh0WRuOcfF7rQDWOg6CnbF
DJxOoH6M5++YH+oTVoOefSUZ2+BuHyyMKTrvqXGzoWPN1pQo/bzUuNhINjxgb+lo
5TBbjlY8V6g2I5LvS8BpeQ5ehihRZK6sXW46tVBDtvnZJtNl7FV8UVF+VgyOrNLR
lNroHw7lrqmklEwDt/ROTaXqJD5mHLhby5yIeYJwiJYr1qO54yQB4gyIytfJZVR/
wr3iU9RA7jtBWHghx8LxNLjd55xRkyYASDoK5+WWHFaSxU/4zrfpUSUItYFqbuGP
cXpUGLhVedZf6aKhZLRxrUydEWSv8RHpxEeSGWH+adkFd1jS5x2Jd+HMoepeAv1s
oxFi1stlo0Nld/Y6xtsBdYc+VvEkF38+DIcXRU2WXzL9Vz/qUBBbVK0TnrgZRgHD
lazAZ7kmlozyPVm4/GU0eV5IXDhFp5HpWw4mYammaLLd0rfUq9FF0y+1OjW6evrD
+POfutIEO4umt03zz4Cdj7yHfresFle0BcIyd85gvsENJozgk5eZgGehrHuCu/kj
NFcxuH7282rdj31CUhjMZSNFu8RPWS6Pkwn4flV5uybzbqvthuOdjLx2Ea0omtaj
9G92c92f7k1w3ThyTMiyPIMbgM+nnkUmdBmTignryB3d+SlPAo86eSNda+smHpUM
2D9rGyiY7L7o4YCp9PsK6XWddeJpbWdWmdXwHXY9tlBPETLNoKwIXCANuSEjWniJ
f4n4othJYi8hAidwHJBOevfnxHfajR1iLo1JVKoDN1Bzyev3peR7GcuO8gBKCp9F
7erAtOBYmow0VO3ue+7o6zM/hYf9uW0pX5w0A0EDCSDNTaLhoeW8y7fh7D++D+/g
gk1PvR7r/7CbmYEmlozfSrRfWQ0B++YyBSSI5hqw/DL9myAuNqqEa4k6zQ5cGDhu
erGzyz0d8QoHhmIXQO8r9OeG4Wq3DYR/pdp7ZQoty3sgLR68z6iR6/QpcRg4Dexb
+VyxCV5o1Bu+BE1Q+ckpcuEcGb2FmnJxGKS1W574Mzd47/jp8iZGM1gtDZqXxsAW
2BhnGSu98za3OzGW4ETbyomMGQr2qcVysjIBaDiTG7L/pLIGWk08uBbWhBaHiWAH
BajNW4EBzM2G38v58wc2u0861XJyiAGxsdinUxMbLMK0Ojp8rHHa0sQt3dO5RIVj
XX4xLBK7YpMKQGtYNm/0RUJsOBPZCpvHW7poyopiij3zOZSsVAbbpHkE6lWSH9/M
LXSz4p4Rnk122gqFtNTBqLaN0IyIyi6usjCXZ/cmAMtKSf1ohc+qDc6RdbJqnRok
b+/X7o+8s8hEkU+2zzj/TLyKhHTx8WEbFdwc0A3qZP0CKYv4XDSgkqV4t6anf+ax
QbNtHI9llo9qrhpAnpbTpdWHMTGZ6UvdQwkboMfRszSqL2wV+7ZKDK79y7HMvxcJ
ThZxoTs0YczeA6d7EUxGJJotIrURX+sL48wkp6kqx8UiM25nf05wL6hFBX4Bchha
FsMwFj0oCHS1AoOvL8pBH7+waiO7AoP4sqQvl38ymLHw+ZExduRsZay6wY9NNd2J
PaPEFdXjXCL0Mz0Cx6h47JruoXgHCa2YDeNUKx0f+RTPp/YnvLN+JcwLWgwfvYbi
UwpSMiC+c0e64rmbZLVHKtMoAlz1d42PH47m737M9kwFbUiz5lRf10iKw/s5yLhd
zzaUqgqJpHl7dmpb/Rf70oGXk6Ef9JnNWjOtiaRWmyYwjnLkuaPOXk+eDWVv+s6o
ihV/aIDkTPseBF+hPK8Pgigg/8jzwAsKgc/u/bsASUjOnRnMDFlzNQqDmpOgPXMd
LPuzTVIeOTd/cRDl+cvbfRrzHYcnepUM6zsUH9cJCIJtcW8Y8c3toCpXRAJRKH7e
GqhjV2Q8LjnCeITf8kFDRbLw8yXaA7xfkWV2oDXKhic/TAcpbeViMzOYGh/Z430b
/Rjkbxzv40fCbx6OeYywPCqUcjwMuNDlGFRVEiKcQupPnVY1zMwjLhnb3LhA4plj
iROqdchODPaqKnL/UltmVo0JAm0BUqbau8smWUoainzr5HMtflmGdwyPQ/Y9VnQq
i+JOGKEMHf2+xnzTJtNDiuLCGRL6XBEbz50qR/nUDhN7selxFMVtUM/9VXnMuUHn
CL+Zea3dXGo52Mx3j9I9QQeLVwDB9wDma2x/y81963RdDwLGQKER9sKhp8LGxjtS
FEaZzPdDCmrzyR41C+BVZfWUBLjgCdrsYc80q5LOQaNyUQ/PU/ujCL78xzelt9po
CNvIoDCk1IfckubHaxlKClxvLMUVr6jpcz+uasDNcwkSqjQOKUMIVahudMlBW0HS
9kolAyzt7V52wkqrXnW0LbCnN+hpwxgZ9gmuo13MeyzcUJGHBVnfRzvQuQY0GXXS
NvegFbr4nEEYMJWK2+CmVNZ/Xl/G41gScvZovdmm7eUd+/nURrCMcARamwe6HrG+
QaLIQP6sXUeCxoixJrVOFzptqh834oGCW/1aR1L9apKQT86WuKwacm51FaFtrH09
xjvjYALytI5fhk/EqygIzZSgulbRZzkOfsXaADQTs3dyOmV6AZQ9Vbnsf1b4ld+H
497jsWhQ1KgtAhPqK7buC3YrwBcDCocCKlhdHemLIudtJHDugiLfzRvJupvtz3ZT
I1U9PX4kntdNMvnjmRfSg07YTGJaLaesy4Krekr3VJhnPBU8Nvm6iI32YuUE8myr
N0FdlU7LLBMpz8zff76+3vyXwQ+9DIx8UlHa/jKKBweshreWhN2mC1GM/7YoJJO+
Z0z59k4lHL0g6XKsf9651MyO/RESkZTVFg/DBcy6+mppE6ShsTvfX+PegaExcnEI
Paf41YNB4+VWCT/gACYBqdkjqyTtA36YIIwaGgA/fnPEFgsAaYzmLE5LauuB3LyX
uufoQqLhgIrPo5f1yaZbY7h4+qlIaWQw6uPn1tnY9Odv9DabeFoYU+sQqwsIGnx5
hWQdNqiixSb18DRK1jXHq652GUo6xCWxSXtAZaPQrbbdjQgxvXehK8NcwHiOc6Nk
+uPms25XcgkjZPiNrH6l7QZvpw9udRU+8+cFjgeLXWZ6SZ9Is+O6/ZwQkXQ+dqOr
6RMEbvySUyIJgZ80P8/crJUj6EJ5+tipZ+3oOchvHVIzT0oyupx62vbrbxeyDOTp
qUy3DN2cYBZC0J4iKELsPljmMAaH30nmkRt9snaI1Ax53bW7Km3Dq68N6NeoKi/q
2ax3E1kD75Erm2qzxL+BH2OrVQj3iPkJOqAocuTGJyCeEVSvKXx2rsOruGdCP7U9
FLYr1S9T+c+FZOPQjPQDzI1wIcbmEwylJCrAJiERFOyZ3f2g/D0X6rDwzmFGoGPu
mKbMJKsn5kK4Lj2cLu/79CubLw/umSqXLw5RAg78F5Ytnq4xRiyAZndan3eTAeuz
a9hXasBHyCls5BEeN+yDyfisgqzQu1g5zPtCx4hf2OmAw8DDq7g85DwGfoAxT6Pr
e1OBCjfRmtT98DP685BGqnHKnJmfqWb64QZ1sN8U+LrCu+hAZ1TlJKULp4o4NZ6C
2J4u2fXM2EZtjetOPuwAx6q3oUxTXaAYY4S3mWlaUw/FhN6wVwd3stmh1+psivX5
sQZNDbYuXaicNcXtCUg1iaFqns0o1+aLmhwX2QexcPzOEk4nvHfVN5gao0ZuBnvu
lg6sFGviQG3ZG17yYPUm9wwMEk9Kj1CcePWhEKLBPbS53g88HqphUqkS7EQOPt8l
5rfF5ZACa69FiOYCHeZpM0DxKIFXX12QowyFIBBHSUU4NtQj3/D0VcKrTXhls0zV
VO4mszFw4oEC7XYilYG/utHQdpqeETGMAJtihRtC5VrMiFieAJPjQybasDBRXz0M
k59CQu2wAsVk9sjdY7ItPC5lqENtHXWcxmG5VdHg2O30Zrk2Yy5F4Bqdq4y0UvHm
Uw5lDgw1qC4QvCeYlUoH9Z8un972ECH/GKZR+u76K2oVBrj7vGpVvk6c3UWaWdN7
kUp9hgnAZSZ8GGgirJ55K3YZ+geDFZQ1NyE3OreyAhk0NiAPdABLxkR1mE6OKPQC
0iJ2g/8xkPqELR3b4lxAzTZRKJYaVMeWJLapnxXtB5Z772fJNZ9as4g/3AceBp+T
IWX3LctJVMURXVhjDNn0YklF8f7nqdbZiJcwBZ6kjN0gfgn47UOutZtHSBAj4/wi
GTOlsykcfovgiwQNI0e9wGGcCTiXk38OB7R8A3dfyJjo2X8NGgf53MfAuILOy61Y
hGc4ZZPxhHNfaopb+Bm8CYnbGNgbR1Z8CsJ7TOWcDU6SxGeAlpvD4SXp6mZfUP5z
61xV+LL4NM/Qn1iWflGjMJOG+46A+qbv/V77328EDolJVkB3hi2fm4zFtv2CK9lO
ubsH1Zb/7KMWGCIUSi8R5HDfMkUt/VS0r75vvRwuiJs2/twBbtrOelYhTEAnlnZK
V9C40JhWamZEwQo9clG9jhJQGhy2ZXBQGLl10sut154vdikocR31+DaDRMitPD/9
YUJhGh5T7SoKHOZm5B6qUm2p2UJboBdQRwfn8I8DkEX6ePZnyy0ooEk8u5sOEm2f
NCrccSkh5Ic6pYpTzAjLOpZCooPQs/3VOF383glAcEhoTwB83HnsXs3ZtXK4WTtw
`pragma protect end_protected
