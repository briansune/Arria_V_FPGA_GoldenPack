��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t��)���]M���UR몖��/ova �m��߽�ar4P9���3Q��V˥��u�sy!&]�?f�T�G�}Y�2sp�7������9�\�INP��Hp��5���NR���?�.��M�	��,5_|a�Y��2��ۥ�u�z�l�zud��I.�F�=�Z�E_�򟘉/ח�C�E|��Ű�6�����g�����k���5G�(By"�O�T�<����w5�x	����������Z�q�>(rI%}��̥l�
H~۾�9�f��c���fLc��n�qws7XO���m`�Z���ʟ�i�U=�Gܖ�њ��T��H�Xޥ���/�T��D�SqB}O$���I��a�[I4�o�	���a5LG����R�v	5"	������o��`��*�����P+ވ��l}�O��1�Ln�Q!�@D��vZ�rb_�E+�`�����㋹�n�������#x�Fs{�Ǡ���������0O����C��p�����d?�8l=$��OCR�Al\����K��]�HY$X�Q��*Z&fAA����t�Խ�����9�W��&
�3�^�X3zݔX �MM�2U'nw����B�@�����o��U�'0�?����s����Vq)uf�����G@a'�$;+��%_ѵ��uL�ŨPrj]tP6�Ӯ�����]�\9�k,�D:T���]��3��$c�&mfb��H�+�0�u<l�-�����q2%����c{��q>�����c������'1�ᦩ� *Z�tށ~5h�t���暠�Q�4�T��6�g�	^Ó�6�r�k뙉�yl��( �)�v��o�+�@̆��ݩu ��kd�yZ�9��Vp���-m������Ԟ�~(��ـ��k3A-�$���~
�ڔ�����(5X��Ѽ�Q�9v�|���8�U��~�B�y0�V�%];�X����i졄}A��������!�A(=��k�ޯ������� �挎K�9:6�>�?<�	��'e��I��9�#���[6�Sr�cC�vP�����P��B�����NXM�!��	� ���0�w�@nq�56��x3jv���/��l<�Yh�R��>
�2f�~>I魘(�ȭ�$����X$��I�S����qg:��綞G�@�����C���� �E��C��G$AĐ?��O㫃�P���I�;^�i�rj/�v\�_��q(�����+#bG��3���l�<�{O��.k����$�a�N.���%��WE��A�u�9�N/F�(L_JX���S-�U�pa���xlQ���̊�a�^�;>�����!�溔������)��Hj��iq|8k>��ܫKe %���ܓT�X@O���ZF�r�a� J��������w�'�yp~��=�ED|-������U���w�x �$����`8b��`���e�v����H��	����$+{�X%�N�G��v���FpNG��1���_�%;[N/rj�Tz�;`�.e�\��J�%�W����c��_B�l���H��QJ���M~���'�b8�q2P$"�w�V*H�-�6�R���mP	��1ԋ9��L�.�'���hb�~I�	���IMƥ��Q���d��Eݿ�z�{Id%<���%w�'h�5���/���A��|O�KK
M.�ˌ����Wx9��a,�	�6R�*���YP(�b�6�tԘ�B#���8����s�v ���f�o=\����͒]Pޓ����k����a�;�@A¯~)���8ٌnY�!�����G�?��WhӁfL� ��!cϼ9_�k�,]�
s�;U4|���R���[-��v��r�|eO���w��ry}�״��怬%��I՚�І��[��R� ؏$ :���h���g�}��ƸWp$���Bx���qI\=%���K��0��i�IaHƁq(��z������,p��l�eJ+f�LX��̺9�[��=2�����L�f����s���e��y)��z�C�pro�>����j����T9*��q(u���<&���A�X�8�ISOf^�Ox&{���lYh,��9����'�*E��ωܺL�D�	5@ ��3n7�!�����a�S4�#�V[���q4�u>�3��]�+�����9��E��>��
~H��?��;����J�]rը´SeFW�E @�D����(|���jV�a2��.�k{sVK�D>UP��y{4ێ9��)��6�*���ˍ�8ි7z=AZ��������,^�1���v
���2�A���Q��/���5(�jud��ҕO������.��W���D?j��}����.� ����k�o�*ⷪG�_t��G��gN]_��d�<c^~��|H�_��m�:b��4���ɏ�b	�&�I
���z�H)0�^+l�r��6�=IjH!�^%�����C�L��=3A6^�}��܍���.2b���|����~ד���&Ư��՟˹�N5,[p���D�=���K����ꒋ�
K��F96�#I;�� �*�|#����抛~7�0�0 ϯ�87D��Aw	�v�)��Mit	
6�>F�"~R_s4�'ܿ�۔w;[�/d<a�-k�2������Q�@{ϵrk��d�g��ݙq9�@�E�}K0&�(��s�M)��j�V��#.g���Е�yVbb�a'K�v�f7il��U
h@s���'c�} +'ҧ��;����ş�d�H4~�d2�kc=�YT����3�����K����myò%��M�aZxQ�ŋ.��2H�ۡ�E^�?��98�&��)D�ƴn>g�8)��[��0-����Tf(-AV�K��D�uFdF��0<Fۮ&S�Jͱ�X�Uh2��dD�0�ɓ4��fq���&.�{�t9�1���%���y?'Ir�E�a���.(�T���Q�� t^^�ҏ����́���Ӹ=�[I�
�?��7}p�ݧ�'h�w<<���k,(�+l�-����y�Q��<��e���P���+;�!�����7������H\_����h�L݌�%lj�`o�:&_���zGm,��Puv��i/���x�#�aS���,�b2���Z��&=;{8�����7I�D-�������Zn���_B�(���$��NF1�� ����$v�Agr����7$���g��Y�gq!��с(�⪼%N��(e�<��g��С�l�2d��/+�,�ާ̬͉|a�&�
_��u6����v�#6�f!fYw�e��Q��ؚО�M,��d�"�������=�X�7�c�jX�n�7�y����-��h����j2r`"h>�(�y?*�Y�ŭꖌ�)0+�Y�\y��Qʪ�foR�T��WN�j��u����-��7������"�4�X&��ę��?.b$��8���K'����� l�V���)KF�0
#$(`�n7�����#�l�S~
d�{�}��8P(o���c�M�+��b���7
ڊ`Lk��A渮$��Ҿgh7 1{{Vx{���U��A4��M��1+d���HoĊ��J����Z�gF�J���2ɯnY�{,���Oٷ�g �2�/�eޡ㴵O#C[rbf��hs�̷�mm���|�:+m����x�}D��(����]�k1��9D�8��Wt��[B��ʵ沧GtD~�BUZ�e5Ҵ�}R�,,�'�੃8�imGb2殨;ȘStI���O ~7��:�nl��h`|��Hg��hT��T#+�ګ4L�Dx1��kE��FM�D� �[q����'��<���'G���2������.L�&;�=>C2sIʋK"�h�Ǡ��r�cf� �'�m�o���+r�q��{6;�b.���s<�$�����T�bU
��`r�\�Æ˯L�/e�'��C�%�^t]�DRXS��F��v��^�V���W�7"��O�"+���P��=�S�L�����.�.�����jg<K�
l�-�*���'�1`�Gcos�h�D�{�9��f�7�:����V�"�A��ݟ;&��%������`&��v$��P8���؜���D-�#�S���[*d�Oc��_�x�Nr�ݵ�o:�:��N�R~�H��?�w�im���{Z���`VcQEK�0w��`d�D3�nf�j:u;�[�h�;���G���p
�z$扨>u����5{,�Ç*(�Es@�K�`������W� �S�[��c1�]�V"b����i^D��Nf�	o�@�9�#��@�����&vWؚ�G}M�8��(G/�0v�f�3ӥ�q�=�Ы��.y�u ܞ����f���e*ӑ��$�)H"�仇��z�Ğ�[�ij�9�~����`�eQ�/�e�����|��`���a��=�D(�?C�նx�����.�Qf1_�ࡋ�M�Iam�0�ی�1��� /I}���g�kG�O]�{1v�����t�����'Ϯ��z�`|>�>:h}by�O�����1��;����S{B}#>�v"�M��*ΗJ<���R��5u@l$�WU�륰�"��t�����P2UN�q�n��2�����7����y��|p�܆V�C=h}*uO��2��8��	%p`��s���4$P�Lm�Z�ET�Y$�ůD����N���g>��n����&��ȵd�u2�+Q�z{$�L���2�[�pQ���/���*���i�g��C����4��&�]xĢ������*'�ۭ���'��=�h4����ث�/�E�vK�k�*��!��B����d��y��I�OT��ɚ�L�&"�V^N�������ޥ����Qˍ�^B�d�z0��f���z�gP*>��"�5~�L@�����ٛ�Τ�@��}j�!7\�'�> ��m��>�Ga$��*����s���ڰ!���@H���4C�w&�i��������gׄ�e�"FnO����٧#F	���j���"��>J�c��eΎ{S���A�qi���	��� '3��U�ȉa1�/g�PO]!߉��O����'9�P6�>
�/U+y���/)����p0���.3:�J����0�=d ��er�R�@�A{Y�ǒ;M�0q�n�%�^?xAc�H�'}6�|��w�r�"\OJ\n��zJ�K�F�/�^/V����,Eۄ���E[�[��'1h)d�������C�S��f��L <�ʌ��i�ʋ�xB:�Jr�����N����� SEo}n��c,E-_����R���!�P@�`ȢW>�gU�ئ1��B�p�Ԝйw>�\�̣C8�!���J�@W3�Tb�9Ղ�=m��ԕ���+{���u����bp7��B~�*㐏5����:-��8�GK38����0��?���'H��mk�ɜI�ֳ�͔��0�P������e�;�-zb���ḇ�Ez+��P�e8������,P��v\[S��v��[ץ6S
k�tP�2f�
�+�$0��_���I��uT�Ϡ(|<�Q�~�E�5HYb�ߝ��a�IZ�0C	�Ě�d�5����e�K�K�og�~�~��}��4<�%�9�Bs~�I�Y��N��G�z@Y�e
Dُ�u/%M����]�K��$�`4̸���{T��'�rX�jF�f��n��0�O������I��\��V�����[L��~o���=y�K)�Jsׄ�XtX���U��^~�Э�9\|�x�BE�>��v#�
�u^y�+/s���޺ Mup��R��pU{Ǽ���Zq~�i�+���항��m��a��m~-^�bR��JZ��I���e��X�(�v�1��@�$�=�H'y^����ܤ%s�y���F��="ՏΦ�Y"�X�<��,o��l�9qa[Z��_Y�)�r��O���cfxB��ꞧP�m�m�����8l��
� yI͝|��gxLD�,jA�OV�,C�;�p`@�}H�%6��)^	�;�~��3_���z��57��(3l�p���M&��Ġ?��(<,��Fa�sE�u��f��[�@�J���7���@��֑����<���I!f��\-;�N�P�F�;�v���f7X�Z(ڽ���jw�{����D�^K���k: �9V�p[<�y��p���(���L?��yY�w�����1'��DZ��m
i�%e�J7�H�Ù�*D�-��l�uu��x��!�b3�/��y<�����ƥ�Á(m�����Lj�I���*�����)ZB#�	��h��&�*| k~�Q��eۮ�6�x��E�O�����ih�}P�+ �e´+1_�UY�oP�K���7N<�hJ�a���!+h@�,������$L
~ �ł���.���[P����-}o����Xt��9).T��k�",\YU�o���l%�?�ں}�� x�m�ԅL�E�f���	MI
X+ͼ��]�vm��\B�ppPӊe��to���̶�s���sU�L�u�ٟ����3�k�����|�v�趨d%�
F��r/p��[)8��Y��;�;P"�����"xo:>�L^u5,�co%'�*!�������g��3^qrjP��.K���>�[N_A�J��m�f�A�&��(��@xX����M�t�/��( ����I������]���h�_4�V!ZC�3��5�&�ev���𢸰�g������
y�	�W�Cho�S�!{��3 �����%�s8���CE����;��o���ٱ�>�d���y�3B���&p���$D�.`��n����*7|a���[k~��<�љj�	a&�R\�(�n!0�e��,�/��\j�z�[�I'�D
Z���s$Ɇ ��
��o$o��U�,�.�YC��4�a:5%�I_����`���E���h�Z 	$� ܡ䡳M���#ˁt�0N����nǋ+���yR���!(r0���19�o)� '��_��r�1fS�![�H��;��+���&`�