// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:21:15 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oZcUplVuFdpgmIGShjvVUQ/knv39GF+PYl0dIcl1mBF2ugA14nLL5TuPSofBwIcP
3itmgsPEbD4K/MLq03at70FG06fHBpRe+jI8duqKAchfQEZOCxUus5gB2uu6fcvW
sG4hEoCMWbojppro+1c4PillnK7Lm/ueuOoHFJaF6Bk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25088)
wOI5m0n4rKZHISzycmzPx938z+aOE5ArTG5MnCieC8XPO6AsfcYLVUm0SvnLQ+Pu
4pkbaLgelEmHyUhziWS3kwNojLLrO82SRX/+9t9mF2+hzFuq3VITK6MGDUqVKthb
Egwcw1uysgB8/QXlDtR3S2lD38fhdb+GZIYYclbZ/DWObx85k8AEHtPLs+OVZ0Gk
wSzA17cf1O9fbw2npmCCCgtbE9GrJicjRyUqUs+bTXcoft15cCU+GlbIKnUxeuin
qyjuAwTgBrOG7nQwyBx6f5OIBuWnW/bx0NObcbODi9pp0VKgdWb6inJvsJe+kQRJ
pkymT8ZD4eB2aGl5/nt9Xjnj9uWavnUpZTTZxftzV6ZJXeNDsUoonnmhSf54n1I0
qzXxvEAI8ACk31cJlNxKOtvhQQfGB9LEPdCFEDGch8JlAUq/2bBAFa9bzD0/KopJ
1/1pzuxqbkqs1mLO1mYPbLL5Plj6B0ZuBe4eF6ZOUNYYIuBx/s5Ky+4gjvWPIWBl
Y4chnuI+bSRnODR5XVcCIszw4QwKhtmL6G+6gctLZ/dYOXocwc1f1maBRy22abhK
F/Zfzdl3I1SDUI8XzMJc6STAGLJmU5By22sc8M0btIYwX9p8UkHpL4P7O80LuoM/
wWf2+mU7s55QFG+iH9zVY94uRoI1hnpGttYAYRslGxruJoKDQ0t2r6cCKUjzenTP
GvFQazi72PON6uIeggZOoodg/c9E9qIYtbfaH3T4Ikw7x1uuDH8Vm1RDpljjA9s9
7gpoKneUd9c4TIf5xCaQtWrc1mwMPoXdH4D475ekfHqcDQ+vrJ3tOPk/ceXLA4QQ
LjAqaJ1+boKblGRBgSRoa7QLXkTjzPm7q3HZ1gtLpQzp5BkDrHKcOct3g6J3Fk9p
vseBAh8BXJNNKceyhrtO+8B+bdPnhCh8rnHYfHt98pOlUWZxsTx/cEV8CHIWaK/h
p7UnnCuF+fB7XytTWtcG4YC0hoW18bPvvbARN30Jc2fo/vE7wCDqY44XvkDHlwrU
vM0nRs4gslIJpX8Q23azn1ewHDbOqGSeDbcoFmVv7Xb+GuzRbFLf8urpwyt4IDN3
kO5c0tarw57Y1cVcol+0V23nXiwyTpcy2V/aPQ1ZwsfpR8FUt4fsEnFnvJcAAfj3
JJiVmQjg2F0tM6KImyFLBxLPRcQQeJhyDMUAxAJ9JK6fw+78PkmDP37uXu97gQk7
3k0ItVrgmhMNKMbGzKBulg7dM99jsIk+Dp64imDSpvwUeHjHA1sdSWuLW2EYD2E1
M4OOdTYuQIaKBsojnt4GUYAnnots3Q1ASZC1lHkNGhwe3+SsrGKUPs6Z+kTEtNfK
ljotR7+8lpKkeph6dNqrsq+8Z0VPGTSsgG1zwk4tk/LG595HGlxmwJ/wiHWMUlmi
O+jpJaEXD+dwAEEDh7UGbx4uvJHHNJ5nZwExuNVrvdFPxBc+EwB8xodk9LCmXzdR
5YyxxeeB0+Je/hnQmUXmimJVbVsjUwwTitTX1O+ObkBY4KaalOmwOLDBWQW11Wjx
EqH3aoa8qzCXlIZRmeweYrOU9weeLTibaH3I9GICIroPfs8V4+gChcyZx4gxNhhO
5JD2+l4hyB2p3qqW4n0feq1cCA5H3y7nk2fAGByltEYbiZyzoLZVL7lwAdX+Tjgr
4YH6ycrve+k10c2zgvRqaYn20gWVps+pJVmfGwSDbnxizGV4WXqjC/5OGIqG9cs8
L6ID0yxu9AsAXlJL7I33reKK9ZCt3Pgqpo/PmmVqNmrCMnAK7ghf5jfer/I6W5d+
CZPWXRo4772FmHIwJgf4xqcvLuSErGxwIOAq5fR4TaTQylJUArrcZHRqIySsYuzy
L5NIj8FbRQHhaVOeNBjDQQcMQnd+IpJ/spD6VoibkNp16dmmu478ZxE3q1hRHAKt
kRHfwuewU2/FexQW2qo7BKgEtrcKmqdFmxH9X5SCqSq3Uv9rlWEKxLum1pQ1s+xm
zmX7Lk1gT10EAtqeVmIiBIMWnHF4ggH2lYuW9f5mg1ckx+DgFrM6bdB8Q2fv21eL
y8bAZtr7e+JeTwv606/GlNQjq0UlD3ikL3D9X94YSUK1VPjwNUFSi3Ou4aps/9rY
G8fVRtb/u5kyBWcC7FInpmt4MA4uNjlXQn7yhPEV9hPUqxN6+yKyQ7vaegqYco8x
TCMrXqtUGFiEXW7e8aKofjsqC5R4LmgFsjUX4SIpk9EAXJBmEIZKHK0fL4L1sC98
33l7wtm58ynhvZlUD5CFt3vTboX9TDoVQ46xLUoo53pQfJ3qAUOxlpZPIQ5RbEFy
FFJ5gUBXezsMGeg6BsroFkdYH7+/9oIAW8i1sJa9WrQcc88Xow1xQ0pr7Bwo665H
37/GBlglTLzs7/Xe1iTwhBNLCtp65uFenBrBNUdSlll+7dqf19Cjg+UsPBExbRqF
BC24KtoDN6XOKOU2kGgD7ZIkL21r92drkUm0CqGNKt3iXeyscuIU29NyJHz3DsEK
9WRpj74RS/x69OEANlaLrijIdZvT1HCKjCXlOphPRk5yrhSlJ96dW5ShOJdNHQUq
+KR1ePTtNt4q6xUjAy3rYgJAf1JcNOSFjPMjD+eZiW8PxwZEnRbNacPZFHYtmbk5
7s2LB6GqA9D9i4/N+Y1adArhCwP1VideucoHjkbqfDI6SxcNrJH4lBYmQEGR2M3i
vMhArJ+NoQ60cXLu9UxpPcCyR8i+JxXeBOHwURobsxSvxBbQRT4fexpb052ZGTjh
YVC5G+7RMF4326LUupoh4xVDoGiSGTDofQhnC1SvxrGqRXXwh5DOzaKJxLewX0Rf
fZKjWKJfKyadb+yhNr9rLvEHjxLwtRJyh0U4Gcm5R0r7oevVr/Jc+Qm4BJawyZ+n
zhgWOQNYb15F2h40+FT24qBSI7V3L0afygCCijZdyDbz08ksloo/OptKBgdbYQAg
6rWF/Zaad0P2OIRuB2buxXqtcaxN3Y9oa1sA1DzMAk+XCjHgL1NhBmf6VyF/gbSu
P6Fri5wwdVUNVr2VGfNxMtISqwLHu47WPfo+ULyQm8sMIHorU4nPsuVM4CaZHQHE
V1zdZ7CwLeUOvWgeJJCat6uEvx6HwzFrpUYUxKT4NWSJXjJ6bBZdReUWW/e7pMQX
ooYH7Xv8PEu0Wh4neIMlaV2FlTKIphU9GIYj2g4qOKsr79ztObT1uJNnXIm/+jsh
aUButwQi6FsH7U5Ywoh3X4Zh2j0Xp/r8PQmEvORtwYE6rfFqNIUDfFpIrbm/T3CY
a6uEVmjpguFSRiXdU7YDSuksH6k6DymdVI8O6ZnnYyLgPMhtswj13F7ZwEYIeVOg
d2sJegKfZWYXOq3Qxy55CTkFLjGLPFBxfcRrcVMQsCls6PZ9JPW+OAriysqnbwnD
n7zoZUPhzpNq/AjuYd8LdONU1ZTfzvUuapPt8F8QFa7Qx9A/24k+HVizDPhV2rsC
t2qBu+zgYes32sYQ7v7pDSG7hcJ2QqVoNQPhbKsgGtxFtEkiKLrwXSqnMPg0DKen
aF89REg18DuSeokgbewL7141uNe9ijdI1GaiXQIwGn7giytBC4Sy7Ahe1GXbqsZr
sznq0/kg25ozOlkY2xLeH3YPadhQSq26NciVhZef706dWpNBVA19x5HDvDiHZryL
MaC3cWBGmTkqckD3e9ob880c91tfQr9yER+X5uv9B0blLeR3nl/wuWMOEutRVwIl
+bvzrtaz5fGUcNtLcaVPUE3swZ55pWRn137/Y9I9loQhlwum+n/zPeSHL/exDjPX
urhXugEzG2uDKDdvpr4RMiR/1D0sALLetPBR/SaEdZTpea9R6lm44+g0rGTYY4IQ
TFL4N4V+sliXUxGESS6My27m+E/tURZ2n2bZHJ3ejbpMWF0fMdKWNwwF94FAc0z/
EQFtJT2g1f/A51Nv2x5BBjCg2/ILE9TNuF/jkQjGLmyASnp9KXSvEusNTpBWSbsT
ysL09cpMsnxlGn7LPjRlXzTHTQTokKHu1JFXW2OK2/sPJhJQ70nl3DVAKzBCil2H
I3e3jJ8VU+glQCCunMKdZT23UT8VZsbsu37deL/2/KTH9bsZ9OlhV50uJm1V+OB2
JpQN/LuXvW5CejBfJj5GiJBuG2m1voMbOknY2h4Njl8B7jqtdA4VkhvmG/zdHN6X
XpN5RObYGn+pyZqmEx5Ol+i+WtIt/lPxSoXF2m0rC4BYjOl6bBc5pUBIYtrKRgNp
eHOMUxixPHTcmd5aXfJHj3P87H1eRTMpvRYSvIQh7xfLsdFQw/4pVnLY+Ftl0J4P
xxPQsnXdGBt35xFjXSdql5oTGQZVfWCi8tNL1WTcNf96bEl/XEB4iZJkPJfmmSFD
pLV9wN1elKFQHqYgJAQZz7JXVBVFnpTpitD7XwFYYO+RKu81lm3DWVrSFvzQ9iMx
7psw1I4z3JQRGnixUas2ESip45vHN78//slHASHKORFrpjcWoGtBtpj7DXYr4aXo
k1zx6GaOJBADERLc7FZkNGNVeQq9aSgYq0OByObsaw0osDbKtW2DMvyX4UJzYxTa
coSv1nkP/0Ch4o4eF9dkhAqjbB6kEO9ppUx9zOr7SE9zYIceuoc5pTYWrSSgv9Fy
6Zx3OWiNZhd0FV6D8vtTj5ldLzOkOrCRWk4Xbgn3YYxMhW5uhwCxNOrZRGPgjE9+
0Top4zY8UbrBpH5Ac4jzdxrJSdZwmZNzF48yHhc7NO34WqWCorzwvm/HLNt5+4A4
2ZvfsxdYJ9YrEdKad3h+rdQCmU233zT2rrzokirXUeJ0A7kDGfPC7w7+VSF8X/rQ
bzb9wCV5PCM+S/G+VLYBiyLj96W+hCHaFHFLFLHvtAmIjM5WDO2pAMDvCohBGAm4
xHufdBlncvwSZn8o6eiN3qrTHMrAV8gZhYa92y6IwQk6jEsDx7lNPU3eCMLSWsj6
jqRrShsGP48yFtaaAc/5+eLqBkNMCTKg0TrHzfCMRBmObbSZnv0d5AdIYLSUMIGk
Qyrfif/WbtR8ufI9ZFQL9bC5br28a+N9sh2vXoRwust6enYWZ083e3dwWcBR1Si/
5P6d8+pbNBwd6Dp9lHmWN7g9nYYmH9PMo85jLd5RBhLz0Z7YUtH55HliVfrOBGks
P3E+sRfVFNM5x+67IaeT83sXhD87QNQFCLSeiQ9B5MZuc+dFkAdc5RUmxTrr5/hL
vtO7NRnWWATxSxUCnNRhyDKVq4pKRHmBaOvPXvQdLwsQCboWpjP7uURTidHeRc8k
fXGwaROlEEKoTr+Llk7TYHCgVfEeBARSor2nMxXcNJ/9lxxe54FFPs9tqywILkKk
PrdDmgdCKntwDPabK7dO5gD0B54H6e4sXYv8CTGMMcb6Y1czU/L0X/DINx5WpVM6
2/xJcHAIwVDI3kRs2a9hAoY1oo1dRP0U68mxSXSnl/+PYgW9IzsNGNAZbOGhgsmT
p2vV71Urf/2zWA7N+0igXrPcuGsbiuLLfqo+z37LvzCOm3isakYi5DYJ+v9glisX
keJ+YeuYybkyn03nBrM6FKkA2ZXBdkTI/HMiv3OHx+0bOoth4e7hrMgUiszZEZ1O
hnf/I9eHvOog/oW5L4HkqHVq6KGgvjQd9tguSAsdWxOqL5PNVHfVZy6bcgiWR+mX
G4LxKTptuhv+DWSkE7K0pIyP9iNA3Ubbr1GW5LZXPQrECkKcdj61+Zq7OCVSG5mC
xzZJA9VCLrG92B8a1YPey2si3GXB2OT277drmZ82zjr5ZGrZjPaUXfw8CMVM/oil
BKwEQgGUe1xFm7LGp4WssCpM2yFhljrCczqHkyvsm6jMGk+UF8R1dcEGPcEsEkEE
eBQQmmZyalZvI5qJxQgOXm+QzeCb32saeoyD7FPSZaw58NFEGcScJ3mZaiiV59AB
52mHn4kH6+KC8c84csDMFk/bLgQsK0//HOF96+lAO2BHxDuA6odfsqekKW4Zrh7s
DXMvuqmK03XGdC8+kR/0Q77qVgmvl00+gzaAhMRqychMifvzBlf900MHTnWQGHV0
0+i7v9xgpfj4B+K8YgKZK27AatlielSXf7ioC4xDoUQ988/31RRJ3/jnk6//8VmM
I2mkzCzIAjQ7f0x1h/4DBUbM8SZ+mHO1N8qzixXBtFoU1txKhpCagK5o9/Dz4UCO
xLUXdBOy61WvWnbWRpXiXeVfS+oZ70TaAeevn4w1y+ZHbMek2zbIxAtLAIOU390z
miSgrLTZO9OXT/E/O/31EXWMERNt9wmH4z/NQgc4YlwE/nLXYlefhx+PtSbf9Zki
yYPcsrMis1/qheQ+gOrHxh9FBBOpkQGsnhoEjtW0Z4qUuxKM7k9HWJkocpwB23nw
5gKlUwwY5H+5utQEuCeHTPyVQrT4Wk76Z9d0aSdj+vw8wLhMlW/GILTZxGlrw0zZ
nRDHrKokEXPPyyIIZi3HxMvIahvnsGx+AvNOe3AgtP7wBcAlxZGE9ob4YA7cet3A
r04cm+Sww/SKjzwpQMZoh2nbSd9uHBkBVI+wrc3L17zbcbw59YSZEELsFFBWOI0/
L7fphLqhFS7HjvCPXa8W2eg+YzVc0fNQp4hNPt5IC7mU2k0pLy62f1WIy9ZDab0O
yif7O8zGdgWE1NCpvQqvhO8ft62DJehgMRBEC4Ik3kvjiPBLES+TjtjqGU0ev+eh
ln1qnSF1/hJcfmFOq3EIK8UMrgq1bFSizfbDSxyjP2po7UuJPMxIRDcNpIBDcFw5
WvcOs8iuNIniOiV9YYedlSqbco0KCnbfAfmmMM+h0grOhXD05iNzFZTOeGsfOXjb
jhpocL0kFjcaL00JjESMOYDTXgvjbJxdvqerefR5fhqj6iOqlHISIlvn+0Qx3bNl
AGfJHrvBf3mp8g+II5QDrPKW7jx7QDf5aFd5MMET2MW11xbiun+ZQwKteoUCfBMS
D6Cre6ZvkaxoMv4rEEQyFuThXK7S3EyYeodOVt1mypM2AmKNY40jf0b4KE2qEQHH
KLxIp2Gd0XBs+c2SwvTD5MJY4Z8MYirzI0VsqsN9l0VNHFXr7HfgkZidpueH32Y6
9qw3/KQq/zHdAckvvxhdlhrvurqiUE0jgMmQMlTX13YNztmnAC6b9le48hJiCOyK
Wdu6LJRzqx1x+iCq2fy1SCUEtnTmQsGacjoudjr/aA1Y4ZYmO9UkBikbEqX9HURB
aHd/tk3Vn/VJ/A/6CvyFH9FkiRVLie4UkXNSDvw/Ewh6mcHHV8ETvOAQptzMLgnG
UiLS4ZIY99fIZaP64JjMo/cp/+myExtlICDKFcfcXC45YGsI9DUbT9EAyecpr6p7
8gvjVq+yVo76qs3iEm5NEULx0DX1PphseyOHAcucS69Wy3q4rHYiB6A19d2pgdhd
mLyx9LmCY0qpZeB6p8BKiTZfe8RWilgxkWbb5eYpfv80/YtoagcSpG55QI7y4GoJ
wSvVkuBgO7iNEcZImMXPqnT+ez1KMKOsflzhH0TwAIv3By1ewjkEK3S3pVr4z5BR
lTinKMVVYX+Zek2WozMdPqDAh67pEA1dJU5W8beqoEyoVpB63Foomt9tIiXtBY5+
Rt97yn1Aj/jKMGTKruNA23WEtVTGec5Mi5oeZ0EzSOwUnshY20/4o2Aeuq8afgt6
ESfsmShZipNrl5m2G8XHE1LUlrDkk3Qu0pW3Lrwkwq5tXuQiq6vdB7HGw3spMzu6
qKJmreBvXnc3L+PcKlwkhMg6CnMhQfItuGYND9+/o5xEA0u4sWY59IWeKFQMmVDr
ZduqnfJ1Thq/2rpQ+fykqPbhSxZJNFJHYegMfD86b6UKuFsPwajRBdJjK0ZWYd4A
a43TlllV99muDD5JXm56g2WGanpdUJT6Q8IVje261i7enihasPK2Ng1TYbPIjfjl
9woVhYIt/FJ0r/1PQyB3B41bD5aaAhJ7O2hRIuYDQWMXD/IZbZLdqFCeV/CrIEdD
nM37lLDoda/iKHwv925k/XUhuo+y/GuGSJDJ0d4n0jc8xy0xKoVeXUjF2vkTFd1W
S3g9HjGILTn2/ass+KxpIBdaC6BucR3bYE+Fc5sMFke3cCwx8zqzgVbDNRbRwRFx
n9prEMqYdvF/niyf4JnsF7YP/M6CqtEMV/+pkxMnoM5o3bQ5gZAyBB+k9JRaLsFk
8vVlQcjI1k92tPy+RorzfGb4MNcW6dIjHc+La5ziLDfyuGqD3ZqzuIM53pI3dHgS
qdQ/TWa94MpM85KuicZjFOoJX/NMiw2t1BEiZ2oppl387TkOJdbtjYZFeaOomugF
rqR8jFkANxFySypRBuQtHRh4hCTPPa2QO5qouAqIKJg/sAU0yNziz2bHtOKcEKt8
wWtU7H+UwYMn4OusVvAwJuviGqGHIlDji4raoeIyHwZdrXegHFmeXPDMoTpczPG4
xRlHuJukgTonwKoruBXKtRlDMyy7tMg4duDVqMgbRgNJSgWkTzAvrIHuCsLmcA2Q
8X3qdwLz7Wz4QrHtImrD1lYrgFTOhGXR4q4tUegJhoblR1GwDYge1iAyNTWOiswJ
QSGq+OYHre6ISDWP0AD2dKjZsm4/8ybPt5IS6UCmIoK9Hc1LR0IIhdJTfOZekD74
n9W3P5PJ71S2wDMI5A93JrXN2MrmzLBO1eEp/aSaagQHI18+gs6tesjzkCJz71Ch
K7QxyH951tWg+lseLI9dI2GrFf0FFxdMuoQrw0SvbVG44P/iDr1FklYICFFy3spc
e0Rsa1Y3bW1yuwRggGlo96f3b1FFDtYjn5yCz0rLm5Ei28B1kBYUAWm4MDlyJMUE
GnIFnyzWsWruc9MFIZTULaKc7h0ng5BXJMqQ9ZSBm0wEAEMplU9kA1mPhUXdJn3T
i621I0Vp6SrotxcszbpxMpZwClW0eZB7NmtkQY6OfTFGVSRQl2KMJxUbAXDcMua3
q1nCA+7nH90DpTTcf8fg51y4lGaapN5xgPCkLVvj3G07s4XfCUx54y1xyjPAN8tm
E+rTetFBGwWfTdcqPrmwuMV1AHCTie3tt1hk/jbIt1PV+vBfyaSihiS8DCz6JJjc
CY4HWSa+48nJmZqGNNxSC3An7zCfv/wJUn7reoZVOnuhBD5E3K+GbQ2MfwiR2PIS
Bdds3AKdrYjRhDoSk3QBto8t6nC1MV3ma1owbkW1fgybhCAUfHJlabRwBIqdAx1x
8OW/PxZuFFeT7b6E/8pkcO0X41oWv30XCffiULTf0MSbQai1f3Cx/7RDGZ5c+Ur9
+7fIjqW2cGjtniG3PunbJXF4x7HZxGYOvN4CfwECpSkijSQAV9tFlIi1X+YVhsck
vMFPsja1FEbPaJ2hORcvusyQKtTCz6t6fvPXpKqEUMz36fxEk3VPhZYpZQJd5OoD
Rnow0wPS1Q9gsW+3MKFRe+WkMAwT41zdLBbjZttqc6cnLTCFIxPP6/XkdW/op5ZA
5/vgMkkqSxo/yOfi6GyqWlTq4s6TolpPX+FURgIpJPm3EkeHjslgsNWHcdm8TciS
7cRHzsAZ7B/E1VGkQGtB9UTRnf0GV5CGB1hBsl1ng4zjN3fheVDucBHfw5OSWhQs
ML9mfN7w/Vnqof7JMBml/PfzB9JyYV9jT52LoojEWH2d5sM1WdGlR96/9I7k9ZTx
RYqt+FGWrK9TWkzBFI1sXU8wtUOX/jAq3SgyAemy3Dg8o9xgUfxQCkhQWlPdJtkf
nCyaSWoGkHuHXW/QwGrWPYyNao64IUfNaWRYW5bFTy/XvUWMxFO0O9vbczOiDv6U
8KkS9wnzAVmDQFrOJ7TakcxjhnGYmbA2hOIOK7BuLSOv0vA2AlDEdmS26ODoOU+a
JXFoBkudz1NnJWGDMmVuFCJkqXbj7rm2Yd6wg4tnKk3G3ZVQP5ekpOCeyU0o3Yaf
8U/uXw61uu253l5SPqMgE/BhwuHiZq8B23UwEgviWREnI577W5jYbcnBoFHSp1YI
pUlo0MZH78bu/X1ldxtZm4ShsINViG4l9NUSKBlu58htpRepTYa5jrWlK1pgBqd/
qxdhlaF7ZgMfEry83q5gcOEOQw9JesMuqLW466yAFlLdjUvQxnCnNzjfg3FQO26/
UQwpvLdjYFQRb6coHYpr3FtryVm2381DcsV9GnQJmoG34MvyBC82L9Vn1FJpnyHm
NCpg0OXoo54PjDjtYDd2c9Mo2TWd8VTvvFgjCHnqgy+24X2QElBJT0+Z9Dtpme3D
FwLc3xtYYqVRDRAiV4FFqpUYlnxnqwI38CxbbAhCVUExSknQ0oGVXGwqkwP11bjC
KPMgTld2eQrkPlQDTac9tzmqLL2I0GoZwiR5m/JobCpTR8Iy/XmOig5xLXWi8VVx
kIYzNrYumhi2mN6ZKcuQhzovpTHyhrCtv81OJGy06NLrljlBY6VK/oIv4MMw1Wtc
x67EqiotCBHbnVaO7/b6rO21HxkdmaXXO/lWmBiLY0CVbcI7FGGvEAnOPQ1ZB6Oe
cQ48kIaNCBA/X6NW4HsJrkQNICKJRWY8iDJoJ4HXvFaR2ZT8hNbjFNoq597zli9U
0zqqw4qb47rayi/nw9BtMHD2+PGClFyoRRlkMZpz24AMW5bnYOkVQgyJtLvfH+3u
7UXy0qK5MrBsxBMs207Jq7bxNByjWqcYbDLjJiVA8FYFWsm9qNpk/BXeTSsgHAAu
1wdfKxjw3Dolnn8Ub3ihA2utweykrPzv+Dr0FvnPbjBYftYG5PoInMJKUoXEJ9N+
dWmVWhrOTZqqT/2wIys3Lfo3j4EvhrDnvgGAvM9o2Ffg/Ob+9b+DxAL6t2zfk0Si
YGZvpOBoiqFEssxz605wcHucQmPg9fpri2b5pAioWzSbfB8VZTn+TpkAW2hlbRrs
RvHZbITp46gUdW73JcvR7N0yNDFhlnlRoChT1g3cpcrNMisDTct5YyasAVcZh4jz
fO9zTGB+JpeyNQnwMlHmpZAcp2eeF1dRXPAXIdgAiU4hrsDDvqDL5bFlZ7f/M5yj
MKe4CHkm3njDZjt8kBvzToTmE5FQZyIzhHMyxkF8dRlZzquPQQDuepOlP/7dlean
Zpc9lhtdObE6p5YKAieXzmpXxH8FI57O7R2nfBdVB5Gy1HVMksYLLlTeDlUp1/kE
yk8sBzgzUfaWfUdkC0HLE+DrDXKvBkoeJduP4i6wx79MTVVHTQlR8u5Y1DFqq0z0
LsYU6c3weFpqbKN2fSHfAZ0n1OJJpAB2+G1IcHl/jsKKBLXxHhXrjOND8bskx9t9
SOovuY9PyUgrqk315sJZ5++vDONdg/EX1xbg72Qk63VgY1/ZneC5FBzOoGk32RuF
i5sMRudwjm2SS6IxWQSRqFwZK3+xiQU9eqV560v7JyBvcmajzeorX1CeE9JBusom
hp2ffFQWwxj2/8Mj0p4eV6hKKKkPlDLz0dg3x9gLSgJF4pXF9uqIztNrkwJuBUKr
f75W5yjxzDptZPDCecPx17ypGcUH1SSUaJ1vqvbj+FDIuer8J9uOebLhryfqifAT
GP4LkZ4lVPv/yP/bfPDYOl8FsyuWipUj6xD945R7Lzg/gQIcL1Lw9CgEbRPRtGnt
OqVJs3WEx7KQDf4Bc3K7U28w3hBIxsJeb/e94jIr4XLTP51eR9AyroOmzPP2ZuYH
VblM6uTBwVaou7x+seWuRybCzBhUkqA7rve+jlIxAAxE2/oocbQpHmJCrz09H+mb
W/Vui9zaDSldkivKb+zzL5tOS3OV4SIZBMOMbiWsYWFfAh1CaDgr43iZ6fzOfdgq
LFDDaAcWtXSxnnNIqwoQl1ygnUU1OY366BnvHHfj3OGphAJGKnEgugAyaWrlmSj7
YPPsvm6f/xvkvDIwktoeVoByiVOyKyxBDIpLN+rYfmnFIVXO16KP8u05ZKr38PtV
WebSjeYVcePJU6hflGwUwrQBf7hYHbrXkzB7OiMEtbTtrWI61EsMgvyT8YZ9L1hs
b9OlDJRbDdR4mBoRMnEiMIufW/VponPizPO5A6jzX6XekVLMavs3VSLm2lCAz6Db
jVQzgGCfxi2lgHTcwWVpzLrd7WEOtJxm3k4PKtk480TfOwSzhuxzOYK8vR2b8Le+
mIUtaYSJQ18bHqpZcuoE9031kDNEjbBdElxG82yJsRcTRQMMIcSZ02lUytuNeB0h
wK5XquqrdWz0VF3uvCcarSUB+6cNCiK1nUx1XJnxiay2WHxSp80E5pVRFK5m1F1G
IiT2iFjSS6oeNTMfRDFu35KHdqJ6WPXfkpaGmHLTcOMUv0p2qfG9w/hjrvhR4/bA
aoMc3Sh4SJmXSO/VYCU/tghpku3OK8mvMRCwMTKjiuB6iNBuowmiLgNCTvSGd5pZ
mcBAWvyTXVaM2lxmY2R7sztk3MLIVDFjsaSy5nHKZ2eO06n5A+mLXKQH0TW0FOSL
gtcRhF28oSmtx/hO0iDB1ze6zEAmFxVdtMoUrQBHaXqY2g2b+SwGjrlybHIq0yp2
nBkJXmL/fGGM8ntoUtW/nM7xYrfMDrp27cu6Mt8rpSFLlWV/ZM9hJsvJwoIiXyjf
FxBTCgrfbsIGAFAtgT/JsDuVNCX5xF+tA1MNyfWcThDdq3Nbp2+iSxCXjAL+9Hnu
I1BzAozAaykAvVsIj1JqtYO0zyX17HnoEav+5XlJCB2nPxdzIfGAA68dFNa9g5J5
cv+5LTOHnGXVawrl9BmlkF9Ywat1bSD7jB0Fgwqj7PSxcfNImRmx+T/+hyV45zUe
MpAV3kJnUnnrwHsjtPe4UT+tQG+gHQWyplgJ8dRE8ngZJaw18S639ldFkuhjGF/w
GIrvBYw2ATw+GuX5JQNGdTh/2iwyrTxZ4I5hvLSO/Ly8WtXLJBRJ8SqBQnmvTDSM
2y0hoxVhtm7RrXk3NhCOa49nnmBL2DT/ccEyNiadrEXkGo5KlFQoXIUOl4L5Oe6J
M0cQ9YAohbZfVkwBddnufnzw26qL/nSKAwz+wmFFugZ5DnkhcHNG+KSCO7eAVG0Q
avRT2G9Yd3MxJH3N30srbq1dk3UdRxL+iPLse3eHnQ6zK0xuOdFIEVqbG740kzLi
NNiEsC7B0OnLkgtCjDoWw1RXo1oZRF237nvaMvQfLkFPGPV1WvCAq0Jy5bTreih0
T+rQAoCWvfeQrkLNV8Eln0N+XfU07kkNrGP5TiNbmYbVSZRzPduXz9UODBHMZZjp
wlJu1WsF/MV/1Cam1U1/AJhZIm7X5fxmy8Pu4LIto1CoU2V6LcModhWLdALepbab
6u/cAA85/KBMUESRmlKvxyy37dkM7RqwpBV9nJ1jmSBemlYgjCsQWmqGb6CgvSCv
Mb2uiu8+7eDLYvfNdtyiEw6Jj0LNXIsrjbwea2nzEdH/ZwWlpirk+btftehuDs7E
UNfCIpZXYSRbnc0mchycP7g18habymTVu0CqsJXQF1oG1q2TElMoZlVGO4lAFhAA
9AZ9GcCjGCzF68+kbtmy2nRM3Z8I83t+sS4kX7zQB/8mLGI8DigONaWkWEnLnWCt
VM0vqVI0RAfaIloh/zVPHjmhRzI0BlonHdiWyRqenCXQUZ3DdpLlJ4hRY2WPKtg1
pZPMw+ZMXqrakouJ/lR+AGeZP7brHH47qm/7lLeKZjCX7G7+8KLXdkeTfXc7+irs
KAmZQdi6PciA6/jnvMGIP50jSrkIZXTjQ7AGFeCbb4YIPkWZgWhXRnabVgSnK2iy
D2CbqblxGXYMNIE2G6OwV/VlYrlG0HcUi3dCTflR75l2kKG7pUAXF/ziK/PVcCKV
z2o/mBsKF4U2EtmbLVwHsYTBLrZhigFBVfhcO8q1KCE7YHZQ4AFhcVg3SgT2mqGs
r54sZMjc+mpOrM2u1zdi2nZg5D/+BUe8EzumJ/RX1pZMM/yp0mTlXIWLJw67nwC4
VnJ6EJQSBgKfOSxE548KE3kk/lpysqUdpYMAMayHMVtyNvFA+IIZWk+qtbv1B3R4
J4zy8Lfp1QB7I41ZLQNLOwymEeLz6xuj2KK1EAnTuOjLzJaWfH256uVG+LcOurH3
+XGtQwj7A9PDZgs2j2Iwt8/CcCSTSQMNig6lXL7QqmI3CGxygr4tIvqUgwRwQ1YA
Im33II49/m85yIbHl/it6F1K6m9nAhOPbApMi+VhiuNS9HdReGHiNWHm09cHzFTh
oQtLy+2zf3LrrFtp2tVb4tQNb60RNBYuIc/6LrqoMQIkJkmM0JL8Tms79WLUqXiS
kmYpkevvXxcPeiSaIiVS3d7aEpcplridK+/Wxbx+GmHzvxKAYJ4FMOIrI8ZzaXrc
pwAxrC8zmIFCXV1Cxcb0N8Q4ClBm8PkebGxUcYNug9hUGHskHTNO/vgjkvfhWMme
wog6WOBGcIbA8yPj86EwcNhwUbiS8OGuPhbz/QaN4wz+lX4BDtrSYy3C2zSKajLJ
fiulXx/qu7MYECd9KsiLVz7ZgP/O63shSoBJiMygbtBnk+TRKKgs4wyGe1gEzu/I
G0EWs2qyHMNn1eAtaOp2ThLCreSZP4iJKSOTpbJ6yWN5FX5+zVao26sxXnKpgbea
BYv9BMiLOtSiiuInb+TzrTZbf/nOMlnJIjyKqTLRTSAV3F5NcNkgmf/5/lG5U8gU
YWEwEjh+dNFzQOsHzDrMJzMdyIJ/ptKKVEPRuM/XNMsgCMP79e4a9UUHQ4q1yx/+
gX+Uj+87lDVW5GEO3tXfaHHJ9IefOI9LhUyH8NOix4uYzHohC7FKB97BzeCf9mGh
78oqP75uE88C1n9bSrNKRJsaf7xtg6d/lzO6xsSiQxbF8cOomzy3Xvuqd67P1Y6N
l8lXum0m0/vvJ5Y+Jms/Wflagj5z/KKj+BJP9AXckK/IBra/Hd719Ou8bCcR6lrz
CWv5Q/lG2FvVCY3nfxsRcCqkHe63uSbCmcyhRAHFmmcqVKHLkU4AwHSQmqsHctCS
TC4dz+9MO/8Zjosy+KoiKuHDIdgYkNo0/nIVmmAIAwFARsic9kugY0pQ76GyHPy4
mJ1lyfyhCXMIxef0F4gkdnUiWJgncfqb77YrFaCp+Ia0exczATkJf+WzIy/0Cqpm
d68Al2t2rLNUVFrwvJZLBOO0+4APuytlcx/JHGWZ4l7Cnqrd9YFCrbw5w+bufqXk
wyDBlXHfOPXE44WfhjNtIePkr2uHav4Zu5Yg72X+sE+Y7/gQcBKvG5j7RU18ukjj
S3y03toVI+OvB+excEb3wRYrRwhlLyGlpPtd4OYJkItdHg7TISl7Eyv3XSUdhAY4
7KdF9ab6mW/ai0dKZB5jSH1bQuodB7K/P/+BZDBJ9OhPmrYMtipR4OZG3uwecB02
2PzYWf28HU2rpP+xdEr1zFY1tY2Q9LwibzVvi7N5BW8sXPUBCGMRR5mleVpiiWjQ
RXuXotpqdK56fPz6TNhyFVfgYyCaXA/yXMyl+iKBKXLe6Yw8CiWaIpA/qsW4CO7I
fuFWbNc/gW2WUoXZ1qB4ZIP0dtGxuQLXuAxah45+eLYNZ4vBhk4i6S0ob2aFaWR2
uKtN/pDrMQI69cnsKj6APNnYIGnLt1AU/obmPx3Bb6LzdnK/rRDEmWkQ8JDWhuCJ
iU5hu7FJ3iyxhoCONtwI85aIS79E9T0DTxmbnSPayW0tWRVoV4/Z7HAhtyB9j7Iz
6OUg8FRSJVSqlfTLOljKFy0FlMA7lA41G4diFb6OoqrQOSE8wLsRTTEJdz9irjHq
DlSZNNkeF8oI+dCwxtTHWpWg8NOpTg+ayPOR7xj0Hl53huXuf1BAIq8kFTuM4oWI
sGAwBijIo+zyOwf02B46w9NSGX1R/0SXY3XFB7Lwf3aLZVqP+ueLZB67EJrSAGm9
2RHzkwKWCzN8SBsurqodiufOlQWrc6KVK3IIeNDgQ6znPl761WK8m9WqHXgIwCi0
G0Ex8AZbf1onXlkTlQSuv8Z8dJLFF7cSWzfPuSmzlYbvqHHZiDYw8l3Qvh/47IBH
JCK0ger3vOjNS9SPbl9g2cTEMolO+IYVpjMOFRPHR4PlyzGpaUKT1ZUmkkxdBDfY
zWoZaQzqHxRcCUyxeCV7R1MgZj5qf5NPGG9q7a01ltQLiMNXd/vsE2N2Q0rp4TTj
kpRvrZpchqJyx+5KMiX5Zjbk4jh/EUCJq5LQRwjQxPCEXIX1lZqAohv5EmedtV5B
yIEnFcKO7xZVGFcmKEFjte+hnIkVyvevuC7JQMZw2RwI3BISV15bGAx5zWko3jj8
S5DGkq0zh8d+6Ags+0uETWkVLJbnf50nPmenDDJNVyagrRFYUq6oxIQnG4LwEJ82
9KthEhU4bCPeGi0uT1ERQbB67rb+kXse5dwdrY+BUTHz3FKHk0MwqSj71CuI0pGX
ESX6curU+WBhchJfdfCcCWYMH1CnQ5MZhsUQvo391SXLeCCUZPBrbeDCyXyCEEn6
OQU9jzn3rzHXZc6gwUciejjp7XugqLKd9e++xxRHYPPasAb2LWIjHu3H8cBs5kuR
THW0lqufQOBlVrNK+cP+wPXlIgYww9KvIH5afyD9xH0nwY0gZW9lEjZDBT35a2up
YX3pydmZRWiDaNxJW2nGcHlUfi2vtLynJfnCWPoFiapKJzSb8dS9g6tLXs5CorKC
/GrKl6K+iTfN4VRwyT96FQnTnrCD/PcE3zvvg7g+s/lTG9BgTQM7fZktA8CxjwSn
Y7gYFWvxViWHObPopITBaejakZzLhRlQP5vyhoN4sNGKI0l2/pWqv0BX+oINAZzQ
6hsrdHG9ajk30CMFyldr3hxOVAq1O1ZiqKgIiRWgu3BVT2Bpd6g41XOy7tM+5ivi
QClZDOl697Pr8eQL7zuv6mNi3jw7x75xXxYbNBNbQOeLVRUBCQpaFKT8GcwOJrAl
WU3rul2TuwBY8EdpFHou6kH5RGgCgE3fxn6Gnm1Q++NClJT52JT4ORelSbldi1Vc
BAyJ3BUL2Qq/UwdkxUVGKsktBROnylYe+YDEKcVDWSF7ltDgec1a9s2APmt0ZDHh
WSp1vBuRt8bUdAMtCgfik3Ae08Iew6sb55EnbZpzZbU//N73e49j8mO5HoVWKRlB
n6JrjEdhiGR3W1vYdymkHJbXEJDbVJXJwQAqUlwqWl68/vo4vtBCWUEngn6SP4Vr
X8/uB9VNgXnpyyScHBb6Q+xTrG7J5OgvDm9mUxYUHfQYCn8PAaUfBnVcO0LhBF/X
N/2cyOjw/4+MhnVXcrk+gOdV9fuio3DKjH5vKZpQ0y0cgeVcmO3LOFUD1BHonkar
PYPaxrETLZa866ub/sjOWzAMVQRkC/ZdaoN/lszTNr4fLQ1sceH5PWiBLAYD1pKR
BV03eX0qrMm1b/1ZTNmGBsAXmLF1gBSYDwUQ1JzvVQ3ZuIGu0XCStiFKbmCMWHFi
K/odPzNU+mlSSO7hz+GFhN/ivSMgVvOFGMNHVU3HNHTYAl6K50ViF2yKPyO2Z6CA
ZdkZV74FqdoXs0Wsxwm9Q5qwoDqFobAie1vf9NIdPEOa8s9LbcgCR3+VtleU8fRc
bGlN6Ln+mOmoy8SEsHpSVGqChboFUS9NpxWPkABVF36CHVq27OfmUZD4frpsnh5S
DRb5uLJSW4OH5Ae6z0c5YJ/qyYLIZHRDdtjXJEEtVOekI996MpY4hvktLFY77zRr
b3ZwU0yDOqRykryX4D+vdG+gALJzDjEqGNu5SnflO1N9e4q7dvh8H1ubGx3+O2ZW
tIJN5nDwBP2Cha1rd4klsAP0GYbJZrhprZXsPJMMCHdMsqSnzka1qfjt5jW2nKIh
/WPhHN84quoAJz58L5PibePG2kbfbAiIUr6PauMXrJAYQ6PkGiV4eCEmN5p8OFGU
wuJY86gQ9MfhNRW6QMXTmN8Xaf+SBcY1/q9bzyfaUox/9gHGnSv+T3gHGAxmKZtk
a5gqa3JxePTw+SfYxxfkJ5LYgrUbji1V3ePDOztYtrhFekRzXtLQyQiHpp/HK2a/
GqfgIR84s2AjzI9lSwrpdTKtqLz211zBZ+F5NlMRWzD4thJcxn9sQEQvMrGvxtBs
ajtlN4cAYiUmQ7by71mYMAOUKQ2mK0WSs2Hd0gQ37eBvMns+AVE3rrXXV86bcB2e
TjEaaTHTM5BGuJYGycCi6GJHCGJoYVt0oFX4NmirtEcGy/y6kNV13XYkNcBKvO+a
KnWHjQoNgXNXAgXWVVDIaUYutN5Dqt+DT1k2bCZzZod5lvhoTqNln1EVaiN19coe
Obl0CW0ojXH5OnU0GSRQlYZy3IEi7hHgXgOBnaiWgU9LDMkUaGVj2w0CkhbijBn/
heHliYsaootNIG9b6FBoqKHu6HGEqrJHdE4ods1bW8RgPxvHC1R7yeBA+7v73UWp
NUl7YA+NoPswIb4ICFcyrOwSthNBPUBIh86sEDQ9WY4Kx5/LGhoyGdjXCYa9wHgS
MPZ6EY4o8qhPqBJU4pRjFAVz9yqXkIGDFH+8jdaAW/VOisoiJ3ZeeyFf/dRe7f9v
71Xm4oACi2OL1EG5B5LYb6O8GMXXA2kC6OG+8jO/KTbuxsQ1399u1OOJ2vmSo+e6
g7K93T69MWlDClt4jah+0820Hp7oSiKUlFF0JB65dpY1FtYnfIsBWbtlFUgIN7T9
wl8GOqIDPt6iiFAVQE6E1ycKsW7UT6TYlM46rz3FF4VwdUlL1X58N1KK3ittIEo1
64njxN+h0TOYL2q6DlFnGcHEzGe+GlhYDgIUdXoPT09Yy44OH7KnvF8d7EU5VQ2B
nBojfkztOj8nY04lK9uX/DuJdwE1JQvxsGKqjV47vHUP9wdJ2u/i0J0yyjnakFOh
xRYXlOnYsQ+2EuZaKhSvbuOavXm2rRh8YrTJYXfEkRlgnGsy522vmXCEn4MwI7dt
6L4rJnQpzUJdux2ZzRDnmBBrbr27h8zzMEuAN1qlBFMMufN3SKIYWuGOU1ARd5wP
98+8kT4oMQfgbfKceBWlm2a826+efnOe3Kkg4texblkfE3LJpWoy4OYBSMSGH6+A
rO4QRRMFstkhj/nNDCnz4DnJMfkRiAtAgwvXsZ1E5j0lS7kC2xBkr/V76F2L+TA3
78HLtskgHEZg+raYLpXEad7v0IhooHwRKNlfdLOw3PYYLFI4WA2rPEF8sZ6v10Wt
MuUFxN36y2XTfuiIFbfWm7/X++/AIlwUvfttTZg4XnZ1md46IerXsMjb98eI4R6H
cxYMMAlHcqjqPJmLdFnczO2K00d1PFACi8YvyCj43UPJGwZIagLryP8M3d1LBxGC
wJPz4OnGvrnYlNZxt1OFXFL7j865GcglfD85IrbmkXGG7kc6PG5JbiQ3rzLDo+FD
NUBarzKrC3MUiEazLstUAw8BHzOGj3BHh270ZVlXss7Wd7qtJE7XS5mJ5sVsV416
/1evrt4amPJTHJ6e6xe6gT4kcPwyKqrdks7wkk7sFtlrHzAKYG/DaBf8GOUJFcql
vtJhqY5h3kc8fzr6PLkCVwct/COV/9xfmJLvfYs2YFNbQD9S8JIKLgtaba+bKIm2
AwylTFCVBfTwyfxs7/4OMkKdS8VXTGdvtKv4vXrz5EfASxzbjtwt6ghm+pNjYXnV
d6TiXfF4ep7+vwr8XOqZalbwIxwRoSPZ8NrfkA1Ssjq6aqN8XnSz+4H75vEzPXtZ
QOoPrA1Kyua6hlsuyESzjltjs9g0g18GWjCbsOxohmggGLNPJb0T3ieQczR1xDQS
ULxRy7/N5yAgLGTwi3NJdKMUt4I0VDIRe+Fn8C+hFEMOdyJnQ6pUkTMmu6i5oEPj
BPTK6qnPWiOi3Ynf4DndMPfpuM8kWhm42voytrwMKknb+u5taOvNWmNdF2Cd3JTm
9W/739j9CvizteEpZcDhDOeOHIhY5gvazXQReOk6MTZvEWOA5NTrS+60XS1GUN1a
FGCGqXJX4TZ6T2JMeQfo5/eksmbLt/RYH84HDtoZPF7j1Bkl3KRC/6z4wjnyRk+K
gcYunDbWJWFx+Sxx7byXCDH6DG8YVA8aFardaO+zbFbgdxrY9oXadiZOwLCzJOIU
YSwXhfgkZ/KH+8kws8Bd5/i2mv/x3pboKG1XdKmA/IUNJ703P0CDsqznSIGEon4l
8azi6kGZv4l3+owa2Hm0ao5jkov4DAhVBSRrR+YNc4Eg32UaskvRnX/pwNrnIjso
JNurBuokmVZpD9BKgod6qa1qmIG5asauNLIrun5zo1h5OaiUOMZwCQ9LYC8OCkyj
v0R6gczQdFW1Yz/yqS7Ce3nBpXVC805HhkY7BdTmMYNOfmCPhatnSm6WYMMBnhil
P5ho781wiby5uhfn8WL1YMKBYVgBnQcsy4OhV1d3Dm4crwIj9FuE6L3R4dn/j8MF
25NkL8dE40QK454C4dXIWbn1E4r9sVzTWrWqndxofDODGVJRr6dFcrPbMPV062/u
MbZGqrC3LY8MLTSKfjFvgEUEuaSVIhGjyIjxyteByIIF+/CqWMDrqbZL2ihpu+eX
uusJXNqpQHVax0YmPJMnEzZKy9NZtusShvFlNKzqvHvTYeI4i7/d0dut5NbCWDXd
5qsFqRu55FdnW0WiogASTbIxgtubjPvubRzJoFj/ZenBkJkeOGEzIGcjlnwKu/pP
V3JWNywihC73bHFjRkGGFZInso4Rs81b32vqZzHdFt6wixvAsPSsm8evuxO1z6gz
a+Za4DF4VTd7DZ7f08ouag5npPARgjsDiLoQ6IOZXrS2+8BRBJkUoPOI9QTYq3Ae
IdAn1jvSr8FCKFhuv+J6VjCPSgoY37IXKfhnZK1arWdjXS3TpeKexn2pqrnD9C4T
j82d6W9wUYSGvnzSWK6RXwgSxOtc5jlyRgVTjoTNWYo/pIINAHfHlTw82Ygi0H6L
ZixNh6LXEfOOSrXeDiBZpLehCnuY3RwndcA9ISZ/Z7Tgq/ZIEy89hk9xQk6s+YaX
FcU9zCe+X5UbikQ78a7hDU2a9jAw1QyhqO0nGFYAuoPcxNb9HuRvzp8XCyg1Lo6S
J13RL6pNccluJRrrV15Ss/YEgB1Rn+YREcS30pLcq1GZGkgn4O3Sb6UtzB2fg3NP
BBl0UdzZxp7lys5bsFMn3goQjplAwa+CPqfSzXkEYInDK7n92QUhfll4d6246BXY
KDXfkh5qfIb3WlkL+l8I4G578kTFnfSH/RjMpU+dp2yyg+sxGuFRBbcnTuvh7Wn7
zLi7b/TFEZ45RS+PQAC0Ck5e3tc7rkfThCGZLdBAHvY+2Fl3Tt8/bm9V3W+EMUGk
HTS2fasJfgWaJyzWnz1FubboFL4bSE5gtDW4MP43q6iKqG2EL8PjawVJMVN/mgHH
1gK9gM+4dgOFK13RTq2+DEpeJLWPHjKTy/JGdIFhLzWM866LMxVz66+YF6y6OyLT
SYZGqDdUT21yKJvPgNo7+tB8yE25i8Q/Bbch+/tGewU/oILOYtCjmg42uC2GUNMA
ohDU2U2mZ6E26FJq17d2odAbPcvzhurv/pIrSux/XSdPYG24L+yqQi58G0jmR5T9
lp7h44tiVPWQ5hjnhpWSvBsJZRQ8qk3OwYESekRv3hmQ8iiAbDK43HUUWovr+ZNy
X7DH9m/sB3QXgwTxCI8EmCLlbh+waBN3LI0ojzkkNqBKbcNCZ+O+GemS9gssYINn
XEBMPH0AC72+TrFl+b+ju+6L0nSlcq+aZtdhms0AV3bLtbfQ0ETmxIs2JvQFuz1f
Qj+kM/dOX66sydZJQ5SuOukUmgnHYaRar+vwzceUGb5RB+cZEK1px5rlEUCrDHoW
3vq84tYIIw12L//wM47nCN5XkzJMcdEW9VC4jgpkIYjzhO80DcdZUa+019f++lfQ
s+bF32jLRPBTwTi90mblhpuqPq4DuDXfqoLprf7HrMWfIhHDIyeKWAFsnyLFHRyo
+xvys4n6b4XJCPi0kzXN4WX7p8bWUkB7Yf/OyjT0d4RdzKoX56GmU9R6sxejxYKh
BP7kgBVjb4nGLk44nPVbCZZBuafxs4YVvQjFXJIIFzzX2kQxuT/mX4IzScVvN2KM
zBVYcqZ+Zoy/l6HlD9S893I/NsIe5bdTSK8EhUUK58Tv7vDzTpeBJs740iycMBBm
03VKZwEg4d4Ry1qkdWNEgdRc7pF4X2VRlbPY1+GjyaEOxs2G60sYWl60plJA3u9a
D0JKRvrTbaKAweQQEPx9kTXLRHL/d+gvbrq/ojJ/NT/88lPciEq9tQD591BRvqo0
DelNfNFQ0cBlNzkSendmN8wCVWriPkzSMvVwQg6+zqsx3k6lpMXlpqdeWnLEeXDA
udm5ETcBeWWv0OHFcEOIi2TwSXHlCW985tOMegR+QMCPclZCrvEab+8yLk/7ejFr
DjqvGG6uY4+oAb3jbZqxct0bEo45pXNovw13AmQYhROcygpH66WfQ2BJcqX3wcIZ
bJR1o6CsXyWl2rQ2X5XDppR29Yk43yfofriE4PkwTMtbLiwyY+q+/5kxxViTi0Xu
GLPU0fWqYmjUNi8acaBAuWbsGMz0I5iimfWucaqtU8+R/8f3MEg3jOt1a45wUexY
LY7hDkjqgbIG6W+Z1WrBwkp0c+e84c91GYh2dEqJQ30osNt2r0kIq69fd9YeP1a+
edk/5pcQDFTAbTI7ZeHUGvkapm4tu/kZtmebhrK+PsI3HANzGBuAsOuFxrfd+Sr/
HosT6rvMjGXOo6+w2repaf/HD/nFy1fiwrs0NxXPY54b/vGPx6j8yg+ZGJjBDlC9
IGG2iOaeV2sVd1o3jp3qi7bAJFdvZBF4uO8yk92jcQ54Q2/TBGPA8who8VIX5bwf
V4ONMQ2iPfZ4Nqq4i4v0oqjlF3qIaIuoNP2XxUlSviyacfEPwC+kM3Z0kas1Uejz
KHGMPb0u21QpIKJackiXCVXjkqa1TWQxdtGJzWOaIrs+ptmKI/7qfx7rOOLICblW
98hC8awXNS4APHK7ZS8R7Xg4cH2dETCzce2melczbsZYKtqn9LzEzccpcGVOIQnB
LBZQ31HgNoOoQEwFEGm6JRoZqXQpuW+QAFsbrepoJKK/GDTuhwRU/Y+PxCpR2eyW
zlmWb+DgfRPdiBelMDhqKlJFJvwRFGXqlslJq8k3QHjUC45inZSYVBVv9ouLHM+E
sHek5mRiuIj/Bf9SA2JJdfKmrXQQDLcr3DgLHqm4Ku2ITKRC3MuXuH6xpq98S57G
uTzalyBC52142Yc+1hcYES8oKB44SJKeq3Ynf2sa1skL1iA5ygAzNhLJEyFS2zsW
e4Rm6+Hn0v39opGO3FHxMLjmEL/ty7TF0WgBdlG0v73+HLHwSQpT6+drisbNqnfV
+CAXBDdK102ASt+GDbaES4iDa259Wwat5y/86OuTOkVEX3vYO63ubnsv/2oD6IR+
mDxsAjHlqfhJBf5Ai95mZR4hdrxUdOZqHgc3j39Iq6+lZUdLC+28VjwSx3gGuGtg
YzTy8fgmU+bC71c3zfPjGOR+lIrlogCrrY+LINe0yqyEAiAY62Mn+9ccW2nEvtpD
9c9LslvjvKc/rgATfWqH8kF9h0GOnxYQ9fCrXpPv5PrX/0wP+1fW9wOPVGx/jREA
nYxJAeJQong4sTSl+38VU5jpR+5aUqVkmOeRZOUHPmQ1yJyrd7SKa9I6VZLBUXC0
+4pCASMnrSQXEHfNWwu1faU9KTa8+rE4zEohzP0Se/W8LSmjlNFQS66J0P0dJ66n
4sleR8dcJePZGoeoV+Yp1Sz9OyTjhKXxkfLBShfqm0UfIBVta4E6A4s75Ykc14N2
gEsQd9IdJ3pD0FK/OADJK9n0ctfkoQGbuid+opy9NgOdTGKlscNgQdNzITuFm9BT
l07nDvOauY/aaYB4EVuh99lw9rfgMqpYAz1hOVT4MWidEZ8HtDxr+lHh9/L0m8Gr
1D6FqfdeWGJO3wWD18RXrFQbEgnSIhAA2iWWft4T+AnHDi6dATvFJKpBM4f5n/3U
ZAj+7/mwrvqbgTcHHhuMx+Diy+GvaIa+g5s+uotdimbZlnWF6MGAv0yN5a7C9OKT
Jwlu67/EL1J1aM6LG2JIa36QWt3k5EQlAo4d9xUoiNDy8f4bMVLIohQCv0dewiNa
Mo+YX5cl+8JwSKdW059BaYfH6SWTZgevTGUE5mM4Qf3n0VFsRkluEQgfO25uvOlq
QoQUv2l2tlyK2Z0PazMwFHdCIKRgVjT/GGjNXJHs1tJkXJKWLqvP3rm+gOU2ZsfQ
/Y51n9+36JqINrnm+aeHIOdt2AqtEPB90DUF74hgrUrP2u9FHAgagwLDCoMb46/t
H5xBDOesE105GrUu4tyAMbz8sYMNcA+yCf/Mr7N2JHEhycSso/hl8o0e2/q/pk8D
4PhjeH2woaMLVZ5RdplUYTaHvVCuRgBDNvEr2WcLc/61V2ceScNNviUgz43Dc3kV
xhoF1k4MRnGRj6fnaG5HHvMs7yXdRJSSkM1g/HxCmWYQvDHDa/Q/rptH04nHl+99
EZNSNN1M9S5ZhaMG1b2dZAYFv/+ePuOV1yFilah1GTNnXIB4T2rCdjehmbyxXftk
9es0C+jAmDnDC6z8PY4OjnjpwDhOmSQAi9E+091gjjWFJ6W3mgup2uSsKy0dkGhn
3+cXnYZ9CEmVsDOVj0aRJwTbp1UylstUWbDPifd/lCEjY8pVUeXWqqUfECOqn9QV
e94wnNtFb7en55Ux0NiWKjj2z2sXsE3couv64PI2Y2I+2ctzw1pIOBJflYY+qLpg
MVcNQxx4cfkJ1FS61RU7Q7V45TuhkxdsPPghPQCtwA75dP70Mi/TkZcFFFJ7Wfnp
2NBUM3HCWEexLSMk/ZeSrAfNJX+9q8/1v8OOIRyAD5o+p3s7qeHxU7VnA+a0/xzP
jx10FYYfYAC1HP52YoEfPy41/Y/EYU4QEem3OBRgY4kK7NL1epzRVNodHGmj13/F
QqjodDuwQvTUYPUK2JrksgOcaZ++obGQ0M/62r3o0MPAPQRJUIyMdmtTmbibIuic
OCcrZrzrMJxBpW1EGzSUS7bhaTr4ZVDOLX4dsmAnOqVhqkltoPg93LdKYmyvmtC7
/peY7OovwG9N2apMI2Uzh3qFvoNWrY4JrrBHlDTfEvKiuwfErSkihdj4pd9kf5Ne
YU5oUsd8uyJTUrWsY4XmrMYNau+Ai1xYLcr3pEfkiOKp9J7UGAjKDWaoiQOfDIav
odKRJ5bzelSvn09ePZ7HPrWQks4celWpoMfSUioZiWPQFV/zipujt1WynjFVycLp
+vTQ7Q4pwBwvQDkrCmL0j1z9+1nklLkXvriIMOzrPzRAgLWy+hQRpWkMSfBZpUgN
3XKDtJVj/WJ8AZmwF5BqU3lmd1kfOZVXw4BggJweJkzvhO4HdwXIbnk1IlUBLaJm
gOF6mdIp/mctRrD2f/NdHbKZom7GOuHSG4w0BVsXzofElQhxqEgCXO0pk46GnWP7
HyicarAh9YIpumOxAkBNjaou/yXZB2guq0WTPPjNfrhvqHyRrS6eDz0EDGpNg5WE
YwtfEgjkFt4O/CMfxhdyPVkv0vd4pIOrCDyCNBqDywMBbkjSdXCGtTPI5t/T69aO
khXlkGA9qE77jThkmBCTha2EjvHYMiElYjsqJn/xMHn2XzmbDv5GDlu4jStcyYFy
SpowS5R6VuOSUYCKUiUma/ZMkUVvOkZtoG8gfzk1G2NbEeW9Rq20JFMbiN9c/Lma
A2InVZJodLWJBluupVwrrEYCd4egLV4b7bpspYcUUrt/QeT6oKEJDZjFIUObHcU8
uVGZq7JLIH5YTW7lWHgULUQLzSTmVYCBgrW4bcYvt0sksPqitFrpdZfcOOSKZViA
7L6ErF+s63G9wG4t/4YNNVz/UsVllDcM8flO29YHnG6xciaJDFCT3D9yweBXLaNu
4z6BK/VQTdB0XbDJ/abjeK6ECYRp7UNhJz1aYs8e6+70cAS4CLXX5U+s1yZjfvg9
ZALTCSL76wCahd6goJ9V5yzpzjrtJ0HZI/zY1D8GmjHep9jMfJDzm40T5OX+Unlz
fj+69WmgEQeCkDgNkstTS7zT1ZSh9feOTQr90HMs1yPvh+lP7J+wwM3Nx6ALdL7Z
gvQpmHeeWjMX48r/0/w82ENhujxuPvxJvopaWggW956fqlpbDCwDC1K7uaJMYiUz
a3Atq6QqBcL88jjf6vjad4gmaACZ0PGJrMe2ALv9n4sT2gPIkXXUtdM0YKpIumAJ
77G86Ma8Iom0kjfYA3IGM9e5VJ2GjH8eqIFQflSiRr5RIIZWA9egMldHGFLOY1+/
GEKYbtKcuNXhOIumqSngc/V7jB6ArQBbwpTDyiYXcQFk+TYNPvPB37djjsrRdVE1
Xr2CcZNJNj3VWouzlztacgju2OA8VV1qYc8SLSa6CFIL1tgCu/tErpDnHgjGRDAV
ld/lsFnX1/30fTZl+pgm5YzVX/jcjbeig3pmQh+YXH9/fpF6fY9ZQn5gW91NqbFG
2z7kWSF1ovnf0OlVCU5D8oclWAJXAW0X3+lsuIrsh4E9vXQs4cLtbgJZFSjL5PBR
JqNa/8qsiXg0EPIKdGlGyA7GSya10TRXC1kdhnuZDMK8T9R7qMaOJpHYxViNZZ5B
aCu+0nbO08LDGAk2v8oZxTIKKY6wg8/5+bIaQfmDkeMX29HCYU1xqJiD4VYVaIA/
sTWhqdyuKYc+1AxtmF8kCpp4+2XX1M4pQLbx8HuJ6Zoxk2g2Bvpi7TaRUMmS9Ip5
BsWv+O82GN+6Q5uVi6SHnFd3re/hYFZfeMtx0cO+735zGV6fSio5eWuWqzPb6VWi
rKaw45yXexbWsfbBK6uhANqeev/OegUUZEA0DS8ewnIRKG0Q7d3UqCpi1M4mHY19
8T/zdhHZnxBcDP5oQ+98j33rvRhS+P9TUByDlTtuat36mSJpU0vbltgxsyZeX8c1
253gmvgaIBpg4sFPmoGOoHx0Sr2CLI2wN4EmdFt9bWXcB3eR82BW5EYCPPFk5c1t
Ff5Qq4+AmvijfYCGyRNGD+ONjrisx/ciQneBzyZ/3JhsrapOGjJFPfr6ODYnwQYF
FZxDUk+ct8Dfd76jaodt5EHNkF3sMT5YpY6m0W4B25Png2ZdanPTQVtLUnkc+yYY
v3N59DHE0mY21cOqQM44RnwzOu1N6PkzSRLH6EwA1/ZS8COOUCoCWDHo+ujBgcWP
t5COfU7zoKNs+I9/1dSIYE8+/aQTYk0J8uWbWm6hJPxeqkH0Aahz9I2VchH2UAA2
OGyJudEPN4GRBfO9BFGYW6c//ec0+DuCRttTb47I+j4BSZFtGWwOmckxPZH7FDLB
H1a9QDuDnxDL5Tn0hcV3mHvhr/j+/xu44OqNOE7fjxYLmca9NZP44QaLU3Gu12D8
CbLQQofuNLETEljOboENeCbSmtFKtNfwpTWanndV1qvPMm83jIWhTkGJlVgwt7rl
vZWArOFI0hxqqdI0PhoJnrimzg/Qfzgg0w8a919B+ZjTQQF9TwD18A5AwdgB9rzL
WdwgaaVeAKeIL1U4DGuI2eZZrx7Bc5bxd8T/ygKIWWXsA/Ktrd7PkHUvpXSQMwY7
7yKm4dIe3Gc29dvEPwaFD9iCqbVr9bupHzM7zTYO8Yc0TrtP3V8wA+udeUp+7yNN
9I+uMSyhxxScmlB7GdHTRqBpo8ZUlFhCSxBNrQhQC5Qvx1VeTk7tUjwgvLJMhd4W
+PhgBPrQBGeJcbp+ES+3ZNg8SF6SZye0HMzQ0nr+rjtMZcwVTnG97SwTaeDkpi3c
7dOlYnGxqBxJrsTzF11Zs3YDujvCWazSQeAcTW/Ez3ca0xG6H06SMADSk1EYQE41
tzrfXUqXi1OyY1LaERnnoO/nFAl7Q8da28JerQ0eAgchfKN/Rq2sKfSXtypguVbv
aHOGeTaDXG/g688EDuuNVzlFDzzv2sYTdlBWtmCXpE5/D9hQPn9CKtZB5XD+mzH3
hs4UM5jwvHdcJ8/wuE2pc6sAGYq9RMLi5qMO4Jt4WbIZwWJraje8x7PcGprpqVQx
XcM/ddZIfIYqpkA/OP0k7EPJ2SHrJi/SLhFkvrDCB1NPS35Dna2M1iFojrtc2dEt
KObQK84yLrHXC8MR/f0UDDIO6ZRMV45NABduhwScIHSf0mAv6Hwo11K4mWoK4DNN
HWp22eBb8wKkFlv/ZO2jSXBZoiqfKj+oXnNIW5/3M7jV0Xe3wvoThtGx3q/TusJx
CktXlJL2Osu2jyrvlYXiwSx+JBzUKpCZSeSk6uEDjV22yMtuyJ4btLGWR063fucT
T6FaCkcnZATgffBAsM8J25HnA8ExR+tHqXs9c1SmvmQE3AcCJkzGR/0D2A42nYNq
+Ebf9rjZFUFheXU07VKg+wUUikphcstO0TMxUtsUagkNx4mjjCahhnsvlw/feESn
VHg6D7yHPPvqVXJAQUQ+y2GVQiyyFoXevGpIdHaWGyv9MV9/EMpDIygBTx23OX3c
z/bEOeGoteeb2pF1qvpExUaPytMoKy1P/Agzu76lng8lNszhas3S210DVD2nopRt
YkCWcezuw2ZPgUrKAquvKc6cFfLO83fRM8R65EYvWQ+oI2602jHt0IFT4OXdVq9h
kPquJfxjAKjTI67ECk6QTGlk7rFskxkVgLRb1d2SDzL4JAalKr3dxRd9pDoQ5Kdg
M1kM/Ma0qnpBrjLxPM6GPakvvG/WPlmmU+bVF+mOXoh+KkNtBW2IKZ9np3kJ2qZr
Xn2qKwktr6FP4dp2fow0itco83/weBUvaYEhbuRXxaDKDGshtsKuw6biuJGFhtwM
cf8ffU5dkx/dN1+SNi+el9ofDP2NSNcAGqg40FPshlccmpIrsnEudSIYGTkFxiuK
xECZUcYK1WkvjcFEGF6zbOP2CY6iYlrHxwdLjX15zG9mk62NuLhTBmILUpJIdIk7
JTKteSW6+3TX8LtRShn3Vb7+50Mds8V6c+SL6lR+1gW+b8P1qHEDsJOQF8ciZUr1
pYEsvLzTnrvt9hOoymD7o+yP7XmNQFLvmO+UcTo1/XQAYxvvEdVbQOopezb3AZiE
6misxl4LRFSDrDfujI7HHkmNRT3bC0/DOQpuUKZLqpzr3nBzDQnbxS8l/QsSxtJI
4ve0W8DHkLzrSP8KCVXS54VPnOvwvEl9KUJz3LT94D+YDnbfj36pDOxWdewHKkw0
GSyW4ozp/hUdQ7lj5LfmTZjRo+feVG9GqMbDvn+DFFoFCKKoefgCTCrnkn6q891j
phprYj4R18i4hVtWpiN+2+sKHXsrQPz1q3qf7kDGUzXEQOCII03GJdOSS7EUOEKw
ZSzru7AX2LqsshbYM+t6eGygN9tikyRmoyEEt7J2arud9yYFTgVvTh8C4V7PHiDr
2fFp3IoJNL3GE3L76NFRkTEVCVPBr17FOrAVDrAcnOWLQI+qC/bw7od4IAIrbj5g
JufDTt+mk1PdQ8Z+7ZsVoyxNUBSNDrbRhkV88m7XpPspoB8ewTZeLdNzhR3wpf4F
tBt02cSOASFCING5trk/k/FFHbt23FriVTAubsAJiP42dM1innfMqPHa1RTBWebs
S09Gtje0pGLrnju0ObeYa5PSUcGOIw9uqZ2m5vJNbppVlibFbTJ/S2N6fKFdfvmc
IoFxkJUNSXxU2GAtHDpEokW5+tusnVYx+CBj9E3GdhdC6s++YvxVC0Aply4CALqN
NC0pTGZZ2lbnhkDL3vaYB842cIrov01OGQ2Y/Fbbvf73MA8VOB0fB11E4AAw59wz
K1ptbPBxaH56UD0RDhEWosnlHk/Qw0ZEDTV9vfb0XoK4ponnzc8wx3L89ZyPIWn8
7Xy5NrpMdzi3225Vcw8B/jyoMGvcjxUDXTcfSv4pMBJfVWbmPlzycO/9oa6RS5+q
Fb99S9bOKbcKcNnjK44LqF7YAC5UP+qXEI9hJPGC/FtY3zwTFqLlD1cu0oNuh+B7
CqlhufOvIzHPq7MC2UUOG9XW3fIfTFLlJWifym7XCMzhaFc7R7Ph7W/4c25qqQzu
nPqySJQqr9PSO428WU8eA9+MBMF3De7iNuCwq17BGFaxoqo1e1id2O9x8ww9ZkRg
BdnlnlkuFsneQkFfrKz0a7eIL/krERbjeV2T4gASN7wrSz5XL1dVdlSktf9CeMkU
UvN/OMHY37UKgb4HwglQ0YrEy6QmzAMUJD8Hx7yI0P+eaROCgT1yxsp8x2gzQTL0
RmeHBb9JvmdzPElNdCCkgQ/X/AYzU4KAvsa2la3yhHwshZ5DEJuYudtxRbTUghMH
c0u/klwbLJjz5Kc5MhexGRIQn8E8+yy2gT7o86K9uLA395zyhGFWYTj3noA5kcWh
x/xxTXt0e17pvhBSvOYF0KsYgQYB/so5EGjc80SBihQxoChgvHN24FpL6Ad2bOwO
aUjXaX2qNGsViZlC1gVx+8bU4nEAtwMrCZa4rVnQIgyek6EkXe8eFBYsxvjABjiu
QpH8aMmuoH8kZn+R/dcNDnPzDlPqxLmZkn87b7gVhFiek+6B76zrllh7wCM/DGTu
KSjx8KD9A1zzI05SUJ5LVYIffONARB6tStfZJbe0fvxyqladidPrmHsmtjt0urfH
USFaykCVkHjVbCB5ZuGih62oJlY2qvFKIabxWtYlnA2XC4L/ovd+/tUcodMF+NBi
DYFuZMTIeFFPMZUBal7L6mjtsA9Oa4ee5RU58G0c92fhA06+LxJxTlBc9pPZpOsy
6knUjN4p4AGTwjQvlwI997+dlZsU2Cqw2KiY6we1TmP+JsnWj5TpI5F9RSq4fkyv
dyU55xUbS/O0DoZTE0nZ9QbDJzAf9XQ64hVfEuY6Lq0kgcgr0u/2ETOt0oOVLFjm
8MMERBXFdoNpWuOnCy742cZaQMZUovF/2JgQRFxyAiM0JcSodpLBSld3rwo8X1n8
jCxDcCKmf238dq9oCNHnZW3DYdRKIu+rJSjhXT2Qm/J/oWmm3GPnQAh5N8a9uZKC
XFarOsqYQ1I3NgENl/IhQDmFpT8hrxEH5z5XPdaIDRIF4i7tCgXh0Rw+ysAYdP7e
bVYmznz1gGWc9l0Q2vrptXaDH+GL0WwXgEBXsfn0K46JiCg6NWB9nnyfYYNXN9mM
vuvhHTot675gkqI4LN5yQL/9ExFryaC9sY/vBkV2MygHwhGFZXMX1cszPwoPDtcd
HkD7CX0b17hzDFZ+knoIrCoSyyFkxTqOSVj/o1ibs39BRDsrTrtTVjD2XGBF0pLA
3wcucyoptsGV9QVRNObl1LCbDsYm8SOedlTr+SWHYa7uaTL9uiXmhArGOfUrj9Pv
TA2aZxtQqjl740PQr7Xass1jcCAnmMuINlF+iokZdgTNGVsQOD26/DSKKEqmneV6
HIgIANBZS4UgYebnXUCt0qz9sJLHPnmdKm4NrRO9p0pR8aQB/V5TTuazfs+U7ZQi
KLmkQ+05rzQkICqFMo0qIuHVNae8KFIMEJW6X+QpYvvCnyzN0ml4oVLORQIdf9eV
aVZNMnPAFg/MbTcVO9alEwdJ/G9UnEY9ZObm3rWROLKABmx9zwVqxF5XO3pBF83a
g95k9AZrNH3isEqt46aoOC9eRNLWRMik5yPUIoFQlvvUl/I5fJh8yl0D8lX9Y6xy
XGWHJs19C/INQcvXCyGfBEYnE+nv3ILne8H0W2beGgIwuNX2e+vre1YBzy++ZiA3
lea33yvuEkpNCC9NFus9u66FVd0FS6I0GJp5/pYXFiMCPPifyJ5zPtvduhCnR8ij
3ezyy6d5JxPu476MnSd2qPO6kU5PBk70mGtBsIwT5DgE2lB6UpieGYsWZ46TfdnI
4ZCoBifhcmfmFdEloCmn3M4hv4e0EOAFDvBd69V2M0jDiTDTbGJk6cBTir/Nb0yi
Oe+m5+t7h+Tt1vH5lN5cB1vV3/II0dekmLqYapPnrqPYGxBNvBBFaEG3uvfQSDYj
GYzetvV/rXr/RSfkW7P8LgakQb4B4nEx/qcZHA9CQLN1HPtGZBmGoCKSYBXx9N1t
kdnnwQ2YlfwJC6TMpLh6smwfenlysCZNro1eu4DpGACMhSqHg9NJrAjvqykNkSLR
ixAheitd1a/BN3EFblX0L9MLw/hlSscWfSgRwmNq9F4EK9lABMxUVnC7VCnRVuSA
f953fZLLSspLhExvXo19uqtubEjhD3gXOdHxGPPIpGdAPVG+DHUSJUZ24+m334Qy
71XkfQERI86l6E20fNTHZgWNge+pZqLt7BarUftHcUQnASEML+lqExxzBTegXf5w
kw3NnXRvij05qXvCMxPc7ytPX9zrZocIHU9+1n/+DCcw1I22SyUDbJu6TugeDGaX
84nL4r/qmsGrax5ntLFEQ8EhSuzRHvpwV+Ou+/wYg9Ns9dZVPodDKsEgz4IH0FvK
lzKE6PvS1IUJYcGpbCzlb0DWPu/kJqsVec45umAF8cfsMre602IMUVwgZ2MiJRNt
YBmkuEr2SZvdzWH/AJLvDKQ1Lctd9BkgSVFmT8xM8Enq7Enm6kbC2V4jyYcr5VWr
cD9Nh+MS5cX+5kTXI+EZCUhDMcXvgKhtSjLkd61FklEeOliXZAM+kgRM60511imQ
TGaCep6TpKvLpzelD/sgyFX/yXbUFf3v8vQ1B22pmtiM7y+bktMsbj/eLuAh7Bxr
cxJfISmKMlZ7H1AwgbYVW0CrW5MT47d5/yqoevUULkAP+PsukzgYlaJndPjQyPvH
VrKoo/rwtOegkhy3c2HLHnGoyROah3ye+ZAI0MZEy3UYHlcczSDJqtulMExe5WAn
0y5u+NqHcyy3kgxTakix0PCvkqpS27yhjAD+KgdnKSVuJ5bWdjUtkdPuxM10UJoq
Ze3Ft9L5z3RRS0tYhrAqaUyPnikuojZaFi1RK3xmcJLho/qVS/vIhkTq2PVX/b0R
vtwta/SFNfVDljdrEZkn1i7oJzN/3JSRwGNTQPbaU9Ys+0quJhNH3+NHOJt1cVnJ
Z/36VQJz8xVhkYStph3EJENpyfAetg5w3ENd6IWnlllyR34F1wm7R9Si8PRI1lBr
WNiSxDXCj1/+FZSjl3lUCzrANpimjlqTcBgxo3UOZyXu6hdp+N4At5E+qpbkChYu
ZDr9kcg5HrDbeus6gBFZsmUVZ2E+gfdfxfw6K5Ejf03QJ8ruvgUFyKjC8TwqGE7q
LT0aQmcfedTWsqq0MTr1PWBBuCrYqqkxTB3EjCVvTDEP6gTsP0oMkHoSSOOIPAco
dVr+4H1psJWSSa0ryGFhuKMU0W56MweBQmKc+GUiEa4YPIp9tpp6eWl37HGbyNu7
caLH/gKsU/ZFG3R+cGIkk9biOixoK3lhirtQ86g5wKXsJ+jnPByrB1IXtMqKsrq2
Wy1poZsrYcvMLf7LWPAjc91wgN87hjVZ9eAw21OHmPuQ14IUGfRswffi0Wzfbyym
04YksMH7P8rwyM+a/yUP6Vami9jgdJBcSZH5QMs+pAU1NqAnnNhz9+K6Ng2Sj6V4
Q9eopcaJP+Fm0hk2OVjIgMCQ9ocBpTS8zDtMTiln+D4JCvOHhxJU4ojuGSGkrZmP
wAWcnn/dQq44NVXSfP9Fx5PSSc5dnRCUIKS4HfUFmh6jKWbnzKj//iJX2HrfrQuW
kcRSOmzIq3o1pX/OsYcXbJOWryMRYFoExDf8yJX+rmo=
`pragma protect end_protected
