// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:18 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ch6gXPXlr8JyDQ3xQhVbwt2fpv/AsWDylvBPPnWSkwGzE9YXW/u6ELQ9OyZWEVJg
ZDgMQ51OeD13uwGufu9ppcvToWCOZ9OA2pdrx8CJ20QLDkUsvFBHlEq6kBRAX2RI
qTBcJQmt5ykvuDpZC9Mgk2JrAhpzGmcM1VyxMBkqV9U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71088)
0xv83FZCWAFRS9fPV8d2BZuzWePo1xPshmHCrUV44zPt23ANPFusc+HZA57qldQc
q6GgkaP+Zgwa6YYqVanZhm6t/AOfF1AeZAs+nbsmPWpaCGYxl9UFIenTlo1IQx78
zMYhgYG+qPC+3suUiszj11XI2dm734pokBGqPHQilewofGMnvdfF5jWphHUcBu6o
xkuxH4btuhZLXg4OhdLkQXENh9M3UokgcmHfpr9nsrZQn3kAEqr+XseELnlwvF+h
CIowVj8qDa6PWQVujm01zQbWttUTTXRIPg3HTy2KVkrmqrVbh/w/KLoz5N2YUbFP
qQNYAwQtrt9hoZOMkZViG0UqtEH+SqSq90wPVnKm64JYlPTz0Tn5qS7N0WjkLwWZ
aIeyuYzXH6rtTsONPeBYxRDpj7XB0QtPNNLyrhMr1RH/72PSGdyYQD8a1pTf0yVu
+mCKJ5Qv5tY5krVWO6Y81RxpF0T8HHaEXSlT/B0um5aSbjf6ggs1JhRaTp4kzXjT
vM8ctrNaxj2TZwLAyuCrNEyMsL+To5mb77rl4xxTndGbm3DRaH3dh16QJvhGxHZn
W8VFrJhKbZhfe8oZbfWDxkUJC2FtQMQka3OVCCSdRpCL05hUCOvMQzSPMzpgJr6w
pu7/fDr9E2MX2lKOjGGF5gRr5jSMm2kx6Ubsp6bRNjgqKKoMbvbvX0AJU3kd92WK
MzYWWOCFlOODGce13YjFkiWdKNSXu2/1BNZopoBNSdUkIWEBhhBnnNYsoMbctbvb
DTMIx24VbyOWB5wzgDhmVdwz/Eg3SIwzfKNQGCQGcd/BGeLMatG6ushPMXixzNnF
OfQfJT5ELwrqSpxYnDWVB1OnOi5a2IdqLMDi3OgD/X0e+OS6gC4bT/Y+ZbzHK4U3
Z98FlUavbYFbgM+4G9R05iiL75Tmis/QUrU6ITgBEYfUbDl9bZrDeNRqR8V6kqfM
0b1CfYK5/EcnyRdzLgSzP0KPcy8CmuiTh5t2ZWqbYNHuVnLcOt6ADJhV7xaRaRNv
lAOB2ZVTpD0RU+dOJ23bfZK9RMfpsbqUhqOPuOAq6LPkbGk4TyFmP0i+02qlvGyq
8IkFB7Rs3hLWE4Bbws+jqKjVdtxNude0sMLDkjT3QtDBSPRIYwGo4jTZTUsQ4qIq
IymeRXAmkRXzJEtWojAegDXR97/dwqXzZNzMEP5AQ129+io0pR+gxE+oOOVe/77O
WbKUpapDzOFaK/uCzwTADl9IHruELnIb/wJd5NrKr32g5tntFAdJL4xjqnqpav40
RHkRjWY7Y5dExVeMeZzm+2Cjuqs1HzHgDnZ+83BKdH5O8jMNoFUD5ZYbnohhe3Jt
XO1HqDDcvyGmyIb3YEYHZXsLikfD3pIVSII/5aGfn0IFuDOU6f48QHZ/CNj1rLIU
lSLAEV1cnPwtIDitPzgAtupwteyLAaOvvhB8595EmrngRMb5syTpmqKSrwgVgxWM
hBxB/t1l8aYUwhVINzeLWZ0BwC8rKwhq3/IavAgasu1RmFt705R7QolZdxlGN/91
SCdgNHT07XPTfHB2dipRfEPxCqTnygDoVuCxzwAERWS0pPVk2LcpzKLiNwcZAxd9
LfJJJ/5AB5ou+5lMKKTc7TTOflddH6R/pNghIzbI5pK9X4ARIylO1G2BitKYJXxO
2ROHS3t8CYqdOEyWVUixiYx/o+9oQWgRsTsGKFHP1BXNjziKcR/UzAbPRHZmzWYZ
5gjnN+gXqXQyWIkuBE0KWE4P1xiqZmCBm4VXf8xXQ+gaWpNJhHFndfN73Cc46Zpw
H7LqqOF+ucyDuor4H87SkPlLU9ubdb1OujZ2E3vn5q9LTZdiItZTLfo3NCr3SqOx
eEnoRZerXjZOlkgYmW5BtEQUh8p+TCJOBNDK1NIX3u/stIyXOa2aFhUqqWDsaXZA
gWcv4velvdl//CbRq/pZxt3hDl9SMCD9+daycphFv3e4HB9eObMXZT8qMbWGOTTI
KKdXp/PaxvGWDUFPPV9gyBdyxhXPU5SI8fCE2pW2UC28s+aCG1+9rnBKB76iunNw
IfIAbgBODK0hzkvvCPsAXLd2x80+ZRlFGTR7Fx3dimDLA5ZLKdUciIEDl5HmjGgp
ZDazr6UCnzH/uhgsgvGseRn1Lsorn2U6Mw8/1H1g3/F1bg8zQoTwFQGe5ksETGYp
gR3+kSiGSWTBw/IZ7Ncnhs4CWONqX4nLqwjk4RhE6B/96CmrcbOyvwwSDqv6OqNw
3VBVTDk1HPN3V6qLDbG8vBgk1p0818BlduMRYqQ6mqlD/ry5E1RiC3GP8IJ48BGX
t928lAv0WKkeYSRvmlJJkmKV42PfHpvJc9sIq8qcjdFgZd39BalDBV+tMDk48+HS
J0QJ75JlBu76bf7eekqbZXUuf8w55sCqFLpj2kx9UB9ExRo6hVFjL2DAeLtY6BwT
Zqmf3FbQW4oAtdCPfI3BHUoYWa6I7n9oH1FY6ptJHtC184WCd4W2V29D6kHB/0sw
h4PB1Ko9tjxx0IJuxfzwf28fLVqwdIR7ied3wBXve+205x511D0BPbxICdPvdR5b
C84nQL5C6sVK2b0WTHR5x2OSM+iHMnE0KlMvtbzUjZGVftuJeZvjBuU9ExECYZVw
Rni1m6bW8PQh1SmCt2DOtvVcuCm2n0WFhzGEJXLhF4Tx2eghWKWJ+oGZMeVwCI1+
FEqjHdmWOCWzmMu1js4LVcmP8oxvQk+XYSirUSjp5wdk6yt/4K2idvq4yNTxPIAh
B/3YFGBZzPkvFJsOAmM/Kw41kPrWCmvVS6yiHNktkkKR0QH21X7s+faBiuhQKyzy
8TBDYDpZGsJ5nUhbMY1oN0TQYtJmsbl8iaUZOA/S2mv1wqozmnhr9RJx0m8uBMGD
VAcbHBZ8sLrRFDF4SKzftEi7OSPrWlHIH4e1bff4QamdfTL4ZvR9LuTu2mMVW9Fz
dXny9UCj0hSDew7xdjqVcj9QG9nBfUqooQzfZ9t3M2YL/ViHofd3Ay9DZ/8vBgtN
bbEhZGVNVjggCZFkCAsZINnkRnNy5qUHSkt5J5YnW9qCMRJYNsjjWgHsJ05FVX51
cfW2FB4dz6g9g8KnUn7xut+JvqQBOsgjGCx3M74VXszfrwJGApXHhyYHpDsD29Tw
b+6AROE8BpbkfGH4lcr0sVbNBG/XQEZmDIC0WgApjhd+l63K9VGC4rXWR+7U/69a
9dpjXv7M7xE20V/pz4/XHQm3jTrK0nKR9YT/XLIqrF1Rb2ehB4K7i4SXycb1wHua
/fW3GJ0fGZotdTrfdPJFgoxqLrRBiuB4UgmfsLKDazH1c4dgM+TB9MS+ukzRDAbL
TIUCO9FRf26NdTs46la1S4zUnyXYSwQL9irbRfin2hQFlENjLqRpxG6riBvAwue7
2O5Jdhci7rhha4S7zklilve12G0sNPcf69PtORH8Oyg6bs9ssDINx5MSyv7X/l4H
SZAZ1FJ0B9+8hfxsVKvFV405Tbnf05wZsFF/sbSCxZABrJ3KZPcdgMyB2N4iWn38
jG7o7PkAp4WKTI+MNGsvMpPhc3QzD0yfkuedNYUBLFc7E5YudvqSWIpG9/Iv2JF2
+NOxW4d5CTPzfoDIZfavKFUC5TOsgmnY4W9Gw8I619ZACamNu9plo8mWiCawR2h7
ftPEpzaRbIIVDerZ8bgbjVnCFIoCsQhyF72EHhbMoKm/i2ErcVyI6+8jx5xvUmmY
/W2+SjJoUtOSUWfeLa5w9x7Z3LfpAGjQsvyNgj/KwbIU954lyBRbaMNUKeH58gUy
87YxmtjUIIzB/mLeQls/Vsc8S9/c4kDzxQ4ottrFtu7Y0627GIMdkiij2dsDlswr
F5yUePH9sQNxFof6xJ9+tR7os8g1/oOsYbkU6s62+J3ysmexaMsXrUiPqgpuchIq
Y/kUfpc2IK1ZcBn6jizB5DGaH2VD98GcPeb54U8A4Kt0izktyjNdV6mU9llcwCe9
+KSlU3tFT47sXmhXiopy5k9aODc1rt6lv8I4gMSMPtTIO/RN55h27dB1gpX1HLUN
U0BWEtItlkmFsi8vUfIXwLs0/FKJU96AY2ut9lTx0Mjx41ONeOYhccqa9nwELnVy
ZrR7nqunHhqXy/PT0WFpvqT2z5e8fxG60lJhZBmmxCUc7DtKYz5egh0HLlPG39Jr
dRZC8ewF74BX79xLoVGBS2ayF1eM980a5l2UwPjXYMgQPYedqdOXekQMDlpgExob
jNmCHB/MD68eOyXsPeoTMLvVPRvi+qS7d8T8xZyqDO/3xi8oeGAsKyBQaJSHt+M0
v8u1DeOafcL1c/mR4JGnPjgoxf6oFdNKBEReXnQ9rJSOn/CmjwIEYHfmWleHpxep
bPmr+Vb2ljYSm1dTI9G4YBO13BTHbb9novDiU189hnjraoTFFZZCHEPZ/yzXwzS7
B8hOIldEAoVPPJYGV44e+gvhirfF5Za6PsmsAIPI77WsjzKywofOrCBVZpMzUR35
isCNjQYYXfqDD8tisjOAZB8kOgUafDzS5j3TwFXebosS7KLSc/ZVFI8lBxoOipww
Kav8BgKL5UV0mAVb68oOfzoSJRJofKTjd7TubMok8BGyN9KSztpdvgGXTtd3ie3b
S4nZGCy0+19vCvScQqPkNzWSg+R01gMTokQakgEZ83vvPQAM6AV4S8pSzrfLr7/Q
R8Y3SbTDGVoteT0Ou2kZ6Ut7xrEmS+96JGySEmBrB5G0FjrPrRAesPtuCiHHIcRy
Zyhi/g8aamqyW36e4DJIXPQUH01F9BTga7KCoOp6mv0APIzkDwsp8IsaeDZbNEP6
DddMQcQSKC9tQf8KS0A44R7gPs5vM1z6G3q2tBgasjHGlpll6ig8GjyVppxHpewx
yitVyXEa6xULx//VoslnpacntmRo61g8BVU2e39Y0gZkzgDekaiJGZPoF5Z90WR2
T8vlt7mJ7FV0yYtzoDrXV6yBi9HXgj4GpKuOazL0xX1AQC09LEzcPLYIdjXkJa6R
yTofFVLrpt+NdMgYezHwTXa9M3Tfo1PsCYhuls84rxKy0iuVczjk5datiVPuYzV8
PZjYdUN8Owo3wbVnwXKmiDMysMiJdgxWPUWSFqnpbashjvUgm0zT5h0jMhBiYri/
DSsxM++4Et8ruVTxaTn4tT6qtYqzDqrAyuHrTY2oirhnm30Mrx0ySp5S5yiCq4W4
Yy3J41f4zm5lk2siX3BvuEzNFESDw76IalpvpKHjEBPd4q6dNykqbHmBN7KYNi1A
LnA9HAXgb57w0ko474inGvc69t2SGfOK2LBUFL0vc/kQpeGw7GqGfZhOoSoifBDF
ph/AelILLKgdKJ4kDCUlShUh7iQO1MCvqVSOllTRMeqbm8bssJodwQQVeXvDXc1a
BvrfQpMgOWJCVkVytXysfo+588AshONfNWsCCqf8tnMIXH12b8M2Tv63V+K/b1yI
yBnUa+YUm4gIChoPmsA0D/uD4qM2nw9BHKkBYf7My1SAzZef5kCxZnLpnI0XqNaV
DT9zcmLVGZbJHCPXFwRm573KjrD1P2RwQipq8qN/ozTwcqHjd0WZPE4GaTA7stH/
LDyQx/8UIOgJwVQ1kI/22V2Ky/n7flOzSwEucUlHWL1AsG5zuQlRepzaNxUiAzHu
vZ6I/0RPChjiZqOE3E0K0DPSzW7qzEgUAemfmQQt/Ff0BItKWDfqQ1ZglcG9T2sc
Lq4Sv+e8GKV38g+4qRt+DjeM6jFGPIwIjYQVixAcK3emAYv8vhq5hYpC+fCLYDSr
pL5LF42IVX5Z0MOzdbviJSS9mpoN1XTgXY7jObz8dzkh/5ghgh31iKpyDEKumZ3H
iNm55SVxhgQ/EuAqSuujBLbwCL3V50x3d8vPifOlsaKdhu5c/UnFAXu/MMvUuOaz
PmFupHreLn5iFFWskLg05YdNGySPI/ECfQ/C346VNqaPcO9H5azi9ndyUM7coX56
GA/5D4OL6M7hRhYAv7DxmEydctJXOjqLEntfhhEW9hqkWeMSuldngBWEb/DbgIHL
Dqff5JDi5ErQc0O9tRGfu3WZHNPbDaXoXS8MR+8CNehBkpVR28P3FLQdvzrTKqOV
2Y5Owk4JFEpF/ZrzoG1KuAFLI8YfK/IcnSgZ/kErj9hOrBVg5jEORHMnDKxm+yDi
9B3yL87f32it6SAQSLucGt+4uFdmI8Bz7s17yWa7YM2C6AnO8JWGT5t6wMMAwzH3
jXvlTijZgMURVcuZBb9PwjRCRiU916YagCsDoeHrrpwCK2pFS6Gq+fzbc/CsQNCk
GMZe4O2BAwQloDjmy9hnYaFdBXWjcePm0vBR8FWxeszxPqziQp4PcJrsnTF1XJG5
1pYF53HxLpQYjxItUP1I6Qb2klxTUchd6/X0LZ0VvMH3NWjOpbN4o/lniwzFD3cP
aF0/5Vc2ZiaM3ZEouwcVAeztUnN70FqewuCn9BFRnJqxfCl0ZdEHKt+74rBGaImQ
PeEPLwySGluR6bHRvCCntI435IsrOCl3dNjFYkZCuEScndlxVf5bJZZwlka/2Q/F
U/iKXGSKAFZ/7DUHlgmo5KNjE27GGiakCnfalEmEkytPxmvRDOKDitkgKEIiGKYz
yI1ZOhxSaqWBYu7xKUKswjjjjuINzLibnhiHpYDnlZwjGjX0op0RyXNjudDCNkGT
3HEci6Oux//L98AsmgYQb9dL5Rfy7h+g7eQomufiBgzxGHz2EgE17a5UIz1+ND6Z
HqyfS04aIVLXAhzhP+A2IMSs4dwC/0FJLrPy5kb/yq0vYfyRFuw+sxC8mPJVK697
//fckYQdZlijFNJsrePWR0L0FozXNJiToBJ2/EpTr2+7ZRx4OCCUSXf2AafV7rIq
qijyCNpSxz/nbe1x1V9K+rJo64mOIIrfxcoQYc6uMN4Dq8jZIdpVOcikXICOfH3F
I5n6m8Y9BnFw5qEEZCSs2IW62NlJYRB6NxaFmETuIKrH/QTRVqWXSotE6dxD/fH+
xkxgJRiyMc0cjV0MnDRxuDBd+Jtpk/I4T5Jqqsq8mnXrk/6l13l8BfVDUQBW82SJ
dYDK939dxLsFV441t/82AJBqpv6DY5YhzIg9ecH+gA/Ei8YD6jT2LgZi9jmXQN3a
LzV18vNU88nY8bB5yGwWJuLyffRS+JMXnB55UnEYZn/ozWKWoEfFTXq/S9sMYKVK
ut+69w0t3ujTh00OLrWRVZXpm1HA3Cd8Bjl27/vfMSSwyi48CwAsW72l2hHyz3Ns
aHtPDsS88NIicuiEhEsjEmRZZdFawugniTEBH/+Fq4I6EQql1E5pSRH63k+x6nZO
5p3jIO1byO7CFS/DbbyD7EQLHVDCVgkVDD1885SW7+CRiXSQufAp9MZq9ixedVdA
L8hITbMQoILMrhPDKvD+rf8Xx/23gcE22hK3AaAkw/2d9lRKAtzSxrvjfGX8aXP4
WwFCOGtpH/+5aSIWQ8KT8GHtSR6tEnkH7RsHSD3XzCgs6LvQe3yQ6+ZEZPiWsClJ
aufT4iphr121tTIBmckP/96ioZIDLW4KcwP3yYUTvOee6WbluqYC4AgARHDp0p65
VF+OYao38FijHcWmao5XwcG7ynyJ87y3qoNJlkw+tvr360tD0TqqVflisB7sb96i
oXVYwpOIkPnzFIoTMGzthy2/Y6HmMFkDoBmOtAoPWd1ivjVKHYI0VQHrAn6M56e0
TQOx7HjiXCY+SkSksWIljGY71enswDeRs0zTjdTT1yntKu3zD5Q90agW0tj+XLBe
VgBTCiTEe9BlPxAKHwCzATmUbABkqZj/0ihNOB98pV6vGGKukbK97PJSGLNRLI7G
yu1xe8O4dSsBZC4V+zaXcvguaVnbIC7em+KfQtWw95ErfP6FfwDmpR1Ds+usftGr
t9nzgXKe41nlMxryxG82goVLRcD6foQkN1g+IAohtLgGfYKQVuDKUppYHvSymIb7
DiSySby3TTHCcrThp/zKvyTLvltrHKrmv2laWSAuMy8qwanJPBso9JrPL6tND5ij
kBNhwOI5X3IeZ4YkDHOGJ735Gqw8aVC4fQMU4V9X7CSS1eZFvsbZXdFceq6vZ9T3
52ElCM6XX8/0uT5ZwtlE0xK4fkvewJ7Tw0fcRM4ZGMx5IJR0e2WsijgHrLPX6H1l
9E/2JeY1lOFnPU5yurd7F8ium7Cxbl8IabVTUYeopFwPmxrEzVEdUi49j/oYz+xP
1MiOxINU442f9Fm79fgKHCLxQoOPpC8DjW1WaM0w962ZF2TuUaZyz3Q++PjIGATn
l7mpj7QYO+l50PittQVa3XcZHjY5EgBd7sVZ6fhCiDdxPWI/6lTu2RuISMXWl8Wm
/xjLXpjq3epVnECVCNCPWDiH4Oq5+2wxLvbH1LFciPdf6RQZG33u9mJk/bV+fDfB
S6p2X1COg3MRrAC0D2thOCsf1c8XVpMgbQ8YP5ZzCXRXUcC3SKku/Z9xdNFQabUH
aIYtEeWKCIQaeLpWQ1v1hhufA6+C8PlGYWzO6Pd+pXXhQWCuxNoCqHDuEcCVeF5C
LsuIt658c6IELEluwB48sruzr8uf78MSCzVF+p1DYpZ1pMtYQL2vcNYqAYbYWw3z
Ga+YtPypbyQCohAQS08Q4blAT1jzSJCgZnbwUJuT3sR4V00F1J8ikN8peHcwiOs4
moc6q2usoR6l8PlJpk5rJiYApC/fK0L00PPXd2189CrSJS0u/yYMD4u0Bt1bl4oo
PZH8RaG7/kQw0B6F5xyDN2X+CR5WI5YNXv1YNPSxi553huLrrt/IUbNmjOM+WU96
k/lCavdxkD0GHj7VF8huP1tnGn2EhpRC0Ueu6UDBp0g6M8lsD7fyL7zGgaAJl7Kf
ApR41oygbhK/GcWqcDXe/G3PZAkWc6exLVFGe7tyMTVuM9SW4y2zt2s+pWtfMaIS
/uJWWG+DKUje+pwuBPkUqtEnM+925xUrbwzB5PWAP/lGfSivB1Bca+qRZxRGJZnb
waOtmKNJiAUe6vys5fir1H0qqgMvJCLgz/3mOF2xIxqi22JTO0Iau5wxzJoiVvdA
aJekd4GJjX2GRHjU9SNdfIvlPAbhvhqIbXZ+mYW51MpSG1ERUFEH/+XHy3+GdbUI
FpOCv1QIzs5NtvrG0mmbFP4RbSnjmtAG5IOxtSs+HphijDzASJht74AsoyrsOIIB
rlIflMNeIW88jZHZ8gitDa3d/NXpI+WYglp78HlQo9YbzjrivWn5y4JH85Rh3DeD
mzITdIIaYzPLSO6XRZHBDqsjDhoXofzGPdW3WzsZkr/9mFxSbxk09NFbvGuJ+hqb
q93T/+yYfK6xUcqnQdLerOfULrLCrPEwLQr+2iIwd1lKJ5d6VwxCv4GBNqLHRRSo
m+KaR0Lr8g70ch6RnJDYsIeCgfOxeCSQ/o/c18cUziTDiX7QiTHLiu0hGSn7bfbK
KdjZ/N0Z4BGwoB/Ud49TF8q0Dk/THciFgwiCo7CHGdRrgRdOnsFC4KoHjDzRQJhe
c473AOzN83Hc2Z3oMTaKWp9v+pmK6Ks5wOuRz2RvQdxiLdkgBJ6f/GbtyoLnKd7l
C/5aBJYzMN8FYnheg1wHLINSnxqdFNjgjMwWZd8b1JS+heQfhMQzgMAP4Tw8jmeJ
qqm8Q/q01uAPkGL+2aJwNE6/nFVBdlGic7pax2dZ8Tc0vnKOshLCgCLR58h0k24R
ZgfDZxcwSY4zUiUY3Bg9hzfrg+KIKESoDVAiDeQbFsfHlwcqcBwsIvyLpacXWd+m
cyzSpyFdDvvc90L2/AA5li2YAxcj1pv+HrvveqTO1Z1JD7GH+Ur5KKzan3nRnQdL
pD3A+6S5qp7KMPtd4ksQ4lq1Ir+DruvI0CsDTfjhayEZaKdU+mGcaImBF/BDP2wA
avwi6zcyKlk7XonO0E93mEO1GNHMKL8Bhu4OYeALfxUSyy4HKehOE81YwHzea0sp
hnFR7R/fzpjPv32DfqJcpCf8DsNBTrvmQxBgyuiESL4QghFDeNbfo/TY15mPFwVr
52QjPvEJ1o8IGj9RQBtDhNn9JZhi3Vbr4wa8Ts5PE4lMapaZEgW9c58/P1voKkpr
JoJRpya2oZauSwMzkw18Io6kyGvSTVqc8gS+Viu7mHQz3Er+KisDsEj9t8JV0MJp
UsUFG2mXn6rLcnwpsdTWt5ahQge4QYM7ADCW8X+ccd5Jm0rjWOqAk+9DGOlnbZ+R
TzjnAnqLKBNXc6WWJ5SOzQ0QkjxEXwjno/FWpAx6vH2WgrrMzw89oNkIvHHtcgsa
Dti1P13uadqQfKKpQGy/SSMn65gUGg7PCPQJEzAeSKgvuTyvIeO95oqODxQiuHx8
fvaY29bHuWbUH2l74v3fedC3NSGNZbdxlqUao8eqhAy7WYaCGbNzKSScF6VHQo4k
Xm0kdp2ug7P/rUUjkljPGKvTJUQE4lFLtl7JAxQWSd/So82cAHUx4qihq1/x3Ekq
WuaJmPSI+JwALmmknD4Hk0ux85Gs1gOGwrrWzAICLhIoiGlUanRuqJg2BdUALWi0
fqb4UC4EE+6nEcV4nFcmvTlSU6gFLLVoU1KyFaKW0wPrF5stQjZ5W7UxWon0cACX
o2iJmQkawKn/TS1aAO1a+lW4ZkqoeAGZK6DtC/fr762//8k1jS8r2gaRCSIcQ+wU
4puyUMkSdiEtE+DLhO4jKIkmKWKeiEfFZjHaYkRTPa0Pvfv2voPWDvVVZ1xKtuc9
V02PxFfrkbUw08UivexrbmKoo0/JOB5e1fNveD7kpa0DDszZj/MTrQLh69LAvwty
cAkEwFpAemjcY4r/rE8dsrQA61ckZqfUYtkraoi1x3FwvJoRDoqADbtj9P2AmOI6
jA6/8gBJ30pJdZN/c2l5vdayTkp3gDaCdRT/CDNd4XMY+eOgqpJDt34USyKlb16Z
+PXTvYvHzjCOxo3/v9qu2pcPpgJymr7CHSd+J6SaS7KA49HNT9+kicOeSMymKO/k
nqloguA4SLL+u5xBgLLB6Szfrt9oehQTkZ5YvwfxuwTHx7T57t/xwVOqZ0rGwLTs
mIURYd6L7iHGW4qIE3TyKJUJ4UCX9nV6X1IFoJT+lLyDsFwPc6/H1D1MHW0a7052
0t8d/+/CE5nvOi/1PQhdAbOgWN3weeDHn0UxaftEHgjQuDhsM9txZXtvs3l0dvlG
gf0K/HYtEMRgj3fAszfWmSAzP+svNq6pvwQQ0XEb67xpnDhksJID7CL9bnguumJ7
vfPlyYE+uz1Xw8HfTjKqJSy0mnsAi/ymYaDyGC+rBDTKUsRevU+xt9cvss4C3HfD
/JWpqCxpJtDJwKUIJV0em23evGEebc6uFD7QFq8iwqBwhmbiDtYPSB5jEsTbQPQD
AiM/JCqF+Ahb/6k0+sk1fN7M6eNUMrycflYlDhS9le7D7W8BSgEdFMugohNaHPUY
8ZVbKr/Q8IsDd/PFrgyYL15a6i+oi1a+6+0hWOlnQnO1cQXR6lOVO24vOxQiUvgw
0TJiunKlhJBKLwlVaiwgq3m9op1qusgeqPJeqmh6tsRcQcu8VOm4EyIajSqLF2jP
jMuJWXCa4DVtmksYoALUdLb8kTN+dJCAnWklLD0+UaNjtfEvrqrVfkM9h12HTVXr
5HBdNxguPp9+t0LQIpzb4FvF2RNDwWDn186fK1fFdYjYZECiq0nITktepSC/vJFF
V71AqFOlWWQv1dKuirao4JiKMSyDLEaIlAPxv09piu1xVhlUaej/0N5gbSnphJIz
FIdL+/X+wM76Lf4C2K3P+NFwCV5WtiuSOg+wn1sHHBOve3ZG4phDsvv4vjIrdbzb
GvanPyUvJiUzRvmF0JxuqCafUOhimn7YdXXne6nukL3G59JRJXI447KregJKIqzu
qmDfvG7RDkjIZw6Fxy8PWrfYDAK8gSyfIufoFbqvXRn+ycYufgL56mHft+693gMa
IwkE1o01dxmj+x3ZsDA4jznvQXQS6kmj6p4bC7YcfbWHZMhq3pSqXw3OsEHTQ2Kl
8CrnOwM0S+VHceyhtjLZu4TcmYWfChrAaakQOo/aj/yL7zAe7r7uevRbenJ0XImy
/nYXkl2vADb+GklfAsnQQRjW1VKw8ZNAKCAkOr0BkeZxqgQ9yc5eKqdsTSc1RlDV
YUgZKVHH3Yr4oAbpVPxLx3XKJp5jcayCkY0VB9wAbfN7QaSPJlpLrtQMtyp/yNJL
gWNSTFNWOpoPUQh3ftjzDFDx15hgIn8eL4LtmKL1NfUzO7lqzxD6FtakDIj1Or+P
4L5qs3jQomUfN7PTcDvzFaDPBkZ6RkKeVgeMGFBLE4OAVPyg2uOn1Yp7axfzqZoM
jyKKVNgRSRrozWN+SrO2LrnrkvNLcfvvtiBynqjg2c5v3zPs/5aqxxcge8FUMayE
q9ZHK4w7Tri3W3PlMo44GKeHbkFsHJOGqR7fGZCTifRimksqAcRBQsLA7/YTDcdA
97qQssV235mp/CWG1TaLrH5FMPJxWbT2WEbXSAB2QZGL92xTQwHcI3IJhgAst9x7
4cNcNm5SDVhmM3Cq12dIis3YeGFSyIgpN3rXjO7ZAud86QMBdmjhDfHIVmvSId4r
9QIQZ3EtoImvwkJdfDrNafyk9oZSMEQYPIfgfOaDRMc0Tb8nWx1+N1FDbfAOqJbW
okRhiOIlebXqRIfNI1k77kCk9LxVQmXo/zdQZ2pe7fKDK9pWlLJQUz1T1ROi9JZb
HZ3K10EjkkbSTwotN6TC0kOD9eJIzYwamvSc08HfBIDOy/i9gxNcaq3GoLRhox1e
MuGW45uN09c5BPiucnIeiLtxtnGvucxJir1FcUK8Zn0Hl9FyJ4QBOGRrcz+4dExf
cv2NRc0kCxXig8WgGkcmEjHLeE3M+ELrxwJ7Wh+0RgAQS2W7mJiaaB9d/NXoUsLE
u2MJYG/xLMd5jxB7MA9uUubolZyTpD3R3IjoWtYM88qbbtQcsWJZWmlTmu6HzwWb
fvSTdXlB0EEaHm4iHYdyZ4C6DX+mKlbNhH/d01wZylk1OxVXL97xTMtoUkKDtvaf
GuASlpEa3jdr68Hpz36i7uzTMqz6p71/ux0gtQYokdMTd8Fam55uDrVqm4VZluXj
d1TLnKQJN6MlWwL89Q5N3UV1ouFB09a33v4SE0EZ8DfaQQDdZH3xh3ztxLtSxNlT
bIXU0yVooBu6OalFsm3vzo1iJkscJZavD/Ri7ddhAZMnnYbu3xWlDI/0wSYXINDv
FoDJfc2Qu5H5C7XjneH7QJpA/L9Od70kIe9JI1+W2NToS195eTdBYG4MSuvz6SMH
kWKgBNA5IS4pgH8Wjvaaqht9CUTIR4VBoUNUNRqHm9SOuuU5q4G3g95LpTPBC12/
JJFpVpd1AzpbWsgwIldC7D83xXx53l/k2j8+RGEeXwS+QkUp5GeDyRzuKRYJzFV4
Wx9dgQl3yhjROjpGV/2epT/qrbiaWioUmBndG/JpUbi8slgRBLegGj+/EBMBRdCN
QaABYazQfjlYGPo8/n/+qB9eJZbjpLwgeLkSmHPhPKgaKwP5/hdmlPrwal0UtilD
ZFddd6IFHWQnwnfii92Gz8k+fFV5OUEV5Y4yuo8WeDqBjPaCl4WLEQsmm9qnc6de
Y+E9CgvXWdzSfYBXcWSX9zmkdYHIcqK07z7u7Bint6V2DsFHbuazICzY+9IXSoUI
0X+Ra6EyM4iR+kixzIke8V4UphYfsoAwNyY5AHsdfcTepZ729Ws9ZWIKDpqtBmpD
4Yp3fyBgJuW6HfdxMyULMpt1PLMd1wB5CX6ns6tNxo4GqsE8i3G+9Vq0eAJTLWdx
BOLy/kYEabHTb9uaG1/RneFvsFOX+IdJQnqpo+Tx312yjotWkPzcE052oKTerFqn
6WoIUbfCLBt+RExYqqndEQqAClp6Hfo8rRzBiDa61nMRhMYBP98u3Q7T27+yeipC
e8jH8pmInDpOKtmdzf1dP7kSOsZARdEYqQK1mEJKWloRr8m/P8tm5NbQgP8sCrj3
uqRTTr5zQdlCL60qARMa3krDHY2D4zbpFPZNeWVXWqEl4krdQuTww8IcKJM/ilZU
xmw39obcJX8n7zOXkQFCNLD+5U0PQkFq4OrYcfbQZOGW/B+ZmW7vNe3IxZyA9og9
biK0qdeFcfPv3G/1nW6K/pHaEWCAlt/IBstb0+b5BfTZleYABUUmO/biwW7JVxKE
Gm8h2erOTSa5+cJgmFGBpEREVPb0p7fzNcQ0DvGQ77AZokhgTBUC7JoQzrs3gwT3
KUPn6g1qQpagLjUIKswiwGNjIg0LTkZhbBoeMeiY77TmQboaYjbxpOGkbwm57mZh
QT8pCvupB5dnrpDFqIqNX4lweGmILscN1bQWxTkHpKzqhsVPqqV/IAcufaEMhPRU
LVqLCApYPcE8w/gt0Nfj91x+Pv1K8R+H1zNJxxYoxoucvP4YHWUkTdDzf+mNlE8x
aZ5apsSLT/0tMQ04NTHQPWs9BRWDrATtaf2dXYdIarBaasngCbXM2nzBAptvhd/c
9BBIMAqUOwFqLC1Nso7jYcHHsxS2ZzEx6c6k1R4z50bqY4NC+6BFOYm/6A1qQcNw
2n56Ya8voF2CfmQxjXXqMu5JePhApofxmI0AipaQYlvdafoMFMas+Wv9MNHr9ceG
Jw6GI/igrZcfAbqCmzdCZL21SCuhez1m1NiyimFayLxu1N5tdG7TBioV9ByH1eAt
VJidQvhO4Io5B2i4/IMo/tbwZ6l/g6+11DT9T2aVDe/GCqYLBUolukINtNKHHHn4
ouJtLa2E7BlpiOSvufRmlBjuVXNJ3r9X6/nQp0CBC5V8Tj5XHs2Ixfn0Tuj9IFdl
yUFVZeq6pNgyWmK/WBj0I+jIuuhfr9CjolBngtXsWNxNXrnSkCQmGLvEkow8VflP
raQ7fqRXb8bE+zllRXYyBfuT+vkGJf3PrtFPGqeDC5wMNNUtlRFQxGKbTLMw4pMH
4IUW8rKK8OfLQaXAsR3P35/hgQjq6/jvJbxf8aOE3lir/eWURz5/ubX4lyKD5mky
bmDKIDpid+X1s3+GBudQO0r+bx6hi3tzmQIy8IqkyxDBFtdPSXi+VDBshbAoiXyp
4a11tWeCVwYbGfQOY7VkX/Vqe1cBireJk/3aVTFoY7kpWCq8kQCTHij+IGVeLkDb
2VFfOnpdwg6UzpakYgdic6KFXcwV6vyd9x8eWF9mNc8e2F2ywqFMT1VdWSeU4sxc
9GdL04qX0pT9d3MCG4KYh6J6TqMi2bN7IaQBHEiRDfNqQeYiyCeiExZQWqoT++Kr
fT8CyNjnlmRs3BI5CLX2iRfRvPTqPktl0/eHQwPO/gF8EN4JsaQRaqKibVTWiCRb
xBkZNY5RkpXqzmOnOrw1CKP5HyCDKrcwpFG5pdNgALFLNIuZLcRKaGn48ZZHWkFh
i2Ker62jGchqblRwfJf1ARNnAyFfq9FLicBnCXWr21+uu0qudH/xD1H0XcE5+Ph1
ANfIUN1hkodR/q4O5sC2J197kyN3TIKGqqCJ6CxigSJZx6S/AlIG5k7lFZLmaFtI
vEy2AOlTcn6PIsOU20NT4qOJHGhY3ciYwOUokA5djATJfJ2DeeRLQiaKdWyW9b5S
/8847O+fslDjYxFx8MPg0ToGkhx/nRAa9FfZr//ZicGRAKKFPydEm3/6lwVLmpZH
X4tDaM5K6hDDPccg4nUb5Oqz5/HxoO/os4U7RcVHczkODltMr3AUnfBjZ2YIunqd
cqGP/z0iwMkcguKUuzHC/EM+9tZ1LncaLyX1cCQHcL6lZss0sreUpgFzrpp9d6N2
KUXSQiovG0sUwjSNhgXmbA8yJQQCQbVinHVcpUS1/F37cwFnvdMscGOah9hI9vFZ
pJjyVDymBDRSzOQXbiDD5uPeVY2axM6J85nclggdiO101/sy9JlvFPayEju9IZP+
QUIRMnvJR/xNt+nCA9s4WcXP/kbjGliXr8M0cqGT6oyO8uw5A2D+b1a2PGJJNQdf
+LCWHqIFVgfLqRqI0q4UsRb5KDQnhPcKR3qqCmbNzdKvdzTCfN7CD87VqQOsP3+Y
W7/vujdUMCBnrZztjLfDnZvaaeojmXzx5xjScnEjFUW9HV2aLnIRsGY0PovUdv6z
CLfR3od3X2GuKxBZrzndfwbU3Bd499N4mySmZiNR/CMYdv8iK/kAUQDk+3Jg+02S
uY+YkIEO2Zz81ViLu+Q9kQQh8J+vC44JTGxx5cp6fl1xn2GKRruVGtEGEar7PleV
LYEXgQaCU5TF9rcCbmDW+i4Ilzlv1E1ZI5TsVZ8byV44yBCZbWztmt9iye4QeiAu
s6PJDlXf9nI++9fuyOZtresibowx6+AVtvFPdzO2aGvx9hTRUIWziEm5Qln7OnCy
wLpM0yxsIl692TuXuJTHZWOCZKDiR2Dw0lFcni7MRi59UCGJsFq8LcpKd/Sei0Fn
vfpRBxJe7njz8N4AhBuZX1uT26U6VdU1bt5c5HmXb6OOzRAw1mrO9XhahcYmjXYe
II55noxq/To1UIosu3cH9Bjqs/c5hDjJPXXOx6zwniwt0nAaHj+60seqDBaiQe3A
j3nx/YI1qmKmnjGHCVWZrtKMD4xX+Ez4vrNvbe8H9d5cN8rpEwevhQGc6Uwn7V2j
97ZhpxOF+GNZ/uEznEpPSmRvz1TQ/5uFf/FPb+7xCiNHefw1SXZB23rA4GvTyQag
KPHQDxUko8WY3OhD9TZDGb5flV1+EOM5hgeLVe0FuZGOrL2C1YaNCC6FIXZ7hWWH
1BD/2X8eh6e5RrBwlSSCS7beYLc/5O/7WKX0hoZOAbrBwDp7WQ7eX8iepR5kxl3f
aIdUb1a60A0mu4jrvctMsksxEio48iBzeFPVUdi6Wf9VDnU8iweEkZ+nGCLKV0az
AZnfnya5oYgGtTk7Olsfvt5igbCTcQAXQvAHFvTk1pmPuGrg4Cf6RuVULI1ZBtku
O2F2Ykhtzx+hhYQthDYkk/5RrzSGDrSNV/ypfulxdr9kPkWmdJXkH1D5E1iIGAuC
dXXe+xBRjGNYHxq4Q1bXePLqi3JhLivtkijymMcXAmltOxmbz3Bdta+IIudUWMgi
qcw+aZIPav04hBKX0bkoz/rJ8j3JmR2IEwXhAw6q9UCeJLzzM1jkYgX9+r1gTu1y
cVWnMhWFnSMz77rog0nViCeTr1meu4pVG4VsS5gcE6cZK1H6Ns7kOSmZ/WvWX9f/
nqBjCrF0tmBX0HiKfOA7WMc0Y/JdviK2Br8FeYDojHQEb4baWmUAllCHn96S30KD
EqIkAvYpFDocSW12NQ44XgMV6dSUxxDr1Y27i7SRfxOft7AIPtj4fMWseN7fn7oa
LaiwNZJiRNowfa+yyn7B1l+La945QZrwUntX1Cd62CjEAUXm025O/2bgtEpWPOMb
cF44JB6D9SsJAyjF0oMqnfnce/7Xd1T8XQ/O6arT6Ac+ixmuSX8zhPl4Xp4WWWC2
9faYQjPQQNjUI1R3B87CrmyBk7BlPNEpgm/+F9JUNofXpjeSBCf5sjJAihzJGeDB
1kYCuSjjM//oh7h4jvTI4BXl3tRqDyy0B/qNywyeC7TjAMVBhegPk6vOnmWJUKYu
O/yJP4iazzAW/mlMLyWDZeX/uVSzPAsuwYTJAMnRVfuEys7UmG914LQwOz/DtUqV
DKtr9vUioEPv4Le0079mDCtSHnDUeblVktlr2TQYn3ai+bmgjruaXH79Yg8BxhIm
83ibdFQ60elforbKEsmrVdkEFUtKyec5opfj5lECobvbXYRYmPWY2NEywyWZXAc/
z6xV4812UuDE16ADMTjTfupuPSVzIijoylxP/EvFoQWpegJ2tgO3x3eCiydio7yP
nq/JZ73Pj6jDw5pUVAGOPgDvVa9qnHVvScyo2ZTiVMlnqnnguYSxaJDraz0fLsLa
9WhPrw3+usEUHn+UtepywrSyZJ5Wrzj0ycfGDFnGbzqRkeQwrgWD3EGvAKikSAGH
c1fu2QxWyen4XlBYpWlmZuCyDrHf4Mb0MN3H3tSfSr/VmeGNF1TSAnTpmSGk+Ytd
CSBIHB6AUgDdhiELYCb7lB6DuOdii2Z0xAjqbJa5YG8zwbuISZFMv1IsQKnba5g/
zPdbAIcTCyPzc7u+9iSqMLuXH3Bh0x4H0cGOo1QUZMLMLwFPQzHXY5Mg4Lgzv6zf
cX8J58EgJmfh6T7Ott3KgXmQzzl1qBjtexXUaV4maCiQdkibD74rpPfqTDFP9O4l
QSBeX6bLKWRuQIGjYGne8xw9qOMREyulktJ1VN8TSCo/3wwEHNslTI5SIyip1XhP
fIHl/mvPA5eGu2Q63wK7HW9t9+82lyc+ln9ZOSjDkchyTo39BCHNE85ecEmPhDPC
mzKYDz5TZNtJOz+F++CeVsylnGV8DQP78pPmlhXmx/sKYWTBU4wA1OK67ZtpBph0
MwEsyngYRkMFSSUVUal2OOOvhhkoJUovEusjPsR53P6TFbMgElgtN1FwIHr8bvKU
np0qtQApnZabMCBnsgTVq+oNaUkzLN2iVMN9MDUX7hmLxe45o16xkMLS3pHDz+pg
dnM0zMeNnIy1PVXp5wj2PfSPgtUmMfDvK27Ewp9yTvp7KTWeFU4nB8XJFBqA8orY
I6cEzlhSnSx+9MsAIwnEPfNdYLnk6A/6NLJNE21+kvpwAKbo3LKOP4Ov1hw24ahh
Kz1CedCggAIaYt0DDcKy9Gx+tvfZQRlxz0cwiC2OQq2xAU2avrEpnCg9LZJyyKN7
ptru834wCP3/yl6YGFn309xJYVtZH34rBKyAuCIv580CyE0lpAALSHElnxrkvwDa
AQALw1TzFye2j16pewDpBIenBdCvpyxJkYYsXrwb5vIaGpteI9nNcLyKORfO2Qnf
i3KQ1a/lVJOe5zhvMYQmhZmZxqLEI1AX3eNwbZGbEXoYkbPdsEGlnRtZn+J5soLi
WGF1DpBvN+GY5CmFlgMS+01phTiA3Ziy8IieaYaC/Dx3aHHE6GV+tmFqJxMJTDIz
QmyOZpqI2wR4FmFfIu3C/zz+gWHm/l7WE7vgv5Mlh9rl0pAzbijaujCDY33YwEp+
Fu8O48YkalBhl/yQHGiD6a9i+niAubUzeYvbmD6Iv5QeBncmi5zk6qKm34uSpkkO
57cT/NxNHDpJwHztelO/LHJkk6CwGlwrKAUq37dmSzIU1BOQ9quWaaVwI2FlEi5c
PM2zQlZdIQ6AkaW2laTLdNIp0wHBlieu0gJkQ/GhGkGjZ/r3Pv/DLwxuH0rQBrcv
I+t+g/dY+O/DZwIk+cxmM9AoVe2xL+TPQLv0DXAigNC8WyWvRdp2KdY03iJoXBrJ
bQKCBtpqouQGLghW0/SH9tLDtRd8uxg1/QRTZB+KOlHDoL1vrVDUWJ+sm5sFQ64N
/h79nKCICCENtkxOP3JQA8uoOTQGtlYjLJSvmCYxOzYRGMG2MhmCF12CYuK/3ZLx
iNetq0xnTd4xFrDqJFUHFWzLPvcol+fear33HkmqHO94uXwikxskYdzJdPt9mnQ8
bgSkoQHSeYBSWsRXwDW9ckuwGBVek5Ibyx+iYgcWOJgA8xAzRbpj+mVzhls91asz
JbASnDUI468jbo3ah3h7Sd8GpfQ9AOsYdf8zBYb2HwfBwjYzuKrDx5FVOGFZo0gl
MOMQjsaQ2/EwJ4WkvPE+XRjRR/X2NzJL0+Y6FPk60/1LcTirDmFOye2tL2BiZpZd
cMjnT0d6AhrEVgVesDLhzZmtGk4pughpSG4IqfmbkSwNB3TiQpCMhI8DqV+p4WnH
QduE2noL6AeEIbqSnNZVSvKhGWE97pmnI3eLU/1HAXb8eakiIe15qWJ3nODc0Pu9
longYFprkNSGb8oYFl6IYgluI7xHD+FY9FDuK7TdpRYR5sSSSBORXnAwOWZhaS6F
/EoIzJo5d7YJxT54uJPU9aSzt/CCJu5HH5Gi+TocFFcc/amCTgN0evKREIcyFij7
b9YUBwu/VRUJqlWX8LCfhm5R0Gbtk4HK7jp9+dyfxTHXX+/pz3V1AScDw6tHSUDz
notCgORtVAq1bHaNeOYohQObblWM+acI3usdOmRmw/XJo3OetNwyEJ8jLzgMmHWa
tEUo2c7Fg0yR9eRXc+Q7ACTzSMnANnkRnQf9WtmeeewaEFCPBgVgfDN670R2ACG5
OjbTW6SSuXwxnjo9npE8pPmC/i+ZweIiEKpXu8xps7obuDmsKEfCxFbdb7flSEQb
AkKJ+bdFEFb0NOnRa2JFOTz3LILPZ0CxULvLTHerx/3FvXTVXSsem3nSDvimt01e
2BxdqpMBbVI9/tNYSS/hOkya2lrxlOaJHPNKAS0DR0kH5vQfARtM9s1OBXABeas4
NNmw/rOxwgT/hzHwej5z7EuXUKhkcPk9E34UrNQv10ZJ9BOMrjLNKhfl8bjdmWSG
7nuVZb5Pj0z6MtbUfOu4RWaPa23VMcVi/ghhWRHRX1mFvPf8dCI9YU+dCP3HLixC
ptwMqbdAUZn0gPll3yNn8mdGMMV2WTNe+lwwmH0Q+jY0h8bNnqcx5+O5ZZumIKWb
RPlpA3ipo2YdjO5kcxBs2t6Ko6eIdm/eUn4KI8ueANjaNg18BPFX2ocideWxFbTk
aqMn5UGiQVpIOgeYvT50MAobS2Ucy25EFpwbyLsxj2XJMbWbEbkDO1iu180j8Pht
JzqeeDIV0woftNQ7DkjljNFnBLIxvO7V7csO//cf68PbyutRdrDqXRIcOLyV/sCC
Y2SrnkJrNR3zRu693XFgCxuxLjLR8gPgr+0IyQ6h0ewamIf8OV6lQYEGnDqF0vW7
jSTJCKdR3A1xfdqJ6LiR7KZOtHveCCt4FfLwS044WkPPHB+ZlO5aj4Fym76dclna
GE+WRgpSjJkUCtv+xAOJ3/7jwoVGrjzeidS0UrhGlSSfEyubZPHVx/rlOsxXXmRT
ceHnjUxsG8MMVw3eyACjqak7zUpTLEWOUECEc7DhJF1PKU05WN3P+H4DE5CR18ZL
x7wZORQjoQ6JGlDgTObU9sD1lqHY5AWH9d2p+6/vNQ698u00CZbLUx/VeQ2YYcE6
EKgOQE5aq7atQxZ1nUDcbyyXizY7vGuq3krwqn/1OeuQgOv3gm+R5QLP0jf1euWL
9MYO79eFIKgIg6dTsHx67Zk/LHvVFYXBxLiG9sNh/5+uuFjiuPg+gKsoAYA+Emmv
Zr90EZWz6FKQ6kGUqzUFIEYrvNBtK6J91jf46BDycKKkIWnu6Bz/JKS6G783xfPe
OGrRmfmraINrZKfxCabALr55Fs2AuLaZ+Cb1a1K0EwGzUqrUa4yOfyFJMrMIZrci
mHKtIVFtPJ/YMVtMIFGtRr2aeJR3ZUC17qPv+yfvUXpU2o4BNCkNK8d05a5IfEEA
PFuUPRSHpmflLZDIwFVxDfjt9oRCdgJKBJSfUtMHEGPZ2zbQtw5+k+yfBhxFEs4P
y9jFIZbqIiCLiB6R2g6uZWj3lj5uj5/DasUz7oKpqHUGL6JvorZT4qR+NZ1wk54Y
LLB9fub4BxW/lx+uh4bdoUCwEPSRKm7HyQv9uQ5LwLsIExxuhaDVre5xYGmHRoXc
5jBcHJtuteQHoHZK6QkSAcC7CL+lVj6R3xIgyu2kBHWhT/cyx/PD805BOujWqPg1
RFkWP1mH8pnsR2aThwSfRCZdYzRBeIpGbNJZIz0Cu0tGYs+lEoga1JDIQS48paoK
a00f+1UUvsycqeu1L46/VzEp+9TXE0snPLeXoOC79viO3Wga+0eMbIXaZRqNaNHT
tOkdSVbhpR81yI1Tmmcq+pDVYg4zRCgyjDS16RF7EcoRhCCB9/fjEqM9MiSA6iL6
UzEpu89i2FCE7Q7RUi576NuyZFk3JtcYnLFhHgaI0u2fBUYtENggvr4B7eBrp37o
de8LJptTJY82lI5IrOmpLZSTU37bP+nFtDm7ynHIhmO+83r4rxCGlFUnR8brvd9a
Vuoxcicwmicc/uiHnC6zbc0x5DWHFXuaV5Qqkyr18eMhScYwcKzxwhg35Vfth1k4
dAm+hbUB9nQxFgo30iheHxiU3eO+8LoV1FyNME8BlDyRfD9WJLm1XoWn/4hIyNAh
vZ47uBVn1QqIwiJmZQY+h59wfCe2QVkQLXbgxLdQNVU/Josr1MxpCDYtyjlULhV5
F6ZNhkUcXiY5c7v4VhJloqFzlcVCNDOFaE1SOulBXL4Al0vaYA/NUuPhfgGY+K4c
FufFo//Vx2Zh1LY4pSaWlI5KmlOF2uxfMGNgz1k4qhmHAAYXWqgDteHeqmWfR80H
1XhQQDp6ITNSdN/twqXINWoDXACncNOjo/Iu156KalaQfPFFHx5gs7Kvi9Mjkpcb
xqKLUelLkUVzYgv+hLX59lbqVwfNodSJmUagIcpmtDreLKZNXfULXV48EkwQS5yZ
wLagCR8DOo4o8G2K/IOZQ3dve1q8ypgNZpJzVQIcHcm+oHM9YEPdXhCNIl22Q6Nu
IW0RNTiLBaf+fvenq2e0VVTOQNILdJv6SP3Vzm+6ZYCZs0crMD6gQzPdbmJXiOU7
2/BBLG0h3se8xbDNN1IKQ+aKvu/twvknC3KM8iTyaQhavjfDzHr3wn/QJJ6Az/tx
ZiLImENSvUjTm9Q/J1nfy86d7xUylz5ujNHHxxbv++ycAuRHXVgLfwZ01/ScSBOf
yEoDNp+OKB/o8Yq7xiwkdNaDUADPgJoo8eLek3nM8NamMXfzBMCzXffu4y6+fmtb
HVpi2IFa7buXUQDM5CIfZWyfh7S/fleytAVczWiBV/Trr2IUC4yeoiWnHPvrsQlN
Ougkj6JM66ma4bIHAdqcPeBHltdOZn3Dtt8SZR7Yb2/4lMXnBLF7fH8GyAzRGUa/
xsQ8WNpyBHSQOc+nQBLOZ56zJuctN90zFjxQ+sRarBiQ3S6LdhtXhMcOyNPuu6VK
Y7oHG8MHsDoLZGws1lC9Qu+GvlbrL7FmQl4Lj3vDepjs17IuL9Abe5wKMbhhxvhI
Yv4NT97xvbQROOqmttR4zUi2AlvP+wOvnyjsRd50AfVUnVbZnCxWon+G5K/vghdK
7FiocBtFS681zpKPY/fggXfnHJKC1sFoTTxt7IaaKBLT/YtcJdXfLK5vtsSLyn1S
bn35uCSDKvxpeJOhpGGXaID9m/pLd96NQBRZOIWq1AjnIvfUF49xHGReYzE8QGoT
ANe0pqQMlxeRMGTJCPKtd8/GgfL9V6wAMvAGNIeJF5FbCAKDC6Yu0DvDyGc1KxIA
Bduzb2MitJLxKBIt5Tc4++WfJKUJ6vO58F0+qAY1PGhPIlrdT0el8ov61jkHlftj
qDA3ddqDYiQJ62GyYZSfNLKlNMuWHvBxBDtVXXrAIlnYfnFiqn1+FeB05SR09Poo
TSxbkKDiJhZqwnKllReZ6cUd/nuzRF3sTOuVcqc52d+wyY8CZkQozT5X6Pslp1vY
nSMTLjS4jXBPFj3i37CHyH4/06rGucBBM5+GAWdNvvXIgVe+NRZuXnvWUBzgDK6t
ziz3nVL8ot07aVSQn7kQ9rHgDbcNkp9NjX79wiKxo33DAH8HCJSmE54Cz4xxh9xz
5OF31eyknVT45Be1W/g6NL8VYUUAviVm1NdGR9Xs09CrZwK9i1P+xp/HC1tGdjWf
3xnc0EB+AQN98OejCYoR692FsmlREZgJy9v5KF31aPy8QZW7OJCjjsWaX7GPUIp3
errIPOzOG0ApdaQ3WbpWQ00dJaWW/4rIY72uUiTvkvztqXY7udHBzNfGEQz6ZY5S
YgUnkDz+DeRC5Ig80NVGXfBk/nl7lwyC7gzyrryfQu7CDjn5l9Xe4dosPf+1qIGg
taPyt2evehujwaR33ANzQM/Y0w7sNXSPfctUEM1xNFexgNHDx4ziX6NqRwGmSLXn
z4kQIqYCqkNat54mmDwNcOS3DBKpuqKQ9gaec60ZT63Sqr1oTIyDb2vlrnp7zMw0
66EuGDMtQEkJZiq0kd8s0i7zBBHDzGUn+etCl1t3+gaxYn0VEXnlfjSOABwxMdj9
ipvhcdQLLr5oM5Q9wiilmrU6Mz1ujV8OPTYdN6gs3jVgQN8Vel/jeD/85mb6Roi2
u9aoSMeeInQMwlMNNM/fNEe1MuJ8EP97gE55oaKfgAIzpJgDtPJn+N9yFbvMmvFt
vQ7u0qeZgCDppZRBtTzp9l4FII89wPLCgYzWgbm1/iAF7Rt1nZw+PUM+mu4gXEpM
U8oQ4t0nwTdGtKUeOqIrz+d26xCry5aN6vW/UOKcH5WUOEUgH9oveRKSVkp2c1OX
ftmUXubNiohD4S/8rJ5JfvSgq/L6XWHidvIEUs1VgOTjkyCQqlQTMg9gm4a317LC
zPZqc5ny9sCcibXsdPGTZdWDUu3gsMPOEIZzWGRq+NvLjLXrUgilURTzA9xrJVbV
+j0if8z8sMDGFDtIMJNu3yHBdYt9+l76bM1GQyug2yUixzkTHXe3hkLKP3kwnKH3
XkneRySX8YNNokjSfoWOKedTO45TJWpxeL14r/9LiHtacs94S1l3VVedrVAEyr7y
ddii2yYurZupbP+rlY/DfTaLsELx4xe/c2uqHoP5N/AYLIUElWkKWkxL8cBmdhdE
20WOYqr7GmKG03xM2kd5PLrGTfbXOKmrw6Vy76xMvY7lWTD5rNlvdF3GNoQs04Sa
UqH/ya/TaCLcwvRn21vuejAd9e8WYQF0Fg4ZrYiQXfJ0qnycqq4nPpSD3YWxIZEo
rIQiSAIVPxZOnAS9yCaASF4EHde31XshNvj15UjbVN/0ID8axHuVaaKa1kyYhs5J
/d+2GtruH13DcvJcrihhfbWkPb0SdrNgol7NMHeH5qcRiyP0y/gkdmrTTXve1CCU
CIym8BhcCCIRWx/PI/LriwTnyB3WJxqGnBHoD//0GQi4cCqVHmNAfXJxwqHzz1i5
2INZPQ/ZRStVfSQzUqZ5B+m/3eswc5BvvRNE5XufMhAogI6mDGD63Dn6B78PKXJx
GFXl5R+ZvEMX8ZRKTX+QFSIQmwA/5DjdoAfwvSUNl5bOlKXiYl9kyBYBRben81dk
aOlTVov4FRnt7zidF27Zz/g/9YDT1d4ktC0rP7IFPXykjfMucBtH8232E0fhslO+
tWs9450hYo9SN8PZOgJBZEDHzpRj6IcS6SqRyYDV8ai9deEkbYY9F+LjsD/XpjHR
2xvbTJBfO8flB7CofkJsDgOcCkqQtCtNv8BilFxipJ6ZEI2Z4tPwFBSTcYWUftBv
ZZOeEIqgvl82MtcmzG2kl7NBaQZFYSVKtOlVP1Z4x4NtIXAeDKtfU+qD5KWmqlRt
NdwvbxhdrtSstCUh2AdNsxO5TU8NUk1g8o+Dulnl9iDY/2ouVrxR9qB+qiy5Lrlu
ua+c2qpZ+8L2vOVS6H9lQKQY4ISgsipkJwACEDBKEdDEYXYCcB3nMlUAYzD7qqvy
4bdPmNQAO2o8telIs8kVO1SgMdWaT6u+3ipj4rfvn1V3H5tIp/yRe9h6UEpMP7Xz
hKoWYkhcwswq/k4EbPb27ivwxnkuvbrc7zmZhXkuVkWr8dSkLfmM4L5z8tXSSr2b
SvGnpB5khtXsXCU1A+hAMTkI9GXb3v7bzVAHi0waUSUE9atDeGT3yM+hK5NPBjyH
wKV5pIcNO61f9VifcdW2k+wUcNNvWHpEQupyigdcK2r4dcHYFSlB8W9NW7uULlJQ
+MV0T1zyxCFzthCA/7j0/beH+Tp0yIRXHG2z1wYikWiZvM9bMwjGaU49ePdNmklr
c1ySXGfj24xPQ5S/Swa5NefVf+iwCX7O9RbXb23kUCATz8R15t9/Jzc6JYDMhbRN
31z8zP/OmUlWT5OBNZMjiDCG5S2fqCN6tIUAkwaDoKt5iuoeWzFZgF9CkfAHiy6n
GYgrKHhG9lLOoxRDysyCFCF2KDRv7tj4SphhBibH5QMnTh+c5AAxNaltVHPX7Ytf
x3+8x2Li2ySN5L1JtSqhSPdFtocZyiF6d9lgNaMQ+Go881Z/I5X0NNleRkEV17a/
rDV2kpP481IbPgFxFV9vjWpkHmO2O+5JCqmxhCPet+DznDgouqq3zTuh/swcBZKD
p0wUUzC5HZI4zTKOLjQ1Z5UPNTynYj6vQnXAQPnXdUjlARCELHITWghDRcAckmDd
9/qOYM5TS6qtW9SJP6SDZnHK+oZBtyMhA+zkBPIspk/glw6Z21DMz2h/Xk6AmCRM
3MQUJWQbVPy08HrprlZ0jBHAH+eLpDq1bV5RYTSwh0GEx0NoubnV/T78YJG26ffW
TynzSEyzdwKvw6gKpzVR6HlNgIX8nPztTYCXO2d5fJPt5U4nrWZZ/40t7qoAA7Tb
sdEmm3uRizXhj04xHGPb8NP/5d3t3SjaKAbcFgNnShxowm5pUP5WpvtFTp4/59mB
J0qcPuZCQUGd0jIwZNqhvWD043I/EIU21OHNQ3HY8OvJOYZFgn12G+7KTqN69HZO
/lBPB5s9XBULuC7qHp8mSsy0xLYaC3pwZSt5oj9e4iBuSUeHlU+mNFwgOosRcghk
cWuqtzJfUsmgaBHVYbXxIb1+GfRa55fAQHFQ7sFpr1iS/CHOOoVW5u/ezwGrtiR0
EClbf6NDRL6atC6fUL+E3BTgTkaFL87GILcnoB4O3r6Hqx0EwMzQssmMF2uh4sBu
Tp7up22cEcsPSXARq8qKG0GX1L8ZjKrPtHkaQ3FcLWrIBCorHoEmSs1kn/UVpq1o
RLJvih+qgbmrHDES4uhZmEGjL10fCxcPfHPCeFlOAjdy/gZ1IYzE1pYymgCmJuYi
qCVBwlLG/NIGYI7H0jpReYNrmalb4NNpp7JJRjCmikGpDtjgf0e4TbREXQo1SO1u
HIyjukog1pFtqCNw50sN/oOAuFRtcJFzxIIl8VKd5ThxTTiDfi0xNPoa3LIxlSyJ
7sku8Hs+9R/Ki7/9CyDHABBPBkd4IBKdqnuXv+Rw+YCfDq9uAMTlCwADMrc5+2wv
mBn4ehdYYj4dbdLlilAFJc0SJ4vafNxbg6VL+2PZjrFd3CdTo5756Vf0p0Gjqw6s
lXXfzle9eJ4aq3EpOZd6H1gCfOOJXWgxD/xcnFKGLXW4jwn7qrLjDBM2b+fLuE4Z
nZS36rhNMC3I7FDArkmbrWY7xG7WzCtLIC3sn55DFJ99U0PvgguDrd36/2o7dJcZ
UUP7S0XfUdI8yumyGZZLqPYSqAZYCgvdC5S1bJ174XNpipZivyRO7YXiPmRQqJ2l
UA4f0wlegwxF5NWgYsdeAPHQiBAad6sgVgoVTqN+O0Z557/aB/RRkD7aj4Q5AJEn
GwHIVwbfdSp6nOroHe/ihLyIblN7Ga2bjNywmh2kAVOD2N5jfaruhL6bOyZKT8pS
i6Yb211NGxjGgVXZPWojt4Pq0YkEEVp6GNWgKqji6ri2Dn2sh240VNjw7lhf0Q+o
fkZelsITxTYr8cBy309Fk8UNiwZOcfBQZJ8m9/9L5YYNeEydT8NOtUcdr0xXNDKG
/yFh5TqfR/wujBNGPCVpaCjLm0CeMu2XT/9Md0xb4ogZUnjyMOmsnSOFfsF6fyqn
jq47w++a4qc93otkx/xoQmAgHtxIz0acAWcIo/iCwFURmkCHIdyXfiCFqLQNrCF5
8mZLuRyfhiNleAmGRB6pHmsM5ayXf6yVRt3IOQLm9/8bXstMCp+FQReyURaCuS8G
LG70RpIAE3GXS1m+fDsJ9+xD0Cvksm5rSk+uGJv7sYi4q+SEszpe3xZ/JKDP6fiS
qGe/sMsuVyNkO6KOqiwqAeTZjVpChDReqhGRUD8bXeEQ7PJ3wRPMXP0qz8DoqAoa
fzahEnZajo3pmmlu005qpHzMLSqzuhxGjA4XHveDJKrMtr9x9uClXZe96n0DgiKN
SphQVYK1c9qBBg4Venay5ozDA2NN80k7vLF7jW3+SwNh19aw6zcMxhpvq5lmCq7E
irFXP+YLMLG6lLlty80haWYina+D6WHetNmCjvvejMRTs57bgkR7DTM5TD75c56k
oYjSdWuBHijI6i9tv64mvVc8bgMQRrYpJlB/MDU7QbbxHIsKWhjkunuYTyuMOgnn
n3hREG5swJ1SpqTyfoP1pOrZVA7x+5owG1FRp0IBnhQUK+gAnMkw65ncAtWO8TGq
MQ1QR5PG0+2jy+N2q5h3bXKxLuZ++jFb5+IRqKs8ACKqUBO7+3ddXe3VkY4tWafH
gy4lKwZQSNLWpeFGKNVWXf7EEUI+UzcJnBjfHRdHB4v9tzjTa/AP4niwrQH6tIWS
NE0OrxtRoQ2BeNMk3SZoxebkvARjJpYgo4dPJCWizSbwBfRTXjzPyf1/qjWoszlu
RUKKfPyWlAQvbnLNioSiWyjUwDdqzO1+T0EZ7Kf3gN7PXwYfeUuDQ/8qNJV7J1Sd
jlyjHd8vpAbalQH6fKW8UhJPqF9lJi/vqk6hAAv8qq1p2BbngOvqRuJ58ykHHbLy
oEvvXq7yzWGPXksFPTSTJFUTog97JAepmUFLtIwG29txD8REWo20cHTp6WjeSw3c
5tuF4rGj+iks/ckYxvwn+zJLOPKeytEIzQNnXHaJ36RIhGWWzRPwsXdtV6ibSyCv
WkGMaJsvBM63XLZ7BOhOQvBWpKV7RdqfXTPyBaDD/CQatrN4aEfgy7cGlWnTvFvt
cLZrrrity/uyIS3GqR18zQbN6qOADCB3bajQLqSvexFnCMfT1WhVGk1iHbv1yygn
o7bafE1ez6vuo41meN52Q6ABQ+qkv9RsWTcH4ZN0wBkcf6t12dM8W1m/53pQ6Iwv
jN9wPNrUqG6m2/cYCxb5Wf4X5XerqsZcZc9EPlOZHW9P/Y6nSHqCALFiC6qLIzRW
ME5Vfj7uidlEXIj38nv9cF/1wpOH3qNK+c7RYkEzlJ3CRZ4LGSwL8mgrnhKwGgyH
Jjp2TgvfTdTcxOywOUufPlZSOEBGdMVl7yM7yCxeeVgIat6loeSiUxN5OTT85g16
rPP/1WV/FwLhQncMuKNwjUSOO99C7jJhjO2LT+QqPiTVt3zLmOVlcqa2tnV+lPRP
ZbNENZKSX94sjyaSbYMnON8+HZUkKB1jFj6CjgiDbeNRmMNrUqdrW5c4mbYM9Pqw
iNCom00J1gpzYc5LAC4EF5fX2ciTzAu/mu1iV7eWPQEK5KVNzH7OCb5HtsHMfS7O
Ifqh35e6+rdlpZc11Z2jRzXQ6/hXOJieH/ELn0Ir0/LCMOgXqEz2E2OnVSKupwbu
RtwdnobeEF+/Nzq3zH17Rz8dBJ1W+/VzrBo1R8xtp6I3/ivNDKYsy4NNm07xedAJ
184nnykcTLzkMz3o4DYP9LZ7MVbtlKvMPHkdDVKndjrDp+JHUnU0pHW8fSDHsiuI
m4AVE4VFkq4qMBCIbclECm6wvLpE1ij5Tz1vaYdcMAvydLEM7nyATEQ9HaOj5sl4
zijj+vGgg4ClZnr6OI/eVGsFRo08p+XkIuu8HrRioTvGL5RI35lSrg3cKZhwX9ae
6gpm2eid8DYsSFz/kcR5kuT1sya4XBcWUMcX+pZJOtTVJDrY629OG8erWpu0VXhu
E77SSBdjbKj2uCsibt5d9KaqvN+LgHzIkBu/fUwyN7iW1GYrZCBy0cni7Pe//FkT
+TYgJJkQELH1Sr8HKUszBTBwjNj//ndLR3JdujiG7xznFgvKYrmAJ+jw01fOBLAz
LB+xY5gK6RIPBQqPlcK8AhR9qIY3jHj/Lc+shQ5ieoTkoibgDh7tWHy2wzQjV9I0
lttuRTQcl6j0TcEw7UyYj5tRmFx4cs1vM/7vTmVksHYuvfhM23mds1IRPjwFDk9R
yRISvIJAggptT9DwDh7ny6vuffw53BAS9Olqg+AoZSMSyrcIXf2OumaaWoLPmWK5
fqcGucXYVY61OCvRlbOkLxcMh3xD6tXSAUQSYkTxkrUgYLDhoRvwMmSR1N/AW4Za
Nv+mrK0QVYhzc37tWYseVT9DdBD/DKr3E2ZthbUNmokGrvgb8iS1nAhk+Vjva2Cu
fl5M6u5u9mx7nGW6HfsRgv2UUEhp/TjGvPSrLlpC8ouTuO87fytueisDfv/qfdGV
zF7x1+77ZBv1TMMfIKqBlN8r7WtZ9SkTdUKc+sHIEHri7knv+w6HgzFiR4v3rSEu
XLjBUJD9j8mXfCg4V0MRA81gAdElgGgowrhznzit8m9YbVeuYhkZ92tX4C1RTnUF
fdnwWCWiWOK9CAqHgBQW6BoLYwMEHuZA9clCq+Dj+WapkbGEFo2sfzgociUa3ZIj
gL4j9TsjHz1KkACWVnVVc+OlpW+mfoMmpYdEZZVsDYmKe+B0X/Dxk3U6hjGq9w6t
BmzGUTrF//5UNWlczH5/W07C3vTjwjXqxvDgUglcG2jLTxK2MZKoVRZQowiM87wd
yNxJqrZSMSRvWsFY7ZgWfRj+zz14uW1macnwnnz5gNalxzhsjY+5zFNcHP663VLH
D9YZ8oWZTrnbuzpN873q9Q9lSGGN1G07X8s16dVhLQEQjZVbrOjhn7nEaJVBcctH
zRCDzYRs7/z8+ZQxoSlhOpiMay+OnECeJow/hb+IraJJx9zNMltOuHqzjDKkQ2Hw
lDme/YkFSPIQ+lyPqrPosc08W1ktJ3i7JJv/jQdrxax0NEdCukGbI+vmy61K7JDs
d0/CrIE479enFbMnxMUHVeDlVaWQbwr5sVEivsp79wbEcjZjmc7yHiiRsZeyWoo2
9/SaGKdEpPKmookELeWU1dYAo7Qi9/E+BkJM+kWRXPVC+WlLobm3XCoD4rYuY5nM
CH123KJNeKHQ18CsTRw5PBsEyXbf2Yq7pnUjPbiqH9UITcNAeTfEGrqOoeKBmvIl
uETJdUECgFSQp/OQfu15uJ6mN+BUIdK+B2V3xR2/2mKahIZZcU5nUhEsr8Y+qNyh
x7xhDr2FoY+0A612opQTTWnNhIs9pDiWZT1CtZptYrV1MJjLDXn4PIJ8uO4D7wvr
DqwqeU5jUoStN8p2WXgvqAomv7PDYEdAcakcOXgt+B5tOH9dWmuq8gDIdszAfQyP
HKXAuMiSYWmF1vLCOKDq3zcHeD9ReMgRzu1y9ngb44FL6vUaT+/xJIq2kOmZbGiN
TzPlqk5RrjsHcAB/j/JR12dKIGWnLHTvfdvJHmT1gzz2qJvyAoSHvF+w6/zMhl1x
Xo7c5wLBFrif0qtTWpzMPynG7HP0m0Nd4wpDJ+RA2HCSoe4M9lZ6wS9BWe+wJ44p
s+PIwe++6r1ISFNkjKPLSr/gxrEPZ4fRN4ecnhFBG45MeeNAxqqs+NGo4tqKzpPm
JYsVlHwYsa2Dn+5UCf+04rEGA3BdGKhB+x5FxCYUKaUhOASiA0x6KM6VtmaSxas8
Y9GQGJ+eyqve1CaKK3A2TWdfsP9lBK8vh7f0dGudDn9gVBoYU2kfBC92ShYZsRe1
p88T3g2OO31SOI9ZZVBgHUa+6TwyhjujVE7EiQ6pFfOGebkN4uS7oPBRzua/wTdJ
j4Zmvqvy1M9j7wR9hbxuu6UnUlygvNCsWSKfl4p4EPUTGy+Rv465MblVIeEe9kej
vlIp0UcgXtd/sUuS9O8g28J+f6L7JK9NXK3+sOpX/4dFrYCmzQEfwsLGSEwzYHVY
Kri9LM/0/TBYDwEmnjnHlvrsVVyyJjVDZi0hjBWrm2V98n265HU30oNguPRV9KHn
7zdsdJMbLX68rEcSdDZDaOBxES02YID/0AeaFD2rsxfEQuqw/GwYyGuRp1W6YxVP
pv0FxFbVaDPY9Y5GfSPJKm90SlJI/VSSNAhRcE2kJSfLaEtT9UiPqX1anRrF313u
0EbgYlWcbwzwHbstdtEigzZOLSNn4hVetYGBk+TuT+23QXkVXNaueNuY9Ad0kprM
bEOjwZBEGBcHqdDO84UKkI5KyVF+E10ttzeG8lzTUbfiemwf30pB8JeHMhBW26s2
cAi3iH9w+JKSw564bc1uRJCRNJQXWZt3Dz1zyYNc3DztOPcjfTB5LF6hOvEmyqZx
435Um2D15rkYX2vQ5mZvTQUH4g60n5F9zppqM3c5fIchaVDd61eI4MB/l4zg7Qj8
2hg5n/NgPj+BAO6esu7taSiQ+2n1TzSKGrCQKcQeytiTD/u9NfpKAGS2gNCFIwji
7fnghuVUZxEFdGZhsOBSEbCbuftM7UW1oi3j7g/1fcPxi8SizhvHTydklLS9QAqu
7nCxetQ/tzlDpRvoz3Ua4ACUZ3tMdCb/viUTn//IUVOmj5UwROF7x/4m73XH6oAQ
Qrz0RZi8/B7k8mwxrrzL3ngs44ECfvl8g4Br7u2bMcqtnrFf4r/psb8UMIO4mjda
Ll7m6x0jxAvgDeDsJipe+BKsoE0LgvDw4RXSkEcshntus8ps0yLvYOnRQbilg3cG
uAjeIZ++GzT1VQT1OaMkg0pB6s18hnYsi2ggH3HMI1v5wE4BR+NN5pleaZZV9G/G
+ikTZyFVQedY+tqdLB8dPk6Af8TPJR81k0ssosvYbheZkfTNUTXWjTTc7+WgQblh
ffzFnI1cYWaK0Q7xyujju4YJHkKDvfwdxb9qjf819cY4svklMQnBzBCxOkTjOkio
rL5VpwTw0tbvslJbxiXDbqgANKwkxqFIaQJJ60hW0gQXqErhmNhhpUssjYtAnhY5
5FSHeXfR/AUeieF8y6NXF/2CZbOj6ksG2mpmJKsB+WLosS7hyndKj0zCXgjcNGxB
YznqBrwfmMVzn074uYTXtAYt+RJAWggJj51XnY2sv4Y27hf9a8kt1+UPeDa3Hm3T
ZnufN8UKNYx4YutvHYOjYEHL2cU5XhZqrtokhF2R+Q5wYMFUj9YUCIaZ7vVHUTZH
SGEF4d/WHlZqxSonDeuwAoMKK2modiZzIFgT+i25ngyaAqvcDNE+u7mNPpf64Q2Q
h/WTMnMyof8kUM+XyH8EXn4ae6iUdQS0IyB3t/8z8Ow1ObNF2k/F6rUt+vaTcyFE
R8ENijYv6yB6xXqgtsCxl1eNQI6tkrf2OvJj/mgC4M5h2Yc1LND7kfNnT750LHVP
J3DGuh8mXkgY3LbnTHUar0XAjQp+CYO7o3ouK12gkFz4SNZaJzscN+NNd/1p71cF
BTCiScM0fS3k7prBwkecw63SlKiHLXEa8wKyZ7qNcF3MVJjs3EcVJu+tIUJRDZjn
jHAVIfXEwn+tniBh3/Va79KOF7idWTWpdplwwgNwkTO+oJ9jSg85bZRW8fMOFDnx
FGN36N5FxOQ1CD1c05dPFcxxtmwR8wJf7DWVEXtsjoRNygKS+1mk6n0FmZnwuksR
h81Tzn9ks0v5xsellS3FnikMylOLb2+dhIHgLo8n2RPZ91fN+Vf7G6JXAo//1EgU
jOwPc+4X+IVuka/PKhW6C+pnpZuue2lYy5M0JcH3RKYDOD75x4ahGDIulNQf70TQ
1+Zm3KTOSSU5o8UptnxZaKpqHQPllazlHAOkS6OVZcFY77bXrhA5W7744xdxTHho
iSjBiGFoinEMQFqfmsvFNLQCLT97tss+bkBrIMvRQPEz1elTDx4EzCkWq3R48Rb5
5mtzVqH4FKtMGDgLxuwDxMG/bH9jFf7KWkwDbuNvNqChv4QDXIq22/EKgZrKSF4Y
6Fg98DJIdb67UNkGy+sV6eejkcacCOUrQ9IHZyQGLyrRrfVzbMLZqlhlku8uEBfL
9zSQoy1PnbI+UVyKZEwahUuf1u2YThY1x1Sx4hQ6QNJhhQ2grLDUMr3SkYjmR6wu
kQefN78Bb9csxT+GSuIBOC73QgAG4lGDFzeDZ1SRJXd0VPUQzJQqLKNJ6Jonsa/o
wh6utkNtERFu2SuJeS+QUj9iyyVVCtf03fv/yAICkBE2AczbqDWi4g3pYb/hiqem
lndtiDEJVLjXWvZB1HI17xXJkMoDvczD08U/PcaVcuU4tHVe2kBnER136mY9+G89
DRnqcKLwfkIgTwEPixlzTB0SdQDajCEnMO6TXRJZ+60fk3gjRz3XhHjPAUYxYAty
pHrKIj7GUeNSrOPmwJfkKOLA62dxE29XMYtcwGnrSp9csWNNaqC7GB2bd1T6FxNi
yhxbHqQU/fkT/6MRFyrBnBPQZb+a1tPBnkfFyfHuLf5ZW7NUDxSTWdbYHmQBtBQ5
7eQPuXOlrp4VdQADDAFaUSCs7PDqbg56q/ZuaXVplQEQUYSQG/7jYhm8Xz5XcWGD
lBLwibHJQJTzP0aARtsXyIIUcObExVCTPLtwYvfVZy90neWPPR+0CJui0F/T1t6a
3WUszKjm52aDLLmnUNjLzqSuT4EsVvj6fzVbwTU4o4tfecYxmLHf7hipdZlf8DsV
1qU94rLXM1NIGDNRRTsEsJ5bv474WCR69YjGFbS7cS7Pd+G7AlQWtroZguE9F9uv
DLslfdaPtC3QSAP+dtBZxzHMZfnJNvy6XnJ1CJCp3hpeDLFQt/Cp/kOs/L81T+Yz
wYEPOFO4dLpMNsC+9JhGRFHLCb2k11qxUOOn1gz6TpBQO/zR9xhiGDx2m/fGGTVE
FcdmhU0w6BM1i6HGNBs3f1ruu+8XKBUZI3OlnmikotXLuIPR5/BKdTMjH5Zk8geg
T29NvzM5keN9i4hKCE6NcHFCB25pu3tcrG5aP9Rk29S67Q6/0BqkbvcqrYaOr8Jn
DCOHgFHYddW7eG6g8CH+J5dGbubhYF/ZlDCsW1wr4isDLze0JpYd2djs9wUorqAG
pYfpaA1VTfRHoOoPHD8F37ccvT1AhCRBKt3Oqnz02uWEa/y+mhkZuPIVUh2E5AKK
8Mc6YTnBNb7riasKUPSkleaQj0rVQa0Kgs/hGCOSHWvK4LaXVkmk6T84or8c7td9
BT0dDU8y1wz2JcQeXDzIVv0k1XNRwipopaHaGyh5/RDlzRSL+tdy6qj1HG9mUBXf
V3ueoTZWyr24eicCq3q+7JgqXz51Wj5wgY/Dikfo6CcczKvbnEiN56MdqoWuddsw
p8RsLnqStn4ZVodTfuOsjCqkSZD6dpJu35TlftjZU3GR911BlA/5o+rtND/6icDq
XhzDlYlEExcMpNGCXxBU5RP4ZDPNAas+08VE7xmTphRtrtRmIC2qKmsOb9TIdMri
d3PMFb9vvWhAHtgnnAtl0mMWhQIUxbPk0/Phs+3ERlkDw8SW0L4BVb4gV8QAjcgX
KEiUA5bGZxz7IBjY41ldrVPZDIroKJtL2d7faqhl4/E59kRo21qF+FaAhMsy4sMV
eMiBMs/3jCXlaYZ7jldgpv8wJhz6zlI1G62yKKsdyODwgfGBl5ttKexCqin9+fo6
G/VBAEMNplPdf1W1D6TuWzhwt8lMZUQkOQzKF07vVOp9tqNNLNX3SeuYRkwod3/4
ETXg5I7QFU/NIoKGaAQd5oG3NJc3r/q7NxhC4uo9C8fpPZOI/O/1PCOAJNWUio9z
yIR3dSf9bzhci7xM+mNZWlOeSLwtl8+7gNyhR/RazflwHVOwi+bTMPhYRDibVs3u
6UMbCoMSyJ3SFC3EuMTdHqPJzyzYeM2qO0Pv+/wFMhwq3CfRg/Js2fwzqBfYgHlc
bPi8fBfdRsM4SZCEEwZ/w6go9Xe8Rh6AAvQyBhegZgTUfF1sM5Bd1T9UAsDQdrPb
UkfgHHGcSKE6DoWiwiZSyk9aUnvEEIqMLQlDRDCU5YRpNpZh68Gr+fsrFnmAP5D1
t7fGQupWCol1ZAJf+ht7kA2YEUoruFTH6iB7ACZeoBRdlS176Tk1rk9+8f0C+pfZ
wW5T/i3Q9QENUUXH/fkmHXFB7q8La7WwDnpFZ2Igis9ir7ijDvRlPa/BW2RvgCqg
mHvLhOdiOjiQwdj415Hx2ydfYmhEd6Y8neDUafa291TWe07ZaPRPiic9A4nCNl6i
sIPt4onxrg0Fz+LHb8m9M70ZZlh0GdM1C+hamdJVTYFfzkN+sBrC1w5mczHiS1VX
yNnSyoTGpv876xeHmIAvDuAhURtIzGbGB0p7aLdgokQLqpuNG5MXmjDezRwYJejL
jJQDi2+nNtdvSttIQaKzJp2GHhiOY0BwzxEHLARpY/MLygmrBWCP71IKvpZEPuOV
7gtWVrpiVzoliMuaCy4tF/rCQ6G03y6T3/z36YUvdO+oU47GmxmWa6WCUWTa5gYw
jwq/vWyFMubFIgZyIyDWq2Llo58SJk6w625eLGEEvMEkUCsHWQx7soa93fV1meJ1
qVmJisQZSQH0jYod8TVvxnAX95dBoWwc650qIOgS5oXrFCxSLokfwDAeXhMaIeDl
Jl7gqL6bVMTG1F1h9n4rMB874cSj1XYSIERgC1z30XQmkEuz+O+B8fZC9NecJc85
/Ik2WYuV5FBvwIkyZE7vsLAJ7wGuw6vBhdOXjzbSNjDq/SsA3Phc8IH0mNXiqcBd
QZg9pkXKWFbzKGhLYvjRawyZwwiiH2JTvEYcVLLtIV4CNF68IhbgOkpAfj0O/gF6
izT/lO8aVaHfSUBJGfOmUNeyJM4sL5sv+HM2uHQyLO7Qk2mJZMTeKAN75RJoBin1
2OAWA/Fpue6ineTi7eqovQJOBtG5C7yTyIg+4ybiUQXZ9RlSEELDQfBjLoEeXegm
2dv4QZDkXD1bUSgIYwIFu0SKvnx18aE6vbrmeXXJwjpbmHzuqm88CKmy/0bgNu3V
LJ85o5aiNk7IB+Uhwv8XEmXhDeSoCOwY4DB7a4GZS475D0lCtlLByRGoMvgO+c0S
+idLG8+hNE5TWXccjrimQWA/Murc0PTcAoOl52sMzwc+W3Nmo7UD4spcc4D8QVRM
UbHuarZqCvBtWl6B6DCNyy/LflxU4pDrd0WpA6pu6ltlFQHEMmfoR3Tz44fZslVH
HVRIct51kEEP2j0sbVi10WK38V0Iezb6a6TrfOJMDWRGV4vo2Hz/bYcRqLEFDccW
Ocl9HCK96jJZ3ZUQa1zZLF08CGJE1sLmHoloVcIjxjKOwNEN+6+ReZekK3vaSWkJ
Z8+vzSgHadTu35vdyTMUoOICxvYA+hHWElif07oxlIyiwFAcMUCvVkkHLv85I1tE
MnKO8/Bf5L6Cf1z+5IVnux9eehAa96BB4oCUjcMyl27KuKLpMrCr+XJEZuJyQeiz
nQLy5YafuQqKZ+CAtZoyYdxQHty/nFwwoFiOsKPtlTXDw8gesHwmfG/nMtbFfJfs
oHTLyoDk/xIviCnZrxLznGdojBCwwPJMVSNkdwaKZPfkt/QFWkEbWcvIDX7Y6pWl
1H0BUS1QfKHjnnLEt5RmktVgHK4sDFkcbMsKJNNG8jc7lsMItjS4bquy+kq4ivfj
aWIvVtDib5H6EleAOH9iD6AxAAWHyw0KrqWF5BuZ02K0IpIcJbPZuHoJ1gHNF5FI
JYSUm0f9udbeqYK8gPp72he+uW4Iu2R7BSHrBjCPLJ+q+85+2yAiMcUuUSxH9aIE
vJUYNeIOcZGFxr0falOQtNklU4VOMO7Ak+/C8RoxBAbeJNm6Jx8FAkRprANWltTc
YKeeTrwpL39ddYPCI/hmsRPlAEHw8ONLYoZD/5/A9JEdMRgIdWYUWCl8Q31pucec
gItfl8TaFARGbwhs3ezaxpSjwS2WAJ7idbmjDaTO9gA5H5HT3VU05c6od/KibV0W
AGCw0NuEiTdvCOptjeFE8qiDhzToEwiq/z27MqjtmWSpZ/1WCvkYDrol6ZyLr4vF
ooiSBRJ6ogrjCLs3OlckbHwz5vffZDEzPE6a+db1nay5xojDPJejEclwZ8cyC5H1
dnOk3ErUoS5LN5rC5y63xN4dIFRB/iPDg6EKXw2ENTOueiBaIdr6+laxKzCAMwub
cdOb5MwmAnMgAofwp+ooAiVFvu5AHDzzDnj3nfbnTOukb6gk++/ucpyvWbJjSStL
mfEmg0NjEp44Y6mHlkkE8MNtPiA+wRCArEeCq952cYHKObOcr8khBLFamq4xdYD+
MsiaGm13jzvw4TewxoDW8kNcCY7AmMXgI/N6vKxTlDAVEegxfeoB6IisGP1hkvNC
jS883792vBWB80PfEARjAR1S+RiUv5d/3w04B5dj6jviF0xqloXwMojoZ/iXeXwA
Cc459YodgGljEhDRm0zgEWlhPasljAqXiWjgXSxZnvUwY+AcQNX0GJAf5rvSxLQ8
QAzvyLvmsZQhRyjgzJisbUpq/zuQJT6GzBSeCG5ZPXaDYC5c0VmsRGtx3eNRDdWs
EeJ98wQei4vdYZQPS3IljgUUhOlnQwdIB///WpJlEfQ6WUgFY+127VNHOUAA4vMN
/pT8ADml61yip8HPROX4POvkoO9mkzFi6ncciRRCeJvt3FKgL6EPlvDZ5roLy9kF
Uwt1r9uIycnLeQ5ArdmN/yGyoPj0uYWzw0Hdeuz++gHyLd4ypY3UcRa0QzBzSqkl
0EHFRUgYNztJmm4l2b0CVq3wFOPGHu6KFNGIo39gYZJM/yFIANOFiTWBAs9B5uzZ
ZxZ/fRa/vcxHrcYy1POev9oYYRiYlOZ6wtNlF8hE/+abqRl9GRjjGX35srW82vZT
IZgmNPCqC2uInqAy8slyRkieu2+3hlP9knyNEwspIN6WRDFlURqdmTfcKrc44iWL
pDnSH/ZxNQ6qR4m/D2KjYJYr+mK94b2gbAfB7F6zo+doyRBzVDvo7UBL52aBv31u
UzgWZWsQWjC55etDTYAZX4YOV1lPrLqkBP+ZQZyw7Svr+iswnOLuEXGC6H7T+ekU
i7QnqtEiVadBmhPEoy+DSfVILvhvOCBi/Zk7QpnpzbZgXW7Bvj7HPMF0x/RP8N2e
S3zMnCKxPb1F1T7MuC2ZQ2JCB94icGWgkMPVNPs9NpJkPqlNAzA9vfTfV3diTnDh
w/vgp7+uVEfD214YquM/gnxbI502XOtvZx2zo2dqzD/XsM56sLVVHERvFgFM+ZRp
pU4J/D0ERBKjzHRteaVJ8cds3dp3OvWais70lGHBrdvlRVVEM57JWQi03ti+o++q
OCJUaiN3CyA+LR1L10VK1Vb2fwFQGp9cJRnrRG7kPbC2GUzwCAGxMBCqkqwxzQl9
OGB0yS8MKy3CtL+waswHB63SpSBODqU4MOmd8XJKYjUUAjO9s3vGKAIwpGjHpsDX
ui1Va5R3WNTh6XnJRDNtz3P6o0jSugfN81ttZH+rYzbDR/c2jnKw3XOym8Z+C2nR
3RspPsNM/T1TBqrUCeXCNXmkXgS9P9/q+AAjoda6yaeA/ks72Wawnu5FupLTcVcX
qs4mFwGE/LxqnT9RiYmx+MsKR+aWbGFZuuVQDcJXo0YaxBfqeGfHFmoq2mtik1gD
hd0Jb6cuULz4l6YG4SStXozax0Ckx4vXliPYJRbCr/kvhzC63m3ZCrMnCfC2fjJZ
Ln5rNyyTv2KAUrF9fW6VF7fLinTUdd8zA/3PFCuwcjxPIkCQpIiPewG2AzBVC6NP
XPfjFJ3YDQaJitgSBcAejf6VoPm7SjrH6rxa0FowI+Ey0WEz+hk/3JZKkjz6t/8n
zyOJA6mjgWJVrBVA15E2YDTj+G5e8WHnLojjod5CokYtYR/6WorLpH5rrISDYdZ8
DiSnH6fqCk2gSH5dEER4WK+ALUXqpHCy4gtFjMGJKFMMYcwRl2hNf3mNMkQ+Qcpq
guTcCGENUGL7jBg7zC5TT/jpjpHVXfi31iKBgX6TjQ40auHSqQZgnlTZl2K07xcL
snr91moD78cZobjwqc/ESo4JJuuqkmwGZlrqqC3cxK0JagG05dpLsK97MsG/uLP5
BraN9gwPUtXev1JhX1Wdmr4zFVJdNpuqWhlaXJ7G3iGtfJAPb5sGICWjVTOmRgor
nwyFx5Ztc1xqpmOFGMEWaDM5n4jJlWdOlhq9JgjiGurebipzlRnKrTpYcLMC8JgC
QIj+4wguCC2BCwHOfBHZMsYj+ipaERUPpzXNGYRlxbRXl/iwHa9gS1yO70jQLg8H
6YYwK8hzhDlYrbx54V+RHXc+mG9L0mzmwUW084rpAcvRADnPWOOeim6nlDw8bnvW
mzqSIZcAVa8tCiRPRH/eG/PkVeWGF0LXI4OD7Kd15ymxCLOJ1ATUOtfwbIqJteK2
BqCp5MWxdnKtikyPPOdUPzZrEDqqqxoBY6BCTuFKPllpxsQA7kHfmbzW7Pg3O6Qm
mAdKFxUNuFcmuFFMH6TqwkI1Bopy/Amj57rInoYa/qhaqpM3YHmAXXwACRG7YOZT
M+hoBCIM/96qLEqKbtH+0NduWHpiFtHUNN8+ULrglVW+duNn4zdQC03JNAD/Tw7q
gAzA9CaUF7s8eDSomqUDuP4ddWvGZnLe2JLlXpYnqSADmRUPrwfBYcj3vtrSsiwm
xYOnWsYxpGP+/6JW7iZ+mXKeBZFZ1oQ6p28aCeyt6xU/XInI6zE4/HdFOPShBB5N
wZbB0zv0jfBZOzHFfLmjUCKAmVx95iLqhNnKE33jPA1HvPPIT1mHqW8mG45M61Vv
OTngGUEynD3Icjl027pRalD4//plCeTOKSxVqjhW0fV2VJ4LBJ5Qhi4ZuCCTucA2
zrzFIYNyVu8f7b9trT+HUHve7wv2dxYHI8NCdzyN6gd7xMD3mt83/qDBvayD6cCt
tdOJdV7wdZ6XhPwU38BLQmMhOQH2jeXTzeqqI3nDIQ3ox5j3qCaFpC+/OksccDNp
7KfgO7EdK2jaob0+BRGKJYdBAY3shzzloczC7kugCsYr7WlgqPVosQO+jxCHGsHS
BUidP3XC4Q72XDu7aJaw6WB7OMHrXPCOzY2Y91T4xQFWFHUyUeJZg7f1HaljPN09
dXiCi3yLbZCNN4K33lsFz8PheqgEU8IQ27+1oSKmUmv40FmiVXyXtqK9F0pgh/CG
DvzXz+rHdZMoLfShVuVOV9Ve+ITh9lJ6+6K53guP8urhuHR9av4ZupPKbJjes6ak
95m8UTrAxJQXivxuH2w9yNBX4X2ct/GhNqwd+qm8AiRn230HE3TgvB1lTVFMjjp1
KoRnx9177iRPpQODQlsbIjGP8L4tYGm0BHCP22qynSl0z1P8uKVXgRrXGZ+8sFq2
/+42WXTckW5OXoInyBVYJ+2BONCjvwdn2Uamw8UxkAj9cJjkeFUX7tBzYTFLctD5
8MjGVmKJ1KfxUBFbqINq1s+sORn/PDNHmE2PSKmz4UudB3XjwA0D8K/hk2GBPTSe
bDNIpjx4BDuzO00WlARHMBLXtxCjPko9OI4KvYThy0x27OLKGGiHSALSRji26MGR
wGz60tB1QBVf8a+eQ9EzQbpP4ppSNG/Pzr05FGG17gCZ7liDU0CshAx0tMszI0yz
dJ1LRz2Dv2HFODSSZQGnzobGP5BtibPi923UQYTIeeW9CUac7z83WwSyCti4a2+a
XKsUXYIj3vtKF45W1XpWk43xx+xC8Te0Yh474n9St6qpIZ0d3l4mxPLCoHnwnZpp
L7BONa+iifVZO1JMsgw5IQpiUmpnSmbxiiJofJ294xxGuUAUaUCMgr6CO59j8AEJ
Q9prOyPD+LBo5bA6CHh/ThwPqRe37Gl7KcyrrKfNO/zq2kVBMzp/lgLlzTKbsfey
Ic9E2U7U60vOeLiPP0ZAvHoNpRFYjKCiTY2rT3j32bksjP7HG7A7TNFl6N4XNU5r
xK+wrIFM3JajKSn/DDSeoa6bKPV+kyrg4VSpzuiv9r2YF1dU5DXLef+04Q/NX2Yu
cYWXLhOA8dOsOu9snjxOANkhODqwmdpeb55IUNF3UBPFB0e7mpViTwdUYGROf939
wBijcNJHZLHc6BqLBb+apJcVn7Wr6tG6wHapX1L3AK6pq0foFnR9U8HrHzXM1fr3
4128s4Q2MjdJaHJrljtcuNAU09K88XdneibAciML5cVmLBnh7MPZJg2uaw15AtTE
WlC2tpqJ5UI7gRKhloO3RIXKkez6K9n9YAAFVLId3ktI2I7S1wb+2VQUFvHHsBLr
cB0STkX30v4H1ZjWsdd4d2C7m5wkLMUCRtUGriulF8dqm3aQBvkhSW/wbhRJbZq7
Jbp78PCz/Gp7v8LTkbZO/fGwZTzTCe6SVsmoi4LNZ2y1FIgtWGV+KTBPGajEgl8j
n50DTlpxMbkhjV+x/dn+SquLQJe6TSlj7jtUXBv8mbjIPuNX2paYF6WCnM7c+IJ8
PPdyz2SX4Xnb46Vqh2wlld30puySs0NGBTVi2UgErvJ4Rcw3AVsBLeclIvdzN8DR
MqOp6C+h7lb6Hi8vbQUPcTo5kwbJ23RlTaSNA7tcJK4gEPb+wT0bgatX+n9TiAq5
wGylewLjhzCbFnZD/z7RnshfBfPRATd9KP9xR+7/YrGOcuI3u/NK29E1RcciQcNo
hdp2dR2ZdM6I8smeAbE0ScrTzme6hPcTvTYdW1vZQFZlATn2XLFFPQY5VUuMhetQ
nf/4yiBz26mzaCjrM2PFPB9ZT3xBLayz8zXgURWwv8OZJY54EdU7OYeiceqrVdZr
ng+oZFTrFP63j//910Fvd5VcX3k1wQlQ/SHvO55h3LjvqPgHZxv8relQgrH97Rh3
DZ2WGNKVgSgFaqHjwl9S/K1Vptrunx+2nPteWsC84gjNDnMEJ3sqyRYovsTmtJL9
QiCb2Cqkha7L2EUBSFCQb0sj+OFJr5GuxDgKN4IgjWWy5rIbfPT0LAC1+j6hVCJe
yi/nDJ/eDKZ7i8hpaCB+XkoRy4lIfWCgszOaS3aFnRdbhS4ChZzBCYKwzkEevbPc
Aqop8WLpWapuVWCFu4OOLhbMhd14v1x35eVIV62HlSq/xRhiYe2pTo+LJd0h3cZb
jUrhs1zsGz3K8EbcO2LDV/yR+a9YnJyfdn7OEFm+8FsjR4I1S6+Wro5bWx4hFBbQ
7pHHFm1GfzJb/AiiacUPk3r9tJ9DkmdOl2bi+iGlPMtkE15PIc24G7TfgVMyc3c5
Q5eHaxhnIowJbLQ+6B/Sz1RvfraS47aHyWyv/ol4NHzr9pLhtYgizvDJ6qJPW+Wm
w41Kx+2fFFmrOuMZbpWEP/cdMshAZk7rNj6CAVp8bEY3Z9Y9/+RzHNG7IkMevfyY
1flQv2HX1pNAyfYniRX0jTLa+F1IeJMDL4XgpvcMV3rMMgBaVZczGeecfWNKs63i
SZ25dZw2DtI8vrb8jZJxZbHhmSO2o3QYxyVj/e/9z1eCybvtNWW2rP0595RwPbyI
WpmjvFcckxE7uK7zwEFFbDS7es05gvFS4fVd9PYef3/qriyYlDANJ8YmtlEpnZsl
bdvLPrM3lGIQ3vUW4SoRT6elxPxB6nVnaH7roQc3r1cwdC/PfiZZR04e40g5+pdv
ifpqdPkzvifNDDwklqYJK6DcV0Ui5C6Ld4fvv83s6t8SDiTXr7qGlk5KRjBLQG/z
mLnZzqgWoy3raFMQIzhMmmEIZQo6sEwY3BHL1whOZHz1BJ47GZpOWg2fVnquVPm9
PUEFsQwNlDfK3HpYLy3IdDIlZASok3ug/hq831WIIbo0KwcI2WVOv+eWfmdsK/dV
SOH0vqL5C4UkgoQTaw3CLc1ma3Sqn3BDDtevgaJHpQhhHr5B6gL0vcdk6Q716VAF
e+GTiJImgFDY95pzGzwb4CM93k+uo0p1x8UuRJAYdRXC2DYNiMpcgwI8p2SUgcZ1
igg/Eajha9+6rsa2IwCD7TD1SBs2alaAynZAZcTmSFUe4WXtJqWsf9Bvh3eyjb6J
/MlZUiSwp2JOXwlrVFZ/T36O85XbTh7Kk8uen43IvkRCUEy/GaW8ofwk2mMwUVnD
8hpHJ8PKT+qTxVokVSl6/YavwfI8Z9r7z7ahbE5sbyaeOfxHnOf16OUnlimyZspV
J5tQ2iukDQ/ud+bNYG6ZIxynO8g2uLLzV4WKOspfMYCWTZruDbgZVtIBU4rr0FDL
mP3mRzCaq1E22JtGyoVlxrqRtmw+TK3+uPXhq8R8TxqrYWIzpXSAk03UV42vkMZb
PZQRa5r7x3WHMZHHvUlC/uus6ThgPeb2pRLGIu5gjekWqzOKrw2tmheI3K8S/GlB
UVhWRKoPlPGcnGhQOKTXXT6IxYzPc0zCOqbRdvApJ2ePsIsNcHpOD0nSSW0cP3m9
h1irgU3eP8CExPiSjb4vpR4WxkQhMoafqZ7v+KjNlEoQfdMiqs/v77hAp6RhjPMu
OvGo5uuzMOOd0jRq3jy5ci+MYUt/j4/AJOIRtHLdT/kwyDWYQRkYUUmG32Wp3D4g
DED/0ejKBbZQHYUzSenRXLJX1vFEqvp+3N8LRSsNNpmfM5OSU1LWWMkRC8Jy/3Sr
B4gcUacpaSvl8HEUz23KAEQxGkCAqKS3Vw/Vad2eLQXIgSkChWDI2+e8ntihGpK/
HlmgASDZYmB5klRjQp0RuRxuFFY8S/DjnefEVBxDt37MCr50Ln0J24eiT78bF69/
YhfRWhxjxb/mp1OxHczOe52rCpllgQ8gMn3LtLdSJ+yO9QoWdBKeJTjGPmA/cEO8
C00zHKIMpZS19w4uUyE10uUW8zuqRDW9fBAY0vtuWXpiUCxp19qMQJXmHNPeOoEk
7R69blb1T9qdw9pnMqvdHUA00GjhwVE13zdIZ26mz8flhTFjhyl5R9a2WcFGSMWd
HaxUNdRI17EIwsJqTsQav2RdeV1FV816baxdNjDEdgLZF3qGFcwwkQuOT9NQrg37
laE6JVvwEaMJ7kDlMLbN4BUD8r2DocChoLVV1PdqZXpdcNTCzJFbBKxH44qfDkOW
73HJpH6C0ADUu2z1RbU/z0iTbg1Bh2yorZeZAEL9argJ8hfA8TsZaFVCVyKnJfFU
0Tho0YxZNFAoQjGf+caTrzOJIvmvz/BJaeWZX98E1s2Ju2UzmZv+Z7dIivXzIGV1
8/fujh45Im4wn9XZedSRuNp37/BlLq2KySzUfGpPpCGBPHjwq0R6H8ZOqs7zc1Mz
AGIYmZMbl/HF1AnZT3MHTScqdmVx8CEQSisOV1y0LTwi5CLAMUhXiAnCj7+AOnh4
M3vc0z4d4WUqIGZWM7imbqau+MPKwFdd8Dn/5tYRiukV6an0JVq4Gp+uxekv6+VY
iiwug4EqRgROb4k3U6ARf4UQaojmZyAWlUa1JqW+fFtwux+chu1/iCqP8V1HMkXI
UbnSIp1R84uRfg3ZI8cwXxRYyUZvXMWE43TpyTorI6bllvxj/RpE3GrF69ugPkYg
DXjy6+ad28a/r1i6Uwayu0pSLoVyCeQCGVZv2h8VDXch6CKedBU7hcWhXp71Js3T
6sYwoFp36qaQGFUKOwvj0zICKWFFvTHQT+Gwj9onLc2gdR9yKjggd1qOrjsy3DJm
K0f4JGossGBmGnthV3hZlJoswLfPd4YDY0B80s95g/Z0vL+52isuTXJmgoLuhLCM
sRny2zhtbCtJXr3qX/9FonLmp+tFpXC6JqorQoXb6h+AoWGcUrxKekoDyimsXBQ+
Gz4PUlLlOhYXzrvkWHVei6z9ZXvxxyCLS8kL+HZ5SN0pzpn14Ve4Edb+gSIiiBnI
wIHepQkg0TY46VPO9QqtiOvBpVO5lOvEEB2Lf/2b19tis4pPCGR5ZE+/gqVa6psw
BXLoHoKcCyZHn2fZl1siEq5NN9YzBgSW3iY9qwOzTNvlXQfK9R0lzWlzacUvaeld
4j6BLdHsNGTu7cWCLn4KxZqfFDhaurGpSNEYPiK06tE1qvofxLGh0fgSlHOUqNOp
OMF/siAhen8zdm9Ttccje1AYczr/P0ZIMrFkILIJHELtei5vK93wsafleIxPnXSn
eHPh+/Ptew8XyR4zxlkZSBvm3Sb8bxLYk4i35dpqIYOEpXgcQt5sMtuDDnOF7UcK
m9ds6Bf6F9lYtxM4n4MmAm6y7cCIIjYoH3hPODQlyxkVf41abKd/kydxDzv3/9AQ
Gskk3V0s2EKySYTmQkhA6HmQ4+5JKgFUIjib5AC3fq7RddgyJZo8ADIRw0mh1ShD
dQqvirUSLn0ZdtaYqlYGlNRFPowpfhFf5/LDHifhN4mOdcRPAZ2NSbgPufYIrsTi
b+lD5KGRADwZoN6DzNvraFC1kbZjV0toF4nBz+scgLVTDHuRIlBe2qRFZxqGUhYO
OQ/UNu40MPOP+l2Lgza+WEBkAgdiJTNsNq16EY2EK2+nDjmFM6dq6Kqu9QSH6OfL
g+ymmiGL8domogEo0pvAmvY6fp1RkIk2vJGQ8Yh4KLPDd7AchL3Y1PMEIO7AF3uK
LtBlG7A1rAbADEBoGbuXoeV7iy7r4pi4sB+0gwH98dp6j3BppSx/OcM6HMyZUlZ4
EWPsv1BzqzZdeWILvQ7YpcrJ7jSqZ7Z4uF2I7myIjIFtk+qnxobgHaGIe8ITRBZi
WZA064k0TyF8pxE1IasgBMzZkdgY4NcuWMA6g79GTf5LZ3ABcmQO0EG67WDvja2f
6fgcC1di15j03PLOFHfeejkRI27kTUOCELRKCWsDvD9n7gK4sy9l5P5B8paI41BE
7VE2aKjx4pHfARulc/jnWDI7pZb5jA/n0yo173sbSAemmvbu1FwI+r5nnmPHzB7e
hYy/31SpB73oy/BTeLoXh+/LYZ56kvei+exOQnX6y1ox7D8QDTP/ee+rj0W0YfeK
OTk3ENJ8VYAh09qkZiFECNzWyjUwTWsk5F1xF5O8MLOQ3qOT3ARbCRM1SBeqKoG5
FdolOyUrd6tpNbmLEERv/3gkL8+s8Mr5uHCj6U4Q6mLvaA58yOp7GKfHalcPgsWh
UJ+VbqGwNHYzlueHiZWu4J2deJajyfiSdJjI5IAUT9huAW3nbELIhcap7Vxy6gHF
SASgOY3L52THQByePui4Pw/tJT2NxxSJ6ingjU/znlQN46e2nktkVsExVQHbQOwP
LsWR82AAE18DLYyDeE3aRdhuNFJilkIH5J496h/ZWpm9BTEFwXK7cEiduLI8l4zE
39wPqy+IMy0qJRIjIyr1vO5KKZ7ebGvBRFWnKkWizVZaWwr/I6LWb2ncSK8Rx2wP
GX2QP7H+AZJZypkHhFFQMNnPnMGqk2wTpBlMVhB8Q20i2yJT3RsbWjsexyQlPOjf
lcO56QS7Zdg8eq/CK1z8aMbhlOS4/DXKKiC7whCbUfBmByNJMLQGhhECrq6iwhza
H3fxgMHqGVYWJIzBmSVmJFDGFA/cEhvlg/LfUtZ/QrZsqLl+7J9adf95UcFQems6
TB7bH7cW5pTtehW4cYAt+UiSVu+JT6i7nyXDi8KPV2vJlTkKB/zLaVhRddVGSb9W
AtHUj8CfstwRlE8X1KpcKciyfq9036ARvc3mDS8/ugTmcZ/UvuOq3BUTXJ+10m9E
PDc5JScy9p3oJDFvXlLlXrcFS/LTkUMDk1nbAyTMrgkhoA+mvUsFi8vxEHOhukHn
lhgkywEYj6ctA1/QTMt8VPZ4sgsaXTY67G464N9xoI8KURrssbZVB7/Stdwcrabn
zXR46Uu1bOCcNUYGVAx9E1aN1W+tVeqzjZaVYQ+dg+X4aWlCPv9dX5FmA9Ewqix3
HeCB7ZZd6drAipoomu8sNKfSrTpYuSu98d3N7vjtI4tBvrEbDNBRZmgo3qLp/3X9
hsCZNTJerGfy1J/O7kM7r7fsvgJYxTPtyXMV3FrAmFtf9WSmwJ5ZEgww6AbjnvmY
XqcMTwV20pvR5H8FXcq2W590z3whQ3eH01NwtfKtjP51i446yaTNyicKDj1KO9yP
LZB2bw9m/iBuKEus0WcXhqda0DZOgCNwM3qKLU7cMmcNhW0mTpO2j28NSXa430F4
RaHQQ4bbelgXN1SeRygS0OPQbb9BpZW++zK6cHcJrxajAnpEuZAVkLuYh8BrNhIH
9pAxE5XGbSnELReFXUD1KHr+UxbL//lyYeWJlbXphxgkaf9p4LpsgpNsrJbGHDd/
Id6uK3fY+qw8UTZ089UHxBm7bOv3sUyRi9RKqa2Om2Q1+I8TAX3lr4X7QD5p3uFL
+nSfTeEwI2FtsQWB7GoGgMcNzwdOMeeZEyh5J+VJ4h80cNkUjB7MUh8KnIOfCaaK
mBKcm+KShqEejUl2I20qy7bm9FtS+BYn6DtyvZLO8bMyPaS7DFLPgmLg0W2fiVzI
K6HgJ9qRnwp4t2seC8IsGccfPLlbeEBh8jIJGgwZtOzKpka3JGaxTlBl3i/fnbb2
YY8kECXA3DTkbwdHApkaE2ov+GyEXtiwoUiwGSteDy0/dxx7BoZUf2nL+/fhMBrr
pVZTkRKBD+n5F44ZdGbA7DQ3w+VSYp6GeLM7y7ugXlJqeHMxeKVtP6TCoSrVFsh+
Jv2+0QyVwt4LnMgLU/FPBToZ1c0paCdLNgZJ3LH30WaT7/+7B6tHNQstHrQ1poVn
pYseBTgfjHXvNzwrDkwD9bFUSCkMu7vYHzviCVyIWrMpDuoBZ7pjJmOWIqhgdmJa
7/nS15GWpSWEwhOyjlUgosvObGLId5mWmrTwJkUkWxi4umvRRkgMrqoBNNFNi8ty
dpPNSXYiSfvz1pQK038hY9bFDzifsHQYxIfy2aPfyCThUenE3gx9nswaxFgEwjLe
ZLYqOwmRDclFdV+HxyQZ3uxNsIRS5vWSTzCouNaYn8WV6cYzGxj9NEZvIMSt4tFU
AxQMrr1exyJ4Z64h4kwSHZo5alE/Qekhv3iuhK6L+bhjalIpYQSJgfxYkgaY1Kg7
+yoFgOlytoBROf/bK9IQuUyG/loy4rdGkeRJLVPLxHtWm2G/AFEvUoVGod8IQBZ/
vkobkTtoDBTgO02FZO+WvRbMzGjcaTcBMgnLLA64LXYYFslkp0gyS0QATSJxWIJ3
36nicPQRmcglqDXhSJmE/iJs4tx14ae+EBsBD85TJlBOvD+y1d+QyIqkkr9Cfu3B
ptVFKzBh7+ccykEaq3euiN1laOlErXYRYAS2VYX7tGRCyZcEUDMHureo3f/GX/t6
ETACZaEXIgydy/dES454T+HX2Wz/kzV2hUIJrOJLvH/8T3LiLugF2flybVfWVi23
8K5XherU8D7cgcBZE05j+4n6rk9msB6WprT6u0L5Bx8iAYMjMTZm5KhwgEvU5rsT
7uqC6mBpIUt9fSZaeymyXfHtCcjrPFtvlQdfXUwlWvZC5PXcs8MJ/3D+6ElfS29a
sxmiD3X85N526AT5xxeQGSoR0fwGQz33oikyqrXTa5l268sBPEzZ1KC06pePRanN
W3ndAuV9GWYfHKPsh/vsvd7Y+rQ1ofSle5YGmFq6mbjV2Yepj7bGODdLTLbD5W3z
W/YH4MoikLGqRhKZaCOoFz6lRJjnwiPOn5fvB1Guavx+M1kdmCJHTVMJvGav9S3V
omYw1ZsLFpUPxNkSzvdMPrQj+Ip+kqEFEvMorgE7ynR5oq/TnBPCyy9hsYeze0/b
kJYnD+yb64fcbJp+WddZzg4v0o6e3Ejj9cR1gyFL0q6rrs+CPCtY4q1ap7A9bCRp
KX3DGtNao8gdtVqnRtQZZJYhDRJyOIRmfpnB3/hoTL0zsIYYFXa64l0ZoyPKTBPC
S8H0XN5r0q8gtqBimHtl8xpQ5wrlaVR8kyHeZVeW8UqCNLXvtkcII8OwKBVjXbsm
IxilyyVQzUaF2PWPb+6t/aGt4ixPzPRC/qadbs5d9xDR4y3Fj17/zo/FeXNa/sbA
O7hi0o4VqTd6GjeRFs4XXOUZg4KJOt1fEfzXtsPhrFZPtaAf1/uNvgn3zeJS6TZg
k+UUPeR2jNZt7u1aBl26X7MPoJk7pme3LUf11cRAAxjzh7/+R+dikQ7pw8v7PqE1
6a/aTZaAPF9fCyhNvgyrJxaKZ1LmxWjAxMyc7bSmcTHBgNiTe22M9JF+1Gf7x6gN
Saih+Vpevsqr7UyXfNKuBo29xYOP+HWiGmvy7dmuqpTgWVfF5GT57sGzzfBNw1JZ
ZJWqtVT64BTqsZx05aL4v2sEtNYjxLQ3BeRu2+Pv2itzZmvspgerUHihig09beLG
pqzJuntmtACVWPzqjwg/qncbG6BH6UwgXA6MBk9u2wZAX33qdO8ym7q+43VgDunv
mUeStdazPEWuwS8I1AOOpYeGBlvoZt5VYT1sCnddmN+blN4hVX+hKuOAjzw5S2UE
cNM04wgrdRDdP5Ym3aUdApF4L+iFITLWb2QabxOl6S0bpCoiZUWFCf9DBrG/4wrF
fZr4FfYnAU1Ov/BROj3sWbTqh8P0InOhorp4jzkXUJw1PvzR/xlbruXNlrnXKe3m
No693wPnxPGrFhImBwqfruqAXXIl9fQmgQaac++k6mAYlARNVZSCTclHoTLd+Wzk
BEFU6xO+/a646cxDCVnb1vbvXh561b+g6WMnRrt1lQRNlin+rbUdqlT9aN1ClXCx
8mDyTy68hMYIHbkLN8rS2lT0LNrigD3006yWsotwBlxavhFbjTaS0hzU/d8mhSiZ
09WNCWkzSkmCosSvZwpF2n2RAoFZGye6yeNM58bB/quiZJeAIU4fCB94SxAfLi16
GCXiFE5qkzUCsY4OmORJjssrupPIBym3FT8etcOMj2oaESaoNp7bZWDicvIG+Wk1
jK45tLWUbxHs+XCY9f6Yh7VTKrwwSZ25XKVagveEEXy22OGO6Kbr5ZfkcgSStno6
i9jIXv37OT9sdm+KXg1rGlGPsg8jg/ziCl8LGlvwORqHfxvfSFb2GR6AuL0ZsqVq
RcVXvUqCTyugepxmtKHczTzae2Iv2ZLNGjvkstMm4cY6EqizBVkMKGvdY8rtoRrc
4pRfgjQRLg3bEg1Qo7MALYZncWdb/tU8KHxVSbNvJRJUmXAv19wImboBQMxVkrlk
8g4R1C9X6I0tvt2ur3uqSMBNwp+OlOL49rWcCwXg6GRHEzBsFhWUT73ZKvKe0YZi
9oiDFH/b9fHaSym5IBu9uiYl2X0yZBBqrKXf1KFMhWkS7OoH1oafZo/hwPAO5OPT
oDq8ICKSCEpPvc5RCu1hXe/pXYiSFxvIgWQLb6cZpumgS4hJ6S1Gs2H3wQXJkOW6
misth5idXNh4ah5lyiEn7mP0uqjno2HzxWYkfrHyqJzbWxMDiOSMFmleR2Udohwi
yNKPL3VPsriLrAOxHEfMjzrGYx06ytrJ6ROVWWaMz4CNVBWtMF34BA4ETcVZXgC5
Ea3ZUVsCSoNYaEs0iNkVOmhGtzzT1MbO+78pIp31JZMEYHU8zz2TNcFIunIac+0Z
LgDfIleQjkqrEGiIPYQSSVV5CU9hBIWSyddA9K1RqS4FsNRgkcJPlHclAhdyBLb8
TmpEz3BLtdOuYUnzYLEAWD44RXD/dqxTArnl8+7YkB6kO0vMeEc4p5WzG45VZRA6
bgloCIIgUZMVA7h24A1skZJZMjQAxxI0+qKL0h6iQO/Wrj1DsN9Hk1tvMEYhaNIf
S67nut2nu5lJV7hP4WaWIz7SvXtzULSMHLMdXz82yahLcB6gIdQABBj2iIMSehw4
YV0Rnf4YH/xJKV/TZDhUJ00f4n1bI39iyGFmdRU2bcyj0SMJBRQaSRIouXG2TdcU
+ZwyNuNDIeEwYCVzoJQO8HXp/UTPNczcntjXucdH0hzTB0E7KdFSgTCvGIv1PwXJ
YkBHmEuzOy7mE54XNblQ+bIFMy7kH34K21/CQLZg0KZ/uso16nZozA6KwrPHhdMi
3nY/pLEIXDAdmAcere0/XZHCBCtopHtCZ4t7T2DHv1QQjgrkAqB7jZ2jcJJnzqtQ
nZqsHxmK7yN7YUq8zQskb2QLlPHaJzr4Hddb2lTz64A0mSMkHSifQCDkfh+hFe4o
xxM1vxDYFm1wyy5p9G039YjqCMgi/iscXuDwoNwwEsq9KlIjoAFmTndM9YQRI9fh
I07B6aZPDDHEpwoFT1NaHsqYmzJ1x0q36fND85Uh/Myum+q2P6ObxBFNquyJxR/E
UpPifzLA81Rcrj+iduR1SLyRmRmK5Hp/HJ+5ONBjp1wCOiefrhbPELYgDAwLjLtf
tId6XWPrCfBemBUCnP73xix3Ax83Z8hAy9Gl+AcIRkOundzzK6JtX/UtH/n+VM0k
Yvyhvp/KxKW7fLxDXkhojRm0MFzg4h0d8XqUAxkyRu+nua/qMFoWGv3A2L2PRYsK
nKylNdTMSpyk3iI4OLh9Ce5/Dd3J9kOQK2BVpq7q07M6XnwW71iyhpTINGfVG3wL
yMj/6t5KALE18As4NUZh/k5jf12Pr4iXRHEbnr2BetXBs8HGgV/gVyNmsCEG6E5E
o0sk4csjnBlzoAqvlP4vSPq41dZE0BWKUrwx6ugxHxwo+MEKECD9tmmxQAp8jTQ6
fwLVSXe9vjpYLtYFkpCxCLMjUI5/8R1EzoZJDV3V1xhKkaJtAnt7LBSSrklkfbph
r23GrWPvwt7ObNM2IwFoJ488Csd/a8cCWYuXNbHOrRqFwy59e0ZflBZJPIgwXtsr
UzBW9ixFrsmeGt1AiFLVnb05tlY0wd8MmrhyduA+nn149IzWr1EZzPOO/MzCmJTk
306v1NrraB3WEcidWBIcgnTDJaRiURBXk3Hin0x4peO4T33vZxSOLW5CVNtLSCDk
xOpv/eiwUrUTHoXMZpb0oTN8f2iNG0eZMzVZr/3zAmG1gfb37j5VSj6AYicg+cN9
jBBBabRfGY6AbjFP7ww2JN8CiGWfIjZp0LCa9cmMml3XRkGOTBs48j4yw/mEaZNP
g0vhM8kqftYPTOFESCQmHBsLjaupk3N+Ei1GgiJvBuxcMl6vpts/ut112tjAH4VF
rWw4CTD0s6MmwGoCF2qhFQVfFgcR59uHKZcJzEl1HH941t1ME1NsIMYbHGm0a6L+
bNZAIDINrnLwGxq569trIG0ytLDv2JpBGWKO27UlaDg+8ZXMEq1SKA3CB51ICPVi
Y0Pdpwh+0pknS03OLuBoxeB0xfPJ3pEL9QR1BzcilUDBs0Sf4xqJnOjjlescJjcZ
BdgcS6eb8onL2zuvIh4m4toCHi2Ds0tpA2jN+0NfDsZU5NaGOeilL2p6ZWe9+qb9
PQb5ucTp9SrdtuPNiWriksItvIFIKX5pRNlK7AeH9rZeeGcoRKIk0qIISPQq3H7S
QUNFdnBUId1WeeheeM24KzbkBFVT18P3YlNNRyOtHdN7M/m38iw7SzT6wZbQ6tgV
zolewbya2/NMYamJvvt4FOjDHjVaxNw8uhKqsuyHCkK667vhcGyc1ObBavpuurFa
nUzTn+CuWbT73csHSfEBTVz8UFfwz7oLpX3JFmIAjzkkvpG7tsTkzu4wjyapUonE
ZjERyCbj8sGw7D6W53mOd0J9sQtfZIyswQWChm78wh8MvDkpbaNR5aNknDV4AO99
AN+ZfBavj//BDcYVYV8zHp/vxu5YKUeNY15pk2i60Lvu7R1SGOh1DxK0vhKesciI
xckY8SkQfVvURr6BImlhOnOjRfEc1evbJHBjZNTpRBlXpUQqwDFWBfiNH2mJIMIR
fmX3AEiylD36AUCZtBXDU66pk73V0171qYsrnTv6oIjJryhIy5NN8LE1AlBa+WW6
rcIsZ9TtSOINlL2KLIvmIkKDlnCmIEA7Qq6gQIuRdp0yNtpJn51KzCX9rzvrptSs
+bfeer87kHvGN8FTYZDv+00LY43ghj0KGXt36owa8nkNgA7I2Jr+5FglD3eyl+7+
dN7a6RSZa73UroSfVKbD2hvBEJczUseS2/XcpUsO31wMP5R4YffjTT7YahU0uF8F
mYUDUw7GDAHZ1CTpSMfYNG/tb0iWZzDwWj2bsh9jfvX6MvrjoiMvkIt2O/n2YR3v
KAhpQlzT+6LzBb+3a6di+1HUsX3UNDSEfSiIWXGvYad667nWmP/upA6r0Ayq8fON
tixtyuNhT09jetENN4iHu/qBp4lzZdf+1369rhBTay+pf0GKDH0dG8sQMrujF9fz
KX3feWdwpbRhbPbKyhQHT3PyUPK9hutabUNFiNwB9S+wobO0gc9CxON9q2XBv9mz
Yy9oM2qnOK6wdN5iAsJHsesSjNllwHBGclnPKKIyaO3CWNy5mare7D9FX/IJ817o
ERDBh95ro910sPo9oml9l4HSvQcyOUQiFnau+qNz+2bQPd037xfAf45kWjxu9d4k
zwmV6Ksa+P64e3NVb0y1pt983MYBs6UNIdPOr3BefaMW7ryZKoMVI7bXf8Efem8q
lQGGQaoPsoNJ59MHxRfXODRAZ667KTQwcaqXU1KAx26kJFCQEC8z5jFmlDYs3ZaU
vmnOctbLJVw8xErMMiMW27p66N3p0ARhccpPwgfEmABFidkGYxDRhQHbGKr+q8Ti
28J4hLd+OTj49yIfM6sEjig+/eVWdK5XXFdcEiL9EeVGml0BMI4EX6nSgZskK9FQ
beJaSyBMGF++/RBSozmmRyTJY29rmDGYP2re9dG4wKYB1qA33oAzqEYkZZCtGe6f
+NoaL9lpLmrdXKntmv9mI5Fd5etknL1ub2cBvHENYUmXWZEKmSSO4r4PVluIFBOI
MiwfUbKYIrTWfINb2fZEzDCcDih2XRAzD/ZMvUW4oBvHWacVv7G56MLN6piv8koX
ODwXmfOHvMqLkhyN838pIMlbYAKWsegndA/2CSRSDZjGJTXnQIL/KonSM4G7cKmN
ZCxwAk/2j9krwXV248TZS8+mQ42UVgmCfFph8VccsRIC/36Pz1fWtWaPmQadqusP
bj0Jore3I2rgcZI/tjDElxkRsj2DtVUbgw6ILeNM6RYvnhYs4gYXgFtaugFt+6Kc
rZq3Ar7S227W5rtNTt2pkK+r8qzrTgESH1jMN/1H4RB46FaR8hnlGjiHasU882A0
MQsDNvKGzP4IGn8iu3qPdGibEvKUZRMbR3nUbwZ9awlLRTzjdJJcT9gTErXYzy+P
B1+F+E/NkXfQt4tK2WPPQ2UHJ9mbJF25jTbyvif3LMU5Dh9hlHH9NaWFnTuDCw8n
sMEcfvnWQUw3/PD9kBUUbj2rDM6NB68FqPIGdRm2AABRhuHSdaDkEviFE0Nr3dOg
MnNUAfbGMh5O1zsh4OKa7VyYS1SmxGuUxm0Xx1GPinOOP6rOpfagFpZN73Tm00Oo
l59i7Be3/B/DgPhzGM4/AYwbfY1At7fNTEZ7dtTWbLnYV7e4iy9Kue71YMsacb0P
ebK2a2CAu9FIQlw8GFP71MHz81irr7AjdfKBlR3tsqhlK5uzLypLZzF2OzXEU6FW
wHopT24WC65jcTYzolG4voPno4BGw56t0pQuvzbPqH/uCpcgI03jRynWA0GicDJb
LObMQcdSoUS+3KtkCiz76zqOOb9YqDhrILa34KIwlRIYEktj7vcSP7jKmJhwCs6K
G4Pab5q2vFYpPPpNuPqP3r44Uq/Bv7OznXBK+SF8wVphjzBbiU5RpdY1L5D5Qfv1
MOJVHNeTWzbV6NUcqufNOvRtkG3VoOOLFBBP+cV+BXUTNdbwT07QqMnifdjvvMjl
u7VRhry2qrzvKM39kQgLJdxx4J+lXXEf74z5xorKq1vjOMfI4db2csLz+H0acJfI
5V24y7wtrb2z/JKKn27Byzz/3ic+epmR95w31ZqFTsWcz2+APFCvmGtA4nSVyrQj
Cn24FLrR0++JWY4XejqoEHpkyxJgiZOjsBr+T2zHDu2aaKdF5+wFgjYBG0Q/OIz+
1S1+dU7XswL+glDitvl0pCGr6BYWYkrkzo564aiDmjgPr55MLOGMzBw7mAgOWKXG
PS7o/fHuAuF5+Hw+YEE64LgFNQGkT+dP5DDtSf7EN14kHoNPQf29hYvcrij4D0nd
B4/dfqqx49Ad5uXa3m8E3/re8CDt0AzckcERXe42yD1U1jhwHhYSDyuNfdzNV3sD
IoTpgOA+iEmoViW+CgsEbK741WkRQR3F2FhdfnpI1coVRna0RedbwafsvxJOQZTV
SA4eragpLfyaZmSs4sHlPsLPgqGyICWXAIwTz2C5pHjZvjcBE2DIjnmZ5GEJLVwH
NnOJfP5H7okT7D5nh/y24beNGAAO/P/rVe1EA3PNmbRGX221M2llJWYy8q7JQ5Um
omWeu7fItzPkdX1phvD/bIkigJC7IS0NZwdP91Du9bLuVns3IYqkEJGIhPPTcE3j
dBEf/5zRPtCjGECAsIXzov9430zjfwZraasDpsqA5WAM3va8EZDDsdQ8Y+xocI1p
TnA68Rtv5ASfgAISvIWD8b2Br4EkdObg2o+CUQN3VV2/O1M0BPi3jM+vsTZGVq/x
dHLkB/c/HT4OtkXho6wwQfKAVoxjVg6EduYfx1czeWW3M6WuwGiTi/G4uwKEy4pu
amhRaxqr1HOmVWh7QxsFpRW2Rq60hP+I+pZrs5hxTB+emqqBf6spngDFw7r/trum
bKipWRG5sjqXpdx+pNfrO/WVa8pP7w2l9giFhwCvaA5l67awsujM2kutDiBczXcg
jxGZxCaQ3Mt1TDEu/qdT0BN+030PwXnPlYZNlY8g0HLXoY058JIErqIBZhLt1XSe
w/g4ayD5wZIsbV75neZ0iRgvhNFKkIt1KpFH7p/d8aByRYSl0enhSbpeo9i4GNnH
7PWVM5tyxGIyyOhovrbsIiKamjLkqN/yPCCI34kvpfKzovaI2Q3akrB39HFFDvB6
Ob/nD22E/4LA9yYQDBCdFB8iEJrf4N0I11z4mlzSt6jE2qmARpo1MAKD3nELHjvg
0Z5fL2Ll4z9h9W3Sc3+GuA2aA5AKedsCjyC5JaPAXErYjSVLlD97fN44W7Kcs6/O
vihSVm6JLoIjd+LzaPVHby+6y2MBYJo0iFUku/e9ArF6udEGJDpk4eHHIEh+U/5g
w1I1t5dpREcpUZ3ZsBn+P8b7BHSn1VjuJn+RlWx1BpyBLQOQ/J1yrnf5S0APt5Fk
p7gtOJtpJUqtfrq/b97ZsD4a0Zkem7W3ZKp4Zn2J0zoT0bWXt3liZdyhWhkJGZ99
4EVHs7Ii/eL7n5fmWKIt9aLh/ojJxFLcm5thTviPfaz4a9tCCXjdUD0b109KZXvP
gFOccSpIzqtOXE+yfeM6ppHJCHm5sItx/ltvMcTFzzmG77ln+oIdAKUtDBX4ZUxx
xf2RW6vKkfwRXyIZwx1VDqvW9Tyc2SJvZxvF0T/zleCiRNsKLrt1/EZTdKGWHc/J
l0S0shlqmyMij9qU9MnzmDEpFDtQPU2O+A3KqmW3QReoKEcWSwapeFrQQZgUSz3n
fT980K3EaMpdEHUuGJdCETOa64HLO3ATDmzCY0VfFYSXdyKOCK8qOrvIOKcBrIO0
Vu8665LteAg+DmqAVUF8iOvwAdj8jOmaN74W4X1lb/TySFz/b7rFWsWhjJBOdO3t
G2R0J7NQVLHlPi21yVVX4Eg2OD5VrkRThpkGXzsX70fiP3lu5xHFn5TPZ6mRy8BU
zXxkK6FdJpLfsWuyVMC8qzxIqG6W3v2/m/ba/F62h/sjKPWSszbqJvIlbhHAOmOs
DdD/tOtABgD8rE64qGWv16Xkw+kPWMyvbAG8t2AG6zxk1bLdPOgxRHrTBIbuG2GJ
b1G2MBZdYveo6LUKMdgLDdNltPGILnOe/hv7TqsMnmYxybQgtIdoLGkbhiaR/jjP
t0jZ3Noky0hA83DDN1jovC4nHSHx/65ydbc/4gOqkaE+Eg6XO2wbx/TMdS1MAyiB
+qXEXuYhW4r/Mx/4HNAfC8t5p+njFfRZBak42BKN8YcizMCi3VAWxn53ZyC//Puy
9UemDCPx9A1PyQtjOl021dQ9yzRyKXptaIHIBuI7iiAZ0CtItU/ZO4P7QhObQIrH
5carfD9TMb8ZRiB5YLTnHEOKY2gIvKYmTJSmCPeRD/91OrZWEVLJr71oJzkeXNoA
YnutB2nDheTV8cZuVD+TO+LHSXXBrJLc+lA3crc229yk07Fn+b6o1SeteVTabsk+
qoKGNXwfQyRtNM9pl9knqJYB8VfIBV0KXSxmpwXzd3u3Qzh1gxR14uMgZIdtdxJZ
Yuj7axNmfAZUSuY+72OSpj4DkZi2NRDC3u84QFO1IxCPPjbFf7lFfl83fsWl7gKv
1j9h2yFV5Wnfg67RF7FpyHlnPiHz/cPJu+yOhQU/dir7pyTzAesVpFW825zo9W7S
wGeE8rHEpdipvoeDVKPWMsKW3oGXqJCj2wQnyJJE92ayDK59Fu/8mhlUfAXI/u4F
bbHWqn4h7pDEGn3hRwLxowQEICx46B+vyeUDMdG1uewpmtQjZZ3joZHOdFVh2RNK
EnuBSudk50JswyLzVcsaw831VR6LUok1UjeH8cwQbZsdp+wsZ3cu+8TljlXcnwOW
TjiErlrdx5+yDRxHd+hHDyx+jmruE/zO3hEzxAzwkJeqP0lbEWizU5sV5sPfsbhJ
Cz5JVFvoJPLAHkIBFm5dMIky2Z48UrEFGJvVWAt5Ax7min9bL1/SyGqUqak5YHmC
nMXM4qL3zjYaV6+L7ulYF6nbEybPAtZFnZFROc3Q/t9WEzPWOHXLy75Eb2h3CcJ3
OoUFY/xyP6VlJ/oYE0fQ+5BmUDj5+4uUPn81ebelgSJ35Y0IqCdcNfn1zyy/vP/z
5uHu9ZMPJ+aPTCqBdUs79sQe1YKXiBYSJ/ncN7xpKc2tC5ubkg9iOslPnEcpE5Tq
cm0fo/1XzklwPS4OaGoxLYxQ2IWsmQrDgHyhWtpcJr/IXgiUMzyjgjpTSoepo4ix
to7dBXx3KAfA9odODGmTXoTSlkerZW9onz4yN/dw2YdjBEUPR90ZM6Ns+Ajb6Dxk
xKK4tGXqxLfaL9RZhrt9ru3u9Eo7UbkRlNOHr1CgAg7ooJczZs9F6as1+tav9uze
ovaphLVC/j5AvLUqFaJ11RV5FisP7Tgh+GQtWfTbAUgK6dODDGIlecV8hU8n1XLB
D5DhoEQGi8YTwQqnrqOzpnw4YhJQVWV/uoE2njLaqWSIW4TQfBheJnQNorePavzn
Pe8aw7UI0mf+NPZtK8P3+pBwRq00qADZAaBg1hm0sA/LRLJpOCsi14oVHWezHrI3
uYcTCOkHdY2mZIK9Mz8HR4tYmlC6qsGiFZE79Qn0dST5SgNxd0a1f4D8YkXVslDk
7gcT4tCpv6FfMBhkH4OV4iFUjo/0S6GOBlRNSqRdbt+yVfO832eLgCUWwyGwAiig
eMCzFMmKVc3B3SV0EckcY5SNgyG80wuElCk0br2wUeu/F9oAevJwoJtjZqkQW6nA
d4qL2tzWbtkumEFcVRQJAxWkJ6F8Uqb/NK8Ih5+IMXlUS1MjZxXKRrxexOgAN77s
RqI0x/6XSoR4Fsmwnb97o5U8M57gb5cN1NKDvqyQH3pMDxgYYqys2fnyaYFCJsWa
b8MFcISKlCa/EN9C46Ir6NLAMgT9RQlV3ICmyLIvCvREhtnhXNPXVBEEUHHUEgiw
l4OYD4QPpdLIPWWq7JiyXMeu0ooO17XdkwLngYAl5So+W6mdnXADPvpkodGs5bav
tf+0DED26GixB61kiTgbv2tw0sHOsrqBdOe4uGMmfKgV5zUUpKjDoQKhjxR9JRia
xONBZQtQAbz8eR5RC7VyWLp2ydP5lNRnk0okTMufepinPnxXGQk9emO8UluCHW/K
vT2DqvpEEfiE03iDqjG3d1SH/oJv3KR9xR47U3coSbW78BVO9wfv7nn++72NVeVN
YiTONNBziE1TdVaEvnQoVyde3bu7cEGR/nX0F8yARo26VRj34zznvAbQO141Z064
zaXAnBSCHWDimL3PFNFIJeJjNViBpavVjX0vLgUbzPj3YcxekEYVawAQNx1cVxDV
jMB90TQs4R3RanWZar8FNQRe0nM+X8L2uHvOIIFpYS4giDMvOs37Xd46yeSJ7AU0
JJTWPUvliQvvydrnHffZpQ8yznvjUA8KGvlIE7lwVJ9V9DdN/b5JfqA1SQKGS1MY
0okXNQ9QsKHQlmQkRpS8OdiYMsKv2QyswQVe0u5Q6QXNO3V8BKJhuSG4sObMh/In
OZylNNo5Xj4ko0qwPW1IYvLFmHmCwcyGv7tB81b482iQb+xB1K1lzfvJaH5FB+Go
29Effjs4DtOozFJsSn+wCYhoJ2OeNs37PWqfy09JUYVeeLsAsleYA9gTgRFveAHW
sqJVwBjd6P/BOWj9AMq5VJ7fsqzRdL7TXc3VVxTarBfUQEwqyLUX9aXWw3vlOdU4
3F9bQ6zHzxkZcs332BNRQ/77IGPtHVVYptOZ6JG+2/RcTesVtFtrX0SHzthmP8EQ
9EOcgQlIFD+JbcK+PcEpSrQx46Nve6Ylz8mT1FCl8zxKgG2irZMDkpIdB/p+yqBz
qTjhhfg+ilYHfFll9sxqn6FUy8d59rZuSP+i4esfyjmLH7mk62c5SqiJueMhgNbP
+EzLotBzZJlB9hcGQOJa6QlkETgzEQoRczwnDZ90tpjprPQtY2LWavOLUAR7ajS4
FUpfaJgT9P2VbpupWo5QFIDmChdaPqbQo1QqOP3kzJfqrHOSJ/za405UijFbbisV
RsdoXrrkHbaGPRBm77nZQMYf+7jPqvr6xINyeHeryaeQk8uStrhJxYxO5Ba5Bq5K
AhrWTBLVCE2MslX+31YEGxCW2l4lupBDVe9rPgmm29UvYLIHVhd3Bjs617jYfT//
pf08tuQLji5SB/kQaJC5noacqKBm7fXfqcu6isSqdth7XDWYx54hRnRv6UGkS0d2
c0Hfbtuhg0E40f2W3MtANlGBCS5yxMIRHKwJn/9IJJJ/+odphbUUQDppo7Fo1dva
MdX1SHWp1BjBbmxp2cBF6yteaUXTvgy2mBM30C5j06tWCVhV69YawLdpZYiZ7IZf
NAQZ26sYN9xEyWCRYL/bCJVpF5A7bZxY2EVOLaxmmXT4qo+tgXnmFNKOiek2QIsJ
kuef727j9dUhxReUZ++Owigwujiq1wE7v1v4fh7OS7rfyFOIhuyzm1tCrglSWF+q
4rl1znztqMqWlw3rUjBkX+SpyyDUoP6PX51RLfZ8Zt1ehhgDThjFRm1+CM7f/bZR
sqzI4H/UCPcx9YNccQJg9cbhNKXWdL6yOTbRFcxAj/NJFswQNANVHJ1F1nxubU6y
JEdROvNl9vgkoHWz5zal9jrtW2HxdAXOZEnVmHgVwCGEaVtasP/9NCIvJ6y5vlKG
aGfgwOA7oNf60hfIstAFxE+7BlZ51zKmqAoHKd12bPh5QOgWB7akSYBrGKoVM4z6
9bxJWkGwCj/OODY7yo2s0Z+fHWkjkFTk/u+Q9aE1QNu6GRAJQoJgV6mcVnRHNojV
lrTADAORXlgvXof5tk13ZMMXl51D75ZDgStZdMuvjGHdh3mhOlcecktJSF6dv1lh
OjqaFPwJjQ0VxtmGfBiUr9pYlhii4qjkPfh8jS5KO2S41pOIWB/CzjYOmuP/XMkN
oWqj8SG2g5Ftb4qVHxnccxkigH5FQ2yeztySIPQC3WjwzGqHzCl1kItLFSOIvgp8
pXLl4XEyo4THsVo7Gdm2HlgFCId8tBIl/WIhj94da0WiU6NFsK76jV65Ni4Wnos1
Rj5dTCDIdV2nlRJqCrD7E6T9nWYh2TWDfSUXCiqK6hFdQyWHyaVBq4Ew5XinuiwT
HC0U+DAYm/ttcYl1zkf0xysu3Ote9fmoS60UiWAYQWGeqXEmOUuaVNEQy0vH3CvD
mvamFkfBH3JSLr1JHk9f1FAnLSbT5rRYOABTTZUP2JhwQsmEIX9p+C5qI2E9wW//
1oaQ+y1REGoKQ0zS9VM2BLqCgbLPUFfODAJ8MPPD8O1JUbZ/F9bkbixG31bOcDPK
xCjYh+hbGjrgTqkXAn49eeSftzoyCxNEecoYMd5Gk1kXtZR1EkP4uiIuDZsQsf/R
PeBhYIqBvvvs1GFNFw8aSxRiwY2WG+g8zbZwq/Q1ldvEvbvMCmxIHOFlBNbZrCfF
PBc9PT3aXPSCULvCgFc/Jxx0ZaXaZLEJqo8gVY9JygJ5bHpPJuyY8QNTLYJBvjBA
gNyvzrOQkSweqj9AoYbfJbv+pAp6lt8JkrLNFtz949rX6cQK389fNtI0x2XpqGqr
vdWEDdeRgoinkPZP9HHmNpic5bl4PQXDieHqTtmBXP8yqQv0SE4RUX58JR8FTAJF
tI3PVT/zjkqBT5m43t9CSha8+vY8fJemedIGS+dCF3NAcGMRsfEKFyHlFGBm63RB
JdhjVv3bLCDtSHSarzsTW8R/HrdWA/DIRzQCHKa7mExR22e2+xISMSA4kgJzHOWO
1bVD9LKTSiAMJ3djI58JIl/7nGs42lDFIuHQe6tRKP6fElzpHYz5xcjx9bEhM4g5
WQMjBaIEkHAIrQbeEfhoKCt9KTCZr5arr6+NuMzl1Zc0q/zdSCZ4mg0XoHwi1Gxv
9pXMbjSoXvn9M6KRkSlXuGmejG48CzmQR+I345X+7K8f7v5Gnfort6ClEHFHpWTl
7YRFrpghbyIl6JictICpwGcIsgljJ4tDSeaVcxmGS4P14aNtmF5pdp5IYeQMOHGz
5Unq8HI4HKZGsEigJCSlzkhHDm1Mz4oy2CJJaQi1FYfrPbQahEa5AUxsbntd+9S9
EfjTlLZCgrSyPZWwN3Du8VPtU2tv0OcPSP0KgoKWeHWvhAVPWaXwOdopVmjx7jzX
utW5BLnD8Ipm68vAnBtPemYli3q5FD9xSf0RKeO9t5d8gPqtfRbHd5j5Q6/6XF6X
0/DSl7GKlariqKS4i02FPf+aVUUt6MrGP+nH+pQDcHR+mvlljuZtHbhqwIRQPsgl
+vzoS8R3xb/AwvxSoVhoW0FSuR0+B2bsP/Nbdf0jO9aA4WAYYcqmbj8zWzwcCmQk
wJS7Y0CoSkEVKCLWuJ/JVMUhGza2M3DyU+sW3h9bSxxywO24gmlCp0+KvOMSKdtW
OMjRx+Zkm2A16Wx+u1MwC5dQ6FB7nibFnl/HSGR6gao5qXW6zcECxItLctSzMOYs
IodFE98NPC4xx5S7NVwpu2R8qKHb9V5CzMa0f5nCXtZub7//p9wQXgdKhYNgTyXO
xeRZmmDq9ju0sD1f6mFIf470BW3X4fxjh+AwXwFYm7SAt70eESQJGglGVZLfuIJq
jPu62wQbB6HZf6W2dp2Z4jL6NuCi8oi1I4i1VWiQA3EkZChHwdj9m/c7MMJtkiKO
WCBPL2vixgRKk0IS5slF/gzsWCn10VhmVcetDjWmJz6vNwM+e8X4hpXtD1nP1NI8
a7IxSmqYx39TY5TrDPlYuRQMBjbS5b0ZRTO2r9+GxsIRVdVjnlOHf2Y6i+JSUAkP
3hTtAM6bQFMhgdrBRZzSP0lsM9m1Yt4YpBBU+s/uKyzqy1p3tBEDrP0uL1JV63ag
Ii72jrKvrLYO2oBc2LEfz3rPTXW89sQ/DmkHHgR9xGHOzHU+qXG7z2HaZEHlvdz4
D7mWBOghgY6mQuHnfSvuhhKZK0m0bdTq+Fi7SXkZWG/PD//yM2LQCkMwPEuNaPU9
nsskAXmBWcizUGy3ZDcaVVnkR6JILrzgZiuc9/dG4zvWrTdXdr79qDcysiuQeWME
RzxICDNFWk8fgoO3AwtrhRa5WJnx8s/r/dxnG/YxBq/vqRamEmdPnjBbuMUJOGhZ
Q0/MSSlQQHJ1pt4Gpe0+eBasouapZJ+TrovkhlnRW4zgfwEc3nC5LxFk2jZDQo4g
yxYokHfWrH3/dzVm5qHVcFOv+Tl6YWEgqkx567KfNoK7OkI+hw1YeAWP5XFzeF/F
/5jjj7ijEnq60x9Z4VMXyTgEnCrreN5MNuZM/WugBq5OXAKpHh9zKfluvJ9bnbwl
JcvyjnyTeUogzcvflbeQKZRjV81XQbe7sT/C5D55PeOJa1xbEljbS8omDyThkWiW
MCWEkajGK+r8YR31ViyO6QdBoioUYxJEevFF9A1T0HA++MV3eJcdIrzj2cD7jaFo
QJ6Lv7KosaDV/Hzm3X/iRJY8k9UUC6Leqr3r2wFFhyoxCU8et2pTEtZfi4aJz1x+
NNKpYfTxFnoTRSgacZwHDctxBmSTmdVZOv6Axpg0DLWjizAnsbDsHNCymat6Rp7i
E+mkte2yJrnRWGoKNOecYXpVbQhYvbBkr9WJN21pQZPSavkBN54HOnLJ58eYu9Wg
AELStaBOVHxZ/ulVJpCqhybwnCI1Pf7GK3FqcSta/jBWXiNhig9Ahpo512jtxybn
/nlXI+LNl+wkifwFlnMxMhXZYWpXQqOt2KZmTsPeh0QPa+tjaktL9I3dn85H8Rqi
dbUekzfyNzxnv/niR8owkWznriG6yltWPqFE1rKdFs84yl9aIJh1cYnomzD84Jf8
sFxGnb1Rp9oz6FOTfEIkSDTyuPzZbxbs/FsqXAFzsu6AB8iU+nCpIJHlocFlyOOR
6ABhHpn830wmRvRDOc7Gt9KZgwmm1uox2rBCAJ1ibu/MUGxbwQncZOizKMQsrwit
Y9iZiBfISRLUcGBknLVcka+GckTm2n2aHzae/aItMfG6QH0FDTyz9MA9N66qHZyb
M3ATSRRXTmvL8QNmPFnH+egGdj/dnaOtyZv1WiyfYKtCWkZpGk6saqLd56UfYgsi
+6BAH8oFscoi6yMyboRgs98MvpFm14gqSsUEHqPnt39Z08d2dqbN2LiJ8O7q9+P8
lx7jbgXAV00mzqn5mepFWDkS5IeOpuWn9msOB1h7D9l6dRZBKifcn187UyYS5uO9
4++nQkkwO4AsLva08VQmwRuOacVwsJQVXq+U8ksPvoF8KjpAlAgqCLH/jjegxL2L
fjgrHpsftLybQW1GXsQgbo+APcUpz16I3IgKOi8Js980CRHNnzHOxnywCNlPZGWr
Q8Q7d3rHCzF7jWC+WH+ic/zfsbaYHtvhcaZz3cLj0Suh0etrN4cqwnJYx1TWoDit
IL5qNHktywo4AYjGgvTgSLjLZKxCW6a6ajPKvd4pX0Jl2hjpGv0E1o8xEyqqXA55
YLJCgFHZTXGIWpoujbknB5LfCN0OggMQ98YSIA8l26f82NBZjPTvSWCtgXmpTStX
KjuuDTOPBZjHiceX6xMylbnGdfpSCqqhxgvEtETzojeIEivgMvNBMLGJKgn2cg2Y
1frMLENWf6iilZMzeWsQwZgtT+cZjjZlgJ13KFqcKoZp+hIcGLGsNcmDfXNAQ7Eg
VDCpApHVEjsvXCjzXcBsSLeXvtDhbV5nGwXPee/dmN/57jOE1ouZhcjefMJLAOJd
AIgOG3UnyO41n355tF7t8kwR5tIosw6UJILSzGYbikCdpvhSPvfD+ZC3Iey/zM/V
3PAvdHh2fuLEa45nRh+0ZXMpct4xYWE1kjWGM39vKEFATgP0UR6RYBLDMVyqpBXA
PePyANXhvnUFhZ/uZ/P/ZGMAx8tirWgS2XfR25YTcNHKRo0CEF2932dI+/CMQ14n
JCwpyJPysUo7QIFs07a3KHVN15T0urzg6hEW4beL0d9yylml8Ynjfkv8cedJv9qt
FlWC/yVfRES0YxpAc1EIezc7Ke/PhbwPdmj1XYKClOvbNZqVVqAsCUi2esl7+Md5
hSX7Cq6AMbwe9oY2DbzsVYWcwRmhd/TpUUTuJoTSmJFzG+XENJIJBg2nhJrlm44D
S5JhpQdEZiVQyQtQCoFFBQunh0rCw/vjfKecHlmGeK03l98FKDXcMokxccnFeUTd
2M7Fc//B/CmHmWsUj5jIeEabqb13u0QDIEdJ+A0sXEx7D39Bz0xOBKoHhNX6U3Bh
/4dei1DDDIG5jmIPtut6xtgYkLQ7t9QpDgzyws9ysCRVomy7rW8hUPJBVeKk+cNc
fVWeouxyyNXODHY3VUZpQ2FSey8t8o6E2OQonXjDKssE9rCIuQXHvoP7WQid8Pnp
73yUgGml0Clow3bJ09gSPTviMtAvZRvxV5PRsti5+TYMhsZCq4SToRHiaTpWCeHe
YwkROTicllwQRerwSK5yBvyLkFdE1ugewKwBwzlGbj7eAQUnpsxhKz6ucNhT0Bm/
9A1nIjiiE4qWvEPUxyuBDaeb3tBGYQ9ntnYc/j7Di6V4xHkFlCs6/vQVvDFuYUoR
0MoUPTXL+PpPr+GITmtJaPyeRUp9ESnL7zuT5/94fpAAxifMIL9aXE2ROY/pzEoP
f6YUgHJcQvKwfGORx7qz81wRHgk6gDbillqdR97iOa8zy/SOVwgEF4IktVn1Q9Mq
VeftfT9zbDO5ayUx9W0VJ0R+PsRka3qnjsSq2zB4qobIQLWI4T5s+j00G42sCDE7
xD/S7HuO7XpR2PCiRg7rBAeJUea8PeqwSeq4XrQ/Wpop4O+xIxXxc9v3pVxQiW+h
HZgS1leYussASZBmWuWg4X4861PUHLHG965lF0bN+MzQjxQDCzZZUyXgPFQ2MN1Z
RimmeCbVUj6RySdNFPxwRws0DJU6ffnNJTx12DZsrk154eipNRJywB9gHQWF6FoS
UfyryFmFgGP6NFcUMNHAF9NlnXrzP3P70pLh3gIYKLh6cbx3yajuSwJp+xvU0QI3
yAlI065GUT/RdrHSL8w/9JCzF8MMSgZcbTMIvxZsUE4EkbuP/QU+xxrh1x3U3sIh
VyGT6yjvHoqiK3TF5EJHQpodg3G0Yqg5C10yn4n0tsId0yxiqvj/pjrPryAXxS5l
OSZ70/q+xO3Af3cVNeUlWtSxg7PCLzccqsnTFFzKdGWvrQL7tIhX4qpnFMc63AzD
Qptwyh3oLlFnYbzce1SyERa1HIlvLdMEOmrXRlqyzWQDm5ztMaBPEN1RjCvFCtjT
/m7e61ERwMEc+45p/eTmvLYLS2G0cyArUZJCWx3WrWlYbv1GYrM/yD0F3yMMESac
w5PtFQJ6MG+GSM+LLIwl8/ihwhl4EcDCNEXL3PoN5tQM3m26MbntfHf+S/CTTapv
0JNkslypWaLKIMANMDYRi/L+pXvKdeMSMqttbFS73GMMDFD7R7W5rPIoGI4K42yi
rKPhrS+BZxjYq8lodVCpsu7Csem2gmJEzoLIV/5UcY8g+AbMCJi+Wa2TAXaviAoZ
ZPakR7B+snZ1TvIAkCnRZtlSbbSA2ZajIiAwLIiotREVbvrcCdqzHRmIHcYaGNwN
8BDiO9/sae2+8zZ1lDvEakW3Opp2e23atBEGvM5W8qq1ZAK/n7CenGm+vMt3Y1NN
UjxtFXo5DR6b4Jjs1FtxYgKe/n1sy+zJNanzn6hBcQj3tOy7TY5f+KtXLHWIGe/l
bIqsMbFck7Dn1gm+S9bR+AItt/kjKAi1p/l+JlNpsrxfcUIYGY23tsi4M647boMl
Zoa66PTmtODXXV77ywDRusFwu5Xt80PWEqqs8hS1PhZgVKsTdi8NnFko96u71poa
/7Feg6o2td7pK4KNUdVIcSaEMvnzmpc2EnZ5r47Q3zFbrp2nRMDgGBV78upJOL86
rjZTWttV1yC5GHRWemcg/pueHN7P+gjZWO5nJ8XsZ/l1I7K44WSrMCutLK2wfQjA
l8YrZxkQv1GwU6Koy7aTfcwu35Jh8F4OFh4bvYasvfg/n0GPyIf5q3gJFZN5FQ8t
8k/aq4xbj6zYTTR8prx5uaMCBJxuYzI5BDFhfq85OwChZoU56vOaycEDhjM7MzSK
y5duTCTRMtpf+VkMzfrCnXame1p+S155RiFdbdJjxcvo6KkYn0TwQjkcmf0AIrdq
5052kHx7c4S0LnFktb5HRX83Oz71u05Fb5UD5EwhxTLMxBazE8hXRIvp1cQ5UCm8
FkBVfnU9eHtcT9gtFFY+p/afmOfjTqZuj8QMtbhb2uNQXyev5gSk96aGQBjYKqHw
kvZ2SJA6MvASS6UrhK6MhOYjGSzywDRFpVQpL2qc/wMsDx93pJrfen8PZUZLCASl
uYE5TZSyUpUygZT3RjPmAF4K5ojVkoXEkmxD0olKQwOuNmc4z0HRWv+k1r0wqpfj
5pD0hCHGa5pimQmu88QSkrdR8VMvvxoTzywbM2OrR+JOljfBgj/tqWn2uzJk1Gak
G1SqbXug+Vo4iF8TfDkNC624CLpef+55uoOnMX5N4yzYV8YcRZ3xsOKwWEV3W2xv
9eaL9HRjydq6eB8+R3tkm3bXzXFt5HPDquDA7H6Z4EmTMTWE/2d0EA/xb9da3GWe
srSz5lef9x9t8oLF6NlxCRU6dShRuNp0G1F64y2uISY4r5pLTU9/uHeaNcdKZ7EQ
ycZxC3svB3PHnc7TLfjll3vuYCtnXZhlp3AM2IiGjuEn8m9f6SulxtZuvTGguHmo
4NLlZTZtSY1I2jMHPaMEXHF6ezgnT+zwr0Id041ll6EYt3NupjWrD+hDfp4NOlRP
q17b7BRBiW+0cyhd08UEyV5eDvpoVvfNjeD/aPQ6cUa2buQD9XfGn79GqqfPugzf
Gmx/5jlJIGN8G6TS9lGIM4NgPmkL4ddYP4/N7P0VvyfmY98TzyT6PJlBPgRfPczt
bt4WnHxMhAI9UbJOqF8vi2eveHkBYiFsLuEFbwYrxTtPzX6Maf9JqY8Cm60vG48l
JFEacLRjLwyNRzryRdXdHXi5cgDHOMejKk+YsEIaqib9aJFADYgT7P3pGBpPBNau
PMSz//reIgMsFiDarkt1OyKG5NLJuMTmirZg6ItlKZunlqZ0P+3ufcpi3cNCwwOO
G0/5swMdYTIAq59c4LDssPcjXWFNY1G3fun/GA58DzDOPuxIONPzT7oDLAta5UD3
u1q9herdYaFAJCJk9zq7xUm6sZoxK4aNV1QVX80SdsbI3PlLRkN9+w8nZZ37tRYD
wWPIhS7Wj8ZXlL85oQC/4SleLx6vrk4/LRThVcMDELXd125EuBwt4Q4jdnjRaG+Y
mnJeqPuAdo3e51ZgVSMx8uY6mjchwvmHXiR2pUcX3IdZD7OJro7U8qBGIWSPatV/
Vr1KpDncdVv+9cKUSeHjcrVnWSXt/Ixy7U6mqxQgq36DMeovwmSvqb3yLLNxRzlC
rN5emysew0/ykq7l4UIBNXg0rdquOITybvK7xg1i2LbiMlIRnzaTCiuQsFBvag3a
cSv6i5m03E5PYExmr+OGF3nmcxIG0nANMdvAEUFXz4fgBUjdvK54Uh24xIe0A6GP
Ri/1UHnbk/Tgmtz7BZgYWjhTBo8x/eYySf2ihXsi+rPS8CwTynLyeMoTInV82vG5
le34av+AYTwkxx1BboTH30mVuqp1mhLY63LmsBopIr49Vg/+AuRt1yj6EwwtUOuh
1TGncPDGze2m2U7Ti+TdkYzshz8D00k63rgUt9iQt0WkIAXaO3fFsQJycWMwFq8a
B9+KLUJRBJTO1XNzXH0Gfg2uV1w7zeUQp57aSK0ujd8hxt4WCCTsPQcl16omSLti
0VDy+c9FYec1ND3+jaKVvU8SrmBFjbf2Gvzl3zKWRav+Cca6KsfHnpGthAbZaSq/
G2Ay/6gtgmpYUbEEHt53waPyeN8kn0+OdtCuPE2roNQOUPT2MEF/iVC3FSD0HPST
Zdd7jKMk0bh/GS5w2Rk2cI0G8NoH1hQ2HdcJBPSMnf3WzRsNrnoB58tNRKNzs49/
ecx1VJAxFuGL2qz0CZcUBog5UtU9ESsBD4jFWNUDKiveHDY8VGu7nDEoEcN9AAVi
uEw8jaS9JGSx+MY1kd+ytq3zxjEYykY7TxlS5zkpS55WDmJCaA29jTqzn3pDyccQ
w9bfrwMvEtzjw8yltTQVLMZznbjfIULl+Fb7qYRbTaRG8NxslzC3M4B2mxueqLs7
1ClPAko0RxaHANskAxEGkes9JrfgkeuBJnSd+Y3AQv8NK2qkGBU4vUDmsyg1XBV2
B9y5G+iiyNp3vWDUsBI8orU/sE9S0hoTk9IzeI0856bj3ElLQOUxbbzuqP+yt9sC
M6PiXOSjR3iLe3/Llfjz06l1X4sF4nezBLS+Jciwt37b/u1GfgNuySJTGIjarftC
9IOkYOa6IiFfk7zBtRvpGGoCfgLchdQipr837vCntFY50ZkRO+MPA5inMTHkYmeh
V09f1Gca4kkYOVMCdSXJXGkFCpcboRDfPkg65hXuy2TsTEA3NmiKJIlrEM3A6O7B
mwRM5fYh7IlIEYioBYIMRUfvh2YLQZojPLIgX7nQnRAa6kTsBfLZ1/unUrYkHiai
5wsoXbN8481cS7/rynkwa5YRAMBBR2DBDR8kZx+j5eXbxn/o7yLgCjJ0mlaB6akd
jLwFIfGt7aTDGu3op/pJE6lmvnq4yacQ/j731yEe8/c5jI50Qtj9j4ML2i2rK0zs
DZta1QNGUBU751FK/c9hk9E4fgp/DIaTpsXTKEn9en5AJFRB456KWDJXwam3t0pI
uGnmq6DC3WN+w0cVtdQfMcCcr9/rGmEYon+GxKT3NdAem3iROJ9Tsez+Zn0hGHUy
udLP6nbxcNZEG+56pUv7es2tzYv+xLNNS1DLNSASLFO98CF88ZG/d6mwrw1I5fGY
g5RJ01kLkGTdJwg9OVRwKCtftOKzBrZ07PQoyRW+aAgYnhELMrtjZeB9EIoWApxr
cNBaCQPt2Mq1ZiHrs9+DRvkN+ssGCwLB3TSV6rnfN7A0aB0i9I23ybfOYntnYmDS
GIzil+cb8y/8wwVb/hlLdqUKkD2AV7B6Poql7tFqJMSicAlHRnd9t9jCqnlwqXVW
cCwqZUNa0oeQs10YCMGtuhRHsrck95ybo2BFtkwL5fVDswzs8cGP+EuFabmCyhxG
rYhUyX15hg8Rc3SqcudvA7ydhE0FRw1SPN1sdW/0egw+M0tkFpZonGvkGEv7f/Ou
fRKqNkK9o6qbaDQc1lU6t7lc2CFbO3MDSua9nq+Yk0j+mKc/LbaNQU2Yr8oZN4pF
ZKApYIgE+SFu3wlDfNh4ffLU7XKAeStUZ4CpKAIFaVC8W7iNtSrjzPN9KJns85Ma
djrcwxbdsO3+uFsm/W9fT5iSGWnurP82UTGKOR6pg2FFPJfjQcP7vF2PZrFRmYQW
EthF4qgbTq6nAFdmvfhV3B/vUT8Rz6+45OOYbXybINdU2atESZA1b3rax5/4hoAo
c+JR1PuvMMysG4bUNo07xkU1VT2DLZORGf808QuKuZJxHnTLJMyDgTg1v7aOsvgX
5vXWvkdR3moeQ3NdUkoc+1zrBSNo1AI4trAAO7DLP4xonNPupgeps4+tWB171tmZ
+nA1M2rwFWfTHAkCprKiW1Agsmf54iLgbfYT0lCZ4Lb4lDv029stBwmyeabghSnx
092N+8euwnYLewXx8DMukyat7mhEU3/8gkzx3OlMSmw7aQM2/93FBWc9ANSbTQb+
+AhA7u7nzfqdDvyNALoJICK02W5v9tviM/T+OCBPiA4S++e2MnR0TXN5ig3IjIUx
Hv6zlFwpsGHX85mwiyRamsJwEZHBCsf+g3YYN4bBmzmebPs8x6E1KmwzDW6v0/2s
wVZ7RVKeFr9WNWNzkwu3DQ0Ihe2PTuCNjXq59ZzIePlpc7Rtzvi2VY3PMgINEN+e
OV50PhRtJ5GQzkJdrPgmcp2XLEnogWy/maR4WaDDl5vx6MwW3HP60iYeoLju9UU6
GZ9goQLHdnuaQMuXcjJTGdmYJbUUcDpP4NAp10tX9/qhNlDyR/DsXHI/AZJ/feH4
KAfZ424esLuin1cjf8b5K+vXOVseVozT/RUFP2vldKd/z8SP1FMCefHS0i1me/Lh
gz1ELZWIx585UhvOzYto6//25TKsqLFu8/YogBV+G+6lHbiGrzyCRpCxJVAdZRul
jXaYd+Z8KpwtyiCvpCcVSHHaZXl1kLPUg59mqKP6LST7C/tNsheopEyXHQPR5ozd
4eaUcRP8rLCoCFZalSVWrrMqHbJ8THXl7lo1crlIo1Iwx7ILoUZfy0UeewZ16Pc6
xWeB4PuWe52/1YlrS08k2krsKIGWurG91xggupLOOCoB3VXy6m3O/DplC1uL+O79
RhDIgZ30Qcsise7fqtY4N8mOzkzuczPFqWXdraU4I5s7GT9B16C+281MxQYHmzSA
9yAy14Y4hcK8gge4SkJea3nY1KNBI+lX0vQ1eqHNtR5wnWbecdmZz3vDYT2C6R+d
gwqdC/Q30hraRDXhGZ5hQNHqpKRDBB9hnHQElz6rMegg1trNVACIos8zFq/RgGL4
/Da3V8EwoYo9E09dEoCxuq0XnhrMud8ovMtN2JRq5cyFNmnrmI3Fvqqiuo73Dgo9
dxDPNNdJTnziDzn0G/sX4jvL6NyPktmoCtbu7sMUVuVMdyoOFb4Ld9iMxVVDSKdo
y38vypcNeabkSsmP05CSytCppVnFeGrcEteUgv7DPIUl6zo7q8JjcIbQMTGLAsbX
7dWDfuGdXlprJLZLRRuJdC5cCeE4yqnYhtZXLGvuQ3cNZCM+8+CoUv2AW2qsSiaV
mRovDIR6CyAaG0bC04ym8l8uMUhC0nXiQAuzzVscuL2mV+0YhXjfdXc83DSO00RH
OPCQdrGTr0IYPC3URWLmfzjH64SLNtuea96Ki+SYMGMj2cpQdTnBVGPzlay8Zf5M
i85+XABZ7E98WON5I9Zzq7OqKMG68fA+vrMjQARqXwhCQW8UFRybS4HaEGDc2WbO
IuMvFCc4PY4XTvzPjTjoadpZeGGlDw5xhutSJqc/ooJ8CqqqVL4gsdo0OrKQa+1l
yMEnKKlGftRst5ztCFr3RFQDLyOllOhm65CS4IVknyEZ+fz5t9o1aSBWI7fO2c72
xdgzTntLdRP6MDZCVKk7yDgpJ/sOdH3C6wIojLFGMRqQrA1kwIeCudPgub7+EVFy
tvKQvHX9TsKCbdBVRiT/FtP4xJsCKUmG44qhh7dX9Rsu3bVCC32rqk5lJ1ACVzsn
H63xVjy3G3Aiz5xyeoFh/fBIpPxNmNBlBxQJH3XeM26gwx14X36QcNbiHdDP6v2B
g03XSmA1KLjme5Q1jigK1/5lAZWJ+WTiPfBvXn6lOTNdu6sWdYs7u9ew5dtXSh95
EwBqpAx2UYjwBuBtdArC7u5qOseGeN8AhiJnGtbn2hVcgyeRXbD5t3lTY/VfK7zH
lTtc4GIAX1sUmIdwORcuxS5sm1ckjWIbzcxk/omz5ss5jFfFsEVRvTIMdupWIbnS
0tRVVx2rK+F2iYZi8K27r40j9kZGsf1N8Is2FOHtClnYFWKMmjce8lRi+O+2eTA1
2wm6l2zm57ZFE78KFJQ2zadFMgl2UD2McMn+dxdU1w3rVZHYgbYELppRN9mhzYTm
k/cnHWHzQiW1JFqB5czOOeFHe2N98Ak3lFlRIOcXEbiARpDrp8q7VA4B+BaitRSk
damujbGsUp0GE21FXd3K+d8weBr61QWLJ66t5cLaZAzJ6S8vNmrPGlZNG4O4ptfm
6YRWyr9y8VkW1cxWp5W6J03ggjMEjh5XZUq39Jn582Cr7rtJ8NLONOS3Sbm9YWFF
Or0MIkEObgLfHI0HCuLFMJACOpa1Yopvj5KLdZuevvQOKcTFbgpbjyzjmcRYPlNB
hVQescJvq0x8FZV1y3UW4da3xNioueNVEODA4RQv1q4HIiuBNHGoTG8JbgJ+3dWv
maU9jXKYfDShZdzSWlq1bdQ45iqmzcO0BuAr/ufqJdDTzJXFUC1sL2rJC/oFQnoM
tzAs/PiUHjwD/+4u8VXMWf6eVCztZWY1NqcZvg8naaBPsUn7KWKHgma0DNv0h0OX
9t1VPW79jGgKyhybA3Uy6QuQPPOnWNTxUkiv9wRe6Vp5CyZR1UEZn9vDc3cXYiZy
3WWC9Wz+2X1yBftulUszCbA6uSnhWOtXXQ58+Vq1ZIwSaVEtsyyunRGsDGl1SM3j
6JNXYKTEeqQ3e4/AqcEyEszk9pW5D+I3mNVnrGcYbNArBWOIRiQEiTNSwF/HW8vh
v+hw1DyFYgkDIkLEA0ZpAn3KeT440+OmaYHAifaS0xv9EdXM5mF4EvWMOmCJK3p5
oss/i3hN62/ekfhh6oWwdQqeVbFNEXM1wuiki71lgfjoDLkXA4bSrIXSF21+9CQU
jU+c59j2S85CXoMTld7f/nfZFvqM1sMXjK5Tcg+r4sJ/4kCbL8+FvwwdBn/91MII
rj/qKhvy0lIp+0Q/BRC7kNS60U0O9IQTGEn2uHtuC2E95Jd0hlNkNM2CEkZmpstn
urbOZFWUL65Wo+X2g991oVLj0Mxnp0Da1J2ZJyMJUxAj2gUyt7l4RJIQNdm4zX7N
QYD3CkEXHGnOkRAh9sapklPn5+ZM1xt7fa3M7zovu6ykPbgyWsW0aJhl581A8mLp
Jm7v4Mh8gkUA84+3lM8zEfrcMayRzNl9ztACHjEpnXyC1OgGwM4yLWnHcNeDJNft
bCt5V2TG2CoVopibBJFtZcfZ5A37NxlnxKW09en7d/MbNRmyQ41qvZXALFyIbpF4
pXZNKZeSb3gRIbGxRAN4uELapjiCxjxob549GCZ0Dm1IJZCEbr+8l6352H11KkA/
PgUDOp5DpMVIPeukeGhErpn0WHWu6JUUNzA772Km0GraMWh9/dFfYlcb8LU/gxzH
lyRuPs6SvHIydzeZL9iVrrayg0TCZP4dxTEz+GeUmM6qMbiRWE8L7pOyzVCQ08qt
AJO+IWw1X35pjSvuGmx4AMC8R0rf8dSFIVaGOEVlh7NYDsf8teLUHo66L6iRfeyL
g0pK3fDFvUQDIqEC7NTkRmu+aIcQenWUm8E4eGm1nQ3ZMYgp8WpUS1kXar5eebvo
cg4i1Egn9lV13hQRy+LTyTSWdfHBdnlv7NWs55Fp/J3hYFDE93lmnRpIAFWdaf6T
i1XTy3SwipkuStsy0zHMAZhVEUk0SJQ/X7QIo2Ak9kxkI24pD/uUOb6WNAHRXJoW
73skHeF6gSaV65FmdyG/vie7yGuqwDmZ9T6DruXKIbG06fqITLWV9g9ZN1RAjKZz
Obcb+C0MLwrH6SaULJb8ksbIX+Lp1yBgag4e2wFF8WDpD6zhEux0l9qQic9965mc
32knCS1/jzid2sGRXeSCN33vPxPJTvhwj216aEJC3lkAiSlHc/ce5i4LSQiU82HR
Mol4adjvWd5RFVCSVqdY7QJ80CPc+40Mbfq3xog6ycdM6rYb8SX+9zh8gE8Kqgsw
eCLlqR6vt/Vtd+rKYhpCLvvsoiMKp28SrBhWwsEv5mQtcTkAEP3lL1zQ3PB4Gw8c
TlEpIIH7DfZsurhEFnn1+nrl20o8xgRYhpA8TakyGkKYCCbcHdBlE+pob6b4Vu1G
6wxwJee6lUqNsg+f2ZFBF/EWueLokQGaDlEScCbTJgqqD8TYs7QWlp22Z5IQ4Wh/
W0Z5AXThEG8R9IDzwD4smAHqHbXMxoDX++jawJKuENh+4W7huXz/2SG/QKWoKEuj
tEG9bkFhcZ+8StYONnlibo8nvZ/JN9/tCF/J/itWDgMNXEgaeVv82GpF62/25CVu
Kc0zZ9sHS62/4VEwMV/nndiTl6iuiePU/nH3Q3KwJ5QFlMw0TDzccu/pSuDeienf
iiu5cZuDSZ0H+Jj47sur5See4lrNoKE42UXSnX5p6r5zh/4ghWQcLlYvnFSnR03H
bo8BZFAcZCvno09k6RH24IJfQe80ozS7k3dEA56gwoErRl9UUlie6YpTcZvl95sU
dOBjfD0PxAyqZnAjm+XQuDlPm1XxAhNxngOiVnvSum9ozdw5v4tf1blgF48tMKaE
MOrDgKGz6SPWOfjp/SIN8kqewz/b0q0oHoUVkAl4aYSyI1MvKlXG6RFL/O73tjJg
bLzOdWUhPrudLPVstWuwdSe+T7EGGhkGEr4FtiYb3S09du5Nv89GW3/TCksjMfu+
4ASDyWKaCngaCI5ScZUwmWkGyR5YSVWvPz5swdTrXcdCofl6ctB621QRJ8pN7a7R
MLzBhGUVahoqvonD644coyQ9Tm4O7KBsQP5bpaIHku7pVzBdrhjHcQcPJPwhNUr5
6G1uX2WZaPH7bnCFkW4ke+jc/FNjx9NS93H8YrtO/HSk1h/ZNCZpqj/w3kCCiUmB
7KDg9iRLvmRInFPA2VO9MRsREVqtywY8AH1B6T1Ple0PMU4o9VvRm+pue+UF41mJ
jYTtgUxeLmq1ZOei8/g46K/GAcsT4kszDl+Vt4nf+cEGOsbt37MkTXMcGsL8r9Wv
u4Lk6CkRDR6/tmVkTUkvo+OBgQR85uPanoFLxi16YD3qTE2EHywp1y8Hxh1hejOA
sxXHqNnrk8BnTLTkjdk5hNz8bDXbA5QT33xsFhGglqN2k+nGyLZRr15TouqFeSdU
d7ZU7carwopFXtperKkJgu47YXBNvCBdS0cX1YagCgtlfkXnIb9VxJOVrGtjbuc9
6a6DC+8a5tyeODHG+ZW67cPrKPx9E+8QmBMAYhO44Ampn05ZmdLEAKbWHYa/WnlP
Vmokue5FWPh77CVog0xUN28rdcmAIGEinBp2LADrjMjnsxCHrEmVGUeqTK1x0Ng1
4OjIrOv7ZaJ84bQp0SwymPpU4b7/efMQIfEGl1/htrb+yZKzRyXg5Kyq7/3Cfhn9
I09Gfaly5oI0VefH5RFKhXACgLd6zQyvCNDCyNpPwwOy0zeKw4Wkir+3AmE9FdR6
ovgl6EZ3jlpTACJdGmQpAug9lJDMB5GLHVXr7JQM7uLCaBm546XyXN8bhjonCzlg
b12V0ykn1rsM/wf+pBwYLe1GAdSR+dQ/w1+r16mbD3MqhkhWNC7+BYBxmprrSV95
u/NjGjVYoUieEpoGzYFP18RPBTZMhTKQhCP80rQZOW20u+iryWeT5MgSLpv9zevv
AuoAgcH3DmOQNJL90uKok7f1T6M+cF+7nRMu6aa4YF/4XOE37NBd298A0V2TKD4g
iOdru4d7fyHyw70U8mnoTRguNnuikGgdxz9ptCrtGb3DKSFZvFMVF4g+TT+6o5hJ
HhBu3u/AGbjyF1eua+W3O2IwK9+rqRIIQrfGPUCSvcWeBFmHmQXGG4anbFL/cdFU
wxi/uFAycNMVoSLTMY99eqS2Kuk9e8elmV8xjL81GyVxW0uCId98IskIAWINX+wf
vXnwBFeM51SXbEJLzxLpmRIsmKwHHDdqC1TeGok8uqPqjxOe+yQImk1bfUfgR0wr
Qpra762nlRjweeAhEfSX7+O8YvD8GOZe/cTVt06MImap2qhmIkNc5SjQKor5yeUR
PxltG2jRPu0llBqv6+cZeYi8GpxLWuxiQ2OIkJ4eGAHTYos7Ei/qZe7LVpB9jZCY
pHtyxshQ5uS5ez6uAJEMgw/rS++DyvY9ysndoKbmK8EiTkdodPRVlQVu20FI78wv
e/1H+u77wYYyY9fSOFwP//OAuXsxWfZUuGordkv4IV5ozmQP+BzCWOoJR88C7Sym
rOmfOa2e73kfHc1R7XNlrvlz1yxiKCiexg/BmUignj/KnVQWqfwL6JPmogzzOPfM
u2Zs0dA+cz6rFdk4T0JaReWCo8HzghDC3NA5/HN7VbNVgpfrjxfl1uH4rpLUA+1k
R9iC04bLmCr1B8aZfwLgC4ZT6gcyp/wiv8nXL84MUHDf2+PFUnd3k9d0i6EW59eZ
1NvmrWUXWjsKcwZ/ogB03h9co0mf1XOxxpSnv86FUOYVKCXJdukH68W99y6zkQ+p
SH2jUDhd/3VuxztVQoWHnmc+kf5kBlg4M+YMIMIui5HT9cIx4fyQhQTWy1I7caNF
hpLBu52I0OBnm0t1oa8aJ5kYLR7eEWQ4e7jjZzN4GdtxfooKLtCtn2Q/kUfkpjGE
9ZNkyOzK+TEzCM3mIeB/5Rhl7iv5B6jvL3CfUb+EY0/kyMEQ7yFb+Qh7KBj9JquW
xpEFa52sHhoRY7pl6HVbBHErlhMHGTQAmndDcCVDdWA7ejbZJQM5FSf2IjcQ0rLV
hjB2GCymjwCGpNoqa5WLV5AeQlyU3uWQWgwmAKB+6g02LRFYGJSd0jj3xzgsN9SQ
WiB4vJLbeLgMpfKGw0Qc0dk2c9A7xfzWSQiFBcRNOlo9FQDheUfk69Gd9TihGhQp
VvILWogwwRFDcmuitZxkW5zijv5b/SSfaGS3F8NhmPZl8AjSrfhNuGH6vCfvI8Fy
0OwPmpaEO9v5lCw8Dsc0VQ7SWmkfLWSmgpYA2W1THxOsVUPJU5OMUflRhNWb7AN6
iFiWxbBdlmxH3DkY7oYgysfaqWzki1aarNX8tM2TeMz0hWK0F1Fjz04W0uRKMrIs
8/j/FiCo4pJspC5HskSjmhTHLQybpdtJ0jS5vtiFEoNr84KxHhWaAcMK+jDquk8s
1QjJkDWpIT5CrgP5w+OWWRWSwRvEanDucQ0s4YxX9pa6hAmaYq15YbbZ3DLSVcwT
8EMPC4NY3Y4+zQrJ+6pEbjHGHUSnFReiYZoJxU+BqdxuHksKLAaW7G0mSPGXbPWW
vWllGj2ZAP/5r3mencQwGN5FPj3SgtiOwgEh/0BYUJVXf672NmbnoEkHRW6ZWalU
97chbvcOMTgVb7CXrPj26X02uKsKEqtobaalC65I0RnIem4kbGdcxUIDGhVK2BxS
kFK5RSIsT8DrFYxSgLHdOVfX3XX4sPVK+m27y1r1Zd5DbFGAvEZwNevrf932DSjO
DXF0vejlYjrZ/naYRoH8R2wYoQttoHQ6B43SYcMLbiImaHrcR5aXPatEKaZC8DPk
HGDgnT3vlTc9FE4i3iWuGSUCzFRe9ky44iC95mbISeUB+bubW0QYwXOdJc0CoPxw
+5bNd4+fFmRllcdyd8NaCw2e/kdaBBInaf6v5hYhXk9FixeZxAseTvXQ8dgoiBQM
/1fzun7zhAWJcCwAgcZBIDnPcSj5vN4mS2iuvojaWTMcVZYsQP8hQOKiNTthYb+U
CaUOgWjE0EzYQgvbPc33GLxTzG38OetNZZQEVQHvla5Fe9a8EUHxDXXrNyQftL5W
a7TJ0k4RDfYp+dQgnXvYBQjssSE9qF/zm3mYU6DuaEE/M6+WQxWy78RA+pJj50tZ
DqFA1IQBNNYaIRD/9GevOnNh+wooNjRQZtRZLYSfgwaKSow69G+4alM5cOOGMeue
wj6fsvOR6Lxsr3wY3FQhx7tErSQMAeNbQ/jBfdfIiZXS/YH0oxuwQ8yCvuWkKY6K
Or+ceV8HKBw3UOiZVU58oBNqXA0HOnNeg/q7T1efL0/ND9s2svwli/kBsVN86x5p
FnqiQA12x2z2vq4QoMfH2vNTgadrLyp2UbS9JC9ZhdGSmOv3kslm99jG2p9gN58t
Ed7kV8FaNaEgax98pH6YpGLJ8CuBp4aUES07i2JkQqKex6xFeL/27zWlknr3xCoJ
rQx11no6YAk3b88XsKTUTOzIePU/bP54IYUrtfMBXMgtMMiKRy0M355g/ray7Pqc
nqWZo+wr9605ZrdAHqv+Z25uSBcFfM2BsTef+T0MJZ9CW9sEMaXrjFpMbUOIvtwH
JRGmDmNOXvaE7ygD0WpzY4dILskZcuxI29NoqkD7msEHgn2Ex/DSOZhHMN5kGL4o
luKKnuwzqd7lHPV4z7Iep+1Us4RdtlzznXC6YdqsueBSNWbQ3/hW/m7ALetqtJ+z
iIKwUEshVohjs4Ufaf514ztWDTkXbAj4gTqplJ4tMEZti5WYIpwwy929AAr7d9dS
pqhYpTXIav2Od2NwfIrseY7N8UJc1wJu7pQ6MIB8OvMplmFOKndKtOywe96vXDRv
bixvOrLzrS2814F9HtV0Ry+QXJAX1OcNq4M7yr6un00+2JT6J/9uDwcj7BnlrKfi
ZVg1TX1vdBXYX70ku5oOneEuZ1ceuxCk/ZDHuSTiF4l9z+WpXVxEZ6v3PBSdr+cK
POe0cht1sXraJ84epbjqiUzmZze0YX9y6OeOyPHInJl0LbLzM+Q8A1K6V0p6nIeH
w6QVdphnYqr8FxKdbfeSwNg28rontT4sljYZmJzFeZlL88RwzXQoK7Ix5mJ3Xe4O
CDnrhFCcjYwpxg6G9R+at4oq+HtcdiAH+8Fl9SMttONIB5VQKVhv6+9KA/R/MmjB
TGOWQUSBGV08MY+Z3D3hooyRM3grDzEKKG3CdyHNozLEhccATzpE1n1+h9Yv5o5O
0l5Qg+2lrIKDaED41LyVPMOcH1DTFpcH+RGFgzWWny1ezlCPUldbV1QgXmHsa/bE
Nd6Lcq3Vs/2t9PpO9/BKXBh9HasF2FGpoVCEF8EHgqYfpkSxXwcPWp788v9cHJik
ymx/c2llyPZuMgjVl48Q+Xe4MhRu9dX2P5AwCpFIV5bxEKPRcZShdJmeH9VYbKv1
PcYJqw8GcMEHYqw4JGtlxbSCgRvY0OtvWTggydQEr2kabG8ERtYCh8V8cktAeW9I
h3Q5sSlJSybkmZacLHYo7k9Gz89ELqbmV2VBxP5d7+Il8SCgvWYb0rLoZjXYzHRq
/n7LWVl1ESObyYJV35RSoHQwFmEYTKB3KLOtnoMPDyRKH+IteWLI6B9V7q4JAHfP
fAqMt3AgIqIjpKyZOkeFu7kbtCNpGsQUhU3LdoyOH0wUDTPgDmBh7mBIQtS8QXow
pbD/tLqyNj6NSJtaCkVAdJf6CFfrW17ETOF/3j4/o9d6S3kXqg597uVLPtPgpmim
2S0w6YRBsbgesvm+uGeT43VxwHS8Eusb3IlLMlMbmnR7kj7F+r6D0mQNZPhjbzo0
wUiPct36dd8KrrTnvbjYwEUB6JbexjVSfsydhNqDsCH8z8HdQox/eWcOKwM6C1Ed
/2A7Hr4pU5PbEtuQCk2kuXBWJrvF0XiUCPCeWqvyqmNgYVpXmAMu6Z+FRYZLez3k
xRVhScsXqLjksL1K3KTgG9hYVH+YuAEggQgZ6Apowf/wEGnvG4s/rlfWdaghKXvN
/pSat1JA5z9k1gbdTssTOX/PAY6P/5YgxpmZfK5/w49Uqome7Xd/Y8VxfvKYF6ZU
DJHkOGTcmhz1GmcNpD0zVsVmtoivqEIqBfgbXf2XxJ5w0MMpes9ikwW/hKoZonue
HVQcEzGu4kGIYtMf6tfDYWfTrTYcsn47gD9OW1n+e+T6F3Zgwt9o/+mEVZFfJfRA
bcxsHL6SvZNmT+f1R10l3tdkVK6byZH+syeDzpLC8KcAA8mL+CpE2K/VTMtIWKq6
5bnopyMjjcx/QXBQEqrgodBmYe8mpAOGdg7xIdJDxhcoJUwANlfGiNixNNKJOP3p
/QSyuCP9VUGA8x2CX/zH0g0tHJ7M0NSrz/7XyGVT6HmP0LTPmHSKooN0LRdGTKrj
4oReePVuRovCd6S0+QbPGAHhmRJOxMf9bDPPDk0DBFNzFwp6LlWkQol5tZOOgSET
4SMHxgxuTaHlPKdomxFhyubZLIX0uwaVCloWHHQG5F/+5L8d6qZo8rJdviTOcotn
wxK+ICZBljr+bjNzdZkOWFhlRKXWtyfyk+u6zFlLYAV77QyuORAxJjsxuiKoPuNk
MCEXOjI9OTYb78vduVVrJSLwHIJ9xnxOOT/u8uTtrXBC1xO0UY6aSvNVbHyPjPYF
/V/mNygksdPXAjZwClcIZ6pCUhPKvLRk2qL96h39+LbTT/FgYfhqUmaebGJA6v9o
wIUKuhgz+mxMtC7uhRdVyV+imnE9S+LbWGFSgVxTzCpyJ+vecmx2Lcavva5aU93p
s1YAs97DjnJ7pQhb/uIUJS4KxTRqpYW4ZfgCY5kd0QnvtLU4KoLYnl7VpapkZHta
KYDp3C3DhwSPDl6G0T2y1mFCqRjoI6BikVT/TZvFwVy62KPgw01uiTfBvCoj8O+u
GAjQ/mElaNJfqRzN1ohPrPNKrAokpvV4owtKJphAl9JuJg57gcWMDlmP/UMVEtl9
PDK6f3cJMy7CasFqKMnxt7m5X3DedoCoOdVZfk+HZL6CTOGSmQwRiL1Z7pydUi94
cio6W7MkWOCXk/SAdFLAMfGwngtf3oiR9QeA+XQy2nKz6+PcsMSk1NEAwgQs87FK
2NJGXIHWWtDshD/4WlJn1M84wJIqnAevw56prML9v1VVr7lG8q1gfQVvMrNMlf0u
Y7BDrTUE5mzo2PUiyu8Esk+eMTenSluoR1UqbjuUpK2u4a0Eb8qby0i4Jhx11Og9
d13EDzJ9wJiEBAb7oGUiJ+wczZDa3kS+1KkIzBTn7c0KY4m/Qdggh6zATXS+icGb
CO4Irz1Qgbm4JuPDTluc/gyw85yAj1TzrMke8O+k6wjYKKKPwqFc/Fbx5rEx4VN8
VmJtg/2QbzGgMlCZZYEYZWwChHLkVT4EH649EK1/iosi9Ivwbsth/e73xpKxb7mP
zh06Xf2uLkacaNg7S4bkm0LrnL67Mx/BkFZm4XEVI5fHuX03t/89vwe11sKYDCUq
OOBdwLjRqbJgdxUmNyM2nkPOjP4oKypfqAXGRdOKp/GJ7qa0TArUCGPs/xpyWIEV
pWJMs3ow0ySRjIyRDW5DTL7bqm4ch+5lbYSKON6i1vislkhDSWXTkBsY7PuLOhKa
GruxNf6eAQvla7DjNSCNe/DKGySNcl4+EN1zS7tA1wNFSQnDoWASv81nNL0UlcJc
h1y7ZEmoyogzuOh1BbNrBD19Np8sTilDHH/R3IXEpdTheOddNMUXBdwJuXeTKFyX
PhCOK9MffpFH0vdhQDjpPd5Iu5r/X7/ELqQ6PlnO8W6idNYabqX74ODHomHaAIPd
Z2gXH6c9mljDtSS5Kvo9OpTeC4iCPow9SmIXw+W8SL5/oVFMc3YR5QX0fs1j+3s2
bheBHGdikIMPfrLGtAwfTC3zbaMOLNMOcrlmQMwetK7h8+ztX+YpdTOTTjUsMv6X
6ekELNzCpXp436ruFLG7jos3RYS+kprh+qLZZ2mjZmHwlUMjCKk7CDIwGBxar/Ol
55kJ/T6QXh8wlO5ZxprTX3kPhNa10QLE3mcVazpfmEB/YF1aj6JEnPtGU5M9d/yq
i+O+giEo+Wdr2OmzBW289z7fiO20DY9PyXbBAvzuRUmnoqwnYVWTJn0adGkK8MF+
WuzOJ8dbLri2yOlmuZcSjD84jpCYi/hGEL1zC37wd5prITutaKxNWa+W3NcrUGS5
F1lSIsx8dGWspKhfHRGAWqKrgpget+udIhfN7sDeauyDrn7UWLC6C9rg4IH273UE
7/R+aOkX7zjB52BdcKiebY8Ie8cVo/a2pkR3bII06kV+sOBr5f5pVbQh2SaWnT6F
ezCcHOs6iv4s1FwOv44Zw0D+fppKAL/PZei+BvwTfOlEPKayQg/gQgCzX63sFPJF
QA0AGvb6cT+N9YcnUz134ROx4dd99g73e3rgM4ij9SYTSLjrdq2LWyhAqhsSOF0K
Cigdip1QPc7NmKwFdv3YHIPAOoKbBfh1MFmqcZRFnQf1PXvbj5ICf98k9y3jd3xf
suRE1GUsTnQuiRPg10fDlITesmCHmc/jCX/cqB2aGGoXvjAhRni48vrlE46Db22h
cJwMA09cuiPPw0FuZx5kkbXtvGYLSnrPZD6wdbkKUoY1CN6Jmq+CLn3HgFGHk0N9
Sh4Pv4pFPvLtQ+4NwurgWupY1RYpvFzO4M5oknNMPZkeEC7VLPscqFEGTUG7poF7
RMI/HQNIqT0XQEyiKD5AJDDg8Zxhi4NPyIMWxkgn2yPynX8FH7ePuLr4kTnc7p7k
103xdWart5jqwNtxgjkDrUJTOr9tT8Wn3rnK8JMfYjxeONP5XeK3AE21JV5iN2jw
FhZAkfqwr+nrYGdy6e2U3hpERk1gWVrd/MZr8wR5gnTqWkPPpLOuSSz0qGYQ5Mwc
LzB7cys2Tb5NF76G0QM83N11M1uVswwQRoCNIe7qBgDR5XAVMZeILcKihLTtEFPp
kkm8ejRqlCF1B5ccOecy1pzpI4U/x8rABPZXBVlZ9xwqUDmw01QnZaEHt25LALH0
8+duhTB6L0AhjF+Lb/h81HyNc0V3z7qs+bI6lTc142Ch6eNNpowUU+KzhBy9rxkB
j/gjMslsi4Y1dJXaQcN82JUHvmDAtLEfgkav+0wfD07CL+MPaFq9aVhB405UlFSC
S8Iqbp09gsqwGUQ/9Eziw3uFRGx/C08d8/pFJ+dixTzWDdWU83GZ/6cxGQMnQmVI
Hg2WMx8Wdxp9CboiklD+IZ72zj/RLyjCqljFA5IfCQPoL87kbWa+BHIHt/Z/niAp
sb30rcrlDSIw9yLeYJR2kKwnPOwcl4gKojX4vh1oJAKfbMaxEo6vPZ/0lkulxlFU
Uw8sW0zMQaay2+0tfsd+83dhmKB+38d31KpvuF+73utgOamfFCsXp3x1zz7rLucJ
on+9Us+19g8whuDlMQrX49iS9zWtnRTaGGgWSnlPG4LWPIGMPYYhPe+gQ9sPsRBG
wsQcALNCsFGB4Gn8EuCmV+fYNIjZkzCY6KZfbwdDvJDdwZez7OGoZY7rfxN/RDMV
euOR/S0Bg6NK7DnJEykQvpRq3lr7pSxyumjAM94OXDvgzUB9mHsbGmMYI7b9kuXq
rjX0cJE2x4b/vuAOFVGhV3aRCWiWpYPL6fJu/Tdp1GOQFf377L82U8vB62bdCKe9
/D7wLk4YFjjAYIMFG3ZlAcrv5uKNtzEFnTuHKSmXTiLZIoHy6m8IDGk5oy0Jmrij
wKmxweqHQup+oxyzGm8MYnSzhopuPj1RaGL2e5RrplcDLLUMBa8DQ/yu85lI441r
HfU3QFviCVMjbGM0oFI2bPZa63AOvNbWtMYRHJDvtmAE2bBzyUMtwl+9PLRNhHct
74WBRyeTE4lqvVSCx5sMI3ooyHQ2NuVRFIc4V1QwCFF4VnshN8IWRGouwcZCrVxg
dbqRohyXaXajzDoEWG0YWsAbbUlN1+0SuoQtYPsVNPo/IDJZx4fxiBRJ0fG0Y62H
V4caFb1U+o+HAi8NjXWYguPl4JGxZGOHBjs3NWFWxyPpAYV0ecyEcOBeWMQXR+bZ
IaRHAcsj7/b2tC8uoaXXTP/9+jgnjEE+Ob13ey6NRl9MSljtenTk5MJNswPxddci
h2d1c6VsmRD+NnDfu2ZIpBnLfPGpU/SFnQjeNA+tT3sLIxg0WZtxt1lhsEGa0mdB
izji8i517RBPbDz3c8LrjOqZ9idXFfw0OcN81J7HtjC/+GUAh2h53Utkm4VuoBBe
QebUFmJkKf/rGARtvbCaj4xTiM+Ywvadv3HmW7WIZU2KxjSnHTYlNQzpYrjYFG7C
YLb68KeyUBwoDYZ0GYL7dXCnXzJ7/5x2bRINcaocJ32R99i8g+eDhbTxyhMWMqlT
iW3ecKf8jC4tf91s+AIngBFYT8ET8VE1KBdPmQsPT5Xstx60I1srkCm37FFDMc7Q
Wgul3chsn1yz7fqHBNq63MCSzHSyhf/qQaolm4WQFuKFMYa3L/Wp7smyZDPfolNT
YhEB+E7yE8W+sjpqWmTpkI6hLSClyaYjF2rkR2OE+ygEd3C0rxJo6JeNEWFwQ8x4
Gj9Lr2xNJYkUvXaZqaZRIgPRfex6LYJqlZRtJ61h/5VkEhx8Gf/XTyRr+TZL1qmg
PYDZGxZ/+N2UBR+rOJ5tHkdq2bR51ExqmL2C0VHnLL65Y1kiteNuum1kVdbhTfd5
Bc/U51pvusC5sNV6JRxVDhpR2vhku7JIwRrp1bhva29EUJ/dtkiGPX64kcFJKzsc
mD9VvFI/e8/XPZ54W08zDnYD7oqAxrn823lB5JhkzzgRgAMvsvgqUr6v+H7CyCdV
A9jMoltaZ5uH0rX0tzJzi0q6n/D5J3A9/BNnPnrBGjagGA/0vSQAHh+vtxpgXdoX
R2Vx+jDiOdIfwjiPrJFzTvYChEfxfqbxigQThgLn4SRosqBx0oEEi5HntTulHcc1
s1CgbswLIP0YW5sbMfgA0kjXzyOCeaCcPul7jjCakIO8/3UCBB78tfOA8VmAMWy1
cTNOX19gc77ticuJ/FYliGWRPCQjypkQt53R9TLcd7n6ZFETh1fjttuQC83ng4EG
PSBR2n9WuE1ckpeUtCOzU+o6Du7qa1XI0os7yyci9X5KYm1vB8L5dm3YM116RyXp
TI13iS13MZSQ4dRgiS/KGqgUoPEWvfWWWPhyAz/6BxGJCHwc5ly/9Pnb1Ua5UCEr
3YKwbbzzsb98eeGGDYs4Kq/g6Y5S/ZpqfB8EeCe4hrfis4TfjHtYKDs3wREpKZFw
qKlwOaM0EBPVA4U+4I0q0TztwpkxqimQkxwEV6H2r0hAHLS/LdHCJ3cXnWmXHUuP
qesNXTpPaOLZuID1Stv9s0Lzr/mkdBOZIxaRlOC0uTC+ottN0A7YHxpxF6EHtDOr
yw26SPHWcN50TXD/LwEieXEL7UUXnMwc/C4Jyeg4MfTkTUBoWPrmy1/W+KYOVP0j
RzTPohjo6JD/heK8wYBchiSWRPwFdPGStCpLJ2ohLi9uXi7JUAH1YZHVKF9lr5P3
a8nd48UWA0rgRWFloHJfU5vaJr+gjQkoT97MKqZDIj3+Jcc+QdHu0g/a7wmPnN5c
c6AP4osQ/E2+7Abhns+/Td+f06zSuZ3LBr+jW4ODNBevg8AlQLIf/rGUK8puMmDo
umiWkC9Wf9gPxmcXMHyqDHSMJZWRcrfePex0KaUUTFaT3W+qXV3KVa+ZjFjue8QK
M/5yCZSOY0/ZnDKDgKyPfEK9aPrQk+CWRoWG1+g7hZNIv8YHVD8FswsxKQU9dqRo
SRJcBz55D2JTkWWD5ywWIYyuzdGy0nBICUTjbC9LNs+GdMoqFDmrpyT8LWq1ExpG
PuWvoceYAGIyHaLyutdMMT8OcG3mZbkAub0jF0mWwss8J2TkNWTdLcVD/n96T0xf
p/fmzmOF88lcA94FmZzoaWhFlMsIYW0IiubbBruGp1rsLE5eJilKUyRBom8g6bIb
Fhru+jcBLpCXU+lRb3BSSNdjH7YHlHPeIXlFJJhyKnkvb2313NsSDnegDXaN9hS0
qD2d8XlI9UCsu+jdY4Ov4KxYKxWqYo9LrHJ1+7LUevIBJ4sVTiWVvWvswIG8Ptfv
henv767eOXk2HUbTVwb1NJlwPg5Bl/6SHyW+NOHuhbXBvneCyeHifxWMkuzBhw1l
gtcAh4PRFTDd0ItW0DZ1d3F1I4InJvP42qo6wmOFwo2zPVN47jEggxbeDZsn/THZ
MVp0rK4OhercCKGty/ZlQ3Mt3Y4KF85+Lr1tF8sZ01/xAbIJO1J6/OIpA/hz2QrF
9x3cychFchjA7VnxeRellqfQToVITZYyPpYsUZ/zQONQ59hgXiNTDQB5GnDbR5OH
tuEweqb5DVDAjSohOPqY4Cm2Rn6Ecs+WmaK2tud+rttmjEBOgVTH6s8hbZ+m2B53
uIUEtl+e5otOgkP2eLvzxpSFvIzilJfb58xJHupFSiRBvWx3Be/pxcyTwFuWjN2p
ClguED0B3X64305pf06UOfSHOAfrq/QnB1SoREXi2uFmiUebwMLutkcujGh/hWwR
16QMewxcwVHuSrfGVgeVO58zN93IOHi3k+bYr7vZ+Azu3Y5fy6H0eTcfdJaD3MIg
f/7nNiyS/b9jPre4Jybx/3b0H7dkot04KVt/W2Jc4IuobBmm7s6bopIx4zgUyi8Z
aetFACwMBHpBzbvMZI0YA8NBVrwP7DexPWmwl3CsKJIToCzaUP6wbvYdie+vhSjt
+hPUQ1GQFds5UbIT0FCRt9WjfKdAZP5wolWlP/r2mdG9gJdEbpgMiMaQG7Wk0/5u
/98VqegvTYuuSFN+tEwhj3cMP9aBnmAh9EU3FU/MOooKEIVU0OyGjnnlih8oW17S
xtCedRqQUnJjAGSpdmUJfbeVsAMFqXZcNXpvGj2sJ41fMudwx4NcBWWkTwmH2+47
3v+Dj2nH0RXnxcapkysx/77n5E1j4EU5doG+/jJcP03JSCAEh1YjS4A19JS77RQ7
WXFyWsLxlbOIAGukQR8JMl7Zf3HxNUimThRJdt/O2ppQ1NsrTh9bjczJ0bsPOYtK
f53hcU1qAUdqRDaDg+xdUQy9CXkcOAQpklYUGX8DZe4Ilk6H6YYB3lAfwFW3Vxr9
wKI31aB6zuDZYypjcvgr2baXzcKc6WWxw16x2cJBywVpWOENLLXHdBydfIA+7CJG
4udDp9rI0eH4UqESCBUfPxx3ATGzlo/hv6u594bIOzQFrOgceEc+UIpXUN1bM0nL
Eo2NRw4oUDhqRP+sJ8P7jDZI5ja4Wgj+SN558MYaty9dH9kmdzVEAMi9p+A4JjCv
TFxubM+4hHnU+46toko2nqZt2dViV2bU2K2Y3NCRJY/yHzFauokEP/uuxtajmol2
12KATWvudUleGF7+ybUp4B91w8+4fPUnfYD19kM8F63eEMDOOQ0kEQ7kZERHM2Mg
pSgsXAgRx0cUjw/aQ4YSh6rVPouQ87GWeWwoqyBb/FSyqGw3p6hTf2hiPDCwPGxT
gvM6lSo4gycQYIrar0KSrgC9f9+GWpCeFyneet1lLsqdQQzlLeDFF+1UO7hK6Wmc
fA8ss3iyYq4Xd/eP6/RglciFs4SaHGXeI6pd+YIOqDtlZfifEzWh3kLJPqmx9Blj
uz70r/ecT93fsuxI5fWOfNNuJMDrvdWNmblFta3qw3EjS2XYcEbWMeKjxnfO4oRy
QuOdQG6zjjWJfs/SpqNMShcbxpj53Y3PhYYqJ9c7kIIGGK1RZgVWGRO1tmD32zHs
7xO67hvJCBRDPMr0cSVX5LGj4EhHED4W2Tzs+jnhuYGjUjhBGUpu+bITUUwS9qX3
qjL5SKsNyY8d7n+w7OF5R2mOrkJyxGVvwh99ekFGpu/gW/5cAVPUqptjIrlSy3NH
nt1FKHoqVTnfORCiLi3lSUuE/tUGxxbryaZJ/FXrSqbVAgUWO949XDmPOIPZ7iBn
H8qFnghQhUuaYvcbVIwT/9HzA1vcMrEEhpl/S87/ww4zYoS7SpAsgs8JvoJd6tpb
Oe8+tL7eaXW6NusOkwik9c48rGzueOyPLmRv4qAxvGCPso12qmYiwfsFckXi1RY9
HZFGFH8KYE1fEpjURc/hZODEu6HN07fAcS6PpIcgOASqZyu3Yia8ku61URCHI5yB
Tiz30qd6JX2/t6+0G9juGem29Ww1KcD028KkpABmDtF9XzzDV3QDTbuw7oWWdMm8
NRxVIgcTTeVTihajxGwnYKU2ZhrFDu91Eg2sRFHomqa4Cp5GY/y9SzVOujLsPRuf
lQDBuHvjYIdfg6Q9dCcXth76YEHAmlbtBiNWRnGiu3BoBfSsQn3qwaYWaJs08/yb
/us8Dw0ypGhXI3VDpusoyBcxjMdwLjanXW7O9i+c7kj/1FPIJHGU3MjXANgp4DQ4
N6nUbGtl67+b28LV79eHlwDBILjZNopE5AXGiUH2y62X8g0dKMBHChHndamnvlGM
eq4wyKO3P+SqP0XQiY6k5dn5EJTPs6MkiVO2TxKW3e6wbI8KZWwK4jq9swJhVdWb
vcQK03ttk7wM0GzB/NRIJdEIPov3NQL81Xfo/OyoWtDXVAkb6AdO14XoodC6kZSI
RfOz/P8pww1VSpDnt2Ux4zBe45Gs7RkYQaR8JjCTttwgq8lluoXs7VVEhIAK0Nj1
s+Des8QK6ZI0xfd8ZA3Y/iTeCPPkvlJ49TaTPk47nUh3IGKhS1vRSqsc5G2+sYO1
mBNntFmoR9CGWtx2D93+jmff6VkUFU6rnYgtT1r2LGRyneq1thhEK7XZ6utV5wLQ
m3PWSPwREIgCVrzyV2AKsdxjaksBGQAqoaBsSG5eA+NRLljeEJ013D48RcvhjRt2
+m6q7BHJjhXQWIBDkzg2JbFOrmmEfKxmUSCxYUcIFUA/H/swWXHfulyIUg7DVEWO
aN+SwyPw4eh+A6YtFHklFoPOpqNvnbi506pS7umMH6SH7/E4WEnXqiEaToJpnni3
Dyg9gscJrHq0bTdxxvOe44dDVdM6p4tLMcVIBWy4gMYfAEiSziFzvEWfj04+C12X
DVXJbttnSqDl3WLhPskA3M874vq6Ja3N21s+BQdLKjxmHX5QpH8yM61FRxEldAlc
aJt9r6BrG8fNvefy3W4ZwUGDT3z7Q2Baotg+vVsI6F3XkczOwGJ63iglGGmYw3Eg
TUoIQxADtfDCF1ak+NVwWun7/YCXCLZyzcP6nL5JVbrukNmTtNK3Y2zOYKHcE8bv
MEeWHqdN3ih1AWokMthHDGoVqezr1jA6tO7yYnL7eE6otgUmGS+L1e0Fq9p3UX6x
1CAjORXEHjqXEg14iCWEViZV5au1pyo1uE/9L155VImsNyIXWjADQKEDD6Wr0m9j
NwZBf5D4hvXwqxNnnFRupgcoBwPRk+5cJf3TZJgkyh5MsRqouFFk4tlrBkRsdXa8
ZRr9CFJdpUrl9pb65miNvKckY8moCaHgidTtNAtb8w3WnqGrhZW/D7OWcUpIX+B4
+Jo+QyVTEPxJnT6SbW6VJNVmpYWPX46k1QR8tBG2rDjSxhgsS+31FuN0Hh0DTVDE
Zqm+5dnpG6mlGTNi+/kaQf18G6x8OVHMgTQAGVL0JTQdO8FKhv/7QszRXRuNQ3Zh
j+9SPY57ezw36cPKjcznoYW0mtXDFL//3KpJ9InBdhkIerkeJf6VYIiRC4mkK6HU
stmwBpRwiNsXzab7B4sLL1b4MjKl18O1OBTi5yHAzb00MUzpybH4Z3RF/kmCtrPT
gy0FiUdQHelmbHSVP4pbzcBswf9RB6b5uzWr8p0yx1rlcpTgL/H4ttt5pwfEJtwB
PPkxzqtdOhTzki95t/r6Gb+p+XJUZwKAnoADsWPr9Ys1fs3E+nZ2sJtax86BM1Vf
7FcLDODLCdRYkuC4K6Dt8DPn/KgY9WcHhs6UWecBf/GpUPQulQ4QAHBYUuoLIABp
RuaAD/xgC+i8yfc4XBJQZ+h/6c9XzLlPDQFon39WEzB3m2iaAn65nxNaYUcqr3x4
tBQkihDAGtRUEtORF19OFRy4VDOf26OFJhzMzb4+odOAnRk+M0u0SPX1lTuFxWLk
c2NBVM5EqJ0bhH5WiprJMFMMxMirOo+TgcwjhD0kJAHoZZXnwx0SoXQ8YMdrmcF2
O9j+krvETN7ih1IoXqppLtGP7HPZAtxDfViK7+Lxw/gjTSRpY5hHD5acBg2bReg1
wWIDjpCevyXzeUjDZIAR7pjIqk4s1NpnLpMBTiNqiaXLAalwp23F0byb4BPxdfpG
/XzUfjjaE+bj0v1yMBSNKJYJ286FJaBWLQIM6xxGUm851RhDka7X6NoSpL2Kn7py
Kmy1uieRb2QKuqZSbeR8CWQL9iwGl8n8feehBSx/fkXIhh6vtHyUM/4NujqmLZ9i
ROlSRX8AQ+blrBCJlY2FfnnTb518/cbIHVlb2KHRshjRu1o7PvJIop3/fuazT7OH
NgzfJMmWUr7oECjIlqLtheP8K4iCSvhJk3tiXa2akOSztDUGdVeB0PPJxBNk1tzx
k3/jgaac8MVJ6WJkw8YObZUnkhbsT7aemwALMH74+40Dmx3FLckMA5pw6+ameklm
vNojIRaBw5OCxS1sOsSkYQEtZTMhFfagLE2j9QtqKWMpPvHi/QZcYBajfUR72Dcb
AKg0nFz6RN+mUQon9ZDmM6VGgSZQveG2wctC05r5I17myGsoJwbfKc4gG21gJELA
4RE6WyFxsh9uzYZbDJDkaFqHrXncPOeLC786CkYD0IrQiQG50etw9Ht26mMw8A0Z
Xy2dwE5lt1Ga9fmppKGZTG0vFItbcEZbmrRHRtWtuZAczh3y7PHkkW+M0YVkpucM
nkfpV++B5bUPPyo3ebNxrEzDVPyQCI0Rr1myi3d6hv26r/iUN/VqGbE5C026Ihp4
9kFi4bQKAxReZsSUWXVUfOmhQeX29G2MNpcamMclBV2RpZikCseYwApJptScklnJ
bXnDOBvhBSbQ7bT8ADYb/FbWkI6nQFaQqCwDtegkU/iJZHZLJw6ePtBx2cdSgM79
aQYFHd+tP1IBwJ6GayiZDHLTH8k88Opcqs599/knvpR3dzZMojkJviK1Vs2wDdnX
vZpNkbO9Cko7RkqO3BpmOq+R5vzOBhYT7JxcxKQ7Si7mwuuRLrG58bnJ3LrB8nf/
4jQR9Ht3gQi0D+qu9cr+hCS2ICK+pNCd0gI5PjyiFZbIl+TYWeVdam/pIYBWW4OW
Xc5NANHgsUdc+SneHxLxRmxSV3HGPQ7m9RQPiW2cwKSOj8s7cZS3BHtPexnj7K9C
2eBPuVnXepftaGYI5tQE31LrDVUtwHk1exuZHm5yATjjq1dVfSGTklm1h4A2+p59
Wtq1zNEt0MDpX1WLR6fsRNcPXpJZ8uVwbJNXz38jNemxGvzqY1q1nnnK3/K1XO40
Ttm/repCZLm2Vkac+AaMtUaCKgbLtJLhU/iREZBfmax5RTxxk9bnRwcn8PTaMzhE
/r2j2Zse4OQjadzfhhtR6E0dgI/1vgMn9pMYjJ9lD9wnQCg7qQb0XyQFVwFLbKsq
PbWEETdBHjwwy4o3cwEhaL8paDOT2+Mvq+9nKF7RqvVDS96t9j5o12hvzvFPaBeO
dhUnVVfkNUhknMn6slIHvNCFNbcOr1OPr+Wb2rG5NHYFJ6NysPrNhD3+g2TI3K3D
IngKDpdiSGbkXboOopaYlm3Dafu70jxFR1/M4QrQbxgNRQzieYStw3FswyxtJulk
szQ5ZLiU7Bl4NLWJ25rsq2CXFro1UIT/lVFTai+GEPhrtfOu74sawmgWzcx9iQSr
Yi8LAge3s3KW0QiNHPpCIoSlJTcuaH4UyHvsAUL8woiUcQu62SUWqBqMyjHfhlfK
UniRJcNsm/99BgPgoogt+4v688eWObuvQShUcXK/Hz1vzdWOafCEi0VivlP8h1rJ
ais47PFF2iyrClTrS3qA4Setx6FuS0e3Hn99Yc3vkZADvoAQcWWU3l3Umimp2p1j
AQ3epikdv/pgUNbcsF/aVxIhyt0A2CZrYg22T/uPl9Mu46w8zXAc/4Z9T1iL2pJo
aJWf4r5P9QmwdC28zbamoirKdawvWiy+FajNLdxc+ZkFpubiyZ+zFpYACoHvQ5OW
YMxE4nmMfCsyObTekBlDFaof2DldQ1v/X+GoOn3vBmWxuCeHbAWomqaLJgCIWZ/n
SUCuhYZbXhrUj/z3MxdNARH5ONmwZqxqAGKYiuwVat1g616iz76IAxjQPV++EYvB
sVYvgsZLAp6N07yMLquo0m2BTocZCF87OUH6sX00jdb1TNRDOb8gPRWqp+78rIhE
NuM0ds0ClcCl2Lv1NX7fUQMjaivhXw65BNC1Eaf2mknf4WHnj3Ixppc+Zm8bsN6+
Eq2Rh5XNcpLOEzURA9Wpiydn/NVPbxDT6QJ4nmbudZmBsnZqANywnWye+Zn7bKvd
tUe8CP+OsVC0sPbjYxNrRBbS0fY3hwEAJLJBUg0+yYlYEHj66mu986s+idx+bBlV
n4DZRvjKo2keo87Ws8a0x8tFoga/lcYnY6d6kYGoEsejy2lKCrzSIKuFZJmiDhaP
mViDaLOgiPgIZYj8G8IuHJgGZ+2KHvM8fvgxA2OrizDLA0tzqmF3I/zIfHbEY5LX
O6tljBkWBc2I4Ct7Wbfh96/Xkq3W8RnqVQs6LYHPxWUBqC8evUHkTPQQ4zHvbSQ3
+HfkWcFoFyAoPb92UPizzaOIkrsM1Yfuyqlxj0WvHNbEMgETsMUEqcznvkC+xz2C
YFbBRxYpD1GHSpnYJ5viExOa0+5wTXMFr83QJIICuY2KJZqvAEodYQNoinIgdpgK
VQE5Y+AGyIIB+rOpvDYx1ZVgF/LOLd0TcmO+Wm0F74SbrjSNb6SaplMnOhdwuPd6
japus7/CrhkHCc6e3y9JLS6yVWwvkxQgzCNCjgWlC+sv/xJyTJQnBUtbDDiYVEoe
3ystUWNtpTv8zXtnCFNDzIkOcPzBxmoMSI9TDeaLt7fuQALV3Jgm82a7ZKEDJiiY
MtreKdve/XUP/SP8BMu8LEbAO+YjjLBcxn/wpJAGRlr5lPsuxyiI5YTtVc7bJtVy
L9zyhLzYAtqXlRiF3HmBIsIoIs3MFgf8VWQKp0kxcyc9RBrycGtiCUYUz4k7NfsH
BW5jEaD/xYGeqrEEo5pqmnJFWNME37C+AaKZp2rAv/8bbgsh2tuvMBDXHdC2f4Pb
qiaQTIGlq6y7JumYYP5CVlN/5Ifr5jNlp+JNdMclQO3ZnsfemZ9CtUwkBWQIjWxe
Z3riBANj5hob6UnpEiyv4z1tANBlYPoPW/RbR+PmrFy5kDkfMh3QUR0bVRQVRQ23
p6E6xXdwkjhuv3i7EZeuChC61ZvK6f+NkqVVH7tfCKllLnrLx6AvTb0FYFqcywQ0
1zr52ENWSV4AtrihQshROGkLQ3+qNjhu7pa7gXf6dB3LJmbYo9bYR3bUcMI9X6QS
AInwMxmk3wWYYwLRcObJ6ctxgq9L+H5u2DlwXgzqLPD27AzTyHc1vz8qaQ5zs8rk
rjijoaAma+lTnWGfGdaABtNW57pjmJU4V1xeZzWpW0zhQxP6J6e1b/iOBHJOcDE3
ZZDKSes4MuqxWld+fPO2cVjBv4y2FIxnt0NfOZW6lUMScKv0lrJXKmOVIP5qBaOo
0fp4OFndtxXlVawWlyyueHKTNhdBAlrb7/Bj+sNpsWwgzVIkDz6Eh2LfWQ+QFm/k
9RxkzQ8Rj+1TmHmOispXfNkgm0BveJU+L7hLUWPLPa9HFOQKpwgDu8y8cfXYP56I
JJ+ERoQM+V0kKYhqOVKfbUJ9f4/SASD7orisQpnSEvG5Y1ZgeqU2Wlhjg16IS49s
iNX701tpM88krjAIQhA5IBbKfykxfb2B3cizC9dtN0JVLcsdP8L7CcM+gdtPZnhf
aHWL3AYwV4XYZ1qlliGLCwj1v2wD3xR4Kv26j6TPY3k4aXUTUrW1/HKup9Q5dOrH
rKdaGo5zPlJo3goKIsrNLVB6WzmMSIXSBfVYnqADxS97S0HWg6/CXBaxHLq+CGF7
7A0yP4H8pk+4rYvwb00WxijLIpV9XdPOhVq1PwWXLKP42bIic2ID/84FoedbIBGm
aw1A3h1Fg+smRl/omJhSq+pFGOnXWSTIgLFqiNvVdjvGWZJ+N1OSM9L/ntDFp/WH
swh+2mJzlsmgwLm3hCVwyOd1Ol1Amnk+4WM/6w8AHxkg4kq3NGkLEiDfsYtvoBMm
ywfpso3rKUCOGC6Hzoxooww7f69fgMotnJLckSdbGDLhKXqlQ/mO5rx8qyIZ+OTL
7xop+wkgbf63ZQuoRUDkrE9gkKJx6eKuPRpFEmJDmfXaXph7ANrx7dkrgXPena+y
oSXXo2DCIvqW+k7diHjW2xGRj9RYr7JJupIVpzI1zTOS3+vMKjExPu1x+y4oFmT6
s+xTIMYHu4PI0G6F0KyEXE4TVLeiU0+rAMLyTSVWRtaZt6b2OB7bv922Pm2ASv1K
SxEL//dQwrJg3+gEm/mRDWq19WoZaUmfnx9HJoEafRJs/HLjuSFBk7ag8xlkf83G
`pragma protect end_protected
