// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
exDgEUyGmiFc/PE2nlcd0QAJkJGlcfCsHWAGzHuZA+gGRRI4p7stkUKdc4GgjEkU
/+i55bSmRSv+mUzEZR1dcWzrfrYKBS3fL4vzy1ysK2rGsPXxEZl+b77QVYjZvlyy
vwDiOHnCsaLw4NIAX6ibJPd1YEEJa08o7OSSX1m2Ni4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
tMgI/dlYINN5LWDHEzol9fjYIWQcBhLjw6+Nds6+PQ8UcKElQcsdq4r6nso/COjP
ZLPhwI8p2j3L/Jka2GFmMA4efHd5yae2iUuM3dM/Gl1mIkldXEqV7HiVFjIR/miX
bv1UmU6r3Z1Y07yxGv3dPI3LjNXIqkvnOHNsSVK+VBuIJk/+yjYHZri+TkWRlL4R
rOfXRu3ol4G73vXlIV41dvmx0UeMMOIF9xTWKNS28QofjdrWY29yCOAdwnAn9K9Z
fOovkX5v0uZGQBqNp179vufXmcDE2G/vPKm9Bzw0tdwcPlHMYBMRZgi+DvdyAiNV
FAg3/Mwlev+6lZ+j4OSQQqVxRerncyHLv1tsxB7Rz2nIsjVvPC24KUhyEEhleY4f
VhOF/BXEJ0H267FW4JuaG7gpyFLkVHNfMCK+z/AcLw8+OxzxR5eHQpLkEv+QoMOO
JTNrir5EYEQ8VjkGuyQpSyKr4Ihz0Eb0CWC8wC1dz7iXZVCHSLQcmzcbt1N7iYmC
55Hwg9t7aAjxCgbtILBrA26EiYTOOG4leLrtJS0STVpBDLxcfcYCl7zZlP0VZCQU
nNRZW8iyKOviLdf/kCePeAdrX2WrXiXdx0pDyVLvZvPD1fe/nk7QkaH5n7QR4mDm
HrgszuLuB4QSewZQepfoQ3B/Oa1xUAtaF7vlxMUp0aRZtfcOpaYwWOJTExQegWbR
rmLvWDQbzwNuowQ2RxlzD4Z7R690YU40mR3PZ1JUT/7d4RcRO6R1iu04z/fduMn3
9vmtjq83iBy1Oqlu19Fe8vomteKk+5Ju87QEXRIMK/qU+jt2CY5GNEitmJTx4XFj
Y5jNIJzPmJBhLUI8hdGEwrMHBSIr5f3e34dt0CxFuX1SzWWok/tIXC18uwsmvfzO
b2Eq7ywMXJFQQv31Nn+7fRPqiAEa5lthxe7Clu+qbm2FbvpCXdp25gtSccaKepWO
xUHFbu6OOugWFEvsKlmmN+1qRt6OgD9Fp6DJszAG88SJM2H4fqmYii83GqzHQHNk
dn/mei/PW2C3ialHOtKC/cO09rzYiAi+Y4/63Zh7x6QCHlLQBc6DoKWYcE0trTrt
mMudb9nXTdAYPQC25ExGZw6DUtJ/fHPctBhQGLYJgyF2LKxDzLtAIq4V8fBhcBzF
p+e5sYI/aukbURDDr2pdaxdHnUpwtRCq99+ou89zc8IVAR8vQQiA2/4659i/3E5o
eqDYdYsNUJosRjM+n1Zf3D3D2L1tAWOtXKFFVhH3j0Q1dciu2mo4gLFMnfZDBFmd
qkdnFHAsrJnzrYPrqgMYISyAg2pMHjwMIsL3pQ5XOaJOQ2ri42bUEvAfIhTOEZ+e
XPjOURAHZuNc63CqbD5FGTJt3hA0qE5p7MWjG8thTkTSKo76zwXpz3mnmVzN0Sdy
uKjVzjoOPQOKZO5toK015+ZghERhpEFUxJ+yiKZUvZNeqJws+MuACfxQFzH3oTfp
VSwK0VFMvUgxj3mL5+rZ1Yh2ExNklzlJMu4f/6/yO3cLhVfLy5Ed10LJ0ajoZi/7
L4C89tyDsaftyvbTo3DRquoaIhUMZMt0XnXUCVgRS7z3Y4AXU2bWsgDBrVu3d15I
eR2NhAxyt6qM3N9Gt4b3mm7/j0Pky+dIZyiP0NAG7nVUXc4BOsZPDQ/8l+1IP4oa
eGqeu/3ki2rlZCZKLQoRyaHYyhv+MgVycu1Vx022Xy5uBAMEtIPBOxAqYEaCNKWy
qKdBoxGo4wog6R8ZOMlJto0+5wz+wb0vLLIGToDTAl2ckEleM7wGHdFs3S8UVasS
wDFT3ls16kcdcbGqFwLvdKO0OvPapbaWWyEMgVrMoSgqGqL8yJtZkP4wr1qXq05A
9uXUQIpeZ8Lrm6lD4TqhiPhWEGXqgD8m78lEI6Z5d4Df7Xt0wnO7H49hHSghwN5P
HVXL8/jCCZxaZa+jM0bDYl18vEA6sqKyx7dkEY24QVQNpJQAIR4CC9cMrvy421Bl
YxGbj8DvnDbr9c6BvM6Amr1w/OhenJu6YnUbMfzAto4Eo3+VxvHynEyKA2aX6YjX
j7AonegQu/rEfj8ObIpqKdskGYqoiHkrOwQxgM7oAjJkU0MwcNZ4vMFmLyp/V7zG
6jn0D0HsKbArH5atsweU4mb+ETLsLCZ9bT54TEkQ2lfcovJbnVctbRh8a4CntK6E
YWqWxG04/6IE4cll7OxU9AEZNw1NdYmSqwYa7AH441K2hJtqpmcXUjLNEg9LuzN5
gFNrpk54t/fmH7sfi4vbqV+/1JjLIOAMn7ZfHCiX5kE2N4RId47ZePD1FmaoaFof
zG9MfX3wlEKUlrSkPpUcTgdhyI0JJq/kuGk/taDt1IpeGiHN63k6P6u/8qHcH8R7
Tms8c+mzOYNZjIBLsrfvObKfc3V6K1aQWg2fe+EHg2SHiFkT2KiRdBm3hoWtkbG0
jjGJeuO6TO5f2sm3CTk6OHfo50jR+0HSzUrhLeQ/Dj7KTxIsAa/A00JPO6/5A1lv
70RtaiQa0Lq/cC1NR/WZElxl7j5o7tLs4kI5kRVU50W3KkPwo7wnYUAOhmEDgEFs
U7xWiBg4ubLW4QZ3/Xv8XPrd61l0eYzM5tflTmSLJLBH/cyA/WQsEGU7nP61CU4Z
Ncpq+PSnxqK4aZ25JGFY7nDZJqN2PT5ZTYBDoZJgjt8GeJnoBDXMEpTEWCv2Hbmy
R8ExbiQpVqwMNSwL7Mh8OWaJRkMpivIBf0eCzl+3LHH8TxynEGcBxmj/cjTwoiiH
OfSe03N9WmhUEVpghNz80PFAMRyoU3+fQMxMOz51tSBz4CC0hidzmqMOGs2XNEWN
kS9WwEpyNdh1/a/cgwzUJGdq8nR98rrjSQSFiCWAKXndj3Dqu4bdm0sVHTF8oL33
mHEi9MTo5v9U8Njhy1Hg3eWVh9+PzyRmlSvq+4BFGGnMvpIvuDTEjzNi0ClwGJEy
jP1UGMO8YyZqEAKRcYehFg==
`pragma protect end_protected
