// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
k07oKjI4Gz3mIv6kK3++fqt3KqmXez6R+7dpPPXOK/n/4vHorkIo02ulAbP2IiEjElMYY6yXTMW+
Hk+y9AXBIXpmp7AtHf2Zk3ynPbVaHHHhneHpG2Pb1IUtSdd1f19U22FS5Ala/6DdUHqFS2LaNQWE
5HCvkml3hT3SzrDM8YxLdP1A11GyE7n0f7uJdAZXr8MH4hGo/kEcPUD0jcIwnUGkxjb1OgkI7T4p
9leJNpL+d7DXtRn5aEH4DjYEBfEdWu+ULzKuACr/JmBgPOnHQLCmkcl9jc7fbU7uOdGtL5Ij8IMh
MS7KFzCs14OUBQO68XDPOYw3Su7uLSgVd0AFgQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7920)
z6iAWzmQ6bs7ui5DTFa2vqPwDZ0OGMhVqanwasD5ZxQC6hH+49x7qE8T12sdBhk8OxEr/KlD+dmv
igylET29SxdBgcHVfa5fCidVTUNV50aZRPRSMjthBxcduvdEzz7AHmVZL/Q+cUchN2ciE23Gk4/B
Czu0k0wRXanOYaXwNfaFKUspQCByxNrtqHTtBCYMvnm0S8PViwG9iwyurR1xPARMdT7BgrnMN6SE
al1KTeEvcn8ux95lR8aKL5W6cQbLOyT9qhtRD4RXV1YsQSHbJa5bNYCuWrqXlax8RgTGtMLKl981
P+7KNcMoAWdl8rThORi5eeX7AsKqjNmQIYuxy51rX27yfzp4cpn374Equ4w381mo3RqKqiqowCZb
vWON+y3L8M1JtLGjw5+hXLorzTrBCF8UCdDHRKgDqRpLG7bKN8vHJSh3KQbBIGtFnzryMKzsr2Ev
QW5u6O/4Ah29PlvnQK2+8PWcAPAd3386HryutTVDO7K+YLvBxsAVul+5i1a0ODU3F/duITgwicfq
b4cpDzzNQeu/D7IRjbMs5xPNtOV9/cuQ8U2Wg/CCJFhi0IUNXOAYt2MSAuHU8ptNRT2eefNRoYwZ
mLqQrvaOt84PfR4z7gpldWifp2zf4eWxFqLZZ53lfI5eXBK32AXGghThiossa2tzHsnzVRV2hqVG
81ivB991ChMsJvHJD0btWGJdeiXqKLeQiK2W5UyQlzhv236cDrLM2OWouTqd23C7H2SLvw6tpdKo
FRIP4OBdQZcwC/4EZz8VOFTuX6wrvwDRAyvEeOwNrE91abTybkiaWOrHye+CGgG0jYnEdtUJWBmA
1Xt9K/VMHN/1kRY5JT2FByfn2jBBCMgPHBLzjsnu+vKcI5zgIDQY4KAJ20Df/5x9xjGtbQ+R5hrg
+QKA7Jo/t5QVYb/UtpK+X1jyY5YMw0RSN7diGJOUcvB7+pNWrIsbANGcd2Mfr4giaAa9ztUTvnW4
5XOdkfK+YRZvu4BMd0zdpnBojKSi1ylirUNmKUGm6djI62Gmx/clFKHlR2w1O7VwiPRKimKzJY0M
czIK0He03GEt1IvYY1PpHJGJGSFmz8GjpdccyXTZic8vlyLSgFknfH/hdYAATXlGNMYBV6/tvbZ+
adjO9GQ61Fv48OFBjYGDyDuxmYwEjIbR2wfowKDhtBJo7hyaCdGu9d3Q9t4RqlSJgkvS0SBRrc9Y
VfWaun4zatYBv4zJPyvWnI+hconIv2vZiiALsCG+iS01NKF+VHyQb422lrplZgcHYoTxXuYs6z4t
RbEVffTmkoMvELICuxHUaRaplXFQzWN/9UVTTv2rKZ9+Eq/73C1BDVBlFTOfnp/fMmZfSd/mZ5tS
77i0kREn2f+63C9vE2ZIqPFO0Pa14E4vH50eQDp5tntygJJr9pE0KH52QV3IGGaXUcOKrN4qyu1T
F6AyRpMSPBnPVtAqFkU7dxcsvXHqzPbJ6To7CdTQKnIvYE7VtW8bThTVLJD+pi6iv+Xg899Bx5+C
fXhnnDwOONHUPNIN/WerWq7t+oJhpmFG5dFGawdoKK02JfaEdxz+Xr/PtfAnN2i0Ua287x0Z06AK
pLkxoRD1K0T93xI9yECXz1FNl2Ks87+EDhi73hxID1QN0WWEi61iyFtpEU5iKMEX18//rEA/o7dQ
IWeLp+QWYNc6LE8cgydGhNmyY6a+weSLwIiIqCHaPRzF7bv7WzseqEdgR1d5wjHLqA+Lfz87gSIH
jVs5uId/37ViCac514AANN+1fBYJljeiWsVCvbO2gOQzyUDo6KdDvVqmR9fc8t1D3oyzT6OrgqgG
kkVD+N1zcUG/QP7FYV+mnV00TsKuEUK0hPzDOFU812tpIetQhDxFbwirx2vRBaIW+X/aMYv+dzyW
ESUz7wlk+Kr5+wAccIYvztgCuUK93Ry926OWluhyW0/lGCXrEHDKJ9+t7deQb/7xV9QsYLd4r6FS
OV6ZNB44npuF7mK6WvMX0AfRMuDhxQvTzwWrxIVC1rIE4UCusi4ArSPgL2xUyaB7T3iOHJ7/QfxB
poKsozTguphErxtPH51hCxiocrvWrDfvfw6NthP+L1i5r9fhw/x0pw3MG3f+/kvQrGcvDzp6ngay
Z767gaxANukVk7zJdD5iX+JwFbJ4xVdpnXhIZHvIgka7L0cPolP6Ac+5XA9UjEkLok+OxoIrIk9t
jjqNmGUcV5aQFwLMojTrPcjD2jTadUKJuy+urVFh+vI+AaAUDhsuZ2scHuVOewWtiJrDyIQTYWdF
0JVYM1kdjI5bnjkLFrg13PPNlxp5knf5AnDiNb3aibxB8/f4d/rGnPgyieA4AJFwD4Ck2H6RBLEj
DYzWMqnxc1nnHzyVuDmEsInOPFWmmxt9BWyiJD4yLA4rBD6w9j/jVNjV7DbBFTwaR7xHW7zEyH0h
0zIZKscrBL6k47U5zwFNqTpnAJG83HBFAqysinzxUUNr81qPUjliYCzI60S0iUVkxniiOsVu19F+
nGXCwTI6/PlEQpJuxZzEup7H4y5HJhLyE6meF3LpA3IrCBg/OxmFIGZKrFN3BRy5zI5bPiC3MI7V
oXvVgUnxWtEW2PNNIbauauJF4XLTkDuwcjMnM1Pr/NL2cvpTZCFGuDweQ5v7fB0ZGIZ1L+vEGk1M
SUicJJV7b/lCD9YJ/zKO1FRFaSh1OSqjNG0zVhgCHpe+yLnKHJLprW5FuV1zaSEzV+M9gdy5etDM
AuXm19Gzy2q9ZhbP8ncJWRHuMVF4tikTakf9WiMQ+GHjrtbOJYi9vjvjjwti+OgtpS9/xRAe5s1e
NwGmdBlTKRFcUiwsNrx/ysuVjCCw+nyQuxZWqmCsajI3n2f6NccxQDc69twT7nEPSp84BpRjMDTC
ctdthinyC8tfJeGFXlGzy/pWMgkKGiiQb5cC8SBh2gVmCW5X/VU9L1A3GG5K1/H32LTXpmhEUMWc
POvyfYxoAVNPeSsSYmlr9oZrzSjtZ5YmO3F1fz/wTGmZXm52RXakIOlg77znLGsDVHTbAk3LCgBE
JR0VR7EXPIf6Y8UW5gUmEIeVw0OdDCoHeu58yiwq17eEomniMTjivXRLC+Op6FltOLOVaU/dtfcq
zuOp6aXYFycjcAASoJ9eMtANEPJMFjb242VA68HnyZ1JfiS3G4YV9qAW2jDMMgUDgsIELR+KI4ME
+GLPyJPCjPTzLi7Kygfnc6y7Z3/0/hcQNkUAgzmFGt24scUE40QtdE+BO4e9Ui6/AdGL+w80RM8n
XO2hjC+B0J603XWDfvO4LGxRKyXjySYYRBg+N3fDrYDQIP5f+Z2Nk+fOFMMJuKTYGvRJXRdLz+JD
9upajtupIqDQu1RMTef/Xgqa83ODaR2luqGlMIdI3009fTJZCnXBwvWRrmeSQ+auLuAOP53Dlmx6
fxGa/TlJUSz9LrPMSQuzquxCFJWLPVnEifIAu9PGDKG5UNH9D/eqUCwAz939o9URdp+U5zj8Gzpi
lGqCvbqxgSDC/j/PGpKzdE8OB8LPYQ8OI8i6bcEOtS/XXRdUD9kqxTr761X0WfpbaAMLKvX/2LVT
uBc/eATzt+DzTqDrxxe/DcxqidHmt6kDEui+llSkVpxbxxgb25ikePRXEsJ97TMTOo+wJ+HOnW1O
vaaewOesAsJVSS1i0akQIP52hDyu0JdSP8tpfW62sIZPvIlHKLOuTNsOfxsP9w+0HmeqGPTWyoNe
I/yOOnAXhm3Jxjms5w3hzi7a/DB8l8oKrr4cn5W88QQn3pd0U4npVF9by3K6H5Pzf/5H/HllkHq1
649hAZTdit0DIWBSBZNT44RC1wFrjzxSkLONGheYZyIncg78hgCCWqNgZ9IxAlzZkXu9PzIgSGYh
2RBF21q6JDc47NlJjEBl6ezk+I84gXJws35l+PunnYFetuGa3YFn25uzEdzWwiSL8DP6cSBTtZc0
v2nbl04MYCXiEbNc2l66UPde7WT1Cn6qqHS6nGCu1gVkcDM67zHc6cZOHXn62rVYweE6baIKxsqE
Rh/vi6KZVFDXJuHPsotofoGR9gC3uvEfvW3QOYReK9704dzw5ywLxzZyEpLwzIUEOZuPfWdgkhde
atT0c5+RIcx3WTBtBFi6Q/DvcyceWXwQmH3t/dE+SyXCVcFbalYpQfFePje5YTo/mY5ZVqSFa3bY
BqoklPY8S0fUi706KaISBbopYlOFF1BpKxZgBlM0l3pwTzrLYkbWcc2rMRQgXRSYXXNBoI/YiNpf
5jbiT/V8n7p2htprRKnqzdtQYmT+yDbZvkImCOwa/3AeeHtBVEKN6OlfZ4sNvc2jjn9kRia0gJA/
DfCRslkFfhUCEJrWFtRRywLLm3FPfD+jTGtIUY5+BnoUjT3tqLnuhQ+/wpiWpCA8vT6XTzmgLTZp
R/YhfzJbXHDLx9mdX+QpzstUZsrV19hNPq6/V2heAoqvE5ja9J1Qw4iEK1DWy4z3kPYngT3MHNB/
qcBsj6AlQrxfKg0FkDtc8A0rHkKk/y/IKvzknNJIc8cPrvme54iox0vVDp77s/DiKR0OSJKHmW5v
Ndr1X0AluAY4gcpoRzLVlogr6USJodh1J/GEzGVrGl9eetEE98QmKTU5J+TrrV/hbcUmht0PiFdV
E++jrhi5aCo+Q+GC0AZ3IKIZhrqLoFEdOb/MKSZYjuC+lTXuR9a/uk1nZdu+FE4zJe6qJfKZEmzS
ontnWMAHDwL1tM2Wke33tcaSxZTmW2N42tG1XKy8ComQsXb1uI+QbWc+h87snu5N6GVLnhYmsPnv
QYl8KKWYOn2UeW8lpoB7gzoq1OFzLYI5+mC8EOC+uJ5GeIuuDtm1uIImqrn5mThz/cgRK18MLlu5
xbzJwinIf/sYZuhfKecZtPOT0zLpcQWRKoO3e28gfeJWvL0QaUS56NSgcPuCWD3V+RJrHuhyDo36
lrVbpDyXADC3xQEa+TImOY43V9jyL0UIfCN5qEPdYSJGyFZiikDB2JaIwkehVG7e2ndY8w6vovoO
sUOa/GYNxVrjgv1LvHwwDlcqazK8uDAxpGntyBt4ZnGRoY2HR8rJTUkPR3SR9DeVGvBe1/7yHo1+
gFCHD0v/uWjJHrv8m+zIQIC8KIwsow0zDEoM0yy50+H8zCsnn0Nxj62TRJ+sjljmvQRAgdhzyVLL
JkrduVWaKfsmHXpWaxhM8E4cSEmIEdXrktRv1veaXPi3ey5V1SCGbmacYRV3owkk/vLTKtgVkB+W
H7/xuR8WYNHlE6sPbxui8aj+r0wZn0J9TyJayCAJtdl58F/uoh8+hv9S2vbMaczH/ouDh+iVw32s
Jmp+XOrh5C3ihwaH6RkAObuIE2+iIaZtHJePttfbi893bNvlwYp0Oyc4XzrNLwMMY43QavmanaSM
3vqZOyIT8NHu7Ts7CxwOi+UqA0aNZBBVP8O6YVXJprhhZ1DdkC8L7aKsGMxoh734RQlUYeDVtjpT
93CyKWG6+JxL81nnkDzPhNwDjN8/SaPy7qiXdo5I5kSq9ZJSRXpKIQG7VOTzCYn27jnjdgOzKIZp
cD0h0mgFXnCV7YsGFFscDT8fhliy4oT2Us3h4hZ1MslqeKUYOesELbU42PlHxKB3WdrT21DuFbtu
8Rq0DfKXw/GiXBQZwCwUUHB46NvAdTP0hOkeWB8sH8sp/OW2m54Uo+llmPPqXbNMAJbat/v2lydv
+Yjg01j1BVVMPXwMxp0bH7//c8yVsKVNTqgpaVmYyI+uaFiK6hmpYApc5A7rAXeIJ8lYCRrOrtlV
ExaTGDQhJASIlWiZ+U0nBCapEJDI/JPiymDnyPZB7XwK4p0VjAqIJT0IHHrh6Z9OBK5nqCBII3o9
/Mu4F2N/+1bx0zcq9SiUhc1aiV3oHQDtaGjsLh7u3oGCE8B07GlYnSqFOm5wQfuT1JkOuYLRZXHI
lqHIfm3MJEWV43FhFy4BnJD3UOj6P1unu5ty6dMfFxWbbqBfsHA/m60t1R/MfZu2D1wAcnI37flU
R6RSr1R0NsigK0StN8TmM9ojX1fE5RYaWEkQa0CnWTaH+1uho3AVMbn4vEWUoxqkiO7bPuocW3/d
Wkv4b60n5pTVGZRZ8BzU0X4jxdHv82M9Jbv65OsT8+iM04NfR43/9Dgmizpm83ltqSAojtxTHEuj
SXe2GjGeaRO4h1voMaMRGTogouVnmY4maukTBrTRv1spc/01eKJ/b35cakOXVkmDGmeaD7prpj/M
aY3Bd3piOUyRI9bGgeCH3VPR7gwmrgEBNIqHYm/TNDKLdIZm+BDOfm7r8cWkW2+oN6WRb2Z/Yn4/
G9fA6mlBSUYlPlR5eryjD7EsvFgWh1+v4ywxFoeAipqVGEvoiU2Z4gbtpxzqeMlOqKtuhi23LOJV
vqFXJfNmRDNlOdNur6z5xRydjVKvrn0BFNJoY3mUr110c8tbH2BjVUWFhSV8Spn0d7A4TqgipWPu
i7ZGeyVSdYqiikzeQcvjHBskeoh4MYHVwEp+bIzqTYaqgzTnGTuyfoYEjKkZa7q73bfDdAU9JDTP
xuPgoeSxi1w2baR0JcYRCfwDoIXhmH7VTAt+VvMykZyyMtQgGBhzt06qIawfdkRip74P9h6Lz2ZN
kN2xCNw3ke5j33BJyIuXPUiMAFNO7qq4hL45QJ1sM4vMkftBBoczqgpewaokNawifK4rtedji0am
07FZJSpUnkdCSEHw/RKdtTKifW+dlbNF+3tuo2B2xKxs88QmH7Faq9Hmwtg6hUa6z87obp9PV/1Y
JUdat87jxl0D/Fa3UyoAoKg/Bggte0aolKtjOyY4wetff5eGwdrE3JEBJhT3Jp+lWmUJwi0Bpnru
AkNfxYrhAW7FKHACyfxGA8qfuus0Hafp0Tg1FB+Ne8niRjRC3JrmM/5hIU4Ds/JhVuVqa75JWmAu
Zu/JbcYePSP209T3LMu4JFNyms78EeMzUO4xpNkcaijCZcEnGjW/go526r469ptt6iuoMMFwuCWx
nBc1aTgYHPQcjpKs5hCluqZ6Q0rgGefAhHaokOYcDmUBdmab01baiYpgp/TboEL91ThL6pJvgy6X
o0PfUEGvzKOUydlJg0qy3fyCmeT/D6oXa5+YXoKQNc1dqQKAkae9ncZ9IxPZtaM21K1RjRihIp63
anC86uITMd8JcO1mjWQR8hFXwFvaxsmLW1aYP5mssdOE1R1mx4+9C2o2KUceQ2VeV4OgLyCGCJqf
CzIggy7qYQNbsCniG6fZvTlJF5e7a+Wz6AzWKiHV0TTJoRHJLZrjikIvs2Vgakw36IilGxxGLjXm
+clLplB3tiVU2dAViQN6P1K/N3eWFDLLPK4hpN7/z/XOIbfUE4bRGo3sXa8slbbtUXnfMJcjRkgT
pb0/TFG1qzoDKXOpxRkRVNiOUFXYsqVYZOZg2HlDvqpOux/GnXx1O1zwgMh5SrJ0DDdOtPKRC944
c7ZILlDxn5qfOuxzmsb1TlVf0wszkMtIB+MjGwWI9VlA3vy8YzqL/9gUsIqniKhFWHipJ/EjRacJ
pVQfvoFpsCFT1hCTrA3xSbgDpY2/FvpPEXqwkJaNO8Cbfi+h6tEFUK/AAPLnUyIQnszlNKPMiJFT
bkVQrU506S2/og+2iwk+D3mJs4+0tfmW63a5wylIlvblZs2CRAh6G+4//UZkwisBb2MQ/zDO4qLq
IVqHBG9kSU3sKLyCKjQpaceA2UjwOtQ0zKNp6LMpHeJSWnvyg8kOym4Q86CAw2ZoBSk1w5jLMByD
tHdoWwsDowFpr7CIAPa0GSG0ZqT+d2GegrlR/BoGayqVqObzVbyjeJzFs8W8m+cZk7nt+VXBWDIK
ci8VWP9+GJ2Qeezzioajx6GpKxr+LKeQxQwtRSHnMxeJ43Za1bOj8kwFvyPfYy1AlOyau6A3vsko
wKDBWyi9XgJ/4S3GHRW7UmZI5jDOPNFvNAytntgicZ36VFRy5RvOqON+hYmoFFtLYDlvE074BXPg
E3vwKh3Kc2ab4GKxRQ8y3wsKWLab+4xGSYTA4zLipCmAQFXphAIL3MtXmpwJJCJYpyPqucApv7mr
Dhm6z+rB+fA1D1VKitqdKZmPYembQLBvrBe+LzmpF0UhAl+Q+a9zn8XSHd9caKqdJyiafPltfguH
391QzljsfTAItz36RD65CiCEvwRE/RN0uVAGFsn76luob6ctSx2JR9SOpaw5cNK26HO7elfb5u+V
r/Byz0TAziPJ78L6ceNP8Gtihx9rreLw9Jx8d+QpJRMzzkKLswteO0V8n3LZd3iOaiw1vpnM6Y5z
VuN7jSxY2qKRsq5EF7hN4niihyyZBSIXbKoSh8tIxX1nsycJWOFEhXzzM4xrL58AgyRB7jtj4JsY
8dxd7aa9gIsoAslUJ2ChIJOokovG/VrXsFQdyh3Q0ypjCPYeXrifBV1PGESBQ5mvvQMZHDIsjJz2
d1TGlKbwBKLAa/qkMJUihtIQgdH2jtsLZOsw2Dr4SgRfOKt2Bgu2SGggwHscQYc/hL/UVCoWJEcu
AvM9VT4BP9R7nJFLEHgz1TTwcmG6P07GeihzPkqeBWQaL9rQm3AxG2Vf16jbdOsWdGTADpIqBW83
T2x/n8dh6GGzNymmU+FtjFBzF5icTALp32jlCpipWqtjC/PJRRgGFLLJdwIZtZKtr0TqASzQZxmG
8+0jM/1EUIoAtap44u5CQ+dDi9VDDWDAtMuP9DgE2DsA1MW07KrKeUDZn3ArxH4l0ZfUr8obBH3B
1gP/yekCFFnSZ4Xc1Vw1VbrwS8rWJDoAyMh2xt2Y55k2fdJlMxxkOBxJ1mvtoFU7dhM+clja6Dvf
LJXw9u3Avngf6LVj7Ca1xzTXdxQuRnDOLk+aURLuttBe/cVFfHCli4Vy3zwL/Cu6iD4jhWM5/SrW
NOFfqD1QkiNx8n8E6jieHt0S40sa72uMNLogqTv2OpgnikjsuYmZwQA81sZ8icSY4dj9hgL3mNop
xev0JLDYUeRdP2PNVJGyCLTOQZaPFUSfhP7PS/8NbdE8rP4SVbUvuiLbyvhVF/GvSwJspC46Z7Ub
wxq08vjjK7FmdMkNhxH9tyV0SMojO9wOsBX+CBOB5LXMHDSD5zGKQg/TpddlbDl6IUV4q4c8w/Gt
0AsbsytctAGoTXy05BWiV7n/i93SuvZXJgC2xXXAwZEDUUka0I3P3PWjxfj2RIFAbJ2WQ6L4xXVk
ILPwQozLELCIrdPoNbJxFgFxP4gRV77X2oRhhwlm6xnNd6ZnsVEYIsQ9rqOh+9MPoaKidWTYGpNs
wExxvRXZ3KdbzY6gyitiass6pYkRD0YrtQLFTrF+4Az6Pa7IcHrgeZ65WRLk73tKsUVdNBoRXHH/
0WGb6u8Q8DA55Ye3UceD/b8f6dfP9R6Ug8oLR04EHqLvPtPLyRZ6KhZ8wXdJsv0Atvk2HEB5MwmL
dxfek8DKVOS4IcwRCznJKKk8IKV1cv7eeh1zNhKN7HPpMVLoszIHGlJGE2nbI4oW1zO8QmGUjkSY
4UZuPPzwS3vnpgSpXjg5IOulylg9t+5JPs8yOCJ9doACY/Od9SEnR/uU7pmG1pYblp47KMceVxSA
tq6sxp/ut2YACsYxVrucvM+M3i05xfOIm/e6zhYcSh+3ZUYjYAeAA8zSTcM4Pv1Ijs2j0N5ohGEM
4/48bABUnrFluTqOWvMUrM8IPOajF14lYG2kV/0PVlvaBBn/CQHvTxbtLIc7SV0wwaa2jRIbY3eE
JMRk687JWbyhqqLF2OcU/yJW6LDTo4h9VtDiM1aLZ+2SXME2LQLdOT9xDY92gOWgWO/sQejf+eMn
qVoz0ALEXwPgc3u82KHZhb3VMBKHwawBuY/Ksz5dqXG0NwTSmlXl9Op0gu133DCHtn6L/EZKGd7q
JeHpJspfkateRtf4GhqhLzABrTELn1TQuUCX72KcNRn/eb6e/HcojStGSplLzWXzTqzi7XquCItr
xHPvSfDtPXZuGtUEImOFkkZL1b9qggxvJ6BSHqdcVWUSkwkRYYK5alrGb6CSxYu4vJfENR/5WRgf
bEKrpmyT9+e3JAW9J0baPwJMouR/yg327kV6a1q8HP8tqSZoIkAb7Hbl9A6szgYxluAar/X6zVkz
ap6WRExrfUtR4xVuo9v7QGiN0Oj4Fkvpx/QpUkxj6vL0uQ5EOhBLsXfNWp9GYXoqw0xPloR5aBv0
ERZifMcMYcCJsgm/Iyi9CR9M3yNxEAH2PSiXdnyQJ7aMg3JD9aILuontIE2eObT5KCW8Uov8gSrs
anRHEfNo0yPHdCK2JG0Oj63NzTksDQOlSonot/MW1GsxBouhIZTGujQR81tp57+QeplDlO8aDWGa
DlQWrJ4ykQIVn++Rio2cAU8rrJ/V9x8MjXQ4BBkO/gaKirCcfxlhtjXTsQHUXxZQqlAjNqXCI1zD
cusFR0X5abVm8rokD1t5Zbzers597YJCNd2hOUuuQFzZQ5/4R4G+buFOyA9wqVInTqbI2jAuYsXv
GHKc4/SzyA/Iw7DcBVf5qE+5IC0Gbgn+VKmr9LrttcjhGXg5QfXGaPprGOD918fzGSRfGEoR
`pragma protect end_protected
