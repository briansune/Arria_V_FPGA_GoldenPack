// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:26 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FY7vwLBWgVu8OyLchT4eD2/pArqYjaDnv1O1OP0Cs6XTv04yTYTcAcgD5OmHBi+b
vKiR60l6+f+tId9j1aKsZF7hUPbq58hEelWUozYxxTDh0x9jy8d6+SYYsemZc0JR
LxKbgHbOynbIdF/CJxj42qDDu/w3JYfp/rTrAwOtSFk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125456)
p/iQP+V67xjtTT2pNR+excSs+MOjqKzNMoOvYlR9AYPjja62qqqIlpZ3ZjvfPl+o
9PlNjVSy1dzw0udjDadtssPDMg5yTTEMOHq4Kh8vwkZe0xofGWe1grIu+XNQ3LEu
15OBR0tlgux+UPbzr9UwTeYSrVk3EF6uh/xrVrohBSNeNpvPf1w+6UrrEg6eKZEC
AMewcO0/n7JX+cxqkErlAI9LfrbieXPdEpa6c8uW2cgx7GzE6Dj4WqkxFqwT7p2f
1KNiHmc+j6VMo2e+16PEYXkke1Yv9EyJDQ2LVq8quLy8vWBYYlVBroBTbnOC7jiv
ZY053P33lS4U58VK+FCx+Pkjpj+7ZhrvfELGhrhkl2yl2wIagcL19+fYvFipPGLo
WtmGRlG8InAUcSmUYcP1/bw0rClvIcD+AN3Q2jIlqTpWTL7g+3uXBEeN0ROwEdLX
Ww2ePqzSuP9IU+XYIlnl8Y5ERH9TVvHP1aOe8PgGAFJT7BMo4OvOa6T470li2HCK
npun4vnG4a57koOUNj0wsmefX80cnQZsZMZ7EN3J4F4C3Mo3aWlILaLj5+uPczsL
3/x6KMIwbe1fEscqNIyMCVTNZBIMB6VfegOKti7eBP/RdvFU+7TcxlfZUprixbGf
+o8r2dSmQKd37kC1O6aTikhwrkDWIKh2i2/6B5vY8hVskRRt/fxIa+gOuoaqWqzo
qhHJ/f8QtLO1td9jDZn3CszqjD2f+nr6GXUrMMhnxsJvdQea1yriTXgdS6gcb49f
aL0ATg4JpYtTBpeIzp0cIYrFlv/VcPNLbM90dNbGsvU6dolMDIF/FjrzCOSAI+6I
3/4bSVKaoTa5sz9FvWDCdZsoJ77VurtdEb+rwpVlmrzO7Pwi1DIhHxR/yaaOmO6P
gt2vC4f+sK6U66tt503IJGcsZsDNld3P9zKxjYBNXmDAgBYh7mHTVFphAwt2hUAp
eSuhyIjt7Wo+lm6cgc/slI/E2uC/0TV+k4is3JHVhQMTOaBkkpyE2Q5nS1JqOrg/
6MLYtt1B5RPN15T1wRrzpM6zO8U51h/9kgJLhUi+i0Ylepb+IPWb+RNXxeY7lXsF
QkjHgRHSehM62MJxjWvWaDNC6S9bO+ygiwoGtk6WCtgWS2HR4u8eKKfmGGWOEJK/
7CfbwM3faYLlGqhsyLEEmf1Uv07E+/M3fl2g7ykMuf/EwIoaym7JIobTzEEo1n+L
V1ZztFAujXzbCnyAmZLJG69a3k2HS4ShiAFb4595c+zeMIHNS28IGUUxSWgqU4CB
unVSg0Ply+cuomALKjZ5dH0v9hUaNT57Pccb0S8OG4aoU2TmTujEVPoqH4VCRhQZ
yKhEoV5fCA04QG4JAJ4OnSATHmz2y5DBtsycw9kjOy679i7uo0m4/Qs49qWS1+S3
1V0Iu1m4c0Lja6RfrtgA1wngclRHagxbGyZ5FoNRIyORRpaxglaEIXNjyTNTU4gN
KTDaYtr72bJYgJ5EEnNUCwAfgkgWQ5vu5EfwRr1zFKJZZzVAA+cDvLgVdhaFqY6T
4CakTkvev1rJdG80TkZIvpvojNV3IWMzaB10PKq9iH4deeN9TQBHEmUwrr4Tuwzd
6plvDqDOGGVlllcg5u6EGdkC8HSNilRmXF+k0gTctHb/duH6LfQ7j8yKUYnL4hUN
GrSJrIDlw17nvpE4KG4RJ1eX0nbM4KD0aQsuuoSEGE8gDoRhUHMYclXqlFbLY+MQ
iZjEJyNzmU4E+CmNLmuyvkmtPT7bMRVB491qn4roJv7hEw0VBhzfOprVkHdcSVsd
wD+E3G16jV0Z6L89KmtZeoY5zdizc7ruQjmmMue0QzY6z9GKC0ohoMi7BS2kxbCs
XRH6CfOVlM0tka73Ynv7agWVQmaFF3QLXhZ0gG/Wp+3lCBpbRrOFsYgTrO50D532
94J8UCcJ5DW81qPVG0D4g3/mUMwkODbiObnloojlzfIP3NlN2GDkiw66qX32mBh7
9tWJ9dBg3Iu9+4xKBj0YU8j+IIDhzh+0s3xf/L2fMcRmz5rtxMMLbObAHSyCiBFD
92fpAQXnborr7dlpQjVngHbddIKxLGsXgNv3CmfXbRpUlnV3K+DJLDiLhvaawiET
e4IF772JKj9Ra2UlIUxFZ71WxqelkogX3wwKEs3JzOIUUDeEqfaLbLcei2cBlulj
cVFvd2kXnRWnCuoI4PNhpnPlJhiWfY618r3yrtHzJakpaZTrpKie4l8ttxDWQ5lM
QG9rq5O/GYdyym0uEs247vgkF+w60tNW+Euemb/35h/hTHiKlmYY7OatQxQyFCn8
yMZRomQUzRwvSt//d/wHAlU3Z0tMUaJZ5Iu0+n6IYwnAwNbuJcqGvZzN2L3+crOi
4q2XnzVsVWELNx82dQuKHgTtG1fIlQsrO80ESKvou+Ll3cCg9KrVkEG0nooc2sw1
+q88BMFwjwttnvPaG14g0bUwzmOzgtFB4zkuS1H4rqMudZ/sM2LROBqHhH97i1+e
zlBOUg4c9A1OgAWuamjofM/5mWppscPowyg0BjwnOZWNasFMEq6lRS7WL+MnKYWX
FxGXzpfyRGJW7ZZX3QDbkacBcFeP8IQlOsz4vy0oX5CLukxV150DE1l0JHy6+ExI
gUubD0N3WR+WCRVd21NjAztGxG8PwgMBEr31a2XTvufJprINGbnLOgYp7h+/L6rR
fY8roRXCB8vrGicm1vf0jgLW2lCTY4Sjv9Npikw1FDKJLUx9TXrg5pxOeEbps21I
tqkTk5MgS8h3+wONLzgGqGsEr+pO5EgfTDq6+4F1BcV/cwPfk5xc83aD6ZwBKk+o
pd4K68NzJHFABsfC12eySR+hAe458iQ87gBYLQKl1Lav3zmKoPGSWWAkGE50qa/w
meUYuGpI7jG5YNsuOjbln9IOzA0xhG1ASGtagG3nCinX58/6i56l90AKHIKYY9LE
HyLv9cfoErHhw1+h6bIWKTuljnhmVCoVWSfHkklYYMIRV8o2nBlnymZZn+hkYt7F
VoCBRL9LDfbd7nfbTspzpsB7vSSYECcSYgxg/+FxJt4ayLT7N42q8Z3Nav2x8Eki
92i6VYYH7CoUJOD9fYDZsdKADGJrcmA0rSU74N3z15L+P0JkKkvhRy67XTEuHJaG
zew3M4yaljShbZMG+uGxYl4/xJlefGwMBKZP3o8yEo7iL1BEheCZArrjM+CQ1JAy
CWhD4LMquAzJFvVcNaaKi/tx71uQKRdYVEzOPkbA6KY0k82JDijTvU/perHgGN8U
V31z8jn/8XJOK8P9SP8x3nOOOJyYdUnIdkmUSk7MzWr2Li/o/Je4uMr5YbmUTTJV
qTQxOaU1+ViEFOyN6Sr9sSjGBa92gsRadfb3bMXCs36vnqTofdAFhkpcD+NGIa11
ZjAyiwboKTqDBkWF8GhDHSnxu7WSsEdBzKOQMoCMC98zd57dUjWTw1p8C1WMi1qR
rZtexCJhVFBITtxpfp/q1fHzxcHJGI4IbZUUpHQPyevLUsyCGocmpe8jHhRPxrLy
aEeKzdqglfg6rscqNuMOMov1qtjADK1qP7btu9zGTAoDS3Rqo5vgI8Fmp/h51OgV
e85P0KFGHtXsXIUltC4cU/uSMIEwXA831llw3zIKNSgCUTZIwSeDeqyTVcj6/al5
yYaXKvTwY15dSgBIi2uK5jWciwwWlwZMFRL5aeEZVUjnIVcviH4ScF44OXWmL9R6
H6xXcz9LwjeuSoxLX792vMmNOL3u0GlJvEKH7OkGDKsJN4mOckH+YFVVyG1Y0a9L
wS2Tw8Dlz7P39nVXr0Dv1raxzn1r/wj6KS+JYRoEf+KgWleRVoXxf72MVt9DeXf6
vWh9KiuCUud5ORetpP4e6mC7u1kRfiEaO5d0ybT8/qc6DIZsERHGBYgPx1FinXq7
UaEaJG/b8MeIvv0Eb9TIPSrd88KZOv+Ey+gyC+hNyuJH75XXR/LRUlDIeU4n+0uP
28b72fcy5Q4zOz1ky2qNYolD9Bd+OOh3ukVnkISuKZkPL+qLv4vcz04WXuYnH+Pv
/zBooexWbR5uhp7uRkJkqVUyk9+x5VG0hKRKf1kbtgtJMfPVhdaidJV4+Jlqvz9u
fBTVz7J0eGVrCZn4QcSUGCqnqn8hqcvN96bGsvPXDnrZonzRyrnR3pCXCUnQPWwc
FZMkv38pEjaXgP0Gl/BxgyD6KLeg2rN23Sdls5xrTv1I1IjOKUVMRWXwCcu+o7zp
8O++jw+M5HkEIzuqJUVK/y1Ncpe7NMO0oxhK53WQs2unv2RMLbVd3/v6cSG62eKF
Sqd95elOoGXBXV+AaCHPQVllCy/YVIdKlNCmMmG7EfrkCxi7WcknAAnA+WK9PiS7
TNSoayrmEwgrTw6RTUMaLYY3gVC6jAjFTYpMUPSPIgwiYPL+B5nWz65ZbYx4eES+
2HIWHVco2R3E25Ai4o4MpEkK9tYJGhqlffKmiSlZSIytYcWo/0spIbxypESVpH10
1Cmaujcy5sRuiddMPjH7irLELIogc/LSqa7KePMLTA5oqCcPDUUoTwiDzPfwAt7n
icANQoYork3GeuryUveL50QTPdyvk8lvGC629T8dtVXApvNk/d+HIKOPWr/4vk06
/JRY+8BG0JoEIgi/CkhbXANB1PVfZRU6xOHxWS62Oh42tYG9UKNytNL4vJcBUagr
3c6RKGAh8uPkMtMztIF9B/xE140FJgjXAGB0lBkLQaaAtrPNJcb06S59KYc/nDam
g3MCeA6rvkzC9kOmG8H6g7aDowwGHXJxGn1L3i3gpAv1iJg0AhpfNtwy0nOTONx0
luTJtjNI0k+mwXtnQaQ7QCOYI02cWKsb1tRTNxLcSze2dEfgUbhKNIq+6yfC7tXL
aqQMBULLktRE0YOGCndh11Znc39zjIAPiEd1snjagHqzRMNjlURgbfxph/F/wOcY
JDa26xLjn4thwGGodt9QxYWrcwi+6zyyYr8dY5NmuIipbNJEywjuzaeENyDLnMaT
L/P0Tqxh3yETKHhoXZwjFnhFa+mvqaMA+Cj8lWF5jE1CDoAtEcnIBCNV+5F4buWJ
fvoYGYa11HzjoQ88wD3kKtSFVgNNQ+0i0s2jb7DLK9CD7H9236cB46LLh4ExA4ig
086wcaO6Y+fuS/jPNx5XxsW1ccn4rRKyYhg+yJh7AMj9bJLYvXdLQCxChcV8VuOa
akyXbIKoJiTymmxkGUh/+2mtXZWLkOfwwYCKZQEnymrYiQznXsr2l5GY3DB7TLOK
AS3IXs51IE+LLvqJKQZ3vQfc2xguFsAHaV3GtqRC18NUGOThsHopbKVwvF/1D5io
vweQDuJjC91AtTUaTAB/ShraMmgkj+dLaGJixeenA4OmIUWMHavya35pb9GbND9f
iNOEB3/hw5DZhBBZV/Sbw1fKuaK0aIP0Uwrh4AR6TZn1fT6oBQDdn7KNtyp7043+
kChXVIOg1bsUFTCfPl9geWthR1QLjt4opxDyyO88WN9meZh6axXzhDf5flyopFaP
HwlPBsFuR1nu6/GSf7+zouXY/cd+ukyXVE+lQpBjAEyL5AT0Q6rnNhv6TisD4n9f
/lcIowKvBz5zvjBpypPa7yit5TyeqTVA77Eos70w10xcuC96iHtl85Nngr+A3a8E
9lVx5DG39/Lkpfh19TRBV1qh7NQeVuqg+ju2hGIePZ/vx9Z+qT9fqCt10xplsMJh
Hm/Nro8QMDY2kBLSa79a5KG/erZGhIcgTwcGHqiQ+aW4oPSnqWJdBKKIhpg6IA0J
nQfjCzqNpr4EfWZvZWkI3rTaXczs5DemQvoOu4pMVxaGHUV9cc/3Qnzug4t5Ani2
REhCfFzfNunONhDXgKMH2SuTwAnfhnq0xvMfyqI/f6OxOdTGh0KQw72MVkxgMMr6
cc+YB46C1KlKyrmuvZKLUx5E+no2YPCvUENHXMDKXjQE4cQUpuJo4Edc8snWq23v
hyFMHmiwWUPtntJH9MKjbUoAyTWPccCTlgvgvdr3wgGjIp3I3bl4bIDC9DmHflBC
wFTbfRQARMtS/42ZXg/WP1WyMW0yjuDuryJkbsOsLIC6u+dtpSarjJE8Rs03b7nH
C679U+EJ7305b0IE+tO6oDON32NntCuxeI14h8+r4ienCYFMbsfzQtEZwtUuL4av
3djLIk/VuJGL2xgjtP88wtxIpOccYVXVHG8gFFe8SNGPW36TdiFmctXGIqQIVJxG
Fbx8x36TIVgvU4nocQiZ0fwhvFIilMe2WrcF3fcrYbXovnkcZLHwIc+q2UdEnjrT
ZQumF2fIpCrkoDtJwCff8tP1AhxwoUt4T43ysjZtqq0ZEXd+GVKXg0XkjwOYjYgb
0ZJjtRpDwDA2lKsVMrijrsQ3e/xCDW3Ag4GIxa/oqfK/YewPDNjoPBVXuox3qdfP
AssHxVZNsbsBdhzBDrqHdg9ZQ3PQ1R4yN5sbaBxVUD/XCLIJtRVr/EG3gxO80c2Y
izwwWX8XHFWoxZwO9l75ZK3ief3KIaJW8JIUdubvQD6UMP1/IVwe1HzMNv8/lFzx
ilLVBv85/d5mRJ1DQrO+dmnMM/KiOlOtTaBjaOrZ2GjwB6FmzdrH7ezdDE9RmKaK
RXpksXkIqcoY99SPCrYZMODHLKQjyxRpLn7vBLSEYza3hr86brg/rzlCTmysWZBG
Iw7UaMAHP7GMfZiBPtiad+RzFyzeuh1SlrOQjzgrkBPWwfBS+MtOa+I0Ve6rhGXL
Q93NWbNhf/kHuRwUyCBfMSujoZJlWO6VmytKMCQ7KH0iPXq6WTQQsGk1QrUI9Gtd
lw4yvjcagBs0XiszOnQl6JpTtiGfInPzl16pIsgGzdBN7m9xFQnGlY/pLKVfRjWc
MDfwJ5qWTXdM8r1Y9bRICAdEteO3YZvvvInSoI+vb0HHXFJ6zz0Uw2M4MJwkvrlT
3fUB4mH9yOkp2/rQOD9PNit2tnDvmR1zewHYRRUjXReBV1B457mf4iGmkcwuN0Mz
8T+ngMorzPNqwhq+nfC+wf3mGCj/G+o58vZK95UW5yli5vBAPmLSiLecxi8q7DDR
8yoUVSHah9+w2+sFYHsJqbyGS6jppRgzdej2KcvtXRbiqSLUYc3keCTozciqeAEw
g8N40mJNlA6LyXGjiMxW2vdiGmRFDywx/pzCmqM2NDSij+av41LQfse1GYINOTeU
5cTCGckdwMJLXsFjs4H3w+m9scQyCDY3fCUs7vn3hKetUIlAO31XuYICOEsjNn03
3w/vAmQLiYWvEf3vt8Tw1mAXExDS+F1OpsNX6rtcrQ5M5J43XUA0IgxqOpU6v7xd
G2FEoPRb8D14l7ED0azaxYe5GfjkDeWqo4G+HgIWuVyHme4+D52KQ0/j1Ng/4C5l
MO4zyy8boUHgLq4zrWRgZgQtYL3KTyRe5YP6KxqTWhl2TSwGF7gYw1ceh+iRXf/b
CExww2cyKf0IsHiKaAc9zt0HSYAf+fmLcJhLl5ea8IB8tui0TqfWVcwrE8AEaz17
cHRJhFqoV3ZIvY6JfZnCZz2tU35AB/2ydq8rXuFRJKOBIeq4DgQs0zYVpEf71f8r
1SXBufp9Wka2vhsLJHAORFqIr2fIZcheoYfQZvVbM50N0/flxO3B4y7kPqlNIOdb
PIrNTOvAl7MXnpcIMbk749rD+B8hLPLb/mcRMmluOxVtLmPb67adaluv24I+u59e
igEUZDhYU9VEaLchgSFTLqAhGJtKcnRqrTvfNlbDm+xzPplpWJFOr0MeDmBWjFJ0
9lIuKT90E5e6MDxQYprIy/bQb8hwq8PVwd57I65V6DsOpIqCuzghJhr0sFZ6N31l
uoFja8nGj15D5Ayphzb1w2X5Yva3aZYdzWitNKqRyTfTw6gvyd1Rr806BaTTEa8o
VW4JgtYb0QroWwslTTTY9Ys82I0EfaeFnhrBbFoa0XLCdiDllN165F7CovEBYncH
GgIJRTnASx2Aqkbn9bS0AO9DD5E6k6It3LJiH5LKPy8/mmkTpqbB8Vq2czXwpnJv
23a2gUk6rDUTQb1nYtv3e70HpERv1xIoWG0JILeipHVsg5ItGxyLSRM3SAzumsi0
X0fkuzO2SgRj63uid95n5RcCalC0UQauHeNRH/HEjTnYYUuVgxg7z/L5R1iuJpw8
XWNBvW6TFcCKw9urqGu/NjRIYJH9pfKW7+3DRy8KAeTolVP1vR1p5ZlUtUaemb+4
7CPHo8hqZ2uxwNBNwVJgUMSNZmYyzObZFTKPBGzXtNBTKwjxb1dJjyPTFdNWZD2N
qgAfNQvuctodP/HQkD13ctFUfyr2gi37JWISeg6XBB+gej6YNodW22sbUu7J5dZ1
tPGasMdWIoW02QPBOReSQZ8D7mAp4mHpJ2FmcMdRbKgwD1FIvtohJ6KUr4OQVG7I
hX3GlEuNIYZKUO6aha8dOEg4aqxe4TRIsGBkElmiz1FjIYeuQ4NoDlfhQdKAXuv6
jH2jrV3bOLuyE8+J3bAmpaLG+pPEbBRPKbwDMXq8rW8z1aSohSCTM7v+ct5NjohL
Fha/qDO5YZaoOvZo+FjiJV2EZc4A5l56HkyZrMN4ajGQLNtXrwqjPHr6dJ59vtjy
T6MixxNjw3oM+iHMErhh/M3oSHIzFxuveqk7Oz8CT/ZeNVCzMM1BV8/wklpSxToX
BvhKxt/T97NJLJYcVVl3azT1cPy9uMwW1UlvGYk1+k8bhl24H7ZBC2Oxko6Qq1HN
S3y1LF+OE3U2Re+OeVe0pfhiumdlxMx6/b3/qQi3QUyEvKy3cJQSutHDWnZqYp/s
ZMQAXE8+ocvqfzCBc5jI0Xgj6Gqh/JKE2FWUXmoIxs/CYq688/KRfqazIwesDo/g
XFVF7FeSQfVC4DM6XNYHBf0InTPIucj3SzNbxkFjFEeuV8bzLdurkfojsTPIxThH
NLH4YzTV0+oE/czNJXWh4WXR5+T8ePyGw3WeVLD2rLGfxZUO+p8EyowiEEnpqq43
lZNW7sWDCONJ/mdArINHnsQIblvMXLkMKBXTjVXrPhj6tUdcJHTWBpBXdCUUEbYQ
/74A78eiV+NK9FjLc//DofxSQTEUMK1D+Aqjd96m7BVaImrHlytjb9kjfAOo2p+b
nC5UA5HzhnH1xjxy0bRL/RoA3lVGqRtC/lOLj7Uon87vvCZYpUxYH4dIjG+n9vfU
TUTgXDGLuyGkU13I9SW7yfL5Pkf7tzi4KteSyTUoP3KRslctyskwY7zgPpP1MFxc
T9P40nYUrZ2r26FhdJHH2lTx51qZMvRs+vINTcfdjp92ez0zGMh+nrAfl3ivcIlP
EjpyMmU/YBcc7oK/T3bHe2fBENsi5eYJH5s/nqwpKhg8CXbvW+hpn6HdLfOEsmyV
8D0QQ8Yp8gA3nQTjIRBjIesEu2rMjZQkl3MfBDPPbO9Bjf3UQ5SvaM4LH/umFASP
ltRxWNGW5fHKUlW2HU86k2fCXqZ64Ww7Qitho8y2LB9K5hLmtVo39ZvEWwEMUwtw
S/11OyXZTwQZuiyMyjbOmgCflVWJgMFFLWr6lHGHE15WwwE4gWjec4jn9tQrD2Ny
6XyRgPHYcPEqGwvmsNuKDdmvaygEcXGNXpM0qknWkYurG3XZ5X9+giFdXXWdOgG+
JCGZSi0rYcVoXx4h2Flt8baIQlbuR2twuT/A2s7UPjqXM0Dgw5uAT8vt9csculuC
FCwlEx2O/CPCIR+R02FRq1suIIfml/btBm6UWwUySngh666gEWZR0EtY8UTAuzv/
EQQLHSgIq131qWihKvLG6pVFuXgGgq1s7s7ucr/MBSh3UkHNHMFTryAxYSkaeaoR
McS5J7cabyDR+mCQ6s6yxSzx2Nho0MwXW1zCcOe6r31/GcZezDVsUR6Ua9yjihbQ
H51meQfJ+9bS2qEcgTq0rvrr5FEQIa1iCClPcwE8dGoZtUvPbt3HPQ3aKtbLYuXq
HS1LA1NHABT9XyQg4P7eSFzPDEr01mCyrw6GmkTbboR0YZI3ip7qcWMdUzgqDjSB
bt5D3ry9IJEWb4v+IWxRs7cYxFZVUJhtjuakWVnMrgKbRZa33JU+ZXe1m80Lae9s
7Vy6KLTEs7o3MMPkPkHnRmTyZ5/PQDp1CbCA5O8TSUjIfivnkvRXaxS1sjUiqNpr
B0QKBzf168e6nbdswF+VqzYML33fR9yokLeKAK2C1ViJhuNxiQ2rS6FhKWGbZ2cm
CdjbuLav3RzYMZA5tsz1qg8cp8xKRHlgYZZ2mx9B+14v/mlv+3eVKOOSZi2l1kww
XgcNIvZ1RN6hZjA+IjuuZu1pdKfoMg6IpRC4WTmtA//d1Kwk0FVnQJ95djI1KrxB
+tuAV68HCbKtWymsNfDRct5aXz1hznnfR6DvaJJAgKS6jsqdjtZbTG7qyGAIn20l
WtNmktvlLna3Vt9XmSTVwGo2gLjJnDu7zi2jhsYTXUTuAL1Qz66U3d6r95T9phYY
9UBXS59yyaN5wL5QF+TNuJV/zirEbMvFnliRuSBhiYd7n9e4ohlFhT/7bgamUfPF
VmYmeViuTqpDgCTLQEme/xXXet129to8ZODJsj8hk+Yq5YGFZ0Wh4jzsVxrbagVn
IQWw6lJFj3nq4HtQ2IE4vWAWD2PbG02x+WJvKLZPSRCS7o7NHtFCM6mC9ylInwPU
WejXzHH9OUsnHI4m2XmST1zueKlBHgRmlhcGZLjvvBmNkeqX++WSYjU59EKZ2biV
18vzVjvbmn1AM3iy/zO+UYWkwGWF64FgQ5R4q2k+6Xk8RHA+FfCBp4vpzcsfiyC9
tzrMMaP3i+n+pjko2hPxYILdAbWhCEUfBS5DstUcU+VVGattzDauiPFaI8D5SB18
HHzi4sOkRCp88pvIBTwevF591MDdXriTkXfG+cUnuKhsxf8CK1FYhCOs4hWjCExW
ENDi9hs6cAWK19kH40EuujhSjjbKHwjTqEmuehGsfdy+pO1fVIBZ2lJRFS0nZyWy
NDWa5W/RGCpMKcQtAzTtQ9+1pgY/Q7sMO7xJOt+rDrha9gIySY36/XnPHE0yNTs/
mHccVMCv7zOUKTbH+nOp1xfOf9bXTi1OfufoJB+jmsdS7lhBm0jmF4QafnwX4Swz
5dmsgqF7XoJmtaIWTmBAUAqld9v5z0VqBhBa3V7ZNTXFFW7/P9CTytw2pvhL6+/l
8w8y9sa8kHQxZJ6vgBkoy51y/SzyiU/GoZEEsYQicSSHu14uk2h9rXfd0/aoc02w
lraQg0rl/KDB9xfZslT9xsw52qzgFHOfpGjPXA5oENg+3Fp7y2yD4jUlNUEcuSE2
UZNPwMXQDTLsFe9ExT0sVgkrhUKWItThfUmufSg3gys5+po13fOrPn3prtwKbgBx
5gEN7yIZ8CJQ1ML9+Y2nb0YnwUGlXFe5Lqu5f0ooxj+qauJFVFkU0m7BphBWxRyY
8yZ45YNI40UeI8QzEFYIqnocUYcoABvMFPsgd1yBBFVSi219mO74SE0KZKB2b6ya
jpTApEg3KM0JdZoPAzKFlld4/46LZd0VAr0mxcBHVKfFjO0XmlU3ph3IDfIQom9b
wEdo1yEOjthFFYt8zDrUFEJs2PW1IfpHTmSrOjXcQsTkiKopHbUP0h7EKVux7vwj
5druK6WGo3MbUNs011OTpshsikBRESM2yCDZHYlz6OhNhEzvaCVjIK4tvHqIUWBB
cAPG4AfxBxSfoxUXNfKHoe8/Wuby60R20Hjh7EjPpcpNSMogbleX46d2bKEL2Icq
6jdW1rZJUasHm4fNVHnPqDw0ifrqZoyYjwY3SuIH8Ne12LD9L+B8aBZTuM0P+ZUh
VQYTAGt+GUx5bCftA8YaP0ZQLq5VfIaAss0knXULYcFNu0XmnkPnAnvyQ++Nkdus
E57d/6AAPBHAjlVpfEWe9QfyM6BDuEUc29R75Sz/8fZvq6myOjeUFRk8O4PyJZF9
cKnZTmc9kKhPzZ41lLULnDZNTWS6etL/QgYSN0d74kasDA+igbtZzSQPzVVWuZ9O
/e4GG6Zoz7nLH/jCsHGmI2+9VI3LlfeL8hWMDYYJqdx3MReKm9tF2hzEyEDSa1t3
LT4p2CslslazezUdXOTFLh5lT/xrBd1tpDkUh6nPwX0KhLGFfrm390aGJDe9PARU
E5ThUET0BfI1vZGM1kG3uBMHcOnfLeAAlpJAdIlG6rhFOcq7zlHzGO1oQ2cnykZM
jDlcq7BeV8Nr/6Uh+wRZBz1sc/D541jjUpiPuHMSEFYU5am0pljBWWXEKCo3Jh86
ebjjd5jis7uR7cIDosnijFqj0/ZyalEST0NPJT8j6cfrKisIIN93t4InAx/7YnNo
6iaCENz/CNocVQwpkGOxGNYnwgKCttZcsCYp7yzM+eQkO8gb23ffcFD9awpHl8SV
bF7De7zyPms7/2Jy7dDQ5rGdPka1Oo13Z86L6YYcxk+TXAh7Mt8WZyQPLxviIO48
keM8AKn5LAYTV3LmdKXQCbJasf1oPdShQpweXWOtjeuGMrE7dT6BObXlvoyGXO9V
8En3pe6GnD0cL9voFWL3Y6UhfxOInqo0fYbT3s59m9jlHxLtYZMrH2uPP0pAqxHl
PHMYe5MV9PgmpOo5+zQwdpqgk9SJBJ3Dz+/my2AeXXpcPLM8fApeVbTuNFDoeeCc
T/3e8vlIQUDa6pq+fVd0cXv+bsuh+xVWS3OlaFTZSrcf53e8cK0U56Q/+GZxDyRL
MLk15z3maAaN1ZtuqEkH0qAVMkUiHuSYduBtpxNOCr2rVyse9eR+dLgEugWUj7SZ
XXb6doG+hFN7+wnryswgGThqwEOJmLhyMFX6RuGIyYx4uChjhW4ZDx7OVigO5hf0
R5Q7DIqNpAub11FivMWH+s3dZhATcUBuF+Hvknd3JmfXuiJeBYxVPxjSYEyV71Fz
hJDx4ZiwLNLkGDV54jwfneArOBUFBUzv52OqjryFbknIcwtWrueTvUNxSghLMlcL
i53loohN7FkQ0deJVtA6d5qFfUfDc9Sz84kALnY120P3zywwJghvi9pD/OkCCtsO
7n5lLH3nSwJAC8cQhXYwwWK89LzH53PWrj2uDDrPMoR5JowfbIg6BcWJSH5U+FR8
c//HW0HbyaUingf+zlPFbr+U6IQ34BybGv/DfDBBxiHrvjYX1kBa72EAY8PAiRR5
r2IVE1OTzEmf+WKlOifLCyPb7Y0u+mtU/msGShOfUb1Zb67erv+VopmxPHMWRYpW
I1Gzm0UD+K0WZ7hNK0uPQds9DSxqnGPgBuK991jJRXZBE9oOyPWPropYxAI656Fe
ZqQAjOOODvBHt/6sHUd2cpQpc8UF30xf8xH4ENODCmKcD/efOggxR0dTTo6uEE/9
/pc3E4KXH2IhKXoUcyAsAT6WAB34S/e1NYiAkl6W+jhSVUic4A7xNM48xMHInVgw
Sm8ZJYfszgnlKtJU22rMBujvDI2pFgKYayNQBnx+N8AayaByi6g/cyt+20Es74Re
tixORYhaiSEYNizp+PjvB/PrXQ+6ksx9IJ3hJ5udD5Ex9xbiCljNy8977hxyBUvc
zPrFQAjci3MPrmDEmNI+cdq8bPnUVwCNtZbElBNMAhJgWWpw0GovbcHFfW/QOtqG
5COdq0Mw/ep5pOXXAs8qrzGlcOTjDvT/W9LCzSIaI896T8roYy1rhnvGHimhnZMQ
QBcnmAPRJndMsZVPMGO1z7zPAPZrDc+Ck8fhYJOuT/c67LRIUp5uRBBg6AU0Zesd
2fmVc4KVpD8BYjG4VBIFkCxMXpLnYePDxl44sfY5K/qNbDujsDx3TXcPZl93LMYM
hSWvraiMkMW6/vBXTHg92gFhZe2L1OogQyUm/bHo4I2nWZjIxjEx12SNtNlh8UGa
zHJYpDt7lkjrHMSxruPV/eqk6CSjxd4s+N/HeBNbQEi58l/JA5jHaTSh2Z9LpKJ/
tO/xOh5zpSKRWYCFHuC4AdkGHAyQsJmgzwmxU5OXwoxUS7my1tvBvv1ZoStdIlOd
UV6VkEaFu6adULKQCBximuCudaqU1yNmOveRcCQEmhKanooLYeIyfljmjW4PSfJB
nevjJkoWh8TRYKqbGgCLpElpIeaPymMgrXcE/TV31h9Qe19s/lsupt8cAJBy1KeB
OInjD273U15wDVLb1fkGJ712WOVir9ZkCFA6ULtLnefLOViQZYFK9CPz1Y9CZteC
i17MvrF2nwRCdKNweY8BIxDsPJZG3+Ky8VKoe+GHltZYgpLvj21BTMcK6WWTchBx
nSLkuWqh69zVmVvX9BWqv7S9G5+cb6z9o+CNaGX0ViQnUNjmbpGDhjCbxb1DBGjd
474MTfcqXlvUnrnXlr15RMYLzNjjTE4A5QElf4+WwnHIRSKXRPTJ7La3C+JP7Eas
N8alUeSZe6+4Gtr8n7AHBNZtd0BCH9ATcQ6SIZSbaWZtAOFHOFLKXzB6ltgIdCae
BI6S+kkOCkgCWxfsZfkZhQRCT2YY/IXcr/UHA3SPzvfaxEbEwpOVp6u+afghRBY6
F/+BwM7wW7TpY3lrjXUTu05EfD2yvKwaVFuwjLJWAeap8aK8/ISDBj84Yhre/Kmt
2p1GzbolGnuyc6Zx2WvNmqETBuLb4oIP5RbY3iuG0xm/0qy2voRtqoR6n+h9RHGS
bSQGunD9f5/lq8nz3q7w5j5O0T5HFv/f6rpetDC0rhikBgCCymcqnfQYI7nrr5qy
onkwQsek1RLLt/n+urusRNF7ClMkGw6evYFnA041zYhHjeOrbBP+uwfCDMy5SJzW
1cOjvk+eJTe/bhdWzPNQfBeykj9fGUEVPIMYGX3gqxp+DABGWneKS64cRoAXrJJw
nW3zS3oFPfT7yh+r0WKW6UJ1ozus8NPCeOXE07rbW4nIEsEfBoG7vKSJK7ntGBNB
9nPCkhn2iB+WKQcxd57XSdReLAULVntagofIs8hYEhVxb/gW2X6RWeQRnVYBrqwx
/H3oRlPwsLExBdCOcHrRRw7NNLqW0NWX1mAL6PhP2sYMiLUGFA89kV0MIAg48YWl
YKcumy/vh58wJaQ89slwv0va8uO3Dp6t8azAwhyqQsmdFD5vXSXMTF1ylsi7WgK5
GQ8gCuS4Vpwo4iZu6O8S6KwSXA7D1mVMZuw0s/35FfISZEBPknBcpJJF5bFq7ruU
S/Xzq7+dd24OR/cLnSjyw4P/LqMqUA49LsONNEBo6rdCLSq5Pm2EjByhD3vvPFIY
40YCJcvW/zVoV5PcOutkbN3Z5OtTPEMrOXJTng28DbEEt+X1kjA96gJee5hIPZbR
bM63aHK6FvlTbfmfYFX8ZGaHHEc6JWfqP4HB64FYoCcqybKQPvtbOnVp4yzQ5CHS
aiY90Y9DaD5q1QKaJtsil9ajhEg9u3w/DPAsKItWi8qDjM/fLGjrEUJB68tDEA2U
vqSM5YkhFk1EiqxQNtu8orY9kDwL+ktRMR8HxinEl3D+qyi4W2PpO7gQLHT7F7Ab
D7rDmcSMru5/BrRgx/a4NZ35uDvY0J2tc49U+5tA3H63v03oMyOuwt2f7ITz/fU8
R3C835on+FAsyRAT3iYm74yO9kiAyiuGU//hPUDv5UQH8NjaVcGIDAj7OOevX86t
TSXkw7e/+ft1Xz4hfCadCJUFp6fMZ8GqIJ2Twu8ic7TVtH5LgQ28RxNf8s1O6F86
T3MDZ8r+fXf+MlC5/uz5O2Cvlxgm5IX0NSm2arKTm8rv5OwIO7oBLelK9sFEXmQy
CSG1sYDIvAGJN73jDg3J/K39GQE9JVXwB4bmlDO+mlYdlCGnZ+YEtTpIGTm3OCKC
fAZXk6AgGOlcTVCq4DkdKcND6ZYvqxtZFsZbGumdysRafDQZ0TGGbhpCG23z8f2X
oFwEALWI6NfTaGe02t1FSEW2oJwNt44+kLPRVU9AbIFDsNwtgBSMS9fSobwEMdg9
7VAc2F/MH7yiFMWRHsSyRr6SxD0egGCTebQqIiWRT9PGENkyGUN8f0e3CG/YMQWq
pBEgs0rsQ1nx8L7rId64MUQkqDb8Oh0XnGLLts5wKqrUPPINhqUXi5NTyp/slvg+
HRC+tm2bqPGsRPOKafZixAIBUMXR+JMj1BAgYBTqSkC+0S1yXPGNiarr8rWFU38G
4U7PpDh+832RxdQrqvvg3Pd4Uu0DhQzT5ib/kkDrp7l9pmeE0G0v8chTlqHBHDKv
dw6Ydd7POAkPAWfj10+gsWrWqCHDGn9AXfHjgk+5p9rpo+JCFKKL4uMbgWD2g161
doBu5GNwiBBbb3hE2EeoY72ZZ4VSa1TpZqQYfFOi32xQQi9PL2jq+zvnkDnA2877
ef860kMzcdIVDEQ7ep8XyRJlUh00e1ybfbOBudYrzR0MYAjFM9bMgacv+E2OPRmc
ceaKpGpaS11TNO1y0Y68IIyu42z/sRQNbCh1NeWh2X/Vy1uxmNgfMJN4p/86Nhrr
TH/yKCD2xNmHt8RnhhsXlSmozTSEzt83T6ryLR6GTACNq/5bIsMnLSpW+1crOMx6
SGIgs3o4h4HtxVxd7gbIOXiLu5n5FYTXJ4osPGyaQk6EMTi5ZJIKVacsqENOHlBi
F+pffiow7DeE9FF/aSjRq39ueAEo0ux0P5P9F0FifDnsnidO8Kvs0WyvaLnpXBn1
axF8cx2OhEo1alEVMKF7NIM2vvWTH86Tf2/qZ8ccI7SaoeZNT/QzNmDImu37vepj
11O68JR7e128xvl46zAUxXZx5uSnCrBFvVDwjte+PMAlii6CPeunXE/QurBzPG3V
bNhSXAidGOKy7ZOcgiwH+1x82kSUcDjSlQIMGA7f8LXjIAiga88f5xYrnJsIgrsV
YVYF26u2kX9H6UuGLIj7+mXHR9ybFeWLa5BaCyNZ71K+wp8HW8vvG65lO7eZIaM7
1NFvgh4CBTBmdpMa/XnT2UuzbaAispNvP5WGHRitFd5jo+mKYMlGUnv0pDHu3bgj
jkoF01PTgk+Qh87xjXll8int3o4DMcUunU9C9uJIqOpXyaLxDhJTRc2GXr0onudZ
mrOzw2Wq47hfr2K0onXL+fLieYSqe2AqhpRpUAZz0KO/WFqN2tSRhGfVIG2qnP+r
TgLJojUnYzXXmVtONeKfQ++23uvAeCLfjFlrKwOpulwaazYQg64AU0UINJMtQlma
3UUuSSI9omsg8+kbrTXxoCSH0sdNJny6elxf4L4dqbTA1s/PWvbbYVmM6osYdBpj
iuT/+wGbJ2jdp7ijdMHntZEwWmTSgjG4+OmPGSRQum0cSg2aomSk/UbKcCLOKygf
+xCVoQF94EGDJsPc7rLZlcRrNKZQgl4X8M9ohnNc/NuF3MLPBbZf1byMyii5Xl25
IKg8e7FOnVi3eydSxAVj5LMNLbIGWT9PBPFWes4kNl60YZB45a4DQBOYIUAhXkhq
t5NdUifhkJdyknDIIW4MuhSxF+b4+mzCh8UgSgxY8m7Fo0NC0IK33isBB79ga0oh
g0eBszxlYHNwK7K4ZvxyX/asozi/EzlowRwTmCvMc0hjOtcQnPdk5R7Zxvj5Zyg9
0XdJ/9slFBrS2P//A2hkHnK1qSHxk1YHPXxVmWeCFNIqvy79zCSIyFHQZ0Iy53rT
afUtPgI2zsA6ma7s+KsnUwKQTE+0CVDXc3n25HTrCO9vV8JmDH7DwJE9AY70BDFg
v+5t75uLBncV1mO6ecuYZAevSfn4s5j5SrXJpB2j2pM7JS3LheYnLyqmlLYy8Wo/
wQWaixAuI8mqD0CkpaSEPNzbM6MIELvFHMSxCNqP6h9iuf1AppJYsNfHIW/VcQFw
6j3pP2DYsL4Bu8Urw7D1EFa/wvxQDgOqcFhuWrccoH7utcn3VtEFwltIRr6iPOWy
Bb4kGgqaFbJoXVQVpeTLtbamBFpjETHEzNYPOogFXSZRqX5u2YUMheR/YHvji7vx
zfW5f3C0tqZLAbMe7oaQzfYp2XvoS0x2HxN6/Xob9JhwZrkeSOPnwEP3cub4w9nO
2Ae0cPJw3hUYWCO/MlYMuf3eN4b9x/SNe4DOD6QcD+dCh6HWemD9mvx7dZGiOSSP
gmkTYAUJFEPAIowckNZwEiOSgqk2LPGL0/XHJjqteeDBqJbxo2r+5c8HVx/TCpNU
3wSAqr3rrJgWaLMHL9xCI6Fh6uJNrRoeUIb9XQK9j8i+bGkt0QEwQh4XOAN714lj
Gy0YlO+NJMk9ORIQh7OJLA8ZW6f4xs+PNwLxxhIsrURM0XFwvadlD9eqGu2y6OpZ
OaoXFW/rW4IiWLrhXVj14xZHkUaTyCKybNA6sIdP1CN6mZ4HmlZg6lr1mi64IEWJ
YkPQTR4g4udGYa9TspCi9FFZgjQBzuycPJwr4ZXEoVqDut3sGx2dW9OyIRzmsqRj
qRa23PM2VnXHt4GFW69DXT9cjxgVVwCKhd+3oEycExUfIvupEkEcPiyP6K7KQktO
Py/dVVv2eaYG6DUwUxiaZ8Tk62+NmsOCyq4Dngg0nC4UybXWly0kj2VopW1PJA9r
/zTcR+hupZ938SajwoBat20WVmQicH0+8RalKDZVwUEpbc0V39M1AOTbuCJUQpF4
g114rr784p0Kur+Rp3i1xkPK5TcMLfb12lKSoF+JI6uPLOeYAyFNjD9/tXagD6Tv
Jv48v+6f3Wy7MvACBfnzswP5kjmSlpUqL9vcX4G9XSFrxeZ+YnkKcW4Ps20i9uC0
N9uYDS1nYrbrWDsmyodCUTgkeav4ZUd4ibb1q9CeYBxL+9H9CqcdnuEk6z9bR5bG
h8gxLwD49j7Y0d/IlnJVBcezlGyv8semNanL1HZi/DvhlfBiwzIc/55SOIRLRMdP
W49SSIaACGWxjqHG1njBmIG/fPIEdk5pQ+ByBk+3HdmiVOb3PqWOpnvrCkXYrv3L
PGbTPA2DexN2pKO3Ykfekp86ZqEPbarwiIpDJ/yzD5itkMHsIYoufa8ROsIrOwXj
gWsk84dtn3NoGalNu1aEgI+SAbm7V9jnL9I/N/14dkdeFMIaA93kVIhYcdvLlY5T
Xrj4c6NyPDrnJRFwCRlR4bps3ZlMuytQr+Pmo2J1xn/Wp64aKc9GcZ8uNFpSzE0y
9DME7Fq3kj3slHbLLGNrqZ/1x6A5dqdHaCns3aAWaOH8AZ7+G1N9TKWXGuewy4S1
llozfpQERR28NKdWeRV4TbXNLVPyqWBzPvBxqIn5r/e5671r9i6ic+wFKRPH+rdn
Mc67UEG7FZzt52SkZ3sJx1lyjUlHRR3Zgo2Qjb29gUdUpxLVHzgW82YcgN2Hym6h
0ii0f4HSxy4yhP4n0XfWK9yiVcaOCMgdyl2D/RaW96SHTWGTgMBSgd7rjFEB1tEx
NusCutx6K/h+fyOzL0bJemoPEfhYY7FAvGFxwJSLj/9kFnc40GXfpz00239Hz11b
g13HzAyk0X+Oej72vf65LS3jMHcnrBJ4bIMV4+QKALtiD6zMhvUR4mSiW9tj9Jwd
U8I+OAi3NV0yRI7jnBzYiotOLEgABo1uhkAmNvhaISL18iKZi1Su58DT4f4lOCrq
vRdDvRE/PAdK/RoYZmBMCQG+Ql/yxK2j6u7ZO/jHxUbr8J37DZkD7Htkg2U6F6Gp
9wZB+ZWHAl3IVbjbLCGVS7oKBq0QWSdY7OKH9ztrD5jEuhq9vz4EIIGXkfqLPFQj
64OFZLEz4zb1v5IWCIeYAU42aw9NzITc19SkLZ+CBpqAD23F5EgeYn3pykSHs2fA
wLlEd+9cZkPuB8E0cMrXWz1C1e1Iljwbs6z+PRv4aFxYSW/+hYN3zA5Jxj7uSLax
DyU/SkBM9T4AJxFPFsogFNhKF56nyXoATajOHNwpKuPsjh9uJsEIC7rP9FFOJE5n
IvHfzssst1jI0J86utIH6wED3jzAuUgQgfZvxSk1fzkcjXmEsvqD4IbvMAIgxdN9
2aPamuJlvLXOkkJuwi95ToPSlVqwPjRgW0GnuZziFvyNVWqpT8rQcuIM1QpqQnj9
IcpcY/pp2SUThtS7ek9LRoFupDHaHxArohw0J9iLrhA+NNRxdJQAIb142ysLXyqb
XgWCByyCEBtCyBAtTeGef3l0RnNsPbGCvsJpJbjykdNOXtJ7WM2Lwqkk4P7nqlE8
jMA7pLoWM7gOs5eTSWNPLdv4SX1Lze3ITd32Nldzr/B6KrKIZwlep830ObU0FQ/S
uQ+6jDGVuMnl18LSzlgDb5CcVfEE0U1nZv3aNrsanbuQ/ZX3Xo7eSSn+P2tVx8uv
QCdfirdOxvFeUpl8Cg+UKsS5ZWu8oWMPrGZqGXGWNy45+SBA/hPPaJdKPxTOxFkU
buGVWlXjSQt82fGyNYSvVngOcRVJXixXA7jNhTdearfl6+wPTOIf5lbZqzCjCCsy
Iepy78V/BByYXnk2qnQCYN5wV5y5g4vHw4U4l83zW1ZE+Is4sJEo2aTTKv4QlUNl
W3WK42vsJHgaylbXeXYJEXdzTj97QoTYAiTaOV8+fDD4T8bAGkO9rlh3ZsB10xAB
4+OpWlB3lsIolcZ5RYRKZG53/yMEuSe5nKqqtmF7qqzcYizYFxHsmTeLLTIka6UW
FyR+O3rs0R5cWv7KukWDleV/dLI3P6Ej5cjnqNz+lPtpwAJzpoCBvW2BJ8kP3TFi
2qmcVpVBF8BkW4DsRcacKEzLYamiKpHO9hxQctiC1SCkpmjXKR5pmW1Zy6QlgAT0
/UoxiVsnOkTRa5S80/II1NWYN4tjniill9CBZF4AprSoldOEJrqI8HPEe/8QNbei
6t63Z3tebq6xU4sO6NAb5Ar6qQgEYX1MRxPaSlCrj7ZVaQkpn/Z0iIswZGUZ4gCc
0NTIisE2cEFQOGy79LX1wW8i2ZigQPEWKT080QNA+XA8supEwbxttZ4EkQo4dK00
sGWu/bAWKArNX6iDwwBg7RM/pKs5hAA7+CR9updgEnAdjbPhx36c8cVw0chkRINt
4H7C2VyhJPpo9xXYz/PC/o91maagw/eQ1WHJIWzU6UnOkJU/ZVZs41yW3ldHXHQU
lgOMQSCRiFwn+EKgHeFQWxk6EtCn18nC5KLIFR4jjAU4AnebnvNKI8juhxf6UDvr
9bGbBoHc/O7E7t/yb83YI6dhnErFfBwNiVXI9JvhihAG2eoNl8I/MuYEJATFTvBl
C/io63qZ/ayww6Y+3flQQfF/GzTwec7hVI2Sg6ZXDpgQtytrgemPQMgQeQhw/ARM
wqgQq4owkZgcBPx86qc2BAsOY8MTQNvbjUSp0F0vx232+z6EY34AsxRm9tbNlyzB
+bmnX6+g1UohBlY85/okeV2tCpDBUBoUSzuYj+uKMLSPTnu3HKRlJDAi403EtAv3
6SV4B5bYPesovdjGSUzvhHK/vw5SSweTjU8T0xLAcOo75HPmG5qtPmCFA85AM3Uz
ZaUdfJgBJuYA79rOP9XLo0hfyz8/wiwk1l+l+L0mYNsJDt6EfH2p5TLRRnZeuGn5
JDYUruFO1LvyX6wqj1TXqJQcBqtn8xYbPugVM8EUetgKOq2/u7w7ITqXr6aptZ7X
xZOTFBTsIJzq2SNmkv3WZ4UctrwwDza/rmUD1EkUsCr4EOJsNmJZxM0vZO+3r0mB
BHlBbZyzfj1duUkgL8Hsu7OCaboxfnd27+bqjHU3VThNwMwVJ1gOBp9rKNGCwF5I
389AXGusZqE4ZhKGFR7+hGxIaSGcnAdjHFrDVsiI3EsT08HFfp6YPXc7Rev8bIGi
LJZQzVaGKb6ijgM+dbH1aql/9sdnOrxxvWIo4bwvEfwcAoq/D0p2gqKJ3xCfgOQy
Kaue0StzERjBy6WRfv0PUT6dEI5o9AHq7Ua8qj5UbQPNMHe9vWjMCCyzQ0PD5830
XZWYN75PAlrh/t7PKUfuUxDpLIUBm0qGMPe+Y3rC7lyj2ov7RYfmxnGs+qVqjm12
duXFpP0J/gMRySOSCrya9oUUT3+vYdg58lKtPcWuivHDqy+SO5ozuSL3ZheNshji
ZbbGWSchV2kEp0T3G3Q8rUCBGhV+I1KhdUBjk/PBR38jUjzVVHy7sav+C9NhxZXP
pHPbVsBGr68LLAkDAkHnD/qVzneUrIqU4I0zz+lecfDVrbPK4nbTwEEVDBno+Mye
0i+xDVIxEHBoPIBqrvDUqj0WH6XEtjlmILqgoPjOch2O1I2XcmI9VU/WwjpecKQr
PPsP9oj05vo+7PrBsczsgJhlR/PnnXArOQ/pfi8BSUfMk/pG+p8V5A2660mJc+Ib
8nC2bC8KsFDearVlt0K/9Cz+hZrGa1sC3vIlQMU7fCXGrJvfEPy4IRCKjHENGKA5
JzPb2mDFlVSWzc43hvFwAXM5PywJYdWYSEvbCUzAgYJ4iqJa3NQLqZxpJNIwZ4eg
3UiWvt7fwG+G91w7pCm1AaDMnHOHoXsiSL0jHVARXptqmMPHapfwBzbjJXSPYKwq
Wz0CU/r8JaTWWk7Vk5jqSrtfzSEcehMSpZG05CmEcMwbm8Do19YPP8kKUpgCcW8/
yBD8JwzAde0O70rLROtO7JSFlLG0HR2jwA/dUXQ4221XpyIlpUfoOVKrB0PNrYOa
28boYho/YrvLsrgf7Qfq5uXO5ga1tbCLLVas+C2qv2GvM7zWorD0Wa3nOXp6JCnk
5ttOuHgf4nhs01jrqSu5q4EQhKTnaNyNlt5IIhkPG8QIWulHkfQbRKZc1OHiMurT
kfDAES/Y6Xk4PPLCsIRkoCeKWHnJX9qsI+ZRFik9zgkUruYvPCmeZMPtyrXeyKw1
MdcqmZh55CF5BYKyMIsSBh5R4SsOygE6TEynobW71WXguvcaWjgSKiMl8XWLpwJi
xNm0l4bBSjbb9/Bpn1jlCA7UsG62xEH8oCeQva6HVtQPFBdu1DoS7omEl1bpyckw
BYr60nVUOqpFyTgytPydvSdiH4L61P9J3ohnrfpnTJ5ERLZ2l4OJ63Qc/EirqJ1l
M440UKiUgVWOE3goSdT44e9LKNzDwKQxYGy6dHo2nhFMrDF2mLZ2z1kUk25+PG4k
peTJJgqxEWZ57jI+FDML6DBikehscdrsHqNB79Y0XOS5iwW96+7vdBkR8TayBts1
xoBDwWrQsiMwzvlkBcSPY0FN6sRgS7it2ujyuv9FH6hADXKj7ANyvsRM9neuFkMo
iQhkXjb/02VUIOkTNUcjzCP5B5s9CC9R7/dLHS4A05XI7NS3de0zxrhSuEaZmXg8
pSgEgHik/EGYG24QmYOOc0sajJgu2ZN6YiPJFog0NH0WBhpflAbFXVbvryqZR1Yj
Tp3f7kD45wnu9l4+yPIGm/7mSbHf18Lppy7mGZ9eA0UthJ20SFBxHJpaSvvIyY4L
nxFViNux7a0Yem3H90DxlLtGrkvdmGx103jaK3aX2fMueJ7YY0N62hhL3P/o4Mrx
qGQHF7AOVpwnNDGgr6FOv78XoOi62Cth5aFIsZj6SHHRT4tD7XyPbrUesEHzgo02
B5gwoNOnSPJhEqp/Oobh+1PvulvpacEEJiP0/AG/KDBEqNvI5x7cAp4J0bexIaBC
04xWMDxz9izyzqasDmWnZAbukMTVU3/WFGksvytgyhyP740hqz82BvjABKXpWv75
SKxHuS1ehttvZfVAfr4D8zCKo7nkHrpCq8Uf7XPVtswjxISUPxsBNq4hrKSGyim9
jcpv+XvC5pIHYQVrPG6Aw8+KWP27MN4iKk8D4mR1QOheMHM2GL2RN03xjS81NsGf
Ewxg+wAq7h1dmTWCpczzRwgKvW1IYDGbheCUk9ayGwGUNkc1s9Ojb5hW231+2LVZ
PpAC9424Z3lLkFW5HuaEu0AbF22bTkSNCeQw+BwgyeJav5M7fTz8M9bBr8y23Xey
H6iMNiD9QJfC7bMXke+ZJNsttvOyqbik+x/dCUQJKRLX30XhZr8AAWa50VKxzVdC
wD76oaHTHLiZYk+aUrmEJ6rLwtfOnuP+lufEx0wNrF8o3MIML7Z+uWqOMBio9huc
Tco90sPImKZYbvkf+o+YpJ7Lh19Rn8dGNOvNOgpb+Lbo/5oVgWTzaoCu8vYXtmU/
yvJlblAh2xrPMde6mm7vKJTvs4i226i0UjST69oipNXrnXeAOb6V5ID710D611Gs
58VAL0bL8kOQAZUitFlXSVb6e0IHYlPXci0Ae1Id36ksLi+5TrvYUTy1NxUjqSqy
zm9KVm3gy/U5Cb2zlCP/XM0kp7s09k3mcKc7thtYMfUbAKOYDqm/O1z3gWZI2PB5
VwWf28Qwe4DgpEqAvD1/ozzMrD848293xHsLcq9HOizQhJVawhaDpFbQmpOp/7ee
sqjep71OKE5MfgcAW/RYi/bXCkeWdC6bWAKlJI8oJF96Jt5P7QTV68L6mEkbhCtF
YQqEQJgpM7YqVVruX8DPO1iOzRjK1rsmz734Wl5QbiXTLEq9uBBWxYYzBgM9pGA5
LjT4RLBQM59rkH4SC2SYCLx0FV3SP4BOdhM/Lx09dp0vKEVvhVmttH2P5F2IJ2Cp
c1RzOORmP4fY0DdYKFQ7RD2iAo1OkKfZy24H13kiTIiUJeCsXfot3mZ8QhOM49EV
BeZZ6Gs8udSjV3v3l+S1Mkx7djv9UBablJbe1rdSJ3HWeDzS7uJtfyk9/CmvBITg
3jeyUlkS8o9ujAPpqmAnzpPPJQKZ1NCi4J3JcvOskgD0l1hYZAIJmhqLhXLP1mk1
uWt/XeSODRVTgacn/i/wXfR2L+JsyxZTOb85yNobHeYOHgYoI+FSXGthupC2wtfp
EkFVoVGnO7qUucwaG8FMa7HYs/0OOz8b2OzzxQ1K5oWxINHITr65J73J1kfOvUug
ps4diftd1ANUMPYCkmctn0iGTAxuOVo8zmjWbvYvLRucb9Q7ArYWVjhQgsHXGWTp
lLJ3SEYisg3r6nuvME3GXEMW0iVII55AX7GCWyQfKZquR0As2nNMTxsXKlME3br9
gKdOMe/8Xx8MmhatPNihRguCTPs5TKYPbSQf0Bq9maosC/xUr8exnIvUsPV23oHm
nh5UBCjKleqQIK4kDCm+28Pv27d/7CY3IgOIwcejH9LZC7ZqSfaMbLt3O+Mgf435
aSyMZuPc/aiCfQCP4oz2kAXY4dBjUKo/2/QgSPkAf04ymxBsUXehs/a8vFz6I7Vs
bJ6s05+ljUJO4C9CuCv9l47TV1wrJL/1dfYWsCLJweIHYBprT3YZLz6GeBYT9ifs
gttzoWGJmb7RNerWbqQr1IJKK2gDWDhJ1Oip+wd6x11v8dTLlq5SRUyYwXrSML6p
sPo+cmiZUCwbANXnj8Jop1q3gUPEHuJr/40OrVj0+Tao1RbtG4VkRfc+9VXXzS2r
7Fr2h/0b4zjjD0c2CzJykMrPfFzdNq4dQO3MM7Ljqz0JysMcQzo6f9DVOel2VcmT
lEOgoC6aPLDQFtf2O9B/JYbl0nJkxKvCYTA8YRKhwcv8JrOyhll09gMiHV2HQRUr
Y9HPjy4eviCnO6yTZ1ONKKrK6PkN9i3xG0vKglseEB5w5eFNHyIr9YNkBkaOxWK3
re0FEsHVsm0Md5JSrpG+CakyKIL7PV1qGBPggGFNLrB7WL8kTiGc/RsCX70iP5/E
ZEQrCHWWWiRRERTkW/K3GH97nirRa5Kd4Eo/UhYKDRLDeUtGfCRyG0pWpY59VONn
c8/HQ0Q0ccRQf71R8pkkDhisOThdQv4NvTNyfHR8pNQVXLJOLdg8A4N5A8QuViYf
3SdeQjRdDifCPjDu0Sc9wDOrIp8Oa8mv9A/cfj1RE0mGxRsAXtNKdFJ6myfmM8t0
mojwNVj08XaqxOkRALZr95PaQk7eDohLI03lAs0Wy5tzU4quzzDRIwhEZvR583G9
2fU8iJa5tprVNlBvCMyDcMm/FaO5ICvr3DAFGlKqGZH3HtcmYXRA9eCBMPoLFSMX
yEK0UPcP8zZDiN4Szgb4AXFZPYRcObSbAbzgWU0Po5GfocNhadkODrjqreha+EfN
Qnn606WiY55NPJGlN1ueCJMmGhSdtloaoovrsFckvS3Exr94KHP8CX+FaIcSl90n
ETr+p7dsjZqj9zVdztLxLZZ5dMFhylpkPOwiCqFXjcdnT481vyDA6j3oqOqchblu
BKTBFSc9B9PoYY2++PjHaWdCs9JZdhUsAcRdn/n5hmiOnqC+l329Yy5qWN5noWWo
xQamJoOZuC3Z10aNXvhL3yTUrFgBQH6o+WiHT8jXGRdF/ilLeeEuiw/5iW8SwWB6
JOe5nX1I2lY19ffWNfilGKmLaYDwPd70lHrGy2cxWfRyefRX+mSZpGCr4BuHfl8v
0ab1h7lWNGjg/tBW15Jqke4mr8lk7pNKUMyVlXBmI/Nye3HlubPjVCcfJysVeoyN
I5LpldzpLd02IUZpLAKQYmjN1JIe/BV5R2FE+3uz3lE/N3Tufi98dfEmOgHZyJj+
Qi4UeEqSItATyqwmNvHpjTLk+PvPTZVzPyjeTJtXXMPdZ3u9G0DExPM2L9AtrCeX
FZUsw4WkNykCpUposq6Toa8k59bxwgNe85LhwNM5W5Gb499h4xjLIHsJpbQVTyS5
C0I0zURnkkkR2oT130b2ZchM3Rw3t9W7JR3JhWuTnzkJk1nibEdNKISyaf9pLn+r
nkIfgCqzNDTGuZWmLUrZZdJI+hKetMjplaYadJtDnh9WRumFLutmMGi9W9/BPtvM
zl4F/wnqPuod/Y5HYd13LFieKCIG8QDS8usbLp717vhYq8M6EhUaD958NDQrTE7r
h5NwtCYqWfB/S7EYJIt4LYGtIO4tzI9+o94ITTPgpYvHzusKVZAXSv3bv22LUakJ
3sRoQFxuWV6q5ebn/wYYxfzhjhRBb/c5w+P1YIBS+ebVJPHpkOoFo5AzQCVt6VmY
rEuuzEPGO0oXdPL0tR2HtNa31mXatis/D/LWwkGFbR02uTqjMZLEnZUdvKwt5EWB
PAn2HAqG17VSE6fTdo6vxdDlhhD1UoZWOzfQisSReUa2juRiE3qx6xGBOesAMBud
F/wg8FwqChq8/2hnLGzXB3KPCI+aSTOJng7xMMGD4e8bkEPrRPWp8XPJSWtl/Dkt
Z8WrpHEM1lEIxdJKPpilBlT0HJjuLo0hKjmUaoJgPn579oN9AL51Ds7xlq97Fpoe
8jASHJeDi+a41TgFgNAeGuvnrpCo8CavlJtK+7XDVa6DbnPvGS0LZPWzq1vW3LMm
Kmft8ut7DcI+rmzImAGQ4h6gQK2mMzt2IemSdIWojiN7s4T2cbOWdVE6xkOQQ3D8
QIQicoxx0MDcBxn+Yar6fQ3HjWtYEGBb440JKcW/wEJ2rLs90QPqOA5EFbk5oZ9q
hf+zDl31mRulQLdS8TqKzQrc0SPCUveK5LoOz/J4sEBY5erCO3dmBBd/MTmR2XNU
wZJvE+HxvViR+mVAE5oInaiiWfFdwjNXBrSlckYX6MkSkXeMWwGHXxboO1M8eMMU
Y1d7boA+Kwl4U4WSz3UfNapn4XOIceVaLj9ibDgYf7iMaIRbC3p9FIgsqvr8Zb7J
9nEmT58L93St01B6kWYH6VqkvzFJMabSXclXw66PitMVs4VlYFfmM18PYOJzpBxk
D9l0nNlROtiF5dUxDUJ1gT5oOUpZJ/vJIt65PYuUiCHNXhgnj2W+KLM6RzYZv0v9
whDP/BCsRd/+eB2ekTJ5Zhmeo3Rma05jaDgYNEfW9vMClKfdGqY4ZMB6YEi51zq7
l98CnRvMTebM/1kB6zzqsdasoZCLX4/rr8w3C/uBhkzaswV2KwYBk2sCbpPtDr7K
Ruzbh1xvx7lABxtIs3jo6HveiyQ0mdn1sc+AuIB/ae3M89JAeddekyLG+YKD5a4B
ealCNW+2Kyq6SArDhVg1dIPyAEJ78EbBtmroUXwfn4yvi7Bj53vJVsbg1jElcJpu
re10ptRFUUqc29Ye/55c9CkyNqPsCCnYIVuTjd38aKoG92uJ4knrPE6ymmZxM8JR
f9BSgbu2KiFc2v9iGOSILdJCoE0bAqdHpqW/F8x8bG3yGVtGjgofvxT7x7mdUtRe
I2+QwUqfWiwj9DeBwscFfemTnUfek4PllZrfizpJoM6FCWSVMG0iOK6mSxA5XWX9
QINn6jfrjc8gaBu7slPS5D4fuHDR6bcQM8qtEZvt8R1B0lheJCsr8ebgxuYxPdJ/
sFq/KAZCor48kXnt0R95ZoBVNAPEyd6NSk2jC8cU5JEO1r3CHjtL9YF+bxwQfR91
40h/7okxI3H10AgOtBoMV+USUPafpC1LorvSgMUooj8pTY9gEb2r3CNLNqMQ0LAj
MZPlnPXzu5Majtxp47AtGWQxKpkYg5XpPwisFU8+KV4bNk8P3GNsM8XS90uZjKxP
VoSG9whs38VAbCk481KJzzpT+UrUJjd/g7gnfCGhSryUBRa0UAHKrHeoNYYlCAMW
0jfj+2V9xvVkLtoH1CDdQlEsSnLRgf+31lC0THgzl3nKTUB90D8crgJeySdz3C2l
jeYJ+0omC8TQXWl0zFIRIU9pqQLdpnpzWhEqiUZRg+2tRFMxfdWkSsfNSseTVBCT
Z83zleMEXfGt6avVqPLjP4tXjEARVK2rEIskqjeNSFL5D7HtyhGmJEe6nJ7QDjPJ
iPZdc5Tj+xLpZaTDanGm3i5rKVnFbZdzYGbnLZDQ4uUTXCwXwYSqMvLCv/Onv/CM
Lb6QPyyjyZ/nKO1lJcwAqjst/OTeiGWOtno9DHnuo6FjeMoGun4tRDz5Qvsfc6FK
beLoMlNfsMlqVw4G7+DmPt2Ji41s9AzybNYC28AgVXx2Fdb91rXerrt5c2o6tf89
qQdrxT2uWkRM95j11fe/BKU8TSViVluKANs3UgArQJZZ80kBginHM2dt0OEd6ZBc
vQSHr1vhT9EhavzU7jleJuNuxqSD6GriUUr54HWJBn7lTiAN5RyBEnTZO9kLRsQv
vtAyWZWPBUqcEHe6E78WAlWo6ZwQ7GghOubL6kS8JVQDMmtK6kxAQcEmiqrQsxRG
Tb24WqbTInXniuLKySP6GPQYkf5GQAnXCIIkZRKq2vo/VS6d834QDvpeUlWJV8cB
kba8zqLnhJ7maYwnfP+M7kFYMRUJ5laMQ0o9n9+YR7ZiEnqHE23NP5sYPiJMt2CY
NJ8wcmWnNoUcJdPhTRiRdCNZVmWZahhCugT4XRc4hojSronZNFn0O6o6lwmtKhBC
4SQt2fnqJD7t7D4lw/lNWK+toNEvkBdVGseW6P5WAFm9fUC5J5APmomyeE38DcCv
M91YDKHGxErxYxbC2DmC4+FMsYnMR0xzSxT8mX5UfHvucXvmEPOwn967rOcdUi7J
8CXwwjP4jvdV1ihB2DJzMD30emJtuMmRkAqfUEeD3lPZMo/67admDKqYQNuaKck6
6XNWeodgYbW8KD1eAi5OtiDKuJp4hhmNCC8Xi765WL6hOC43uKMCR5/S2s/BhekV
VNZKj7FeTXnmbFFEYitscLZkfcBF+WXxJZD7q+cTw78ZOPQdxdYxSw+4MOa/s5Iu
uMhbvHyEo9qYYUNSgtEFGgahBPcNi48XFYGhOJEmE7pfOkXp8gT0IfhWP0h1/Upl
JHV0vYIMzaJqsmxkvhkkBKxfRxoj6GpoFxveuLhlKy81J8ch8VT9wVeahDLHIhYd
TjWjc6Yz3z8K7AGuwvOiSAwSIbFGVipS97DUwSVR5Y+cqEG0SfV0z2FFJENgGeTS
DwdEcVMBKzgykod8KPPcLzWFjDju5cOOFI/rdAbqgsVlfILprHorVetGXAOrmlN9
VxWrI55e6uIpzogEvXJ9N3ggz9OCyW8TcM8CiARbWTixJP+A9OcTWciS6GUqFIdT
OmBZ1vYGG4GBpLrSC8QYyZoqRilaJsHbBj3KxRjhxtXUSu60y6+jirmeHYjKUvUM
XWi4HX88rzsyBnPeQ8hQYj65jekIDVDEKKKoAXxLPBgbx41Gg2sKqnXyRx5Q34GV
ycJQ3AIMIWhhCwejsaCDyQ+NXgrqRQUKKcH3gKdZq9WG/IPlQfpuEaZ+uJy5dPJH
GmD25mJFTD3IKYDEUCyxh8EOb+1L+n8fV9uJ7vhY9gm9J+YzJ1jhMDuNmwxjSn/9
xfmzdY9JKAXvoSM/k9RdK0pcf8ZCZ6J0v+HwapRMB7HkV6WqDOgVUE/2cNar/uAB
Z10IQGjNSskgZZ0Udqu094bh9VV7ecwPZA58gefkmVzELo/kkrIG9KSW1RMjnMPw
dxb7NTk3VgDeCk+a+ee94ZFZfNFSmmXh51+JfeeeqxIpc1C1OnnMEgJVVDT6vPeO
KCM1svKy9FDhtCx0/90DCR6Ewr8nGsjnTLNSocuqzb5eVCxEvt229CEOjMVTPXrq
lfbk6qH0NDAHH0VLrAaXFYafDBIJ+wd4CRHgP9LKphR2L67tHfaPMmTZCQpu2ofn
c/SGh9xCv71kRtgPR+wmPPHTkcXye7y1Y3Y7hMu9AXma+e7KzcUvkcMStAhaxQz+
JYcq1lFFwqaz7dgAN80xv40YEcF7CnguSd5kiGDBiJapUpJL8HQadG0x18acFQnL
eURKNIe1TtX2HGnIPc94IqtbvIdC6PSE01obEVZVKNSUi0xGh+nVsCvRmO8sRMYG
KdLqtIusMHz3+njl6vQW2FgGK6hXZiXMt+vYw1DcGeisKwpN3E8YqG+jzz/R42bJ
wwMsz11PUiwJj8kyzxjFCxeO5cyNO0JS8+3netFhpe0vo2WhXQNohrwW6HE98RKy
cZ2X+Vhn/p68OS4G8zPVpKyn3CRJFExnSI4xOquGlRO8NFvsejeV/ItpAnNlTtTi
/kqvTh83z39T2a3GnW/VVlj+FNB+8UlH/mWFQKtSJgDxcsKplLX1fCzNtk/BQIyu
236Xxuzj/9ViGAqc9XEh+vdepJEitvehZoozh9ppyRL84NSTID57MW0wJ39Xj4mP
sj4sUO3Sawjm8iGriRKanP+aN4DhxFCN/yTInASyHWGa9ePdCzLuZhi1FubFdDZo
v9Kr08fHufu32Fv42uNvzbdyYN8pWBw6qcZclh6P297WVu8KGzf488lJ+YoQdb7T
hvFfXEeDQBk0Am6aCkb3eh92ejam37MjUQBvfhNXJzpwaQIQzSHEh3rpaKGGLEMc
Etka4VdlQn3rgmZeR8uIJHzFB2xltPVmDQY5BcGIQBKOZe5jUc+JNwYDYVt+0jj1
K8wNjuDnaMkZ/ZcKkCZBGMcidiICnuTtgSjxDQgsjBO31VA7LI6CNgQ7WbQ1HyGH
/aFDKh9o2Fc8Qu2ShUssjVYfo/6HfZEos4e82ifAJ+QzJXO/UNNRu9iO57O9otpf
7YbivCB9Ojf7d6BuTmMoZZz0UAxjEqL/KEPD3p76+4vFxZKhnJPA6mV1wgFpic1+
OFu938ebXNf7WYqAhGschSWkDzc+UnnW/s5gzbinRH1MRJcLIfTMVHXhwBxJXyUo
XieYbWLCDKihi2ZZVikrMDA6Ni9LnbmfXUU8E6EKK0IxQ983xI4lsdgwv9bsDZv3
8IzeCxUDRi5VCa/R7lx7g+dDeOOCb/grVHXtvHx7eLMyLj+IFNEoncJovKWk24N5
y/nKl8ud4tPTjs/WvM4sY2zYnrITbYE/QB+7ZSzPmS6KSzvhC4k5AfPzM107dNse
1PCIUmhmKQx+T+L6kJRricvkYA+5QcYfTvd3uDquuMUgNWaQDw92GEGboneymL/1
O62nWn3cI4QXvGzhWU8Fz8XOhPwjwRYgk7dkV2xMKbRyc5kU5q2xHXPQmqnBlr3U
wVhbZdCV7eKQKknlc0BV7CmsOAmgx0NU5sJ8A75WBEX1ZwbCwztJrIoC1RB9418G
Xfkse2P+S+gIx5HUw7ENB0AsSH5HGmukCOPQnSRhkxr0u2SOD6rOE5TY1fDia6Ag
S+3gkEZ+UidY+TK+y+cKjMz8aAmcZHn06qntjVZMbr/g5W6e10T0YuxwN2MMKVvA
CjGScNGWSpKZj+9JrsEL91bBegBN6s6APR41azD/tmKoqjn6OXXizr1WHwqQe+TF
3R436ykARBWqZwdEToPaFe3N8JcPFiA/Yqq6prJBHTrtPpTPaVhOUU/U+u+9unUq
Q/lKfdmby6FbWzyMLFAzNLY+VY8kJ1MBEc+x/DiYU8+uYR1p0MHl4qnd6gxOx05H
mckzxJFG41Sv74uRlx1ptoXnxZdXV03uVydbOHEYpxJ1YNryXbrl43cBD300xNOA
9j89wQiCJ9ljdYaKGrIQUN1wA24Tu/LTva6ZLkUZc9NP2Oe0kWV5KCt8tygV/pTG
ri0+nTGk9zdpSwZ+kAuEp54WdT2XjFsuDlyCTpp5Mep3ewe+BzWJ0HRl70oISYeq
J6wtshxzxCEOIABCZ4usvRq8saUBmiv5MRcAfFTsUL1J1SGN0ncsjoVta6lk88EE
/erqY0McdOZ1xgLKWLkgOucLQwIrB/UwUTmAOn3jlXdYMxkgiABYhBkR0FrPATbg
mbmuL/5Rp7A+4ZJtzE+JH1gl9vsot5HQAMF3ONUlB5fv4Ig+sIQdclHkhGhqPcwT
ib3bwxxc28PiQBzWpkNvrh6dN+zFfOaL4x8o7H5ZHjrhSl38JFLGguGpDdYB9XIc
eYfFMY7Weoz+eMkt2ynyUz7NmuVDRzBW9rHzQ3gDqWPOezzJCKGBxEugrWMqbEBt
YyJwiNpmgO06iyN4//oohi4+5M54Vs1hls6XPsmOmHzsHIh0ZBYkWh/mtf9NVmiW
8NdOH/BBlrDFPy+FpKDOPsbYgYNnKMlqZ04zqfZX4A7mSd8a8xcJp2Kl3gi4qNMF
MgsfHDB/WIZG0j23hMsuNNXgFUE5TtPYwDMXnHQpWqV+U+6+M8VJ/j61MbkGoLcI
XPPhVZ3PoR9YeeQ3wOxBN9sP5zdZUCrzsJ59b4wcPBD567iHBxOV2vxnaqn75pnY
2KfvaNz01OvIob9mRuVLrI64CGsjFutrGMp8Tvv5nWw+1hOzGI7wKxDI8vX75+mL
Hr+o8Q7vJWgpKL9Qm2IyA7mufJJsqYRFlSyMmOFMzTRAHaV0ZcKYJb+ELz+TpTjq
GbF6TIiedoyiMeuVg0zNVqI/JY9/NuTgivWCyejtHJXfHTszAE82s5StelX4CXeO
6dqAXORY84pWbL73OZy0rLANdHlmwnN8v2D62hCNPUqXgoPPm0aYrhaznsTaBtP1
fDIQjNC3CLL2UmHv/0HClONh3rE/d55eF51kEkQLmr3icInxVgHzfjZDeT9I+Pkh
00bmD3m3GvwwVZ7ubeYkfplZDsxx2yNZeHfsCZXOGsv9ovbc1FskAm+mBp3c/IFP
O1naTakIPRXSk7QBjTy5ZToSFRb4qji4avanktkBo1zjoNPDi3eN5kFFg7Gcnpgv
nJv9YzcmMxpK1jC6AajJ7nCJ8bfN8frflGkqqhzbRGJUDesce/BujEU/y69ymPJq
BPF6KgkkPYO4Z+PGeSXQq27ER/sqCbcXW1Dlu38w5fQUgXga7kznxKNJaBx7ucTw
9jlf/eFzEAqegylAwXwiuWXZE4u53/cooe8X7Oci+XyyKZlDP42ujCcX2njVFtxZ
/3RPRCpJqMYBYiEsULJCbjBG4pX4ufPmOyW5+NQZy0DmYSqkGTyvokP+56Zqi91j
FlgLjEcR3+jKhtdrAuQsL3ne3tGkgYLGPl4anp5XObGhm2sQdGYOH0QnWyO0dyg0
/BNE3rnAPevaiIPeImVYsgz+yZnoNgMZ97M3x1IuNmsaRJeg/EJ4oSzsvDhQopWN
L8zewPNRH+YK808bIN+v0BIkgzM3hg31bL2FpcWlVOr8pSXSTcRvC2BQqRTzFt9c
8NPgdhMCoHDfQae5Xo4JOSo5dK0gGBK1/eQ7awlWJ+ZDTPL8Lihn0NGX6CVbvXuG
feA602UCH/HtKmjD9F7G53bJ7QWcRUEofkOSFA82dGQQuhrYWR/l+xBFvhmNg5Ba
PpdTn7Mu+WPFKKAAZTOxj/mJbbjSjrBzGZThsjI+jcPwQL8LJV61x6WcyvCky9vS
lS6JW0uvcSSP8RCx6LDOot88duMkb6MWV1kECXgNbwOP1V8rTAStyaFG3e9A7Mmm
nPLAZxtc5gZzok91lQB6GaVbJFZQIL56TBeCaVH7pikzUSrQUjX4T97hIW2YDHI5
3aRJxrJjVggKh1/KMngpRO4sVI6FWFNlRk8nbzNj0CHbNibkoh9lPN9tK9JNlcgb
dHz2AkGU/IVf6foEtdry9maozs/FTW8vB1XYbpRtQmmsvsPj2JKUlga/ZiKo/zPa
zxK9trDjtZBAsNToIPwRwlhpiIfpjbiQ4YokSnoggfVAQ1A+g5/dufMf/8hn3abS
RSbp29T7OMuYRwtwJHcsuzwYdrrJGB2klQoZijIvsPmY8nYWuj48b1QP6dLj2Tiq
Ws1CpZg/UnuULw80kLY3QTNAPEEd4+Lezq8s8FnpBsr0bREIkFxse+p5gXWTEBc7
C0DpDpx2+NY41vEEs7yQku8BhpbL7BZDkYDH8N2alC02Q+7wgHSkJ/5Amin8kiop
nROZLnUDM/rXULRFOYOjaSWxJPc+aKVjwsPLsAJ0q3FpuYqISwve9pm5qvfxb3dB
oNzd11ruD+KOiZ3Av1hDVGoooQ+j6ZPWEcNuQPUE8Nqpk4JVbzhX2r6qBhN6jBC1
LQ2/yBWhDWpTXSKR50uyTSwBqVN2wWNjjbeOSmw3syu8m2DLQIpmKs9NbNEBINBq
tTIkNQPAT6Q92KgcI3RtNK2c8M0F9HpKrnH7Qx0WMt19icFiHuMoxvn5WO9A1gnE
bobF3cG+5EfakYSEX3z+wUFeHehbgGVwnY9M5zdXTHhoB+mteGXiy8uihznb5ObU
oFfYOOx9o884IH48fUY1H4ZcCYZ1FKUT3HGyrqleRc6HrGd+moyq1mRJtej7cv6O
Ghfo+bO5CT336uvenfDDaqLz2f2Lw/Vo2qUdYNyvuCMX1X+eTG7I5Zkb9AzIM48G
j7CwDNXxR9wxGTWZqYXDYZa0q5J+9fq89x2yM4UXruxjBs37dmsXc3fTSxXDiySV
KBFWSUBlFvzoBehn+ZTra0EW+RlhWQ+aUUd3WiGXmur5ExTjjKgArz8ktYQSFmz4
FE7iIF9/abufDtttWeGvjiQwITQ/XxBQzRCQlmKUBnVhGgeQoqQ1Qp8u+ZiLCEsV
pvWfM/HJ1uuN5bbOvq6SdktbZIVan6Hf67HJYFHTuVldnUuJNVk5AZjew1QncYAk
SIbwleAoytI9ecWC6N8d0EZRNrp/ZS7f/7YVW+2oaG3/lznYfCdh9Iac3leQi63A
k4usR754hwtag/8Q+ZaRrY04bNMWx8rhVZQLqbrotxuMKM70Ai8fBZwmk4IOw/Sj
r+PvYHILJKXoCtb87UeV5dlrmUaBJbmrAxQxZewuxrxKWFqJfuj7faX/zTLAUlMt
ZFboNLTQ4ZKwcsJWREtpR7wQO19Z6oy/caEuo16evc9FuA0CgD8UwDV49R+IRbvp
DlbQuwBUDEChen61BeTswB1ezXCYzpNV0R8EapoylOAfgy+sOzDUZzUoRt5dhjsF
OUbAonSb013leD66T5sYJdmwIrrkYcsUvcURdhMSd41lFhdnlcLJle/B6idiTdxM
t1hWDEoxJvBcB35YJp5vusR7TkJ7EGaeyEbIg8Uur4jlBexgbwwoTkDnAlcIz4Av
mDqXY6xBgNx4zAYJVBFrDZrIOxgTuWPg6WX4vlahk41RMZW5j/PFIuq38rYFLFUq
cOdLXk5R37sYPMBDCyg3i7sHhULGFXtx+PAEzqqwDoI1kczb04mbt8jS5w/HCMn/
6hmWp9Rsg7LjFD1vt0swwa3QfN21Y24uSLsYMQaPXIPUsbg7YQeApjIs7UEaavOx
+dGkQLldo4vv7Cg9VaUX8ZLN6Db4TGPmr1z6bX+E20fdSqIJQC6P34RQOXHG/TRK
PAow5SHsIygX1aWp7GzZ9KVandCIdaW/rNv+Z9XtruS+nnm3X+EifXb40hXQSnAZ
PMM3XMJpRUbhwSEiNaTcj3r47VU2Vn/ZVTcB29yCglnxJAryLiwuATkHcYEBc64f
VoGfmAiCS8h4W8UhxQS6mORKI7VmHM5k4iQCRh52+HhNqDloNMHty3R11uWXWVR9
UWNkagx0tJQgK44yhPc0dcOJ9pI5eqGZjI9eUCDRU7JcMnDzig0Fxmv2VsHenIS6
ix5bKl5Q6+/ZqHyMRNinBUszqpN4+iy96KcdXpP3F37DljBwO/uf8+OZRjJoNxjD
AGp+Wm7jQleEqeaL6t7jhsSCqcchxDGD2rrC896O+kNIWuMukTKzdFL4stwt2qSm
iIRUhFSLIoSfIyHqIdpKzvBEj85hif04AopKDfjYL1/HxrXRFepWbIb9kphmxJo+
vKEdE/SsJXA60h2zY4huQ3uPa+NK0m0Ir8tSFITZkp2aUXws51EehMBrZoGsCKAd
60tAEyKsX7pr/EiIAqt1CjDlrSkbEJd4pmt0pebtgPqcHX8LG8awWArs8XVuId6X
J8XB1LCSXrJW57f5GvG4mi9rsIi+pw4L42tMb6Yz80Zw8u5LjbTlIfBw3e59tPBX
iZShlZEuuQWM9kNOhppCEpqwwfnpBJPvPj6wZBOao7oPttzNkmkj2SX8QKZ/aXbk
KBP38SgkcFH7OaK0tN7sw4LEtJnaYn8kbn8jbFOdpdolTBQDPx3lUtU8nvabNmoK
CK162p+BmxWzYDGDqDvYBFzJrTgvivpde5RqpvTlk7HZ9u8yQ25OFpQiISlE8SRs
o+s4/mDbwnlktOCFH/9QA66Kq4qdRkLBlOPz+QA14qSytb6X98dWJyrkRsZnlqHv
5G3WEgcnYgwzJiApdENERb3dBjZ0pq+DhuL7WZxrQs55UCW8e/Qc24sNS+N+eO/5
J13uNdn3Dlv/3JUtThP4gX0pp2lBXQNzX6OzQ0C+5Ve6eCJjmLZPH35fRCOyo8zW
BDJoAq3xYIbmEeQLJxooHaVidRB4VyFXlSqhQ+dHAlRHmGZHQ9qu7C8p9yXyICDG
1xBlnFumPL7KYBQJDSjUuj4lKyMudsMzcfkYXF9zxcydJOGjK8JGO7T14EHFNZIT
6ewfkOvDR/7uMgepRaR+qDIG82Gjl46QBQV7EoRbf08bv513VR09j9AXHTELPXsi
nrIEzA1yHyP9Zw+r6j+MPs6e8sJu4k25m9d6T+UAAS213shwQbzqDyGH7bRsuYd/
zFj00Bu7L5ZnRxulZy7PILo3AFKMW3rz/3WD9FeMu4M/Hb5Q2KsCR269b+njgNTA
yyFB7yOHZdLGk/Nc3QjHG/jFxMR5nPcJlbwbHL4ZQeazNesMkWBRw5PbkA36WvhJ
anGE4uOViEKKBcZHeXDlX4yfmtSb/rbYSAyMnxhu5yqaD2YWXyHvTWglNQPNXMAQ
9HspbhxpP9dw6+i0h8pce45pOkr4TqVX6z/qatgCLVocGPX0ONVTGWePoRTxY1tH
ZZLErx4XOul7KWOZgfkrJNA0w8OgTULaAmJYsDppuLRcylF0MCtAoTuQTpQBoDn+
jbT9fgrD1zQ4PSuLj2030PxFjdcyajrFOVmn2weEGIxeDgTJAuytZdKZJlZ6gb7D
T1lVA6RNpvnbjgjEbZEtc1TcNo9iR+OBs7xAMhKOFQ9C4YJ4OjnA+5u5q2TIdxVJ
1hBM7kO7Mxvchy88BZ5FPL102yGyaAuQPEic7PD8wXuHW9B7pSkj0UjVXE6oER9Y
rjE7PbYWU6DdXY5qzfbl29DVx4ERSqkbwsAoVSrGoxFU7wp94Wv5TEh4IUQhGZlj
qzJcAaBQNFSlZK6L/5bdOlzUE6AIMMKxmReOqzmycpXQSaR3KjIg77gQZE+Ze1PL
aAM2Grcxq9I4baFp57/8+K8qHH5vmQg+08gy+4vSxdni8RaV9mlhh0Xkvo1hSqxC
oGZuOUGKBD3sBQTiCnC9llPj50Mwj2bNo5LmZM5YEjNhwNPaBL3wOE7jpy5A6QjV
YJhyYIBtMIQ40y8smzR2qZ5QzWS8pHd8UVH2YVw5tZMEdp/x6QIk345n1wQHrHo/
VdIFiYOLRcD8LhnuWOY49YXhLxL0CSRvBbdP0/3VUN8dM37Bidx6h/GRzJ9Pgt8F
1t7N3spfMyoB6+ReIoFv2KDoSZZtuzBuqdwQWxuXOVFaxEA14jEZK81TXCCvMq84
/xDoHsFx0fi9F8WEpICvi45r9O3ghhWHG9h9mKAesVC9tG/cLIE6lukDKd+2UKfv
6yIl2JbkEgLg+uzymjd68ANnXwjXknBSQ8uD1VptzaTvOAgypB0Uuji5WU2LzlIs
NffDwBnfXJQgHzbWZ212D/DJuxj3evVOZ6btbbMjY8BALngJlRN9d6ZUO6yhQ/A+
zP6VTZYlg0mQ2ZBJR134lGvszrKIBfNjE/MuEKH9woT+6T3RRfs9quglQ21K/gpn
vWNIF7AHPP5TK9jQNFTvwtetptq48HNNY0JNnHCBsNBPVpt5fQtsISftpr2EwPWc
wK57A3j5t9amNFHtc46XCIfqf2tGopo//p5Rx1Opqdw2zuHXlGdMln7ASzmho6DF
ADiyvvwHrXiPwzbHarQt6NfuaHo46/248HXPm5Ir8kasE52D4tyPCMAkz8pabg3d
dS6btdmZCJMsNvVJmROUzUtvc3Fmz3OvQpHD0whqVu8fi0Z5FeVzdF1jiZTxdsV/
y0EQU07lerAYxFjVfrs0BzMdqSwvwJ17M0ebuq4lD1iCOmired4Tjdm9d6XfArCQ
bKZoS+YX58A4ihI+mBOAM8zu2OIRRRtg3sl5AdMXRuFCC5Df0gRRGr+njmN93tas
/KHoOe5vhBcJlr40UV6Q0Jbrb07IuB0apF8Ak992K6OcMQC/zmdwAHCXZkjkZ2SO
f0UGs2dTRmUoQENUbq5eKMGE1W3YhpOobCMX/x7wkfgz4H1SA5mi2KsEET2Pp53u
/ouqq8BFshl3xI6KdmyWogQZDTaYNIpYtgD5UUCTqxSrzqBkWSu4UJPXJXmFtnA1
Me/Da199xSk6zD32FExpAvAHb7MB9R8BzVRN6ODAXedijd7s6agM6/4ltyCRAy9W
U68RBubVnPc7/PAmbvREvKi7sQtgdPuJefxD0RNjbLrN4ToWyrKe/Jhu5eu5WsTT
VzEsntzqARWL4rxSeBTh45MSqtaUd4tTGNrkEBjhSuIqU6+yEXxcGuqJquS6LYFr
9ogRKJbpc3y1QpEHk/duYBffBOa+lM7YxlXh4n4ot+K1r8MtbBIW8m7zldN8op2m
jQQ0Il0FQvA8dA0mzv0DSnQ3Fu/PvR1qg482NszHBKHjscGAx8N7GjuXLGN42n9s
aYJDBUp8RZlljdHHEO8IFB4Acng9mwlOzGrHZXpfL03/o8R8xjSsSPtHG4mZ3nbP
khKzI0MoRv0rMHh29+Gs3xUZf1+H8gU/hyAXe140K8pPJw/1WBkDOLGECe7t5Zo/
Z7g7i9iW3pP04GpDKXuOfgye5lm4e3t2ZoUNr6dvE1e+S8ercCcTklUJSyZknJQf
2eacte1r8cSHE2AT2KBpuecnlnH1EZ+KvKMC21c0F4Iql9BOVw3asKESb3siEmSq
nWe+2GCrOWGV5LET4HQo7i1WpyDksrNGGm0KiHyjIGzEs0qDzH9EV+HfjtagISvr
Kt+hB7sDgKbMW7ozZaGsQFSkgtTu6/W746EUrzGw12e6cXkqKlowm6NRwhm5Be2Q
/jeIS/KVyR1nsdYvp70ofQfsf5OirhSEYEIP79TjtVz73Lw2ChZWW6j9uFJ4Ek69
y1T5Exdju0/3QdN6wNPXBwZL1WOAP7TbL7a+GZNUjHnTA5n6xslR3bHy2eJPkT8f
PHsCrdFcIPv5N6QZa691jCYvC2prVWg0BuXbTZrLy05/z2wrjtRKEkTGHWbXT8sd
aF07bDnAEHu2Z0Wh//mYFHC+52aKKzt1Nv95nlYxByR2OeZCdVOZzsn5fzMzRThp
x6CrQ+CV4i92DMk773rh1351jDJVpKKppWyeWBNe59clUVaLkDxGw8MMbyZ3rcr9
EK7g+kjoIkIYMCAj9XS5Xs/7R9yT4an8OfWfFxFw1qsLa9MTOeMru9W75xPI+Qy+
vud0VzyFEY0s2OZx01GnhEWQ6a9nWsnxYjFfuhcYv17YlYErnr8kniCvES5x3yiM
8LTWL28bosCGpOQLPE87lrgW7GOS8vW9heFLifph2krq0K/Fjt8GJFgQe2tcT2R+
QUJwOLMHFt/047CpHux8slJygQRrR6Cln/KaXOJhZOaTnRf62oPJ9ohzc/3Z3sGq
/1UmHZ7RkDStrUyn/yzuruxL90CWMlfGY2eROn4O43XBUTVqOB3Sscmg9ZcDpjgD
GuyyXDY5iWefftzZ3pVRL0UpnGYdalq89+1VGyVrOlBhXcCILsfVyHAjDqi2+m2D
udYu8owrPwhnE4gDY9lydte00eLoT0pbIsbanMD5JWDzWobNClipLoRcMxtwJ8KR
1yQpvru/ZI+awzV55e4RdaAYKzcr42bG5wKHvBcrhCwhGTNZTnjrMESRWLNw/N7Z
4D7kR0f4V7TCWdx7K0ZaI6iKYcNxM33qxr7a0K70FCbP+ivYSwLjPtQqelshXu44
tbtLm6gDii9Fg7XcJlh3r4bPKoYrfCT50mZi7juqm9b9CHzHYvSmo28Ng9XX1078
c0gK3ElwhCs8j+ZmWn07Wxwyr/hjsPHv2Yecp9cTiHt478CWA1XpHdboE5efkhzK
lwcG5fsHbcGKkO+48BGMdyTEVjXZ4x8T94XkE79zfIsC84/2z7UwBFJtPT9erMtG
vbPhM72o3rKazo3ZZkgyJx/nCXzGeNMqTr0Wjo32C7dR5MycWvAvOdtLZd6rax8K
t8ITNygRM1uzmszEjByrTQgTPf93Z0F2mwCDtHUMP2p40P3CGljlvYhIXeuBFmqN
tDVLpTEA/oNHlgA65chBOmXbk0HOQLh72+DJ9xCXR3Xi/oHz8KN5uWWEQWQcjvdk
D09Jw5ivrrVfnUYwZXTB3Z/P9BTK19ji8IPEdIHpFwsiduW0P6U2VMO3/jyYnWv0
wBWEVFOEbmKUSihlFOo0dALsmtOwM+MXa4ZF2KZNEaH+GMsjdzkf3nCUjDl7AF51
3eD4fatTxBt38B8ttOqrSrPF8XzV9RH5hIz1Fn1SRszwAjgvoB3Hnr7AnSJTvtwd
HIPtWgQrEIl7rlzLBrXkiQD9Z7IhJrzGE5nx5vAs6aFSMw/KD+wEtywrOmQdjJGJ
jqUFWqIuUHIWkbxgXKeEo9gDiuo3hUXFqlQLaQsQcc2TyAb6XV0DyNNW7WXa034V
Op0u/ZMZK4H0NKGFShOXXwh6UoplEwy4jqKHNZVYuObaAnjcbqb7df8cA0dDBnN0
OUmmvcUAaI55MyKpia3Qp6EPx1KvsYHtGOWM3Pts++nNEgrAJBfJJ5J22tBF6AUP
p61JGiP+2rrMamACvL+MMpjV/hj+xZiLo4Ram7dtEQF+ldRRsuVYX8hrGWTmrYK/
AbmcBg5IUKbZ9mxpFrQCeDOqLN5d4xRHqgDhEvk54/XFFixgcmhXUpMREelH52Wv
23tHrWRuHxdxm/3Poll0/sFJWn6ZvU3Md+O5I9xY1aMRNiUKHMeBxDwVRxXRmSYY
jgltRpCyR+TVMiUFXgs/4c0PibXv7e0/zWbeOZda+BQ5PpeU6zN03U55eXaQHSL6
YbGywY1+kXYacOiRKawY1mfingqoBebZuXYvbeqYAiISe/VwvEKvBefozkjcFREO
EzzSFkNnF23VAoi5DsRQ3ApF60xo0wDUdRA/nNCz3VAnVpnMVggipXZpFZC4ifUt
zNbUZmT4dn3Y7SccT7bgOuJ0DDXWXb1lpmtgGV1f4k3EMtp+ZSZhErfK3f8Qi0+8
XSrzMy4NQ8jap6I+czwgOyqMxBIIbnkeNS2qmxgZ/D3VCpBo3qilElX+c4RA5eBj
GufBUPm9wpen5KxqrgYdE+7StJjDbu64GqHX1O6kg602dZrpSbs+5OeK3loe8sjd
Me5CCTtAj2jOFmk+yWM7YZchTsf3UOWLsDKwA2ceMr8i8Ak+zxgq9iscos/eaB5Y
TsX/18T6HmmVZ6GBRuvMHBeHyHO9wPBeeZtbwH1P46Ri6ZHDGw6iYbAcUU6SOc6W
4rxISVApOmzdPf/+6U2z33N6q6Y0zJ3e/YJQawN0dOV3klUaSkYQ1PMK3/JhHxXV
89KhW4nqRawgJPLrwpt3afvIOw+8aR0JIyLSc5St7ikgBeVvVFtALNnfLUmpw3PX
TxCDy/xkul67izV0vqYMfDnd182MfhpZYfDEKOPj9MV6XmcWbFMboDf5T43gmnZF
boMvrdsS+OZRJuctJlQ9FK4SyeBMyowoZxAufqzz2gTYBlvxZfhDzFHM29k+d+fA
5W8y+kD23ST092NI8PR5LOuk5OWAberxnLEYmCNwYR7l4mfZ53nbbpkhx7E8lGtw
HbCuRylsSGaHSExJD/Go28065DuoMO0q2b3sdpxk7EzI8yDuGpxMtIPFgLSzmFu6
tHJoPzAubXthlL7XNEE65ahCBEz3jDljIt602lgGGrHCWEa4QqCrAtHjauu9IGI0
U2Wfu0t6LqZdOwnDBWAcZyL13wHEMEIuInj9LD4cSaJ5DhQwTUhZT8QhKscH9jTG
YcEbDy7QIRcOogZhkXDdNeCxN/R33L6hjE0TojYUxMlvuv/8F4nMB7tCBMxWXBl9
so6bb+rqPdeOqR+Z8czQuwbXa9lrV6KfS1GwIvv/Hrio1q49dOZCXOESphjFXGKH
pJ4uGagE5rBBqiZ0Oao7KpoU374r01lRpzptT1O7M8YMWD7knF3Ci8vc/AoCREA1
KijgZ7hatpX3+iDlJtpwFhJgOv0mSiF2s7Byi7EvbRMcjTT0Vy/+vhZHyLljcfXD
nKXzZKIw7/bKCHV0jQe/usYzk9Dt5IYOv/5ac04mRdcnoMwONS+e0YS9HTkix7+1
5jwD4y7crsuFB0UyfEqNr5mHvO8vIx9w2zGEZqhW+cfZnsKCrFghM1ied9YfthtM
LZy5jTz7R7Voxvgrj3E1UUGN03/NoZz2CscH9vUu9goVmAwyXp7NWpta33XCMzob
4WwqztgphibuDn1t2F8eO/yF0gccB17Cbteyd6uQklo6Oc/+3aukhK5r3AY8yxi8
UmGaKnBBHk3iqwwOuF7qBM/+uZuhXGEW7Zbe6U0uvRD92Rz1K5+cZo9Zjl1xipDW
kOMm+F2lw+RAIvkkf73MaGHjvCpv2mxXyey2emayySkLlBlSxNqk+Deyc5M0a0sM
P/pajL/E/sAcwYt2EFfpiZ0HfrEooCIMm8gdjrRlsj7zRZec82o7RStVt9Hrqm4D
ixsy26gUlWL06euBbWaZQErk46l3cwpN/pLV6JySDJGOFAyFomMyZQ3joPI5JSP+
U4Nf7WP4GjSRwGiQK3txZIX21MtAjO+/2Yqk/F/3FAWZwlr5VXIMwW2lVza8YY3Q
03uksV1Cs1B4k6y0oV9C61z1HXW923GlwvtNIktCoqqINlZWEs8Ri02dzLPpgDWT
S5WgeV3VdwwxZu2HDrLZCVj773lIrIeMQgHY8kMt0PIpmi4GDbjTMOOdol2LrT6C
ioFpY+YimnG2Y+3Sb6qcBGV4yF+suzzBNc3dWuMetHBhrGuuQk9gLmRE18vkPltP
65mBu0PcCsCQgnEMqr1GzDm2uCqxBXVKd+C1sdf0kBNDcpRmWu73MnSR4GdA/H1l
bgTGXIurCeYHBaTOzk+/Jkb/2mB/rnu6zGyaq+iOlmvWbIwBLeTac5Oiz7hCTwyR
x/n3A4b2qubp3n4tHzaWp4xIw/jJhquWSjBFXzfNExG+0/sTyepTfUdtu41O8GUc
NnAroiM9C0l2KN/sCASiNTFsKwSHjfSADovYuB2g+Yoyyjy4jdlOJCN6kncTdkH+
j9Dy3hi9A8QAZPgDh4zd3F+82fsAWkYrtZj4e5R4mM3z9Qdnm1LH3JvLA4s4jg7C
coXuZJj9TTH5VL9bVBRiO6YxOgm0jYV0zqTQu2rim9JBg4WbFizf/AY9Bt7TR7Qm
Ejz2QE6d79L+uM1iEp5dm2LqeI5i1E4FkmHk8WZxDsC68KF+w1jQJTwiqocizPMC
BF7vrB/cOILy6bbxEYfFNTUnE+TPM+E/gtxQxPSACb+g6kddk/VjWSeu8auvbmPx
IQbGYddfTaCBSXF0+VR/8c/TXZ0J5C0ynjK+Ipd9rfQtamz+63M20d4xP3LIZPeb
hQy1E+DKrmRj/t9k5uteVLpRTteb9CjtJPmOArHaI826jHKB0wiornROMJNUR+/e
Es3eNoS1eaFANTD0+epN9g1PiNKJosjgzDmtatfPye8VOBwGMCJcUNWxEwDkZi9V
/bm3NHz6PXdPMu1fTZhNjlQv5/uxDwxic5xy3gBxmsAw9hIzn+0tPvbaKOyemlDw
4sCWK/AjTAJ404Jb5MxpNsq/slzia1qxjVww11hJkbvHTGF+vogvM2CoH2QGzacp
v9AcpB8f9jnEb7EwdYhMUejMkI+phKsbipbtpFpods1DpREaGUUFOIt7DRO1ftG0
fjxvmsZAoLxqNfhZpfyeqQoydh+aE1iCWCb+Tmts66tyEoUsvs/E5mAGBcxjTeAI
V1BcXAAAPnAcCN9MQirZ1A6H1VYTnMWS8LKhI3aeIjjx25iJLEfFaIxUDvOGabyc
xQc1uvB085njo3m47cDs1jbKrYFIAd9dMd5PVmx6cUs1Yx3Ckaja2cK0HpChRxyS
59Ct+nupVIbZVqDPmG5+35WtfKIIel7sDyQLgjpKROXgnkNiJZ4tg3SVVq7txycL
N46lawSy0A6KCB64EgHzkS9woU9ksjP+E4MlIEXL24cpwDYl0bCB1b+6W9Hi1Z16
DZ/DWCXW9VxWP1vWffko3Z71WjXfTo0q1yaECmjjEHSmRGZARsgYcrYNddj1Zqbq
2F0hHsmPUpWygk3ZuvKrTQy1wOZKlR5az63jD1+k2P1Y2JCzz/aKfShzmqLBDbh3
b1TROuosnbev4xgfoqAXyRjSRRatLjWAxg7JI7f0sErW3MunimrmaSJ71l5M7DUL
y8RYO77JHxY4aJODWrtdskTwt5WD8Uop7NNU4YOZaCz2+uUtZgOyki1Chizp+evk
PHxzxTNubVu5UKTtM0U3NO16StePzpflvtn23+PRXbxCo25czh+gE4UpeGrjupv/
PS6m88d6COFZyqLur3aQldAmKZlpCsYbEI7xLg4ubbcYnN1TNR+PSEsgAHemzPys
snD+AYbRi8A+Y1V5kUY5m/uZCnCrTf6rHcUWXxi0yULUwESE/ex4yoEPQK9alZH4
7sJPuGB6opGug9OcE0f7tDJFH8IJPsxv8GNicDfgdgez4rIwi2tZ/OMjewWu8K0m
7dNbjE6NPDThoXnzSVNVgq3R9yo78tmXazxoPQ3tROSSfoACg3FT8ubo/8/Hy9Tx
ho3wX2vIJlDG/TDl0eMrNXGQ3SzzDNZxySHVrbvtiSUT+KpoaXzOC78q6pJWt4/Y
dkYhVCe+FeeZEdY+Su5TcKV/GAPYh59jmDUIC0nZtWh8+PkoKnLtNMptTSNsqj2R
BDKTQYVz8AEKMxUci7Tk0Ltw5M2yAzcv9bYOaPA/xCHT2B57T0fhK27Y+Yu/lSVy
1xeSrHbjXmILqJxism+BIvMRD7bB1Hp47MhRNnxv8FeVvq+rmC0s7tjqrk7M154a
jD57XDUMIiEOEyUECmJE+eJrFksF9Q5bU+HbpsWvx05dc9FDtB0sbGFWWB6CXLlc
vVes+ZDxrh51OAFn/S0xiYnQVgLCIngq5x3c6XyNVm7vcNWaWQbCVw4HccaqWQCZ
f/BdmDL6nPJjQa2DPQMjyCoivuGjFvgT6DOYsj/9Ozq99vB4lnyn23iLIOMdh86u
Lj8399RMLbJxc5W18qfqQa9Iy1Wz9hqXBnYsq3y/TeUMcoc218ih7SHLQTzcgFaw
L+xl401gJW19Lf14AAjlgPQbuXNGvkLIK7bDmzAnR50HJBYmleyNI4Avg4KhGrSi
Cntd0dYAiJhRVPhvK2L5WUnyuL0CpBVwuqM3/mG2XIH8FUkrHSqpLZb8jnVnQVs/
M2u21sVkw8nT9Xwvai3M6r8F7ESAlhr7jxWwz9Eb5iU7llbEZvedKaLS9ilT1rNo
Ti3Fe9DhQWD3grkZlGZ+2Cu91ohGUbEiVUQdx0eqhpQCwaTNd9QaeqMvgUcByP3r
OYpR1DSXjUX87xSiL3c6/Py3BF8FPxLYfx8oWnNe7qGjVenHO9T2UdReH9Ce4lI0
moALFczQrBNG1jRVwN+rwTRk3CWGxgHKg8yICHd9aLN+FE7IC0tK6XeStwNsveCR
dqwBcwZ4El8NzZNlF96nFlGCEwP0H449IE06pyRWqirL/aTfA7QBMKLdnIsaP5t+
5yaroNTx+gTLHNfSpI8Ft21YU22bavm3cwKieAbdvMsySbKxVsgu+0ifANluYHTU
+0CRKc7xOb5LOXEytEJ3vbkFE0yqtY9O1LI89pIh/lJKuR8DQ4VMrWy2k5LQ5oqV
dkvxzxgLh+Pz5g0X8njS39eIHUzlFJRN/ee0CUvaklssgsc/sgWPI27CMATgXOLJ
vNDoIpidxSATdXNIO0WS8574ptx6ZTaN+KWAFdn6w3ACP9dUAaWhMQt79cO6aDCO
PXXhDfwtJnwrtjkCRIbYDVWGopdrtseO/n5W332CUMD1I9dMBXJt/i0wqtOv+37g
bnDh2d3NuiTdmtI99Jzqy1+wxc6o2K9wiJALX32Fvmq8DXa+tWA5fjSYAEsX59MO
AgSZOXEEPnYkwP3nwEQ6/7pVTRqBiXTBPdF82BGWQMn1DAzVBe9KYEaJ5KDKvna+
dmVy8FntUYOrf3YRJjb5Koaq2Uc0DePriEuGe8N+yPRTBO8jzCPQ8QxoBkIp2EYV
QQUYmw3wd4t9FpZDCHXt41zLA/99TKNc6FxHn+P9PP6an5PLsr0novNcE2cVVd5q
3rLpyH+8mGM0SY0IBBYdeWJm4eCnSxiptgxpcBWtKUaqK3RN8Wisr4cqp4/X3i3G
LGX8pV3WbQG5OfgA9mzMa32dQmZ/5wjcYzhj9gAVcGc5a2UOilydcscl1TRQ0xud
o+BQIa3R1eihjafN2FWHvDmAYB8oGn5kzYFKZH60FisIbBmg8O9/3d0KOFcJPAMX
DxzzeR14pKR4QM60PXeedKMSlfvb/1uWg79y+Q13qrSFlg3T5Xp6Vxi1V6Uncsg6
qfbXqVSGpR2jpUmD8z+54y/3LsgNgAJMBU+bpGdSP4+5ey5X9RlP93KVP/nJhRgJ
y9EDMLTuJor5IagDY10KydvIihG9NR5yqQ+IL+Yr/GTCGlpgkyUkSGx/bGdI+76s
s+G67JS0PR4EU5OTcOpfb7IKSTTGFzT2wRgoLcT7WwV6Is5HX/t105OjDVRUNi2o
3zpq9QXdauzbSUA9Ch4+h3JCJT5s0KIOVB2my0uUiYTQX4/k/cEtsiFhGRmfo8IN
BmGi9O1AitibUo4VNS1bsyf9e1yuK+WE4SG8b6VbckGO7b3cSOGnRzAo0DWN3Pec
NQgjy6Q05oRqVKitHyNZazmbuk5RsXNbxqdqfFozKK8QP+k3DIAggiHxBmRkhH5a
YyE944rHb45CWcoEDEfGICtBswae5Ts5ihINnWAj9ZOClpkwR+BatFoOXtuwTYIK
T8ThUC8OX0ZqtNVtuPyo6L0ZG2nNGNEgtlRDwJXccrzexb9IuyyZkmzq6/0tpLLz
S2Oi5GH3tkeVxVaIm4otKbq729zLiQYPGvB8cvvKiJQTGJ/oEn/gfgvKOBWTZRzV
Rir5osL6dig7y311aDbJjN39sx7B6g1ZAPbLeGMjBlD/ZeoC6nG+TuoC6s1/FvHj
fg7U9f4P8ncs4hFhhb0mSH6ChZbsyeNO1FFybZVxF3Q1Z7mx7rVc5+QLhiX05u8w
UEgZ/zDuZ++easpzEIW2lHjyfwxb0dQUwDm7vf8KtcEqTnKuil8PYzGtmfDJ7VTF
yyULJQHq5S3MmiSPcVvvBKrvOIoOeFzgfNeQRaxQ3Hh/WrSK5B5y4jmnJAs7hLpI
LzG94jxp6DJOEqOLHkd9kEIsIfIUH/LhADOPp47Ycn2VnAHCrz2i07N73grvnbiD
E3wyDYIePWdPpBuX1+UTvVjuZqpJy6nptADa0vba+a16vlGc2hM1/A1GxrXKGGJX
TcPlScwK3gUOjvSyYmNOWzulUEeqUqIEzb9Ys6lmu0SLsnaNDZCyT1rToDwS8RFW
TW/bxyqgkwcLzu0BFUHm9h9tBYnaomg3vUxBrLUh4+D6bOmNsVPtifD/Tb5tba6A
gwUW4NP+Rd0115gEEIfrEsIhPl6WRvrxtz2+W4nqoIv0R0HMtON195STcMYAQLaK
o/tRxV2tH87miasmvzftF7Egz0gb591w5zSRsUN9Qxw4Eg2go30qR4+jzvOsnw0l
/IXOlobBwyCpv03u0B/vUEUFsziKqQS7PVKNndjbfbUrzoPXN8Jhl1BDhpeXAQyX
ljdJhX1yYrjo63PNFvozImOUtu9vj4oQEImHRBSd9COkFLVtE1rZ7s+upWhj1/ig
YXGrh8YibKzNpiqeY2LvXsOJnvJylnrPNzyTxj34fmBqcfi4sODLkPmK/e8D0Eax
hHLWMxaicAEA98k18XECP8DEhDCBOkJhXBBz47bbO3UYPMWAxWnk2/WJnW5IVG7s
axMYPshguq8uKvHkYvvyBICgBBZm86rh/aBMZzq6iQCXUgzie9amLawglwGrXO05
QbYmwpSVYFEbrMf5VVGKyvhZq+xZdJtHL0Za0Jd1GB5ib8ARUdQlz+Bwv1snQgJ8
LsAy/CnzCgx0sNMuCNAvv9BGSH3+svnw3QRftgSB/vOEO1m7xsmp8VJ+3MFRU26Z
nuJkU1LqdKeX88Lm6YRTJ5TQU/K9+bj33LrA8maVBzjjmP22eTT3hd0CLkeXML0x
tTL8Rw5JUnXiGJ7K/usVKe8c22b9wqetk6SeHNN7RC0E7YESuj1LO+VBnyQCdyLt
C9BBs1LTCmIN64E/bHwi2troBGFx5a0svBWqdaFWObraGL2KWQuDKdCRSOJTvYj9
oCEobopH9pjMrEcq7SV1BrSwALXgg5ullhXKxKgEA4PuTd2ZmQd6YAqgIxzjCh+T
cD+g39mMTMNK30w/fStlpdLT1MVOkwTjTorzFgPBRUTBcCf9IFbje9A9AdfAVNdj
ZdfafkuFXbRfprn230IKx8RxAmOXqMrU/aiE+beIXDuAKu4uderNygSlzVHt8s/d
nO4Dgt1cnv/twApOThzyLx5aDSuSKT7AnCiW2eTL2+55hofPe7bQiBmlPOEuJPWW
qJRd0SxrnQ7akx1Ii5JjfJ56gBlyGfW7UupilEPxEc8SJlglKMKHzPjPCOB2mz36
kLaGdVieYbl04Wx1l0A+TXp5yXHPZJTExXr7Q7WdgzDzcbR/c6Nol8YRq4LquyFq
Ti4lVfIDitilBYKjs2WaACKMJyMwDAkcsS6jaWNOqn7GFc+OuDegve+b5vzIQoJS
dTtPKyncV5aIMEqC489VsjdOidZuEK7gN4HjazBa4RGNpcWE2rPa0aUOolekBYio
+KmeagPJwiTI8awuPcUS6+MbGoas1dEq7+mGj3XmKgtJgiG3GKIzR1QLbpKilNdy
FXCdRSASVwUlhTzNiSo0MRwGjHYHXdK63Jq6SEgKvlS16BawSD6JWoA7Up9tsYr1
XjqiDPR+/l1LmnZCL5kDXQNBGEdzoov1LjxmAQfM2jTfvWMC57djev2IvZ9XDDpz
3FcT3hqkIRRGuAUfq+JeS0R5ORByIpLkEnFpIgNWmsA7+XKfFuYnZGZpboCQBicU
aFVgpKfvlfopmCbvV5MkHC6S2AQWNDP/9X4E0qRu8No6JfutjTIb7YEdNfwUyKJu
CXpLcYvaC9qYR461Lj8X/0t2wt7ZOEfzsuZN7ijn+G/zxUerQ+k9mimPetJ3z3k4
TjCgT3RVbKegkvdwXuikpxJV9f0whRcF6lGGO50y610CLfhYJXPx28rA7fIUFebV
SRGKWkV5alW74VWxcyqwqJ2b3xjR7nv9+6lKP8ARVB7rVio8K7kLxEzQ9EAOPfjb
sQEaPqVMJ9eK3yL9JjYVhXRQKJtdNtrFe5YIAZpz5U9/t3lAJRhr7udD5PjTkJEr
NKktO8ooQARHpo/oOCIjVFwlSGsmGJ4HRF9o71Dn8+5ct1UpKflV+T6WdY+efJXx
kOQB4frS4hNwzKpWHI3gIVgmNsmgtnVOLq05Qpm+KhUFK+dywjFybbVMluh01mq1
qGkTh7T3cd7//IEnVYwZGXbatB3jtkce9NQEHoanb6Zbr0gaT2AvpLk3c7pwRdrV
+J0qzeVqWD/qU6WmlpA5oT8P9e4tVYKQ5xhee01i+qPqiygPt9R9SaMpwyqALvcs
e0SG/xlmPH0ieajhB5bCKaBYIxVRIzHIlw2qhO+MPQmXfsEVljL3QtQiEMRYYN1m
fzWWDGUgotHGMF+ljqVbB3M6FdhBDKXyf3hDj2M0zaCjKi/g+EVYbrdDkDKt0b46
sCVIi7eWcAktIFCX5HtUtRtuYEss1ueWUR1LVcCjYjYWaDzidLLyTWHk1qNK+xvh
iFsIoambK8sd4jNwdqDEaD1/cAP3/MbLfQiVOwcpmGIHYAgMDBFUcxE149NM7ai3
A3Fp7Ytsd33bb4TKwrkWuLyUEd/4FAZ+YwSxJtyeUaG5M9DFEVOM8SWJ3wgkwbFV
8E7wTESpHcbUR16dmIIsrRgBEdh9NW8XCOo16613k7QMpkLX/FdNqE4ofwrw1Dl8
qfXfJwDmBruFsW56gn0hRH84v9Z1B4BorB57Wbujz8FbU2/wlP+xaOozGKbtgTNd
HPp+qhy01h3hBdQ8yv2uzSsWjvaBhDdyVPkRQW0Qox2A1C2YbLaF66Fnz9afIz2O
YMEVP0xUFEsRac2GKVSIFtun4O5rLudh+imlBZnFR50mcUzInFr9fhr6cGw0/yoa
XMwsnhAgk4SvBr7QKjdFSw89k+L5kzD6X18LqRrrEo96VFiPuve92gIYKI2538bK
hatv9XgAs1AVVmJyfuQv3KwZAhA3GECjhl2AGEO1Z8qNuupgclPCC+oORlnDOce1
vHNBqjwnKsc//pF6P526IJ6G52qoW8FKgyL04gDOP7+Ke521quCyf9T+EYFMLPuk
a8PewXX1FthGmIsomGGVB6+rlwxGk30XGMAJwF3vsEx6u1UZXCakPYz867hzNal9
j+ynGnAZTN4YglHf9ahjDwYJ0q0lmY2F2YiW1jEqQOLmeuOIsZWvbkbubXF3I+mp
ZJyopTTavbriglj1YfqIl80pajI7IawRf6+HeLBkdiP07DZTmbEqphXfN1KjbGI9
VcepjiX+j3DsGZ4SvrErC/QuFobuQ1ZsGC9Z9DG5a2BPEx0sbnzT397nDdtxFcFF
AQ7m+S2MGve9tRN3E0NfCbfbsdYB5esTVnxdrc/YFLbwyOYtqkoqPDtqmu41dwU4
bSaujAwN27VcI8qOu6U1QCuEruRp2gq1KhvTcXKaP4KFcVSXzCjOpsWdlaVOlJYj
JU9/GGedy4mHOMDGpXtDTGkT7GA3JPQhGH5C0o2z5hP4H8b9xNXQiynHAJBqRNGw
hhMcKIhf62fZcDS5K1uQe9HWNuAKR8fHAXethcVW1au1W8zNVYV9CgWF9NX+kZbQ
+LUz2+xtha6YxrBsFFDpLyWQEFZ2C5zneY4hXsTrR57szQVAV0+j8uBBjf4iGu4+
4E2C9LwPnpSpClBDjS+BNISGNUVSS1Bewfk5vbSUZRMAsqqpxFo5L/fnxSFkF7ds
WqRIPkqCxJeUAJgplTgOKbBqsTWzoFdMtc4haAhiJGZtcV1Obn3KAFmfXVHwUBqL
joHDXZsRU6AX3WkkH68cmovhi8jZOS2cO8F4CtUJDscIHki0zvi2hxHdBeTDyi7H
mLplpQD2ruiB3jFwKrATiiuS/WRmSQu68jhUdV2Jq3uQIYtiWrFAbL9ycCw7Hat1
B9rpGrmaoS84HqeyYs+eE9XLoodgQqyOOJmc/3U1dM22gc0XmgLQQVY/Kzubr8/m
Q3czCNZzDbCBraANbA956EdVJZJ9YarJljUD+vRom913flX6eN3+I/NHVjW3tTUF
2cKL/GYlfdwQUVWR4UdYVGE75Zt+FmSVS9lK2AinCMGGes2pc4yKcUZchYP0oeeI
ygqZfUSTVsWMuvdoKWnzicVKX93l53oaagx5qZqs5fwDr5X5XnRc8bqc5VPO5iUb
C8v+6l2z97bcANJtkPMx5juF4/Xl/9aVMcpRUp4FcXeMndtVPbOS7071RExZtGAZ
kraMHohngtkwEZy8jW1jriM0DXs90e2nxsr5OqI1mWuvujbM88VDgKu/hU3J7BOJ
oVw4vRhcglewNo2c+mGQr+kkQjmn4BBLqcJHDudElyEZfwrC/oy+JwZFgHBVEfZ5
tdma+p4D6nxi5u8xQCMle0yobYhcgxe2PDrBfdjgrPSEqSYW17sY1sbm6vlT/Z9j
zoFsF5cWzyBrqgNxpu4vnfcMg0UdhmiHlsxkrOAK0OHtIarn2KZX0nBwcZcoWOE2
u1ICM+S/d66R4xhpYDty/CqwOxxgXIOqxq2lOH4Td/ooq5Cl+MN0JBRwJxyyfZ3p
51PMjlNKQY1X7eh7r+CadB0Pur/Aa4251+njCIVacVfPxXoI7xUGB4a5UTVxqZ15
1cxnYU4QfGZe2Nivc4AMAKY194zJuC9AdcA54WV7BWkQ8XJjmhof5LMgHXs0U4we
8WTt3ClLgKVxZG9boodfeOxe4FjEofP0m2csh9IQkL8oHQRo0CdU3StYGNiJ5Fhe
VI58kXc2kXzXfGvjP5bhpUXZONxXxonbpSvygzWajfSSi1szf3Vl0seIo9KEJH8z
KhTJSFWZIub4+ye3/FI4T//ho1rNTL7Ig6BvIzG1S5AhTaJp7EbraQfDB0BM/OdQ
jkhXCqIctlLNWoRAmKrhAxhN+IRcnGXkN6OOWl/0cefjd6dGthOsIUDO97b3SiFZ
T1Lq+sqtURjWKjvBT2ZLUUFg/BQHu4jDQ9oVSEqjc9OquK/vrY754Sqz9ZIWwLt5
wVEizat93DWHYU35nkMSfyCQQLYzO59n1018p5Ej5cYJv1wWc5AxtDFJK18Un1iV
eNyhjj87XroKgiXsRuZ6BBq98kfeXcBNwV0VpgHtv+JY1e10dzJBeqpkptdixTv+
bXcvuPOAG8JZ2g46EsVJcBkNFkrhmLM/+kJLqOf8QQ8XeO8xW0fF4aeIAeaeU3+N
AmnxbX4snfHzIm4e6mxuhgOS6EbImBryNvQZ/Uy3vrj0+XDj1e2skKaVm2NIYWfG
f5GVJ08z6MMq6+FSIHFEGmkyvQRCbP5Q6wmCAXq1XN4m9zS3wf/cL6+Bu5sCKctN
MKqvBOS5ybfLMDuL0/q9s/ZnigH+KIMF6Loiw/odZr+d3v4j8u8OnUpCbrKF1UHE
3DXCr3L7b55D4Q56d7rEovD7jBsSrZDKpJDctmQNSYaQRwDPoYYca5kXQvOwx7E5
FJe8YmZ8bsQfdSQjF1pwVTeyyBcIVk+xzFqLORO2EF9BnthnNy1LOJE+4nGz+JSL
EuLBBGURForLUAEOgpDbPg1R+BuQzzIs/fVEXedsGNvv0NSr5GXzn3FxdWMWIivh
neUpujkUzrV6f+mDZNMH2iJZ9YWj4ApZ80ZoOFpoG3iWH8gr8Ar0BVrpFAU5eRNJ
/N9pxzND8Di537mOv96WoZON6oJtJzjBK+nuUW/a7SnfLJyuxMwDjmeHHFGsCM0h
sikKvI3am2xRlj5H+/VlqxVMmlplihwjKrSgzntmKDNgEoXwSXB24J5XLGr28L41
SK2wPMTNHJdSNTVz/BZrw/QSiyzc+i6pyV3KpxSi4BbrTSCisJL1TG1dkMdVwLy5
LyV5pZa8xjLmeqG9M2N7xAyzXvZNAFM84rAtgErAO63Z37OgbLYTw55zGquRY8En
GM1dKEFPpKia73+Wk3fEv6HncClM0jY/CiBSJlE97KjY8pNfFD4yGf5T6XbnGL87
HDq74nEHFa4VCSdyCrFCdzXnMCq7M3gPpKcJw86VSJl0Q9x1tlwYUV1RdsuCNGbQ
paWTdhrtD8eqKi71mysioaModh11jUOS9B5jE/qMZncH1gZ+rRONczTWOjfvrNc6
ebDdCyxkW5Oy/x9toXPBjdzEu96wudI/Kf2+FOZ2kVLbDoDmJZxhqmyFuarG2T5Y
i3MkagElQsHO+MBDdjFVObsLRPnzLy5zxXnU4/uVBWtDu3b6eM8/pJJJqC4Dpuqr
2MFBaf1C5gEjcVrTqh0Z4ODBvafLbJYtSygc7I8RnOVfn1iwEezBGKGJ8P+k8pEV
wCOPGW6HEk170z3wC+BMWZccb/8f53niRyWTt/atKpUs4V8STjrB6z6zWSi1Qd4R
28Rme/SithtrkXL80X27mywHhaYqSSp2aRRnhRji7pTsJgU/AzIXM9lIt8UqoKJL
QAbTvcvRbozNDX3dq6BvjVne58gchnfrT0OfhjxvfEFaS+1RgSpkWk7cSD2ODvGm
lkBCBJct+TuVxH04PZMyTsjGN3pzxOEBgMGWTkMWNm9Ik9MgnxbhepIObroFFVcd
xfFw6GuZcsW6UjO3oGYF8znvfllgor1PF1fF6c9GaFadpB9BWzvfKkHEGF5Eqa7c
PeA8j9HtLqj3xtVCp/1j4tmw19D8o5c/HMjwnyEq57LJHv1GRr1uYV0HPUERKmG6
6J/UCUbodX1e+uKLB53uyUvjFFOIRzxFZDKqlPIDKv4Thq/wag7udIU4CfdbFu5Z
d2IgwTNe4bgsUd2Om0l9HNAnq1sI9s8nWos8lPc3H2SURXnmUMG09R18/0uxBaej
ZeeUv6gSTWGt0E9IUdV6HNnsd/EeJPadSwiQDGlAWHwkWSHeHKpSZ7u9d3Z6/gi2
rcKk+8+N6idfZZ6iXzUcyjXnSq6z481wQeZX+zdCQRDDhhve7b66i39vtNcYnwCc
pNdd93iyjVZWNyPJdCYvh9taXq+Hgv7fLJzxL395lE8o4Yd9K9T0sXgxOkx0ZUOD
ZoOgrx1htTo6pQ+GbB/ACaFeDhPtl4h5llnS3J3cOpDmosVyFZCbzVbl1RmiLM4q
JZnRv3kr6rldWOwZvHhyHNTU9rIUl2jL3If5IyG1j0hacvpABuAnidZvz5mnE8cZ
fq+AHKYEV0lQx+bznrpNS60dptMBHXppxbt8mtKwctMGqMWRz47a+8gNLBmovpmP
IUuUMv8R/Ba7r/W8LIs8q8+HJpNu8aE2V9xzGlwhAcqmti5kACax2PSprGhZsr6k
PrA6CK5eA/7MlO6xpcKC2/KnJ4kps26orM+zqtvVmXdlioedDHnG3Vc6k8O5+YkR
XJMPvIxn1SkBdIN0Z6zFgj67PXPm3G3m8z8hMNXcbftSeSplsvkaNYcVlELiLoiU
ni4Rd4kcWZIO0ZBhu+WMaWJO64VWRfhyfSr/H7ORfaEgnERKP4+MIkr/qv0RLHMT
LIVUjV1FwjXrxqh1w9Nr/JJezDOFAZLcIgaGcoq09zMLwHcJaVFpgOgfz6Y3G7NE
e92BuAEWiluxwBXGH4SlBUwpKztM9t+ihewmZHHfw6n/8rLBcS+gnVWH0X07MeaW
CrX+KhyL1dOdW029Qvwl2vhBDcJa/8EJqXzukwCJHzu19WNZs+shovfIACLNibxh
GeY4W45SvzwKRv8TGaXBwqsh+djAlACGhZYeOW/PjLi9uDUPqUH5uXScFPO+gBuG
fx7Xfkw7seqRXFjHuIy2egmOUg88wTNAbbrmjdaniLDX7+aOBzVEMJR2RqeufWP2
ezPidGmFDaG/5iCimUv+v2pP80n84HKk71clrP8EySE5UMaahW9FVRzkFOBAGHhA
gXhHpfOiTM5SvjUqN5nKZU2GTQv8sngGO4mKzmdfPV5SQOYWOeRqA1ZvpAIsXvd3
Urj8PgsWim4jbvabvLjmmaOP1dy2j4Sna49Lmo1KUGCJEJcKmeB1Cu5E2KM7Qr8Z
CNq5vijBFJQllzYzyYeGJxgxLq3RV2kOkOwEIoM8vm3ZFp0Nd3DPm7X3GWwGeqkA
tJhNd4gT9wFEwIAKa56NHo7pYUid/HocQGmHGZlJW7PGGT/++45X7GitUWx/IKLd
+dZs/0+nGcNVcXwFhM7pi7/FTNwWbuTdFIdwq0ysFFqIpd4fMDViHCuDV5t5TSgS
xJuYpBvugiDDmbBrU5Dl6l7RoDTKa8XdcTTaOVcKnNKDH/oj+ZqB/CdeFNRF2cqj
pEDzoAQWICyGqf469L3b45JjWNsNd/I6F3/5Fuo0FgDFbD1SoqC265SneQip52n/
5G4Zuk8bC06Ftvyvd2lz/Z2uTHwUEBA4Asr5xzTgTR+mYfsEBKlaL39o/hwckb6C
ph97H3tfa6ryopYdiAYj3lVWHb8+OWeBP+36YYAIFBCyni1sqvvKV5UPgHGql8E6
TXhE53vTnntu/jVCmVh8g/zgqVAJAgySvRxdfwkiY0wACq2n3wo1MMIc5wORj7Kt
yD2i8JwZVQ1ePAuSAMxsEu4g9U8Ta8z9TshkkFIYskKSvE82JV2FpVFmclb5racy
xKwpen5Qn/61gvq+vegSNhmDB5EGr+jJe7bOKY7A9ykqOlG24d42G5VfrIDoXLA7
VYxy11iE8ifd4Q6yTrJP5iwSk3Y4n311EIIhfEkN+/m008X/RmpXaK/kg9027nn+
FA2L5nQ4+XSo18C9A+bkELJlpzyYzW4mHZ5PZls+J16VfhidRFNyxR03JAvo8WZR
6oz1jy4t5mbIM3epIovorGIi8hJBh7fGoiorjKB8p38JQcnOmUKXTmVeg10YBgGp
alRnJxy2RMZ7TInZ8a/fQcmup3ogDujyCARa8SYexgN13tURWbw70k8iEn+Smgzh
vN9bh0BViVqiTegysjHgIu+AZ8NftZuRneO7JACfJ2njyjmFJBjMYZp2M5mRUi9/
Cd1EZqR1EXfYsj9QrY9pujxxY05M9ZScaZt4KKUQY9LLwXwmEY8oVf3HrcDUhuFo
bOT8vbpjAztwoSmE20Yx9QXIrfgpGOMDxob8e/Rfz+GFNmP/WatDMtbCaonG8wU+
jSrg3m7s2F8gyQ8TpS8kj6v+vTKv9ZDVQKHOIB5eMMfyJVjH62LOWeYOnhjlYacX
pLiFXvpM1kH+jQpgoFd+mJYw9jc+flU+v5CXvui15lRFcecWju+wbsAuip6u+juw
5MpvIi6a9L52JLi6u3tsYDq1c93UmnpxHNj52VA+2ebPi6c+QP3wIWWlZ09yFf2p
2I0YFVbB084t7aqETRkvGDa09yX9syAswhzSKgu6HjFydWZH93mS61uepoUfc56J
HdR+ReMQvqVGP25y7OEEjQyPPmcwbu7xUINbd8VIszhqy47oaWiSSCsB4LaNKM0w
cyxIaSnpfXtGa7EsvdCQM5NLkMYZlJ2aqf3HWtgL/kJYM3Mfcqq7kY5xrSx0REzL
PPzmc0zFizmfvUICohh7lPC6/zN7FLGt+EcDCZnwuWwkR06yMcNR91mxOS1H3uDY
r+SzV9eulB319TUNscn9kQmZ8HzMYLbads4mGAn6xibo4jPI/zTgRzNw7RpzjzK4
2MxXHVQfZMXgro28vzROuWrDvZya0FpfaNgaanxEQvQeLuXj0YAEpsrpkpuCWK40
lhUYNuKPYXEVVcfCXFJ+zNz7twRWBG/ztopaZfonVyJWk623Fq5gryx9Ll/DE3+t
cKYHi5U4SYF4+33xrs0rBNxIOh2JU94uv3tpPfBmsiEJxgvzaymmxTgs7zysRc5o
GKzvi/hz45w9duePDRbMOu9ByNtvI3WPDIePpu+3T/QQzq6KvPFf5IQR8zQHDIFv
kIiHP6enyyPwfM2+8j3AJoOvuNdd65be3D5TlEmX5e7FBv7+I+NFRzfNj4pkoFeJ
JYUBRkq0Rm50myv363TZxDiyUCQppY1ZT2rtg+hMryLxHDpL8KdAasqF3uA5lLzI
y/5tUgAu/7RNg15Jbs8N2D5+IZIE2GLRnKzqj+bB14/N/O/AgiEkCarL3hPSOaZ8
Dv9g68ADNdI+8dk8xUmhwAM+XPOA5eTXnI93Suwyx4dQPqbKWGvdnbtGQpoBghSv
VdrA7W+BVQ8qKKZ38FOFsb7DtXcm6GU6srsyWFyFoyLbtbvfmig+6+zdcjeJmY6g
86jsN7WPyjuXpuCqkuDuFZj0l+OoFHDV6/Rs47ZAi3xJJBGGo36DrVKx0WkEAvzh
eLAI1v/M43KN6iZ5h3Z9fEr6+RbA52HKIxhO6lzz/WNq+8YOcYnWYyZ/Rnyw3gig
oX3D6NPlkR6xaOjWZvhTkIeSegWYAwLvGib7EPJJK4IbArZ8zvJ2ptqSSZ6VVqYa
nZWxnwoU2hGhqoCe2TTjivh6abUpzOlBERVVPu8KtznKllgvitu8cotJUSsjeB3/
DxKCTxPtMPAGluIe9wKZG7Cmy00AFoP6ecDJAu2l4ONkvLI7RX49elWsJYByrkfm
AGv5aH3F9pZ6Jj+ghS/NQUka6gL8yCj8FEDI5La2P8+zXkZQwwoSIHInKl53CoSj
LraOC+/co+4d4Qj/x5uxKrwjIznotn4xTuSFSiZB/4UURvy1dG/HZXhmj8NqxthS
zHjUypIxd0Cq6LjB0WDCKCrY1spZ1UN+6w3iHpWkBBtEoSJNH01f7hWqUSgHmkTI
IVepMYkYz9VC6yqAxAkfYwd26iD1yy4EIe1Xfh7p0K/2zZa+GbF5yNJmU6XFv2uu
hO2OyQRaPhIxqg4m6UqrfO2mUewd/LoLJ2LEGyJJ/EJpZStRJ+nMKklyH+FfSuf8
XJATn5oO4nTK1ARZmq9nEuezaVIyE8zAhUMEHJbh7Gv+Cjzx4eLqJgJ8UjROXGOV
2dtABCJ8fAJhrbnYMEXbfhiyhH6T/6UgXQZQwX0tIu1nCjAkxIUmQ3QSxPFZGRUL
Skn3FYhhh3bbomatLBJOADMEHSf69uitQraPb4Cy+gEbz4x6knOonPsgTFanDvGO
Z3FHjTSZJcbl2nqzpn5a8kPU6osNIGUY/GBbX+mtPSaqOeebwEDBcMDPZ4NyCH7X
Artx8i+K5T93swnfaHXJskd6Xds1k7/W+McvqZpzZCimPGqq1RjMqv9HuyyI4Jju
nm5k1NLUFBtpYItpnDvGH1D67uzlE7byfpegHUVTsNABsVVv7h81nTBUhIfo05XU
Ksvp5VuwPzCkgFJycVOgVq+9ygvQ4DZ6/SuVYt+Em7VOOjD9xIXrMJR6/ZooC8zJ
OU2k/MA1CdCuNEsJ9+X/Gy2MxGktYL+1p/szNjEiddIpWOq7GR/IOmH/3wQTZQ5x
ZbNNBBU0PWbPUOQGhxDEIeHOe+iSMmoQml90B6MGN5iVkvxYkb4j01IZ6cJCMYfF
41ccRO6ITDcOTU8Vcmo6vuy7dOXgdgWE3MiR0VsmkpW1qXFbDCJIWvKpqpp44e9k
Jk65ckMmNhAjRsi2ACiErSLIxvRvhMfZKEWYUuOM//7wWT3tpvusJWcF8ftRR6GZ
vfgckxre0ASH30DPCWb9/JC+k4pmFV5lFg0gSh9AKPzH7ufC9ZMBkkzgKtNFItYi
cdaWKiaJrn+DnHtugUXnX6zOGNxp434DgrFpi0nfLUOJoPcOef7nfyon40cVOXuM
F8XPknMUybNis44ZLswjniAJ6ISYgWaw2+NMukuefcc4VMFYgV66bao/yZMFe7sn
XWqIsnvdcAOwx5UyD1303ihiMaj7m6hSkVtg5wsIBniawnCIYVNlttvKTVvmxjUa
XO1rp7mZQGfT+MYX0AzgDc6uxQ9c/kEX0NQxiPWLYPJnTMIVNEdJT3B7YXDDXxzP
aZg2HfoBQYWSrubmj12+I9wwZRIsU9oIa/MLUSSuQcstLEuIlPFoC3dm4uMmR6K0
23j6XivlFRR6YI2rO77crr8gBkOUrwqCoEs6oWU+NxXjSR40i6vK8w1/lBL1Je3P
gWsJQ1eqniKfNNRKyo2jXKfC1WlcgAIO6xIc5nFnk0KqHARJLs3ugMosanAtJ16a
cdBpWTFz7SHmup2yL5BYC78h1AWzEH/4Bz++ahdtz1v76H3pMhXqxmTwbaqKalGF
UV3kSwGbJoRZVVXa3rrwre996q9cli6OSi3qOHzZUdlGh93AdTUY1imcYaIBGP3z
KfM46of2hXAlMqjQqp5GNeMiwHn1NEzz7WRkzdj1VvDqkOx/rwpsS5f0T8rH/IWS
qFge+V0QGqvZu5OrtXMPmvcyliQZzev0D/1CGneCE94vLhhPbJp1mHsC1BDC5uz6
LzQBx3JU5g+AmrQ2xAGH19NoqCjzWjSOyEhfpGudXsxlVdLOqII/Mny9cm8tH2iS
N5HVQH9Xq9R/wI+zcH/H3mFcUZZ8eTXCdZDIZenMANMx7gJof5AhJH0pdef47cmz
tYV0N+8wVQ+33/Hqg0eiKCHqwO1iwyqSBo8lr5H34ny0Z0LUY9YTHWcCIz9S5Tr8
2FONPvn+22wyub95Atu5h/RG2j8tp1IKqtpc2rEfkAFygG6S5kjCD6ulMmzdbXCX
06q3Cbcm57Yh+g3+h8MSIJqh4LQw01B1czYExeS3tkenQHTSsXupjruYoyLL99Ex
i+cV4TUEy2xXJeOEBnz8MtFIBDMZtqRCB8xeZDZqrR035EBl9SjzgDZvmi7vT19P
1222+daWbmIv5X5JSR4PRKQD+YcY8FLO5LyiwHKDSKhsugXattFiUVLRM6ZM7rfB
NWTaxXzd7OCcsZj9/40Et6JgP7bFOkXWoRn8rfMieVwrB0Cd06mPpKGLOhSSes8j
fWfyToK5Ye8eZOJP8GzjYM+7PHYY3h1CeCMwAx+QA93oqjI9DUROCo2JeApUHjXL
cgbvOeaZ0r/IjeXuftsuLOPlYu8+kW8WpS5bi+ATXZyQhUuD6vpyZXyIo6JvNDVB
rPONVfr2ANibh5fBobHlNnMEyvA3NxV3/Kc8m+Tv5zvOIH8oZqt3H2B0d7ruqQjo
isE9xfUxNctIqetdYTXdkq2RQMKtZSQZckA/xsG94ilc+SGn52ecSVpRnjlBI1XR
UrMkdh1N0ArFg3gvaBWz7966gy0sxBaVVy/TMsYY/0teIsQBRW+QEDVY/anVhXEB
RqYvTYwqbfXfG9tH80/nf9aVSbdL1rE8sA2yc051rDKFxpd6DZUk2IzkBTzRAzx2
Muq1D/oizRb68xjqVsyYi8r2MYrBdiGsPALlDCkmSZ90QWAuyASHY30qz9m2X85O
q1Ly42wzK9enC0x4uBQeLzM1yz/oQjmkkOFjqrtjn5L4ZNja2Fbs+UhG8p16UGHX
E89j4ZDOogV9W/4lNFVRzdUKfac8pcv3u2umlMop9g+H2QRsok7xzZF6iAlFb3SY
TcjEYOHKGoLCeArnJry1pmGpgswxRGr+7rnopl+EJkJDrf98EJ0hCK9js62vkj8z
W38Qx8rXdRhRvCS5xsRV7UwXT+6j4U2iE+0OgvM0T+XG49lpWLCptE3Cwz5O+o2t
Ems0dHxiOeCzox8Am2LHZxK0mPeesZRR5Y0b2ABUN/cAA1T+xUPtEhU9EWCtpr/5
axaiQ+dY0mWTMXIETNk5wrzD1nhISAs71esBJp8lDLn9uQ6Pk8mxBSeqcerwsqn9
1hDk326UuSD6av+4YJiZFS+lgnBToGbReLn6SxQU9d6l4xUWqFw40VHjFySua/sv
2uwK/ZgbDeJKwXU4qnVgIJIEGk0lS/Q7Behba5xoVSFzqdNCfb4nt0ku75sYbhGl
Ms4bTMqNCIwD9psQIK6syfN84L2pr+lq0TeVqmgofyYkVZ030skVS/zOEYCm5NSd
0Ll+Erlci7WVkczV0zQO2KlEWKPqkP8TyTTXBEYQZ2UyOfGytvN+831ZxP3JQ0Wd
6cJio3BhzoERvwHQ/LETXQNCvJ5aaZnnuyp97RdWJXdC6Q+wN9cyt4+oeYWea84Z
df1j+OnxniTu/RZ2OXzGBreiAEsNt62WiUjLrQWSQbbOy25HeCLQyZOyACjf7OQt
HdnzIX+ejYhSto2B05a9U4pC7uxAqgTObKBCR68E43KB3LTwEyp/2gejf0Zd6R4K
t4X5+MYMqy3vFB3iOWS/MxtNn58uj6BFn8R5AI9LvjDrtRn7LCD4dSwX/aTtKPlG
A+mFA/MkOoVuK8fh5wxMBBhPJlNaB+n18XkVAamFkRxrY/gsEIi5v69gDtdhYjnr
6TmUYOk6XSAz2zCVaI6iXYynm8EQILyh67aEsHsgZYajPvPTFPes0KzCyT4lPwyi
Nk9Ha68HCLZuPeCNX9hxoLNM6Dt5z8xeczqqcEPl5zh/OuorDYHMmr4Dtt91rCiH
9JfWM3vKWtsgKsrxRgqck420cJSX0mkxX9VWkdWTfu8fxhPjsIlZ+I+tCq1BG8ux
ILyRoEZEjQoJM1Ye+IWvQiK+zaUS1NhiGVOxbD+fqoby7pZ9DqNC0Z3GV859aZpY
ZPsaNBVnDdxRaw1eN1LRW7FpqPj9KD/wQ/sAl2QO5rE6w0cRKFFc5ImpFd/dbZ6K
cdRgCxA7Mq3XmCCBU6wE2sZv33knSbqtaCVm+n5ykWaQ1Z7r44+VJ1pK2tljZALV
5JYWX2PFoC1ur+cI9flkhM+jFThu7bYVND8cyns+C2XNgx3QpQs/4wDvXjNaZeif
cDuYL620BYiuZHEWBmh6YQy6/+uyREUkiKYpF7XkkErJ/4P4xBKXT3xyl2dMxlth
abDflTm5Emv1vKn4w8RkDei4f7ibpbrfV45/CejDO7dvEqRvBwBYIp5ZbWX+nr/N
To2ZnVxFkDWN9fmLfRxSTlmvTxHNEHnd78EN/f2d3axs1xL2FUk8S/JovzuplWb5
VfBOwcnF0uqHRqkitXR62NYccASj57v2rA0E9I+3nUqA3WcooXXgZ56jlxjad8RJ
f634klhX8tXUpucgsrEvQACZQ4e/ncONQyW5vgEfb4CmZnOggDiGITtZ/miHPsdk
TF+h3Pu/LabAdGI2HTRQOCSnTGfOiqwqaFvX38SA6onjgv0Ke8zajqBlEPv9aHmN
Jh50f4eRo4r7P7k9/ItHlVB4xe9bkVZXqKVDo7CZyH6n1MUZsl9RFzFgHJbT0kdH
Td/t0w/lH9dA0vhLBCaMYlggR3vm2Lmd5V3shDDiGlDzk3zFiLoHGxYHVuyRTglO
y8BvWUSFwLwF+KSqfucB/hSgaGAYtJw4z3WpbDFSuqCjbs/8osyrnpg5GbHAWtr7
MQGy21Fi34Mh9XIzgI6QaWh0Xed4Z5WJZ8FDTM/IKBC2YdpriZhMu9aXJkAcqfCi
HNsb7IqPDSsEnha3BKhtPzWRClyInYUOipc3iUB7ED78dwtKmg0CPPV8ZXBw/X6N
o+/6bSXM0C7X/CZfAKV7ywUFjplYJfxEXpq+6LTQZjgglXIS3MMGE5CaPw5r/wrR
Hyqxs/0WQGq9lF07a76Ar9MamrwY3BF6r400gKJ2mHc8XDO3cI90e9D7ODPmI5Ds
k+rbit3IALbXBe5VJ4MedIJ1htqd1m/MPu9Emt4vhnwEgPnxKrLEGHsAQyLhlV7d
36ZJuyM/jqYPwJmD4AunY393bMb9v1Y72K0IoCNR9Jn6Ol6fFvqgPAJSoVGhaOvH
VZylpU8kMVf6egWWq9CQ0LrHQgqZmli41oGl4nwNRSdaLjL+hG5Md2PG/B2vHhmO
f44h7IS8C3zvofMCogf5pBI4HrH8Hh+VdSRPMrGecejm1TSGb6af0N59L4y6T50f
W+iIVtiHfYcQI5m/6z8yw+fz2bb+ocZYvn9p7bv0NGR989xy3xsr2De4Jx49RHrk
LfkyFS7st5VIOSv/YjZFib02BJK/qzS6le7D+EcG8qC80ck2MtSJZxV+QpIALiaX
Im/bidANjY9NSjwpiF3soJFLC6LVlE1Fsml34K/cpkCx2TidfyBGQdHlJ+hK6gHz
YGuRq3y7X0laUBHcI0J/1R4sfHZrktw382JgKGrOZzyda5sMGE5yQ64zyVZ7Tmoh
Cb0XR4PBqHzT1eNGqJxsJukNQYIJN9kFon1pxo+jAYUkRFq6ERWitgAAvUwG4FIq
CXn23RsWywo9V4JHfnRcwk2ohN9C03P+ic+S38tar0k7dd+Ic/EyomaSq83ij+D4
4m6CPSxPKzezsXqSOURn8ihRse2yYIZ+8Iemqjwq+wDoU+qn/HuY8wdAxkEgWbR8
60eJM/kbAMUJSsjdVdYGjIMEnKQr2E6/bcxDYj4mSG7AFhSyWruOQvh1cQvQFJ+0
0rxmXgBZFeQChhbkHXfcvFSR9IyFAqPVw3kGBv7Ztrfjpks6uOA7ODoUJ++yXWuL
iL54eC4joexgesai5g9R/pWTf6sW/1jkvCOsyuSdNXNs1wH0imVg7weoF/GTG0Tz
Cai9TMWpmKkiq14P4u111D1LPQSgXxe2SaO4Z0mD9THD4DtaFL0cHxQPMwiaCGej
HvkQt1bQ2oQBiL+1Dxj08X9fs6Zwwpfo6Jaclv08XqkSVj5Mx3HQ9Z++rz8uzFdu
tq0+WKjl4HjAJJ1DPRpwieUIMe6lYfwha7KYazg8qyhnOQq9W8W1bvjoxqIXqy0B
PCxS1hMfsqw0ODLxY3TUEhgjnjN5DzHwuhcGRiTwBXaVjlaDa0BLKK2WBinNpHXy
eeEXrslZeTLN7rF5XbVc9F4677GugzueTz/13BJ76gI5qW/zCbjb1Jp2XWmbq+8o
8YnauTW102uYj0+b/a/cnlmVZNwwhOWKX//yy2+9NfwbJcfNqm4eZ2N9/nfvEaTc
YwTo/YFBHC+eQWfpcln8ZiwqgxuvuBRk4e69+vYoD97dJTWFtdJSeN3+YyyY1FN7
T74NN8QGxQU6s3GpNAhUhUoUDQNwU+DAytM5pR2dHG5EMcT27o7Yn2Z1btWqmk0g
8NTtJkpSRs4lnrfqQpOB4TLZpGpGOMlMCX+IfRfvyQHhg4OqtXtRytLgRP9EzhCA
hqXZO+UvIjssT6zsjiA3TgDMV0Zusqsd9ORiuPifvI7V0eHjbYaTySUG5SO1zdX7
5/+IpA6FFvnFgGqU3r+Aw8FMjYu1HV8ddMU5rJOhq094LQsXa1YlQHBR71FbKCmA
vaoOTsho15EZKZEPgjjCqRpiVYg28W/yECLMrBMIUKSr7MTAZHVy4jtl3Li2OU6S
+7cCLt3H5tBvgyZDpgcQCm00ziwie3hHJjjeWOQCG8F+o/wDsGP+teRDqabVrQNe
2CEuMF4ftwn8XzQU6S95A2VBDQCZPjiAEj78Kq3QiMtw0zybaEWqb9VmkPR4EylN
aeboCPM9WRkMsWSAHYOgyZR2L5B7XnXki3W5lMs/wXnXVUvEvX6A60NZTmfBWgKa
LwXtPHYsjp/mg2mbs5pyZCITmSjAbbFUB7miZs9SQZkKvdDY1eqZpBrIemnmh4Y7
rekcLxBohdAnpz7ngMqFE1njJjkEJPbEqcG4xWLtRLof8RRtK1ZWQHSGA57S1CYB
Hl4fD57nqBcup9P+8ZeQsdkSW+dQSToga5S+XA4VFYOg6pMen32fd4qvg5SHb7uw
1riwkoJwh9lBb7yuvf3g0y/gsnbxXaG+1MV1MCpKsgVN1WwI2dd9/kRtM+YgVwcE
wAzar2HuIdQRv5mhJ3leeOpZMgCW9u9v/p8ZGyCvIqp/2phWbI8Meu7lKa7Ua55I
my1ZadEOSwN2IF8io6kHH0+mpylZxy57g+57oK4J50NQi65soPh/Us8lhZGL/nhJ
m4UlhbEH/+AR7L12g23YbA0mMCqYeklmuwlWiVB41E1SdTL6AMqGxzykoFv3Qftd
iFvJH7lHtRoWUOO3IexSX+SONFeyGMYfdv5wnqs3jeOcyDttGVI3cvTrsoXiasfO
vV+wnVQ5Xt7sumiJk1KCwWiegaUA0QW/Tv92rcXPknzrGiHp3VEGlr55mxud6MHb
jXZsZiMokYYnVddiNcsnT3f+nzou7xa8yEoCAuxoHlVi5t5qfnXjOaN6z/hLBvOE
uFe60mQR9B+snnEJycKHqUn3zXQuSmg+MkRgxo0KBOioYAzEJNkgTemfD2yYBs9G
KYOKru9cOm//vc5JrkUdUz34Rc4iXM432CwK5eDlQeIOyGBO3WJDY7Ccnt+wxIN+
NYgqjovfr6MlK28+9bVHfeM/tMOcfxw9ERkkEGTU1yhprjnbx8rzwV4d4VlXXqa7
KaEs/WKwFvnToFGSZKXtLMuQZ28LHbu4OcfwcOIMmCVEcgMS/ViZ6UIBkW5SamiH
Owmuow1TNuwkJ9nVBs8ZXv5vfybU8P1iCXDpEuDDrIYqCh61sGLBNVzYKm4XaOIY
0a/dd1qGGde2Ium5H+df0yatRZVO7RUpfNvXbXlT/AR9ViAktetDEYMWXHlbI3eo
N6wDjJY0eZwybtx6kRiCcUOeuTZVIt1FpxnkCsMsyTEhpx6QnGmyxzeG+FbBqvQG
D2qC5FHSbJtqsHScfeTEEVcXfdPRDz6TERc+bJJbu1pRdtUV+z9N5nB5g13qWeRt
79DUbPIV8Toc2E5UZ/nBoz0X98ljHYUKZPIntuuTDQ/hnNw2/G6oq0boyhKZYWQU
QiRYv0zh2K75c1A/rteJufCA72SKEK6mrVUpgc3cEWEhPtfhKKQ/WeLC3X1xVd2z
86WzgKhPmPBToqjJUFnhOnnQz4uOx6Jccyy5t5o9ptGOU/VmNC2TJ+JyMpiEIKyA
61bZAWStwlurAjkAzG4jZTgC+YG3ArxOXDnGcseXBRJuAiNrp3SqsI7CB7lGufzm
Nn8nh5LZSRI4R1YmoqSbbJpQiwplmPhNIzkF1MsgL5fjxiv5vU0ec4Slqr2D5KmA
kztyJpul40tKOk1IASy6+BVHCKCL4D9M5bhAHNkHBuf6Eaek0yjFaCQg0NhqoYoG
VjhPY1jEgcnRiH/XwgwiO50D640+xLqLJQk9qZ+JTm7sGzKMq+Hq6JS1toFwxp85
epuAdT323BeFt2euc1MgBs1w5yp6LlIn0pgvEi+b4cX1P0P8e8FzCkaAHWpnxMew
wqu7mArPHwYR9Mi9Mten/LM6cfJjotd5ZaNhBbgOE9Igechy9U9XHkv0wdnKB4Pp
QxOFdC+ufHrAZriTWdZ8G4eaS1avplhuNLeQs6sEfjg6UhIORiNkHbmcnqufUkPd
g+zZecj1jntYo6i+/Ihe6SSUyIHiGAWUOG4RHFct55098F8sPL5SYOO+Bw6KQZc2
ca8MMVKB4OBNmaQeJDEm9Tm381sFgLKDgU7peTkybKXkpX7AsUGwNIzfck2dANVZ
pPvjuJOTlIuA6U3ZJanYqfiXoxyxU9Dba5fXtCAL8QU0z0gVh40drM4mU34Oxq8P
AsX1yTctSQhKS9nuSd2x7dPlnJRYRFL0MqBZ6yVrlfylkJoawFtPqyJdCfNZEJiL
aLmqPvW7CKdTSdyHfmY1OHDcnyQlBzCi+yCytw9GM4mizNpgLd0rlBbldA8vvNV3
d/ECAqyOcJknaLQW/M3iPjea6Ct7bV+EIetsXTXJ0FUKB4CR+wFHDEs85+1MpL17
zeUcVeknzxFHcsDyaoixbu6XvODZ+/8RctAWR9y5xagK50ygkOrynWtUJm1qJIus
gw06C2/6E1dWHj5zZQA9j4Uahmf8wHAs2jnP4YnLiV8d9Eqz0lpwChHAa1VbbGg+
ZJjFIU9r8MUPwgOkotvYKDleJQqFHapcI3PvacJ3ofgfvorBbz810HeFAUfv4I7d
8/cWNG0rnKdLniQ66bEnpVzTUH+EdXvKATuRLkC4YWqXGTTwyUnIe7sDEU8ULD2v
f/Q3qwbHSV5xMmf9mE0K006zoCMwPaH/Lnayj++7mikbfCzjV8g3U7X7qgQ13CTp
jI8F5GK+d/qN3ZdJ/TjRxeWGOzSrk75WQRlQinoTjsfjyHKfw06raV7qdE3O8vQw
y3dhluDH95+BoTo5y+8nu09hckNyn5/c5FgYNZKKLq5kh5oyS13Y2IG6iB9A/Y7Y
B1SpiRq8n0DqfbPVHUbVIN86YIujUq0uaQkmljZmmMZ49+2g7Y87qi58/tTePbCj
PBZ9F5YaNzYbzjeIdb9SwZdBJ9jSQVs1BWuAW9hyA/LHuWzZ2Y4eJ8Ml6oPL6V+b
nv1dwPAjEmKhWodUzxQG8pzWqcLFgX0w/iDVGOEsKkpycTNfkAoYJVoybsZV/MT/
AlAmuPBMzI8/0eVOP19FbKovd2buyZ74FQQ5jkP0tB8b3KL1x8KEWBTuX0EFYBFq
BaDxres2v7hDZsy6jeOFL6ZUj/09GhnkSmCdLZsVAAG9BzCjDoYDoU+oNZZFpn/i
ESzOoNMtR8c/ZaypYlZTD/tS2YtXVEACy3RCs67TYRfKRb08DvQKym5fMhhl9Zs8
7GDJICHOwEJ57MAsp4Tmy/ysp+agITi6hS6cV3pxBkcRCk3568S15Gk+VKNm/uki
SVrRQmaBrHn4qAE7BX1Qtptz2M4CIRcCWfhHWPOR4kxz/qD4HHoSwaJRpG9ZqX5O
el9IkBQ25cBDL6hIQe9AWmgrVxzZs+VFpqtAnpvEvoeZiwZ8goMiTgE3YYgtz1hQ
YU39HdAbeRDYuq1NF910ihAJ1SYl35X/dHxL2IL4SiKDA9W1eE3DBKn6WjW4sQQ7
NSk9zT57pQizCGqX2c333JIfWNkyx4yQNybUV0TmNqUA96tqaX7AJoQSMpAQxp2E
W9itqVJ8UTd63klOdLvkCvJSMKr1hJEuOXIEwhW5JVhEpbcHBnKiVI/qYnM0ITr4
j5DlTRa+iv9aYH+ERk+2D6ho62c5WXI8FTo3HSJPTq+N/Jgqb6Ek9epZvthPh8aD
4aRFrai/LbVR5ZiLinxtjxAuC/Mn1uJ3csioqB08CkfKWU5YVeMZQAPmNe3haxvg
KYrVVPj2F0rXP+EBMlsTOFkGZ5j91LYIveSVGdu99IZxJnw3Jc1NX53px1kRuI8V
OvjNZ/LtW8fAKeKRB+YIs0z3f79w5CpwXBOw5ucJlNO3/RkF0dgQQTz6juyugRvt
z7dBjUp/DXpIT6wphHCgSS6ufr4KVJ37Iiw+65b5UF8SlltgrD3xIA2e0U/7jp0s
kQHj/Jh72XNVhP/jsAs5jthyCPTrC4mXnRfO56aa13snaxnOTXQj3yFtOIt+9qE4
z5op39ieak4MYIBtUwvOdZm/6OrIGfLCk1mt2WJDacMZ/3tZ9dqPn72zQz1fdJlG
r8YZeZgZpp+Ny43wDTWlvpgy3BoY5VYghRaROiKVAVEXctfsB+BjdeEN+MorDsec
A58sdVywxTRt0p1kp3rHb82FYC3MYlmUe+q98F9B49FFGS9Kh8FXIPmn5DqqDufN
QHF+OAzN4XHdvC0LkN9GOtWaW5MY+8ChV/8i23XpC71/SIS8eVubOVY296sB9C/a
RmyYNrhTYwJy4tLElEwLXhdB+hhG2gv5hgXqrkMFz/ZfgKD9dDjs5rsM9mmi2fwu
2GIFlSIyS4NHzz/NfjoQiV23TUhAm0UnKvR/lAa5qEBWXoaZu8aPkETdPmZMGGR3
sB4zF5kyQDrTNgcHFdWNXRhfwBpHCtBKK9Ell0vHFvcXSIQuTe1M14gm45NXB7xh
aSEIVrue/Qc18NOFS5lC1F7Rha/CMFv+3wKVLVhPSRAYqMxCxAufnqNLihrbYzkN
g/9M3mpHgXoO4plEoMOwXqP29zz6OqsLRzKjzVjUKMggK9ma+FPUOK04uWUgdkvQ
fVdeYxEqWkcuJSRsqbjMveSMLXY8n2uiBfUX1Dl0uttAguXz2O/sfl2Q+57xaTuS
5u4uFsqT/+t+TJnoWDQDszugaR92BOko6z68CUkeydKYd8/awpXgDKzBlGT/85Tx
M8eC3p/QgaVk8c9kAasD6976L/Ep/b351QpzpIS3EvcoMmgScATUcX9EIjZYsxnL
87oDWECwgZXxmk1ddXLjdro+TjBGoEK/seQ+iW2K5nCKnE2vHgWKmCdZCHwouPBK
OH0vQAnAz57YVXA+Arh94djRY28bENppNJR85Gwl9H+hKbpxlFuLygtL6V4o8fYo
pjDotqEbNp+APMvMRujYe+WFlI2SklZs+Z856ydpoJ1nDcLG1UoWBbu97IWWcj6H
OjMtH5Dw4SoEWQAfx2cW1/4FVmUcIeZFINXgOxxO5OsdeuK0yPuo6pKLoUQBImow
ffTbHDVh+bkmnjThWmg2B1PB2wGmmSYWb2qyYLOVwnQMI9zadfXl+AAiHq2N1HQ7
vRKvUKNrAX9Rfrt/cMTvaxAammsRIVOOR9A8F8Atre2ogvBVWuw+OkbuTj5YOCeX
viCcG+p2N0XokGtApeMu8hdN7en5+RBp9g/Ri/2GKf4sTX+RJvWboQBpHsjZinB0
Z7UzsJefItfE2VDhPvz3f4FCjdCR48Hio4KJMIurObUlZ4HuBno5wwYalZpieQx1
EIyoDOW1lzAM9Q6mgS58CY32tnLXsxomndMJfnFXxj4rBJdH+aNHazAGowRKiPdf
ueH3iNca10MYbpSuQO1ET3VDokRK8L9fjsu14XcYopnM6MPIUvJYDsyZdgl6iHOB
YrsSGAyX10rPqy021UO1wxUFA/0cQoRMz1QdZebdQ1xW0W4KSLcopQ105ARfZXYE
a0/mPBEy1X6wDqnbfxL9X6sNxB9UINUk9ZEi5OgAO2KlPabPJKJhc2DpBHgdOIps
/C0zp5qbomI/9QrRPgm2XQtLWrCONXgs4RWuuqPt4H0Oo29h6JlN2+KIUOHP9IYq
zvLVZIL2hjNYMGa/drxkQAwL3aFeZ9et8k1Bolym4ZvyyK9MWUySi7E+JZ/+G0+X
QpdjOEzdYCmQwCwajRqjy6aoVRl/Gs6rHuRMR9z/jfX4Xg/ilFafccfDJxo3HskC
v6Y31aTZW5qmxbLA81p30LfGE6SRl0XZma7MlBRUyFfqcSZNnkX5MXuNj+rg36C4
9PZnkeTVZnX3KONIraR/vqLkzo6TPo41lY8Ja3Pnh6jlWP+1eMgzA0PRpf+UEl7a
B7DCUotOG4Vtm0kJXB4BzN4Ysu6YXJ6eBwAWslFVkqTPnz+iX3wW0lFrVKP2PHGd
TXIEopzIZrSAdKugFxaUHdWPhFnELb5eFvk7u6sLbYgi3y1Rlv+SjxISm3jfEFgv
xTH/1EpiHSWrdvASvItIjJmgylrWTNtO/eq9DgkV4LXkofuxAFMy7T+KR0XOaBBs
encRxtkr94q2H4UbfvLNloPmXjG1SZ/a7R3rhZ8kT8nbRtXWwJ+SFRiNlpKiHhKi
l83sV2PvrbLniZlKBMb343axXMy1ZDb7nUWGrmI7cEU0HIvSPVjIl2H/Q/EXSDwz
ybQHrebBnrju+Vr9qRMPfQC4ZbZ6Wzsm/UlS5nexU1kCnJ9zegYZtjb7P3cVqp8f
MzJOfHVShkdv3ObJIMaxsuqJK9J60GwBgRsFv/mexBA/cBfhFRqLYTop/NhZxmHG
0JyFkPB0iEe1IeTrcz8ihTlOcy1MtCBBLzcysmjBUQLM5ZqhvXWZGOKk6uZO5KXC
2I7FoIQ5RqumLFqLHrYyRpWMdHnLA5yJjrlk7n4SQMzff8+yrNxZo+q4+tQ4Xu85
DXbPsmejSkC5g+H7LyhsDCTInhfSbU5AU3/ahLUBz+gw/Srob/goxgx59ZkbMQTu
10qbWDz3B5m5nMEww/Y1WB25fk0h/yvLvW0ZGpcPWBas8JAwO5t65hhrAlEjxhzO
lf1+UFGv5qKRV4lU5ubbBUPSv+Djrw+wZ3vg8kWzyz7G1wC3vOlOXWr51F1daOY8
vEdgj4Zz44Hsbq67LjpV/t9ZnbCOWIdBV6tdMUg78DyyO4FeWYU8gDjFmfDTS1kc
FJIj9Hfp6HCh3UYZsieCXVSNWSczJYvKoVoWVNeABpSMRLmG1PxRXrlubg9XpMVY
qeCmUaChQMJA46SvrHo1DuSyD7qPyStjPQQAhsmyPwS2BixtB6vrwXypog1JGCoa
opHk7gTyuhgZvYkhFS5DxCuY5IGSTxzvVc9QOm4kToZU/5fCAQ19zHPHuzj7apTm
kld8ZJHxRykuqvrtaqqn6b0OIVwdXdnXtiDBPGrqwvxzApcpbWYs2Zd9OAV2rnL2
psIA758ujKIKBmoUK90mUO2afe1oPSjxuGRaK8a6XQ/eHWF/UM5tPNogl99PPz5S
kh/BshPryXgxOe7XBbTHinqvVHXEuieo9pf82AM9+O9BIEmwX4UpkPT/X/ysxwA4
AmjcNnpSVTrHQBA87kyUNW/7vN9lV9i7cBxU9o/dyJtWqPi+eK5gOJ+i6w8Gs0D2
EDwwQOlJYKHFyxwraYVoeBR/y1x4bSiD7E5rRqD8588I8B70zbQWXtDzF58KnAZp
8ZlncBHsm2mQFBvX5CTZgD4xtNo/bBTvIViHJMdOkaIT4GStX1lmVoavyrUedc1A
3D5AlH9ZVbYxN9P7TrRqECm93nb+7k49Au2xxlAjkyJOVwqyk/nlgOc3INPUkUtX
lbMaE0PoMrMc/CdfiFhUqHx6/q4pUJk7G5ECupPusSvWUdOcRXFD44JQLMxGiZTo
XfCZUnNdE4iJxO2unodwb0ehE8f611+tG/lovSq7TMcn6BJD6y/pgqAggHh88UyA
ud/Bzex/SMhAJTHEV0cjW0C46UtLKFJGyuABleNCxjK3O1L2lBPCD1Avcx8DzAcI
dFxNUXm0Lc+i3IwYcJi9lXoKBUdBT8MfeR4upGS+gHdRCGNTRTPID9Qi5HCb1Hix
UxvWnKdyeFzU0xaxmEcvDm3HiXrRYrvX3VBi9o7jXjeZqllmoIJkhaRt7za+xCO1
m/khWRSvIZ4eQao/7A7UOcS1h+x34CS47sFTBli2DylO5x6C/9mwpDL1cON8FWg0
7Y+Yaa92I/0C9cMmnw4W/iL8JJxqBdS4obQMAbly3luYb17g4IeXqtrUUjSsLfMp
bpVnXXARGGCMvx3Fof82z53oC7SN/WHUncpQE3YX1N8pw7HFP7wMN+ky+0XoRfsA
z6FuG996yMkgQha+5a6BOxiuTfqgpWzzO6XiCVZK/YP+jrIk7Acy0OgIbbxB6v06
YAWAEKV7TV2riidCw4gNbRkDRkozJw7TRaDpMfwGS5QDMv5hihq9QD30WxtIKNDB
/NzXlu4/10PH/MFkYQvWnDLcXYzXvZk1BpgG+c5CM6UHcoWcd2WTIZ0QVkTVI/+s
7ldvwb29bZNwUY4NbXB4uVfsXjBeVWogKHvSkcTXIyf5l18LwQdC4yPYfBSGhkc5
VkY8ocBOJdHhEGn9Qe4NSt9/aCzBe+1ndMtpCfvlNR6LHMy7L3HK9/pOmSk0QrJ4
yZOIQYrrYohL+ywefbJKmxYBFFZjMLoKTicsg8+7rn78U7VCqs4eVFtnEZ8b5OAX
SrT9jRYQug3qkN2iiydkor4UzH0EfCrBP7Zcxc0wA7WSPwSvrkmD6sR8uvxDXNSg
pE8xTVZ8++IBs/510a5InDArITi/S8CbCuAJYCPm/KbwzMI2dXMFHCPvuP11U77m
KopqwneX7RHuJskyxy5DdVxVbfga9hsGoAexbHoIkA2wmtcIlVCMsmijWNyWfrcO
kbkV+UwOQSMwYeQ4jX6W+dfyaptubzU+lwZ/jtOVazF/JXpwWlG3iYGjWNTP13gI
g7jWaWFkgLSupRvFTATMNDkJZTm+WVjLqTEPYF9s/odiZ78WvtzOo9o7Z6xQD0Ql
hUJTDigJoCb/w5b1+os4WA9WVvYD56n70taagyXmncX5jl/vFZP74iPUen3AQX6F
/Z0b22fQ9Jem/LVF61P29z1ir8BLcy4KSiTM1BamxqhBgNLL+4O8jJe5n5NJwzkM
ck122ZU8vYcUfshwoN02GxRrU5YKwYTGuq8za4eeq6++F7mQXztU/+UFY6PPGuWX
l06mOC5+fTcBvXbpVJOWwDVLLFUZfCjJ5ZQ4+Gk+iiFJDOVonqhUUkRJYZCo/cRY
9O4WQmag8Dnu4IezCRCqrvMgksWCdO/cGV5Ei4ga0YsdtQciwbFic+zusQreZ4BJ
FoB2Q7/A06KRUnY9zskopZHt39owQlUXrrayzCpyyDl8n9azyENnh9zEflLhvMIG
EnYhF89eDpPY5bPe3QLro8dWaloOPDGw0ddpP2nK60cCP4K0jt5xjAxXV+n7Fvzr
UsFIPe/YoiVzG8UefY8amTDV60MjQxwJyzXJ+xFzhHC5MP7ZluD551Vryy2tDkGo
JNSxIa+thconvADkz7mwfgQEQ6ozlNBkhK/wel8TwHUNB5Vf8b7Ij+iToWPN04by
/poNz0ugD3OF1h5pO3iynO3ELtZHPCUw5ktH4uE/Tg04l1PZJ0Y1c8FjAvohA0rg
MrNDQpebSOZp9M2zOIksqWqVU+S7//ETCKUzaWKpU4R1B9u3iu+vdbzbLyDAbkaB
HSVJEsdrFZ38dEXn4QJBALCu/+ccfBzozTxvvlFnHoymClkHpJcr0lCP90pX7fnc
jU87T84dKuBHjNymxHkyKD6EyXXGD8NhK16M+9tIK8sYlEoEtAXEWonejYf3bJTr
AoZ4B746ZD7UqAsNdvjrCDI51QhMLNYixTZd0zN4DHCRzN3AywpGtAcmkDPedxDi
Tt+BDpV7UeEq6iFSvr5USkZnFCtDZHj1+AwhRR6xppKYgHKQjh4ftF3rsPhp2FKP
rK8H3xuPrOkZZ0HSnspvpsC5cYSgvChbJE8pzQqxh9MR1a7y85IVCKXvpcBrC6tn
GiHr0q/Va03k0cvHfeMQxs7F9CKXtjZsREj3xvSQyc2bKDqjp7FkTPyNSv+KQJyR
ElPR/q5joxN9skoMX5dbZMZpiftLbWk6bwjMWdV6/WQSdsvvTVC+fBW7A0crMnTr
tPx4tLQPCM5h/PaFUHejEbU0umWKEH0BdI8P2AbVbuoXCobzC9Ii7LnmuG+AGQRc
z2GynBiqR6xutBixJFlLTHFfm0QzB+M0R3yzGHFyv6DJcizfGit4J4dkHIpZczjI
hfoeDCfsMLHeuwajlFNCNpcZIwO6ir10SlzWeXeSt2C/e3Gb1DfiBEUQHvDiJUsh
PY6LO0sPRXBZAY6TYABvolVOY0NHHO8IS/Fq763LnvXZltqMS6HL5540solyiywV
/CAa+gbTZRB+ihNTRaYMtiggOAdPiMRfkHts1bPZdQK0unRp02rtZY6eiD1/zX85
/r0LSe0WBBR+WfbvLuGIY9hlJ7HrRuZY3bfC4Zb/kj7oMG0DCxtXZLb2hB5Rv3GG
MaGXxQiyUTqbUDuPaqbj4HcfEAD4u9AUesz8F76DyncQlBzGNAkHHiyOtFah7lCo
LfIPODJM0ntMsK8OvOG1K/0N8lnSDf7hmIel5rd27oJMD8gvwHztZUYT5hinxKqQ
DZtA8E5DXGB29y8/AkfDX0aWzFVkvCHvKstB98RPUClc2IbsrUYW9rB5tkfD/2lm
b6K1kn1/U6d82JtQduG+DmGVYApDY6KhtUY9sqIECjoPIIPF2VUkIf39ZacFEEH9
52gWnLC1I+tjzSfasa4XpwzQ68ap0UjT/PveBbmuOb1w5sHUDxwgKBjjGy/FQbJB
/gbMcvq2CJpOjIG93QoQB4DzQbS8kff13VZLAvpvLEAo5pLfjshk6Vs2WoP5M9KP
zk9dPNMu+db1k1SyrX/zHTNUl+T/A/lb0BOYRwBZEzPL/OxKf+65xYzWfZZD55xc
AkxkaQ1nMJRPbqO+5Q0n7+cGWWZ9lpGFeSzG3y9kHt72AFsZydDKANBeJVHs8DKc
EFL7OxvQBl3Q/v68BOurfnFu38dkiUkoNvPdQShx06CNlKRqpCeThUsFUWsnWW11
g1xc8UJccuKId0M81X/BdxL7qJjz/qM+iJTyJg4vuMIO/hHIRGSzgSLJw0/gSNJ7
cCXj+6+hpO+n3kTCJGVef5LzT6cpuuCKiwcqt1F8HjevZDYzL+by9WnCflVkRmIt
PIjLzY0K/rvsV0y8fRFy6ktTB7bIIXzKw2FhB5p7OyUDPnE/4/CM5twZIPsDadZA
0hFL3xeNvZIV9s7JFYe0tTnjQtI1pu2KXNHcT8NnYyTZW9VqKadYpam0gP2A0kbB
i8aIcFIe1V5rIOyIcrQG3GswnjDr5MmgPTCSdtvFpCbpEIlP6RbMRFqUsHAVPzJB
glXWT4SEW2DtorGGLh23AOOXL3fZ9gleUnako0jFWqrWKiEAMPBL2OV3Ed/9AKSi
lV6fCThprc15fEN/krYrDZ+UUO+nbj9OsJt5PQbCn5WHpPVJsT98zVo5wViFyjNs
EE3EcZL1AtLXQT0yeqGkA0dBCUOoQPtIc62YtwxjaPoLpno3obbaBhC32BQW3gYa
j4VQa/IVppv3a1QgJrXcLFDhyapAcf2NhrDP9hIxIQNzFq5ZvOYZvW6q/xC3rL4K
VVGTxB4tiZzV11e8fEAwXYg5FhbBzhfMYThuhcMVZQZy9jozoIg+5bKlXv4ioYop
cGSGYOz+Uar5lY0flc2bDMLRnntGBkOaGS6QAXitYmVax1YNof3EiH2YSbKM3HQB
lM+cR0qk5LeFVBGzybjW6uG3Cnu7x8TB7SfeRGLniZ/YmU2C7/9HoaVRygtRqoZR
88A5bppP2Dzsco/d4uH1POBXfvwW2EF0dRV+meY2ZWuIVROBloDrYFt+otl+47EE
VJPPp39ZWTScD1uCfjTgZOBDKJ+UFLKu0KNuRkV7zpaOxnKBxE+fP5AO9faGeHoL
8gQun4en0aimaD0/fQS74MuxVsKJXHv2p4RLg/nHzgOjFHKoZJQq2ojN7+V7dSvc
3n40rLR7fa7ofpFOsa35HX+izCH6h6YNaAeTlilrw4v/bvunzURWrZCSOl9XqnzM
33mko1hz+HocpRt+65YAKFrEMd+oRc2xRC7tcueqNEVaHPcu0vqKCv4be5iEU3BR
3qRjh7GfD2hhP7dChFdgA0tSJvjwtJpTynr4VwN8I0niLzRAzQDbEjLa13iUqjaX
JVN/gc9oavI6F5oiSF/IefJLXl1eLlgTbzp9n4XLOIgXfgjl/INdrt4n90Dd0fvL
SwKv88oRoh3mKc4ubYoFtzYVboQoenACJQXAj7IV6Isjygn3Wc4wwgztE39r0Pjb
A6oLvczGiz6bSIUf/V1+N37XyoS4WeNQ05/7L+D0SZUno9Ctwaq9EOKZQ5C4h2YB
+dgXGBsQxUZ9egWee9hH8sFIg3Xaadt/GbRaVxJWA9tnsvSh195UQSP1E6/2Uw/J
fDXitaU96zAMu3y3un52kZOVk0e3O65FbOV2WZZiSueC/E3ha0H5C4sEjPNwFJLD
Be1EXLfshekrT4zS9PzCkyojbx6ukZx05rbqkDz2R1FNtNKQiIk29cTxAjBntImV
feaGjZRSQMinIBw2qirJYnBsEyvZZiIOT/sDY8nWrtHjBrvRBxkSKFWplbT7y7JR
295L0QObEKRr4fmosWExV4MNnDUqgNqivsmY6rOryfqq8QFbUasveJOLUpV1Qkf4
jIelUtCdVzjRNPPGLz4sdsZbD266RHzWKCsOhQp0xPTYyNSPa39xOfhKyo/4Qjf+
g10te5Ocq2GkGuzV/wozjE6+x9MessaDLnibmIBbLkf8Fx1itHouRFXi57Tey0vI
R2s3MgQ38x+KopN2ecTAaNjtZUM4Lizlq+ItVBYSKxR8qwQ/HaSiq7zCdYuDHhcx
qHjlexxO8IRU9RpMtbWmBNu/Oj+2H8NS9/XUu29GeVHa91GO/8CmGC+nMJNdgJdl
zEjMCwpgsgrcdWexcZNnibLXmXEPwPQP3SAHJeal0oWT7BQZ01ja7q3g/6Vu1cHh
jGhzVmc5PUHb8fEmR4vBgkQQ3v5FXCtcTcsHaBbKVwY52jAFhRluX4N4Khrcx0M/
cWLZ562S2dtw3uICbvRvrRQKXgS+HMfoFCK5yeA8Pqm7VIuwysnSNyfXVVsNIYA4
RMTso5ClJfLsFDEjR50ZlZ2QxyD+I/vNoGbOCQQYwqICMEoMB2c6sDFUwMrwMD1D
An0EPuDtZhgWiNTTYRuB9r/iWoglOP1XUY9oooN8vAFR4lDs9Z8dGhuKRx6wweeH
CKoZ+dXb2t0Vy0YsX86Io9TX+1W2uLKGg/Ipc4/o6qB6NB/JYfmwfXKBRh7/seOU
IVH2qapxWH9/oUcDeYLxul6SfHhs8Lf4QWZd7Qu88hO0wx1acXQ5q/VzXdgdF4Tj
QowUHUkgWwBMW37gSmhaANxaO8/e6PwV676iNbE75P1y65X97nsMPYSgb7zNdhpm
XoylKOkYcBbzgFysr2LskP3wkHBbsrhXv8qDlpxWZPXiTZR1jQbFinp4VyrIdRXG
Tk8ILWBaxQ9jDn6xBv2NXLdi8+3kYyQzaEu2SO12L5RCdicFjFLmZpgJh5oobRI6
DV2uRe85N51oq3ky2BkLLt7j5wH4BFX/HQD3iuVJfCrGLp5jmQEznMi10DWH5BX3
3jmRw+6SbDcNkNX1kcFQ2trzsiN9sSVZui1XjDurMzUd5iZ9GBWgWH8v9KY6yu1Q
D+PWVi3jgXEyuWnXeku0nBgBWqe7XegPfV2Hu4AoQkfTO+kDeMK4hR+u1Ty83Qfa
NPUNcZjmmJiiXMu8LGwAZWnEXMq1F+eIyk6shDoWChkLBvZaYMNWcaz4ZbzOgDfI
jEqiHT3X7ErUVkux9p9IyqtnPgmhBhi5VfwjJTqMjappurmxnnGPXukw4cMEbw/4
T+QyEHUsNumVPA9A9vrb3Ilze91HEhRVF74+cZ7EIpcr2G7Hgt5rvQRZPQW3da/A
4i5meLY8hH7c/lL6W3hzaUO03ZaPzjBoRa8/dSBl3C2gaK5TcqZ5PzuQra80zIfg
IWW3QRqosmV42DXSf+WTxP75PyJaf2NCjfhHsHPJGY85e6/x+OAwgvxsGouyVwTy
QfFM4WbaywFd+zx4OTr99z7Mt7mGI8yuQbpcDDa25GNDX5ZuwLR9PVfvAcTmG0QG
a6nCTwg5j8A1mUdWAO8TNjcf4Pao06ANu9fvdU9Cp2N6+9+TyJlg353TAPNERFf5
lTpgkJZ3OYzhbU1C7Cvqtpm1WYA62PE96zBF2NdgKbHE6RTHGNPn2QQCrDSADisM
qfkcxSbeVoryDXf69cpyco0KlZT0mphJ1qRPWiwgZAnbYWTFtebItRAApW+IU6/9
65EfmWFZ+ZKG7l481UOXjy+2JHM0ouRZbs4EUqrN8sl8hj7ZRoywNMqUz74LVb/K
dg7FraS32gz4jlog1K9IjoP8/k40j/CCjga6a4klvoMVMZzY94hxJtZDrp42gFmt
skJK+yDhBZCS7NkKuKwISHnaNo3VKfcx5FTwSp9tUPjUONmirbmad9YAdcFDkEfB
BgeCC8d+5lPFbfJsetsPv8HlnmZ8VnKz3wbjqzYVPwZtRU9NiTPWBB+18AnU8HgI
lRRc8JEccM717rv0tKYQSVgZsS3X0sKq5kz8YIsRe+niUC6truC2dxxepqTqXAph
TkshtT8R7dKWsTQArnZYiGIPo9zgFz44oWLhX6q4Aonai7g0UWm2bkoMkJwMlZBy
1A+8YJ+LDYDLXSLbs2qvp0Vgzd4eSgQI4I3FgiGdla8YnnbuZFKyqExpEDClEo3W
tnjPJm6ZLxH6ftHGNSxI7vBldKP+NF0qPjrhgUh8Pupt0qnB2CMFACzYWeHDsOoa
QWGUvg5iLqHwsVw8AbfuukWnqoKMAbAYBMvC+pe0yNWs0+KsaYw1toVbepy0w7FD
5wt8LXIikB8tUWk/NmXNxEgDbeGAPzFTXJjWMViQIPjE0hmGievqenYk5diBNRMp
6mr/bspyblV/+9fcDmwMuDy/GeYdbuQw3Ww74Jk5CoseMEXo2Yjq25xa52UZ4NWC
3OVWZauIh7Be7J4nspNaOeyjloWi+5/qRjYf2dy598j0a8ztKLVhnFo2XNii33hr
sXntyuF5SIh34gXG9QI1x/RbDtPPMviHTr0kJOBvtPGAoSRyWQDrkpoFmRuYazhC
bXxezeiMMAhMw0ole5Z1rm/jak2+TTHyVZVtbQBX6ItJyHf0VX3y+LKp8DCq3e+O
/SX0+IiXlKlwEP3hVbwIllmbqbLR5hg6/tHqi6CBHVU5qkVxMBt1fiUHB8YaQ/vb
hZVmcZLsW0uZUK92lJbQ1sEmx2GbZinSdPFDLUf1pXbf73drJb34UgLO4cpY7lW5
ktMDGdEcvzvkpgouhQEERkczLR+6ztrMCX1bjCrhwq1ax6qJlS5XPgyfu3s9mwV1
pxosI8wXwRtjfGp5dbf2mrctAcTf4G1duwAVYhGoW7HgdQqAW8IYxSzdVtyiCEZn
CAR0vm6sSPtxxm3zk0ABEtFHMoa+m0S7MZGzd5OqkPYx5B4WDgvFFU9A3mSZfm80
0A5w0s9YmDgTNuXrVzCIqWT2bwKV1zoAUnMVc53M8+7r8KHKdjY+iJjmpUkA0JTt
BO6LTBytY2F8YXCdX6szleddt3NJjr2jU8SMmp5+tbI4FgO590RkBjYozn/64a3d
hnAt8b8UTDGvOE+FjNpUbahO5NHhw91J5swAbG2q1/3Jy94h+0/PuqUJLyjYWw+1
I/tzC0itO8NW9HFFRDMMNBlOIMl9+YBCScVIosANyr4fcTVrXOqIPBoxasqD+Jfx
gOr3+ldhdI2/LpMoz4h+m7TqbB2Fm3WjjsQRFoVV8xDx7PQOifLiuQBTmzKpxgak
TuAs10XH47DL8HJ7G2OtLlGjKy2jwsd3g8agBtGijgZ6OzxY2jRPZw5IhhJ9ebzh
sLRcZfhSrDcMLqDI4J9kDbZyTAwJZCRL5f5HKSBLXetvwYopMp+nPr3BEn050ncR
qcsaiuLg+UpWc352UgvIyRETz10B8IIQPX3IspL3CLcPFKRPc4bqJMiVF0N5BQt/
/x+TityL5DkEomUuQBzM+/6tnI7HnIHxsVZORWxKpdDVg3DzUk0sHneE42ZAnJcV
mp5amD8aKZVJFSetysYNzCdswJM9uWgyoCQs2IjCjipP0LC8z8TL4h5cgC1hnvuY
C0qbK8eUYe/lH8iAi8M0ApffFp1ZsVWurLLa+HlOjxn82LwMNGh+mjK0gDopMZ8g
gQJqkzG7+UvS08Urc6Zs7P9mABqgpJ5WPvod2CMDs9YHmUQNRUOhKflDQpiRshLK
vF2FZZDn6KIuck9hso+AAezWaG+bv1PjfgDHh2Fb1v8k3RmOgINrExjHTBzeBC/y
p6iAIAAZDvyPiGzt6MJp4B/CdKEKd5uD15RTNivpzu/Cu1rK5LXyaiKow5f10dPW
EpMU1gXpViuXW2TvWeQixL3hFJVw2cZy1sYUJtSY9HZ8VkaZlLjNUMucaYx8QWhY
eywsRr5W6CPztiA1+pZmvDkT5L+DbqGxvfJsHDju65hdMY36xnRcQliZsCE80fNM
H87DvKhoKZznNSFI3eBqsAjI2cv5/BgKDCJM/ycIuDZd0GI7mMor0QTRj+ya3sGs
jMcs0IdJQW3MmuHNknU8kyDotC9865wBVbd0wtC/80rZYnkG9xNSKsdoBZ2MkTq6
5RvwDUIvWvX7P3EmO66JIET6KNnSGkFL2BedVshvvXuvqh/Xblh6uV6prvBAVHTo
oNDZB4ILnGl+xQ9Alo6HJx7UVML0uLF655RAmofLfVGbhopO027fPxP1QHi001xa
vey7up+lA/vFLWbsK5PtcTmKsGii1v2poyhhk+cpkopUOjc+YIm6GmI5/tpev5tK
PX15zwgOJwhqjaZxbwrm5m85+/kTHLTiZgioNteCf3n9vEl0BaF8aOk1Jk35Coby
znHctma/P5nlbmgiP9jBSTZ7ilkgDHtmPXkuzZeJBCN0q7t7CkrrG/W0dXQ0BVnw
IfTAyQIphgNLvTGYr+EeX3Gnx/eR5YsiU8kpBkdA2+O8n97IsTmTLp/RDL2nH6Pq
BcssZIo1fUOsEJVBTTw1vOuPp+CL31YJBARaTSldDwY8uQ0q0FVf6sDiWBFEtl0z
lTHG2MIV5hDAv+rtGevGRb6X1KnFpoZWHyFZiSpm3iEoBl3f77PQDq4wb79XTWTC
OnhhkGHT4QlQyAVnWVxK7niI9S6HVtbH+9pE4v1CsOsTRmurLibFmjf5VelmTTa4
vZcn3aayXwHEnrqQE5dAqs2Dub7LfeH4YLAWVqYX4wsrZIq8lHLW9F1aHiklWkGa
ocTYkKZ2Xil+2kvepaCwKmDhPIAL5j0I0HXSvwvIgHoFm9GZSbAc+v8fMg6KgppP
nf6AfhY2UTZqZBEHvVaTYd23bwWX9IRcq7aUXoR1N4nh4AYYXregvVh5NKEhkE2T
8hcgrsBjjmT7S3OKIYSdW2eBgNZQNVGLWqKnoIdmsxv8gwisWaLHntoxCKPfO9UL
VFM9o9UOv6M0fysyg+9klalaeWTb8e1tanOvX+AR1W2ESwwFPMNPGC6E+IVS7yQ5
E82DWgW7XB+s/FjW7bIXiBfcJqA5bMbKp2s86fctmMFvFyKaAwfbcgr9McRB2G5g
rWpASEwj9aVfLL/XKC8LUwIL9ZmVAZEu2NG7DKyH5biZwZyQhQ374hjzM3ELEW3K
XlYM+0BbocilHWlnTq/jEKtEcOT+O0RRfF5tLkuNAPIMbPKJMClEk5D7LlEkRpaz
vGQUZ+nUgLMklAhqJ7GIEQ7vvqcPS9M44CGAj4dAVYwZ06UTp5YOj68uX6iDKqR6
TXntjeNWdPdwPU4XOL1czj+SSdge7x2SqL64uiiV4QKAinPMfN9iDEHtDNMPhaOT
t9NadTt7Q370FAM/uYMRlGnVYZZ7uxI4qu7+XFh5Eu5xgr6BpW+kuwwgrxETgGdu
0oHmbcnS7D5egKHS1dPfDoe6oOEDiONlWblRTGBB8PDEY9wl/5YirmI+W5nmwO17
C2SEeU82QGaV3gqfcODuImRAv2QhFSgQnVFsqmPcz0H4Y0he5zsEJEQIMic5pg6D
NAFIxvOdrtlemZI2t4cyblHjFe/ABJM25pfD0DikxVEN8/jsmrmJy4QipEVpuMif
JwFEc2pTYomK21qA7rGy7T+rFSIUZ7k4tp83IxiGTExPxY4hROgTmxg8r0KqY3FX
aG3QgnUrEbqGRWVq5/IwaZk8nPQUBjG79swg3dWELYcdOr+hvwNqy+T7iFZN2dBv
bGKeXJvKaYSQGzV4XFVubKrRn4uUAudaiqCBZVYAmS5qjJv5ZdT2pTIeKJ7caD4P
WagRJPDJ6YjE/XMcgvfQSUZJQ5yQJJzTQQu8ZKGomAnDrBn/zpZL9miUnnbN34wR
xIIudLisXCU0CW/qgs7wwdEpAE23I/f/Pe6GBmg7GRKjqlH7EFed9+JFggUKArTk
jUhryqb5jGzDOCcBiMHEvnxyvkkcbPzED43/kvbHACNRjpYrby7jzYxuyR/YF/3S
LQsbi6T2ZOSxA98BKiPsaLLFt3e+ZAp8F5xTNucVuQ5T5OLeZbtBOVZ34CMeOmO/
JvMiJ8YkZOzXZlNDV4+3J9N59CJmsliSmO3AQH5oQs2CrHT8tRyUn5IcHbzSkt7k
RNHJ0j7F5ylITA/xVKQlu4bV198fokaBckMKZCdHG2tTmS/H5jJc7Qjd1oJXOusH
M+AUaPvEdj0c758+33XSggH2uMuWaVqbcb319quqCRdXBQbIioYjQKt+kdIZA5oI
10OS1A9gNLESN5nNqfCuXiR9I0JfXWe/efgZljUP8RbKrGguQzcm9o5UgCAIxRce
JAQtc3q1Z1uAKX+vAblVlni5qG0ALDR1EWGoscPykxnGcwFsZKr5HY7laJdzF8Jb
7TZBTkev/P/pY9RVJWfdQfKF/sbVpAD0sXQAQj/q+zbVTzNS5EJbWnEemaVx7o0Y
YDrAaJdnYPCggfs03H4L/up+dWUaLzGDJHX+7KLB/5XHuVAef93/Id/OFYLif67Y
YFsHUsz6TH1+NY77lit5flERpmhWWZiK3GRz7mHCJNzGpcar9F0Yx/qoCWkk0KdL
37IBDI34zmXroUUXyuIHphaIpJ024k4b/B3s9lQgZ4O1mVTgqIiWMyNQNXJPubpG
mUmad4AKXVux41CNnOax42hxHZ6YYnfilBGmq/IMl3S+00WYJ0hgkfQRxydFG5KS
eXmwJm3TqzHGYya4sGZ2VGVHUHRlcb0F2gxcF13DX2lablIjcdHeAzdJ1RUL02kU
egY4LS2tCKlfwjqZNFieFdniYuzfCpXLY8/Q5iw0tdINbci3/6NnxDJux6RorL2Z
/n3dmnG/sM0c3P6ub/9Ymwf464tZ4seJJp7Z0Bgizb6dnwXESUgZaEvM2QZYV8RI
kduXyqvkFGHpxyFB1/9PuFYz7j1b4Ly9BDaO4ZVhUlf45LIztrMiVakCqBf5ZEWF
NUtKIBOCNSIN9nzb7Iq8ubY7wPnM908iIeDxGZ9tuhgCOqQWKHJxOCBlDfj8aw60
9Qb0SdYh6iNTacSG1pdR+1/mWSzsKMjsOVqrPAV0gfualIMLnKvJwmMzXrCPXDzU
tb6d8zkEGZcyLGqQHeg8DCMCrmcoAAR8cmsyTTdgtOPtYmvGKa6sHZM89XJztaUO
p6WYaUzjM+7VpgRVzzket6kgAIDMr9aYfTI+sd9jvzH1itE312orpWokwOv4oGi1
boPgQbIfZoKmFRleC0uS3P611rEFN9dhfiqT97nXUXJizejx1W1v3WoYVEsUOOz8
a+5cHrrfdnDVx/cFQr4QlAgFKUqBydR+YguuJSCi5WsT6p2Wa7sf2oJx6TbHcVP+
9zuX77pcoLZ6fOzPGBDiZsJAdiek+rf1khXOMRbEdfBPCF11FCXRqWxE6bG99MUH
2HfcW0TBIxNRIZlERqvfRxia1ylBS6xag7NNU0vzBpJEgo0fpnMU2z05Xzg8kRgL
XwJu0GgkBNy2NRpJzvFFsl261hK8LoIgqlvDgPtlMh97hLyRh/311w2Td8LA4M8j
X8vvMFiiKC9mBUB+y01wleGJ2VlZV+zbcyRWe/+5DRqR72pemwfnKmo0O4wQsPWA
2EG4pLOvUcbqXXq+g/PuK4I6XPe6CeVYjPmtyJxVgZxA4EiIpE1JELdvuD2Du4zJ
jlgrwsWH+F/s6XdzfS3oOuleVX7I/T2ake1zZZE7nx3pW0w/Oq7C9qmABlZvSu2n
cpGtRtvoFyDwlKWTjM9oNUe9uL2Ix/8WNu0cqo0X0eIlZGcHSNreVhHqe0Nap5Ow
9W1tpkKeVae2yk3ANWHpLSas9+tNwZUyu7CFH6uFW7bssj1h22RO1n01U64anjmB
0MJ35HlWb4hEaldZumqjSFmDuoa9EDO/qR4VRvx4MZmV1C6e0FDQ2lKHAnhKHAVk
p2usCnansCYK6Jfe8a60C/sIuE+v+ZDwxXC1P1vJjAMhxJ7Zb+0SQdrhQBB1tckQ
Uy2RfNrtkrHZ0x/fVkIh4J5YR39ks/KwuIbvmE2uX01uZExf2SVJv0vYfop2z00A
wGY2wdoqnIHMWvw3/1PQyg6ibKGzGt9TyGhtS6iY8BR9VCTHJ13JKNRpctSo5vyb
D8MClir5toG14dbA52v2pkDzKa0zGB7weN5DHtRX9C+IEY6n5VLAizki6OV362nn
XL0//UYJdQ8abXpBSIPpaSn4h6FS0I9qdzW+QRr9HPwb2tEx6MKPBLH0MWX+DJuM
K6xMLfzLqP4njiiW6iXwtUWEGladm8iri2XSVuOZeIRnkL2EOQkDKDDg2WFWw+Pd
5HOthfBoknS4ButPi5fEH6XgJrmjww31Z9uE+sQn4LI+2usGudk2d1ps9JWkucN7
TcZuVOL3BHnuQB1W1YIoJTm89/KJ7Y0lKnu67fIVLRpH29ApQ7doBV4nsvoFbtj+
+Ho5MBr743+3DqqYDH/0NuGz1GcobITmxjvqvHlve43KGTMQ7htS0tFGn3vee+f3
TcJOhBO8+qirC/pYsnpq3HS4K29WyZpt00Kx/LlPX/wipo+WRhdOnP7lNTdfa2FN
6mrCfRHw15euuL8x0coIC6n9jlOqnv1lS2d1JRo6i1XROnCJEvyfl/Z2QyBhLOLQ
2D/SsvDbl33PqTZGaGWagoaKr2ORFO95TVTbk/d+B86zYpalBJZq4vMiHurCAwK0
LdKsG96RSTMJR8UPd2J+xnFDOTNVXn1oqDdv54iG/5ObX0nk/6cS+wI/mBDplUUM
MML/Azzo4r5ydgwqyVlJKKbJw3i3OIAgbVfGnfNFAowTnN+SNjRe7HWAKcXABSrq
6L/8xEGiS416xfgbhUcTph2LFiJH2Ybd1YOwm96HP93jziTXGTjm9G8jw3BJ4S7u
R0ifTBDbXxllesp2FCApYyByPRFONxYmQdtApVuhup35ssa4SEnMFMi+nTUguj2Z
RrmScfzjmOCavfxYxh3+WI2FxDP4tbzPIGmfkFSYp1XS850szdsilphofZmt9EpR
H36E+eBSsZAOYEyi7Ftxu3cGY8OO1V4JyWlSBTz5nJyozenD9ztlJtnVxWSmXDKH
AGUfLGgIqj0QrEN1yYggk6ue0PjxJ8z7kW/oi0OZYl4ppnyEKl2jIMeovgd4kyYh
CFt5jWZ8zEAgJ2NFmIUDBwx8GrYj0CgoOttO01kdqU6UMlEzsUhzeYwZnfyvSOIN
TxS+eRDm+Mfn5dlBeQ2k9IJ8JtUkQNw+ZiOyE08K2mI5CtxkAbsFzGai2NavXRmg
aUccesj+JdRW1v6i6ATZ4LkyySkQRbM371RfoPxaKpS28nriz8Zq5aY6yoYVh5UV
06C4t7AO/lBkdzYnq9u1kjjHIuCREYDmrcwdsY3qKUyDqcDnEOVPWz3SyKcu0+zh
6E0+W6/2W6/m6uPfA2xpi80jrFaVT7cd1Zn4KCTVk2741stNGfCUiuITpYloooZr
LJ0CxwnV3Wn+Ho9RzQVsEZpCD7sUyG0hBdT09rLjYMjrYdQU3+KfswNayYjNYphk
XLe67eXEDiiW3u9RsXAfrENT/xWQggPjZjO98cAS5pM3xZ4lXXs1HQkjTrcgDchg
mdC76E2hUFZFT3sjtMd3HQY0cRRvE+uwWys0KBA0302G+/IEXsD8Ll+liKs31zdJ
USWGVaTnrtv5cMDkvE8/pr7WivDF4GTzem996QgX89x1nDmQVZ3BJB6WXBQjuaos
JBtlP5vBgI9wslDV01KXL/B5AZ11no9fT1uIOa7sK+oaZRnReSfaTCDCDOtpeqj+
1K1/O6ej3cacBSoFkTfb6U0zRPsotBibQGSVnVJt2xhf+mJ8jL+EIkVOUK1hdWNW
vCaHGHZswRXoHfZNp9qpsfIssDLsJkUw4ZDAg5XqDTxg3XhHHUtnrcd4WlPI42B/
LkDB/2GOZQAorDDpkeG2KpwntihrZk3cUahLffoE/n/N2QiW+i3NSeWhQHywM3SP
1F9mX+I2N/qpAWZmHBQ4QKLC3Cc/qEYBaZcOMPQE+y10UPEbEUOAw6T/TZZfjDQN
8HQqdlDs1hoiaMw39PXjxkIlumoCb2mHxszcWdVq9IcZoFbWjCn6bp27uyvDAVLg
4jhosZfxA9t2/UCR1sSGHLZQCXRHe04JVtYS1GulcQokeibv2Ft6yzglPq+jq4KO
I61ZWp6KTkXHgY9/M6dtBNV4SBBgE8fL32d59h8L391pjOfjfuSzXzyEWujGKj+F
/lQNi0ECDVtpUd69/koG+JPwMct3CKCb49gL5J9Du4p2j4cdbuF4y39YI/bOxWA4
aHltIaIkr8ZPXMwWEEBBTEEhUTIN/N8lxCLV/JNGXCYc0SZ3OPJB4DQdokMnJXsB
vsn/bzKpcYN8usWDn6lODNKF5oA7NzZv48W8oGbVBypip3FtF9lc0xeeVeNt/87E
WJki5VwAh7oa1sdVeqOXI1y8CyWhMtDDFerHNlpzV22ssfimzlSQ1nGtkNbOURBw
hQ+J87ES64YGw/T99HBYwhmNsKMM65E68xLSyIxzIPxqQ/Y4C9Z6gutblMa5BcL7
u9DVmXYydiUe9Ifhfrd/NEATpNW1gKVyZafBu+Eti4HGqA8tJQpiNAatQp/4DYMD
hjWVpZYP5IOvmuD9IVaykDxfzwzRQZO2CFoYomZy9mxBW6coY1L7KeThzKMl9ApT
wbPht4knM6XNeF8QhbjYpIMQM1iX+azoyyaBv/c1mLoIDxdnXnOxUiu8gtFxWp6B
tAypsGR9t/E4Uo3U4NTLP60kMz/+6jxscvENlwPVicuMDSnqnVLOlLw1hCIEe7ss
55YrPRw2Ow3toBw/cIP2w4i9bDWO+JRmNjepHKzFgBgxVJBa8M3mdPQvGD+WrhjG
j0KxQwW5dp4IeAXduuD7hnhDiLqULeFCT9zJczTstj+hh4lmtMnjw0yk5In6vENu
VyQDSBpSgcPzpM0UWbSfHQ0oaXpcbH0JCuRCYMI8BtlbfYiz3NExok/V9tnu69dZ
UHVt9XJccnxJyHoRv/cnKahDOkmq2fGv0fR0Z36W70qKQcHe/Wa7uYnSS6qUfmVU
YBJwk/6TOjdz0fZS0dhmi6Pg3od5KF38msm9ynT0VT+l8d6QQfONS+CYZ054xGdB
hmNpPjIIYU5qX9LBqBOCTCrHFtnlITuupKU9/R+SsYjhBNPTYIxlCnWR80AQKPey
DKh7gH2m3hGNxhilK/cT50hC/6hjHNt3vovbdwIyxRlGtOHjsyXWeRj9X7VOI11Y
54htLEE4kDtrH3IO3VL4f2SMGn1+HwAHSm3xoPrmLMgpv4l67INXeZfhHh7qLdhO
T9WLbczfXlEPtoMwhIonGwr9kZuT8ht9hgRO6XFgdvzyDQqmRkvReg/al3ULeDTv
FFmw5vUC4MAmgHGMctFDm8ely3yhBbJ1rJrfqrmJOET6U4lny5tYmSVw7W2NTwkq
53cGtQm30Ys2HsOTxdW7uzzCbtS9/TV+b1S4OFemDqW4JWbZHF4JkIqi3kxaW6W4
X2Q5dExAQ6GraaErXIn9qyUVmyFCFAXSl+dIvE2VKGLdpBKdMV1PM3k792G/OLJd
F+ZpWEePt07LwOFkPSoWPjSBTs9lMmNF1OG6RwVN7D5Eg5DnVS3z38DRv020QhqL
PLi/fV0xNswKD/5LjsOHptOsi0ieesQr7ERQQ9TiOGKhRFd5dMdGy73DA1sBtqUS
qlTkaTVSUhvUTTQzIfdm8ITh6WXlCaXcHXwucTFmCn5hO7p0AFsia3gcxjHhrWWK
3TDHwAFhrAo7imEcf9PgcXtMeWd9zHSYS2l6ls+FKbAJF2m3i9wu+253YD3nh7yU
E30C6eRQZkAGSmwgXP7y48x9MEaw5huYyTzjR9g+8z0IGUQ0AYSogNdFmwKoWt9p
IFmBWaGteewT6cZNbVI9a4H6LGcr9pc4t4NcveuK9p9H1rUCUrRA6u8HL91L/Hl8
wJaMdIo5KHmNdAztHo/8q3QAzJpbQDoNZSubv8Di0a/hKtY/gWoB0bvGPfB03lSY
IgNEPCsqJlOd/f9GyeqtLDNd9yS9moV15hWpggKWdL31S4XYFiCBJXi9DO3rVZxh
sN3ltJAHIHZSk3fEm8ynahvMi88l8Fq9OkTiZvPVoi8ZwkmWx+nr0TtTeWoyFlzY
vZjqr5+Xo6RA8itCcriMwitob0gDvCUl1itP1WHWDSKN4bOUtK1vbuM0KRdbCVl7
jf+I4HdsmWmA/6J7FVnHMZt2yCpozFjhZZqi5JS/ebEWySOJnz3dc6G5b6qujw0k
IeP11sha+Eso8Jzs5bY5zt+rGBkSVhBMZhFNli/BM2oJVVQYTA3GGw+y3rN/+Hk2
dorjj5tFjYOW3QPBUP62MlEWvO3YRByk8VlaF7pGnK0tKXZ8zknr+yJyEhBALOg8
UMtILdgdRVEZX5mJErVu0vQrlPcMNRqHqEaXdu8qmvTICUlp+6D+3wPDzhUTN5JO
jhg39RR8XtYzgP/vq3SyPhrFLMsmZw1KVzoCUePWSikNbIABnnigpfEPlztXALzo
wP1kk99d5tdIiZscT3DsEAAASIjnQ/JDtfcjp0UUEvUR3HfM2Hc5/7Vrh/5uJ6kq
l3aU+zH+pkaanXiOyVI05vNlQHH07S+VkB+18zNHF9420mKMmQiyicaFI/sJ9WD7
nCawHQdw30VNGl15BxjDLPls80m3MypRqjYSBf4LM474kn+RLHUiQvcujxU/AFoG
sgxloRxbig7oXcdiuytvH4GAZj38nVuLe9FmNDuA90uOxxPz/X01bWKQJfhby0gl
MuHmrjvH+2Vn6zRecBISRh5VGzXENop4rOOD/bgsqK4cZPLtHVi8wG/790mJ9Tv2
xDgLmOwcmK6OLm33f6wGatFxl7+/d4J6RT8xHgBB3BlnHMMN1a8MszJ04BWo/85s
6EzDlo0pyfwODDAAq8uJj2bZIuj6X1rPDWpyXHo2TK7FAo10qxnsi9GAGb830hMz
B1T6Kd/205g6N6WfHwZ+YmgG3i0FsmTe//Jw/Eukcbj2Rt4jgcb1QQr02KOhOUnJ
gK7fkAr/XfWT3waDppTnQLuzOzTdIodcVNkumOg2oHVa24gs8qYvpZTUPqc2WZg2
b6khalo6hZEPJSawUP8jcgcnS5SUrNUPFld7HYeexatOMVslxgX+Jxgl+OWmPtXJ
7MZHT6LRl91OgS26oHGM2oq4wHcE0cl0xQXa5w0uBqmBAjVqtNJBF2KrmyPg0cS8
rMnPzI2p/uafMQ1BQHHvCAlZl0zgeE4AXVHIb0EZFJi17TbM60txFIFCnNzvFhG7
VaJj5UQhnZaZkjox8uAJhr3KyKVakfsysuZoJ1BEMA6yK5txQQWPofGYhyyVNNfc
3I6Fi9FsEHG71VQyTK3QUDO5e0PrSRNRFqB3zgV1ZD76n7wEfpc7zOOnDlMN6gGS
M1Zc/wTp1LApXCPQccp0M73OgLdrfk2aIoz+6vVqvc8d5l1u1qcELpp4FFN8mGOd
om1BrPtH81sYGFttqWcrM3JVnwv/z6KQZsZdDnBJVvm9eog/LMVXvXASGIcfWiK8
gxo826N2D1/LKlpP+uuZCN4bN8I5D0Pt4ZLE3tnPtZWJAW6KPWL3nSEGnWC2QaLV
E2+HnQ6MO8KPer9oAqXCNmf4X97JEbss95SLGdKXqAZCdX7uavD4ZJL7z4pYyVrE
RD3QrIyBifGBxmgtkb7RNA08bnshfErwi/7XaHAsIc3in1PzlBN9sLM0/hGf7vxX
z48bJxNlFEi8XANpWdkt3iKY1Vq7nuWCluSdCZgCft8mG9IX+OSSmlWBz3BJrPus
Ng9bRLoBGK2d6ZwwbNws36dQOBIbC4YL8tCiYj3GrFd7ULRa39YIEkkxDJWmGe5h
5CUDp0bdnU21JodBeUz2C4ktG+QNsKmV1SlrQaZFftS+g7W0X76f9aNCrHPO07Cq
mRxWcS7+4tbVp6tffN5jIkHC8tSdWjqniwTlyUq5DxK600Gs8KbXGtOvfIT7RBtj
ZXIzxoVTwue9lOr3xTOxZ1hmbK6WEU2h+0o0p5EhVJhvryzgANPXLcGlwz662Cjp
w0yad/OPSYemj0U3V/dN1Wnl6+xoPoxxBdUuROJZaYZwQHCKGst2IhEH9VNRTj0L
ObYJFK0BE+18G/NY3RR+AlopdOoNlK1kr7uERumvfIzEXZvR12DB5swWrUAE7eRw
0+aCu1Ks5e5T6Hha+3VtuCAEDauVbu9WO/kyvaq0xS+WLZn14IBLEZbI4PW0s60f
Mr6iOKAiECEdUU53lDMpPpm93cchMPmBLjhjNJ5lkPbFJYPhy1VsxzU3hVs5evp5
0rVFBdVNVPLR4qdF458U4LycKyTuxT/FU88IOeQP4KJ9RMgr9sPl9UInWQJRyGAq
nW9cXAS0exmPWhHVWk5UezuWrZeev9dL5CLvmCWuLFaXZPSbU0ptvJQFKShKi/eO
HKbfI8TrVSABkRxplFvz9mHaTplPvsI8ML+Lixr5OboMeTKu/Gx9k4qLDakY8IqT
FvIm9e//QPbzb/ShQAPFb8oLvIP4Su9B66zscFK5x3/UA6cZizsyhwKYCwQAkPxw
u0PCoyzElX0McvcJzS5gbPphndrrvpvCr8AvEWLMoGXD7+AbILmsU06Jjv4Wq3AY
rn9Rzmihb2Er02uZUzfSqDiVsvRtcs8HvrFJDpBJQBRukNEECUDZ6KQxAHzPZQwm
WpYcyJxqgmjA3Qv9+9YiNJidJ5i9U8vXcJiH8cDBH7WLEoaDKQKOVd+GPvnQXrVe
3Oq9voFID8labOqKAvWXHEmYyopat0KJT1FFLlmi4HAAcSGR5+v+w//SCzAOcoD+
IoSUbooGEszbt9shc1oa74ao++5K+L/VTVQ7e4tKkZGAjhaesAbpVIyII7ndCiUp
QIxhYl2k/hgArSdZp75lSs21e9xneUXw071cV6FnVI1T0qjNIuzlrJjjRmVYvn3z
QbuAkwhskRnb4XwfuDrjMxpA8EHNH6S8+1NU+pMk096pwnb8DQ8Rf9Y4lQASLgIn
JvUdyIX+qZczV4eCbyFlG9jRrzK8uKyHuhU54BSPHRXPqrALRfMZ9zlzEqbrEUQy
y1JSoHhuDHW6WCEfNQU24unWUYeg7TgfHO3K3/W1BI3AlFDeQ7d4pw26JpPbpk+p
ufutBsl5hmOrkjCW7hgN4oZfjTET8EGH7ID7mxWVCRdRF4WbIOreIJbUnNq9stB8
PFvJvJOZp5+EpJV38A9KXolVFVPZKcqtM93vLWIGh9icB0CVr5lq+6Si9JKNJ8aN
VzG4ZEmiogDVbHw1oaatGBysj0+Wh3m4dZtSB986ItdhlQA+MtPtAIv2c+n66G+8
hVEsotOH46o2cRJHvqnIxDDdhAlC+a4S3BZ0fBAo0kBJJl7dzlupei7RoZ+PFChf
QE4h8DjOw07PYTE/ogxveJ8vxNr8Kny/YE9fo7zZaZ543xlYsYh1lLEa773xNYb4
hhzbBtVKap0krA0cNsvO9vH/i0obUEGIHuIGxn7RJ3NRN9Ya49a5II3ijamZUWd7
bL5lEg/SHv72huMjbVNXjxec8a6KWG23QWGaXcxgEesUqNQYhLnDDWuzmrVV7Ufo
knHd0u3k4nkPsQJsoipv8bXXZNL+cVKglFm1AS7tfpnzdrHBgqj3Pi2N1G8zuI56
XpnkkyAWCl0RwxB5BB33zZWwXktBeUvwiJySkBqGIbwiMSLFHgS9d8at3GD5YGvB
8JHcobovI7Dc4zdUm6cG3BOLTcB/K+HtVZjPND3sQwbdt17gcQeiMXzEvYRp3Sdj
xk8chkJADuOLrFwxShoYtUzgYBTt2Dh++OYx3OmPrv8Zm2z5aEpegTAeqfoQC5FC
i5CFCliaV998qg6u7sljEIJ2JCZo+X9qcQb4/FdBByniOS/ecbusndhQAL/y/znr
yFkyC6LY615dIparUkLha+cZuEBS4wr8z9A2s5rpLQVE5xOFRfcVSyeuwy8clYU4
JQQI0uqpRzfgZksC3N7/I/XqGoR81yfARnngbnKtbGwUOJxFQy0rs2ZxQZuPSsuE
W37qIw+g3GKqZgJWcguhEIsbvlTVI5GS0LfSK+p99s6h76Ui583B1HqhQ/9z9u6+
ieyXczepncmLkdVM0GBQR/te6iByiR980J2hNVayLtjrRA7VjIasp/VkMPl8qjG0
vPEo3hvUveE56x2DXl0zq1N1le+4Bl8rQirCB+WRN6nsslVRRqX3rxF0fzre+t+D
mnbUL8vq2VGc/tYlI23Bm8x1dYarKOwcetHc9R8hdYNiFPmwJDBxaoIoymF10Asc
kw5UMceqK39neqgBhzi27veBzS23fTd0UQqcsFxjmzRLqBxksiiZTJ0I350t8YQ0
apnrSTpb2yk2XbGUsVnxk5ifY4sIs9nfnqul3z75pbblgDzRSFmK7KvjtVnADnrI
BjXT9CWBNr1dPCpNMSjUmhvzi7d7AHEzqIApR8sz48n+EXeBqVhvM0Yw7lPNGLcD
ziMlhhOMPEsy1IeSaQ6T8r967eOxWDR2+kocupDKCXF1Z2FZNLG5+jIy3m5oGyZl
za1CwQR6ylpJ6MXgcQz+5X8R8V67+yk+12fD5RAwsvX30/rnlu5UqV4kAhD00nW0
RpZjK3RWWo4wpM0yVBTUDOZad8QC4ZHnOgS5uG7juBDzmkHA81PlTKVY03RDkU9N
W5VbhOCY/5IrU+VZQsoAKhgx2x1dq/To29MY1O4j6YHqCzK2zze6FRQz+dAN3+lq
sxN4KjCMmaBt5b/0una3C/xzdOFdFDdZeEkk61vEs76WxTxL4iKMqtWZGqkvPVhJ
KXalqDltOTKIhFDWFhoEBxaeFCjaalGofmAr4Nb7+jASwexQmSbNUtMkzz7hlPoc
LYbxgwx5tgTXw7XBP+mBiKkEjoQi2J2p8YnVr8qkF2D+t0wbmAe0Gc+74WtNG2P/
eFqCTR4vd6VnLDnbmgQiW2Aqs8eoIpeZAy4JLIM9Ym3sKcFAuiLxBFE7uVtSK5yU
uEbXxWe5tSH9DPOGyEZMgzonosc+rh6orzcr7O1rrfPS8FjMp08yrdoqHB+Fgq7c
FdImWZvUVSTl9/zadcWCcuDBR/FVMDzMCX/v271GABVdQMGcxnwmzqazN/7n8+cD
oYf9E3WQH5QhEWbAgV2rd4icz6nLvgBau9iLf/PH8Mlk38LS5qG4zZSIt5qj2Mf/
gj0buLZqoEGF7ui0t450dMHbuLLRBBklgxnUehNBjbTfrOws1+2VgK42LA2yrha8
FptMn0gbEWnHCCAUXMOwSafMP4CQ7NGA2wYAhul+x1nexcFx/kdK8gpxy7b5l5x2
HS3Wq3cFy8EBJuNOxmWpvexfT5SNHEZvB531dzqlnrRhB8lqcXy/ziQixAjuN+LL
aLjKjf1NZ3KJh8bw0M/K2knU4cE98jtAwDw/JGwjOg9MsUMrQeJum09YI44sYNzS
RSX9P92vNJJpTp8RSQX0Ac1P+aIpMK1I8nNMOuOZ3J8y2Vwy/kqDzL4OO1y2kpb/
QAAJ4j+F50Xv/KtTaBSC15n/qbmRAPOtTUTFoFzi/pvfleu74oGkbbuxuPECKCEr
g3s41liEneApntZapX5imrkVltURpFzuLaEFSzcQmVbfLv5usRj+ys/6AENVqsM+
Xyqege2Z3TS2/I0/qEFdo6sJwxAGlAkckpZRBIGQ5nRZFhu7STCc6jD6dRHPMrqn
gicUQn1cZNoh88xxy7W4hFFPksSbz6Iew8pnn5pUVVl4TuGA03pE9dgKLb9IpGmb
WCNLod8aiqjrWE5tfIfFkJxhOwJT4jpzLPvf+ZFTK3XufxipRimtnrTaz7quH/dY
f3dvsbhnWkXRY//7Zksf2+wcP2tg5WldlGMGfKFcMoT7bBlJgXnn6NcinWkq4jnK
Zhi0P1BoVx3PNqHB0BwVcUHlpf6ydy71nkYaAeZF8K6IFRDzhZLCoTVfWCzl88vM
BW7lU6yeMx2lhKiwIlYl47pl3KWqc3BYGRP7pbEAyAIp6t3grfQH3XUCXZJt9C9q
oVIFm4kUUMXsswtQ8E7pdighHa4jWs2b15fPLVT2odPe1bL/Y6n4+4QtIRdoA98o
A/+72VWP4jHoL6AXzCyIGxmxvfRA64aJgLg4UklqwFx1F2OkILGbedMwo1vZGFYw
NTMMwGl8EV5AQZkHa9n5eAF8S90os+IMt2qRtK+JkcvAxHBa9WRJ5VtNjoBetebd
cNPDCggzcv6mslc64CBsD3BFWlv+s1RizGymt6S31hbpaCEhUomjIjYAQtDr+4zi
2UE9L8LcjjCgAQFoYO54egLSspI75Xnc1mI10TBotuzHlHAs8Ccllx1LBIc2/jIf
O21woYqS9WUxhmDz9MQOQni7UQFLylcevAuHN62BBi7aj2gP192REODdXVQ8AuYV
EPB3odyvqwnG0UUwIKNUy1z63BW9e6Ja75Xvjq6kCO2X1lhsdFfwhZV7u4Ms2yBB
SAQjLT0HB5b3QcbJjZ3Z8SLDZVObzT81Wa/b1u36ajrqOYkCmXG6S9KjFP7K/FrO
rDnilsptgPvBcY7anZwK5dyOIANOsYaYj5Q9Ep59Urg5eZEnolWn1/Aqbsl/Jlg6
T1yQjWX1BESEm0Xyn+JszpgASSMK19bNE07aYzprE3SS8AbK0QfjEDW6BGPytWt4
+TrLLwIGYy5nZ/UI0m4nj1WIv3shVW8tnoSMcEeEd25J4QuK1zeiUQk/6IDU0UcB
czpvDbTAth2t0HfKf5mJvbwQ5nl7DB6wUa68YmRHyBVRUuReLaDOmp6Qzf/nYCFz
44owUV1nP5Y+4weteqUjn4j1SaMOhXzxi7xhUIVQKK1Ef7rGT+tUT4BnT6DsW9ig
DKeXGn2aoXwcF04ybYV98QSl9BEhUU+Rkxq8RN3ONXhgpiru3BDCh1V6Nvd+hMZC
JKs8m6v9oZ9U3EgdT7woN1Y/flUe9Nh9z5a2L5yUkTgREX0FQRDUDeUYAm5stVlP
b3aosPbLUlFRAT0wEM47AVC8F/uJgWKxegMuVcoy/yZgbLFt9Wh+bSRxVx83LnWL
nOm+cjNLLrCxTcpeHRGd7cpnwMGG3EpN5+W7m8cVEjzNMS4+v8+Dp9gmPGUhdcCM
PayLQilEQWFMIm/vNYyBu1USFvMO2n0gDGVwurTalKIoo9EyfwEBsx6Q6BGzddDs
DoNyT+TvNRRaHVPdAS6L+L2qVsDPQQQwOVinZyniHFkVKsIOcB+XuLYGKqT/Ysnd
0tynxFC9hqjkXthDXrT3Vy807qXYNue8Sn8CkJSrLBmoU5oTkGLw0wg9lQ2BOm7Z
SQytX4igVtzR3MJvwiLY0kT65/RrQf66020bQBBg+d6KgBf7gPAwa8ufGz4rZp0E
MB4XhIEGvUxTw0O3O0qLZowv4pz2eC4wGRdSV5/qMux3Y/kQRByZJqbmpfXYf1D5
b2sBYneh+TiPbwfAgCr/lcgO0fdY+yOC9aQKUD7QVm9Kms+E0Vh0NSFf09PZd49+
hIFIWJj3W3oTCLnkAr2kinXXin+rPrCM2MBcS7a2wDy4HzHamjW/IYygBaJaRm3B
MbvX/SxgsDofijNb+c6Pd49QwulJude9dGz1mIRAZP6N0VQRi9RjlGhD17BaapiE
Lu4qeO92mCERETfgmP6u5AZ7cmIV30Yp1QXQKU6FFypBq/E/Mnm5NY0V8xoPtBGi
k2p/IMDn09C1FUkZZ1TJKQerTavVW3jSvY8hQtHjFxvPfYnxfUdY/q3aHws6OJF2
roIk98Le6h4dzG7C2G0Vlv3uMuusJ09+qIiSlCp4xP24SNxQJNOFelGifG3uuB8c
AOdSs3FKgFmDwH4RbefAwh3KBLoxinXNiwSxN02fjH+adkhmTH0ttCh3dcWwaA32
nD3OF+1unh8pns6rStVpRls9qemsI1O8TUbhtvzAZ9necDb+u0LagTnpejDDM7Xr
JwwgKGkYayPp0GbqBtt1/6UyNL6ONfrVkfYmbJFH+SZ2zqbszvSKXUFbA+Sq0YAr
1Ez67nn3VbP/Uh2ftg9x07YK6OJqkVQaMt8FvKyZqT203VVEdUdH5JKurfahdlmm
r+fQbZMnGRDMtQvuWfx9+XDu9/VPBdjmGbzf3/BzgJtlnNRWwO6dZdcNeaBjV8XI
JOouYZeQHEpv6xuTnbwQ9InVM2r5gh8+jhv0IkNwk1oDXcQCEMGoyl/1BogWJ9Np
wjlLcZVOz+vxiHev0NbxtW0cm5HSvE+auw7C2j5XLg4ESWxKKcvT+CYARatwKRSD
Prw9a7JNjW0k7p84o/RN/HoZfqH1x52RO9BIQrW0cAcrDYoHQv17dUXTwp230xX0
Ehhc6PzxwfGOdPPLTGL62CHEqQQZa0KCokauYqGDviL1KsvH16RCxeZILcPBpNwk
4ZAAU5O6g4VCd5lKfyfhlPRZ7M5RuLyZzHS+ewoaqmJuw29xLl5umHLcav9nJ1KC
jNQasHLrzFBI9F01zCSnaouXBFKFCiJGbQbE0KayH4N1ee6t8GIifdYFAqmCZUs8
n4CNF7ifml8y1K1xrzzaT0h5Vm8jozW/u+8zoEyBn4h7+a6qYtgMKeNe2K454VOq
ymYa/N3fR3h6Sji4QonbjL+TmI1xv9FTtX+Y1Zw6z51t5r2ZOdrQb67m2n2X7FYK
0nXYrbYEhDrdJKzGnhKZ9AqL/RpFMz2A039cYZsKTHkm0Hd5PN67GUPY40rcaOrv
fAvmgBEzLlhsp00mAjb6UObNiM9YZyilleYm4tIvF+2T1FsZhawAkPIp/AzLfHOn
B3sS1IUuuJRWDW98t4c1OF8SYyxtnK9S2GfCbY0Q1kkPPZfXKHga/SKkAQnbj59j
iSPVxhZVpnnUFqaCfpIpKkr8ZY+B524yO8G9R7a6AUC200lfUNiGhVouJQ/NKqjr
HHlZlKG+IJf04aCcpPLBl/V73BboLRucPZbXTcTYx/3JLQdzQKiLpZaq9zP/f1LE
udpamTVv1PSdA3P8048EIfh7YgoogocrG4WtQZHf8KtaLq/MBMCYCB2NRhoDl/fe
wKZ6ppXRWCzAb8zfoyWzgy8gUX4At7/pMP+Ee5WkLblcS+lfyamqla/6WQHIGKb8
/lFOdyeyJuurymOy4iov+wPs40InCjUqYp00MVfFCERaKJrRljf7HumXHEdXT7xh
t0mogW9iFI8GM0jgmCvi/qEYcS3LeUsdX8UzzAPsmCKyiCaufBzt2vfBOJPWEieQ
K1GbHM7+4bYkw9kLQtcj3FqVV4HjCocovmBXFgTGSdr/nZOm9YFqkc8FwsgwrKbQ
RkXqnBFPuHmcQTtyWXRhLDjtiPhiGvBT1m2XjRVVwVsV7C7THwggUpQoIgpmttsF
vRfjX5WgPgGp9L7ZzvnxorN+0njkdsVGpg7PQscRsxrSJ3eSktoAPxovQiZaTx5K
3tr9dSkno0A3Pt7EXL++/HdGEHZCvvub+WBZl5J2Fb1WHoPpBXLwwdvKEGAldVS4
4RhNbwXho6uXpwpfSw2yG1QYqHvcgBFNqF54oCyKEFDqYrOXtoCEHuA/Qsie1MY5
6Q6fUbneCu8SzBfiYP4/twxtOZb81bCwCP7RfMRHIxVGrxP/mVw5/vDs3xSjeM9L
48repEb80vAnAIroNRl3Kp49ap3TRVlA4OhpWzvcgbp+7A2BagjrRYvKuurF+qRy
ZbvJ//v+a4jiy05SlD9X47Vu1s4PX6INIBshThJojnX+q4e8IrE3V5+1wl9pGrnT
fOAZermj3/GEaqcf+fa1ZfpGIGWiUkgPweYhAOsjXIkn2Va636ABchFJjp8PcshW
rj06dimND1Q1CfFdTDOdDRuE7b1ppzNRNbd75DTYwOcFLED/CGuvNOH4LzGX3FYa
EMRRO4AoqM93VlRPTo2b6WeCsacundRNTK+1AX5It/xR0LaC+mNInIdpZP8pDDoF
i63nuSfcdnTKC2SeyZJgOZUSQguJRCCrzvuy/shnaYLDMFl+Mjn8DDaR3I3jznEm
kXyHA8B812mBiSuAVdmIlgf0iw4HaZ+/hdFPo+6Rt+vbgLPPiAzDzQtU1r9YDp3z
eh4/vHGAlEvniHNqJ19hevpAJXxJIRTVfPB1hzmcOGOL0szcRhfU9QbvMgJ7sj8A
F1ze/62fHThJqoNxxqjRyCyEKnE3hQ5oATF2S/EdTBps4N9ZNtekZOOPyYI+3At/
zAoUfalKdw5pC1na1vFmffUfpZmMrKoQPSMuveWd0+2OP1XkIFkGdtYsIHpdIsHV
TUL5u1ynNIUIgVxtZjqCkMC+2a69MssmFq6vZwr7q/VmtreX5aj/9cJw2COliEND
EytmSvh/eVwaxkBZWzotDGj+WBkUB+s9rM0QBmkSA/yDYhaKRm+CXfyS0FX1GULJ
2R8GfJ7T8YFjZBiBdgYun8ZMsLl2Ge4c/n05+I9kc51dm0yj+XIsP6Nlg832PuHa
US4x7s0sItW2bJscZDirH4oF2q+goM2Y52qY6ON824hGxkCJdgFhYQXH8cHt7sfP
h6TZZO7VHCgjKf3DarRC+ufAocR9Gi0uHTfr447ZUUeQIrjxlPDGYMrvh4unA1vI
q1yk82gSMOmIR+BZFFolF/guSd9vpRPdmzAkZatqcI7ys3R2HuRmB4ScqHAlnT0n
ztRJdcPDmU4wX+ryyQEsvZO+fuwG4uDgtHgi71Dm0PJddOQgDdT8BkUKu/IUR97B
EavjG9cCoCcsy65R7vVg12uvgSCSFk40nME0SGvZtlPlxy2ikvHiti7Jy6N3KUk2
GzDIP1JLqbsZKDDEIIBIGTKync/zVFjXJwaZCFDWfRNA+eq3O4XHoU5Dou9BkRJl
JAepAjaG3OGbzF8SBJQ5j4wZ3FwDCXG9ZcWb7k31inr8U+EEGH8+Aqsv7oCKMS3G
ttOzKwFJpOrh+UW1AmV61KO/L1i2SREhTXe+pWp/fLyvM2BdPnojJgMKPPktY4ef
OcXJw6+f8MKTun+GS1tZa+2DqNmlDDIC/bvHkTLgXgyOdaCmT8ANzNl9CuBIvGxl
aL45J4eiQqt31zVhHPb/ltg0VX4dD3O7wTioDg8Qkix/JeZTcz6YCITp8a6wAe+5
YGOHBalUufiAp8F6HFoPE9UjdaE7bWGZe39tIFB6Uf1mykFDi4c6DT9UOv8vKWme
g384k9vQFU7s6lmYRgu4P/zLO/K4Bx8OBAIYbyofjUpXr+L3rjcb7OAM1dQ+yQ8M
ScB+MESoYKpUe5XU7Q310gVXlmZr8axkcOkRAaYrcP4cG9IHNmtEiDHu0ZJ6FiPj
hWOc2O8WAfJnFpeOKJg5GNYGT2PpH1gf8crqIM/fb2pcAa4iViAi4biUnNtogpQc
Shu4FIOuLPoeYYofUWoEhHsJiw+jGZZuwkpLoX0T/RkCJk7UnG1MFUHT+2YLVDtq
RwSnYU323Gf4FfhqRTihJtH8fs41O63DHseFIJk31/mCV91IdY7UQSLRlU4BQfth
LerA4wTvMAoVLlCuq2doU8Y/m+drZvHCnPiH+raqZs4pryrTLWLXbxYid5BBYtUC
/6VQY4UT/RgD3NmZDDZLVYwKiiY7ZOIPxTUB5Q+nKmjBQw0CrqP58bjLnBhYaW1w
7KOOp7alCnE6WrnvLdlCvvvi+beem+PO1DzVTSF8gnvXqC5BYGi//V1JmJoVI0T/
PJ+rbA2gL+zQF7EQn3vYeW/kn1Kqn60iEMMohEgczlQlvVqJD241Ang/NevVWuk1
nBb3aZGWQ91jKKUrb/Hp5c22zWbHq5iLMQWOloB0X6sJFHUne9h8v/HA9HvY/kEd
y6d42RoMmZeac16F6Zvu/Wqj0LHYS+5SHgAXdYhSdHJa8TcDljVWWuLwvWHuCgyq
BWQfOs5dDMvW0zrpT8nX2JxqViI262otsK+hqTibzfEvn28iAW38MPW8gS5QjSh/
lWcaEF7b1uxPiRf/oe2Weab3xGDDPn6Kv19WpI4SWvueVbQ6moryBWvOXG5kSTO9
tibvz8y5ByIBrHOar/zat0Xt9l6agTYIgDOimwyNQVqKXgXnN+zL6raVzCva5t2u
NfLTseCSjBvkyFtBLP2FAPGmCvjPFcdpjGDZ0iWu3bqDfIyqEcgGpmP3zCBOTefC
Sz5i8XBmaQaa5ymPzLPnlNihoFPf7wYwTMaCBAJeumLqNqmBGcO7GPsWMDSJBEhJ
aOppr0LefDAlO+TYFO+4YxiBdsdNjjtTnsHp7DAHH5EO1IVc9qJElLipPdfg8kk/
AZABpdG9vzpsSA9uuV6heQ/VAgapOnPz3VRvaMEDKcPfB2bEwbZ3cIRG8YvmnEP/
qbWs886ywoHIKj6HrUXntR7M5chLpV44Z3opUiFhpwrmeHlFeXz5JRBzWxNkwotj
Rj4ybIDj26+SGrvjz4d0C3tj2fi0pGY7VS4KfPJJOnp7irgzBQeV1IsqH5Fk7Kjt
o5M7d7PgjeSA2Mmya1J/br+ww1HqbCHt9AbQN+15D8L1qb5xJKbPEScWqUfAcccr
3m/dXxzR02EkaBETtb2AOK3hDR2ZXFHC+pMPAH1JYAxmb72MTUdrQQ+j8s1Q8CZK
r4VUOl1oIgCVw7IDTegtEREdDrgsC3I2YOq3RFKcgUJakn/uu5hiFE75fqFwcB2d
9nA8IwuIkxu5OUFoPr9wz3QbOzYiynduh8PGzpyj/OMq/gATA2WWvjj5TRKhtBI8
4AnG6Ds+MBBOGyjwZsShLtpt1eqCD9li7cJ32mNTfwG3KGx8qG5dstlMZRZvWxaE
JxOcm9bC4FwRbH1+q9CWK55DANquPUyMTayIWs1qC/RQuE8LSaSfMGexN5XoNJSd
6sFDN6IQGBYprjyw6JQ3ktOJS40E5Aj3C6mhlZusT8ThxCFl7k3fVWKWxvlsqSH/
FVuFzRBmQEF+ECixpl73ZXws8ZpSy89RlRCHT3gRJ+NT8UoKpeCgLPSHNdsdg4jd
TW2Hf16NV59DAu+8SFFOoeG6YGg3FAdekeePPCC0+1IyfNnbyRD03GEAOgYBI57o
BvI6Z1FvqHGRnT3fEIcws4/EYeRLpjnTWUbK8Bu6IE4vdXHNVyzStont4iYXpLBM
6QIn8TwKeoOfqToC/aHmCcLOlHNpWBoM7F/OAY3Prw6NrKEzxD9LFAzQk1h6x7S9
pFpYGaEq7cCHXJJpbLM97k1NhS254K/k+UAzwcsoBomyr2EIbaAzscQitJGEO9sP
BxplZgv+UnFcy8h639UNY+uA0VyU08EiuuAdw8EfGRzi/JboxIEq0r9CMdwgXKwk
aPZx8uUqfwAxcu0e3W0mxorqXal5bneRBJI1ZZ47jj6d3nez59i8xzHxCj6VTbHY
g3S5zPsdASYTZ25H4oHNBHxOp+RsaRFWC84NaZ+QUgMLY/Rc2AjImLxAm5oVGcrV
mUPwzjZhhVFj1c9rLCGbt6pZoXuR8HNiNnGly9FsSWBY+CK3QKvMAUbooun5axw9
aICHmyUjReGjSX2f6nKqGrzh6ruLfNE3W3QAQokaJMDEfXwQ8y0SlBFafm3HdzWn
ZQv+EWUYSTv+ypnhtVFf6hcznkEAOJYoBBQJfFeT77BS//8rRRaDC75rgy/MC+bz
ICaKOixCjKagJYN4uUoXNs/qsZbB//oFgE4Ix2YcR+MjqoT1g7znkJzCQyb7Ofbg
1Ib/8SEbHbb0MSCQhdo4l3sku9WEY+JQ25kFNahPK5PXj8AiEGhyA1jWIng1y9o1
mFv1F3OnxIxW9xnt4GiyL7J8EOCaRGKlcnJhZoWP4mgFAX92+8snxihlIzZ6EY2J
X1bD9UOv4bzEOJwNVXVzDF73x6QAPXANZNxpP7Dl38q8NzXILhEapW0BgfRhInUW
z/vUt6f+VfkeHnFqsUcM+Wz6AuYJEbQ8bO0CBCZqyAiOg6Js8mdVIG51PAmI9TXO
XUAP71gG13z1KrhVKjbj99AroBxBS6sT/8Mmy1WUflQ4qa5GKg6oGgBegJItThtm
nj0EFv8dKUNoxM0dkaXYof7qyWPf6BF60lBqfdmXUJ20Sx/42BFtv/P6g7bszyg5
WMGAXEfNxpfKReXXuIAIt39eTjgPqdWzoLp7lg8VmE+Cz2PoTwtxo/XNLhfeQc4p
cYOFiP/HBRes2ois+zkONFcUtEU5eB+wCf/YUR0eDVvP27P9zCdkTLeESXsT7zX5
52IRbkgkNgM07ie1E6FmlLj4T84oHOdD36CHiymoMegO93KRru+KjFBQPPhAlEEb
WjnUjPrKAvZ8W6nYqDwGkmT8GMFviZ3W/E/ULbqKvq8Os2Oi4R1IDCKBk4HTrQb2
jBEXEfv9udBItcFdVKmEeZFZbgaSr8k0bStzLdD4StfCZX5fOHTUWOAgngXJMq67
+Il54H4b7dcpr1y01Eb2WFI1IDjPFthle4ViW5IQcGHaLp9vXeqLH4MZ6rOLLBf4
5VMdP7gp8XtV4u85Ms8hdMdzU5tD29Gm/VtpQr5pSPXTOU5qwjBjKenhvq51NEm4
+4OhVEksfncOnIHqN7MY1sl1dlbcfRlA6Ea1ENSsofcfcsZZukgKLlguzl+wNwIN
XZXbNHq9krEDCjy7jyLBntX/RlyBFz6bdyze5TwQ6OeLpGoU28gLrnaFogg6BHe1
4aQ7/65rbIQK8EvPEDz4sRw5gonynAZNev/2/QMDzjTut/Rsr10llHSjwddsAT3H
fQPG0U7KxMxZd2FguwDA6jxIZdvymvpM451SQQ80oqQX2KrqXhCBqbu5NHR8+EHB
GAlvPmJHXCjT+BsytjPl14807rrxPvIiFOy38/mIjT5wfpmeujikpf4T2NLc+Had
lVMm1HwnNQBpVGwp6g6w83luXScs3kp1LsyWCQcczyL8yi9cwQEXzZDeoq2NFzap
6EqT25LQkImyoByDVEDHTZ4U7PtmFmVKDDx5eARjPQIYXvtz5skett85DFNFK07J
IiIEOpsUgz3a5Q1VADr8oShhFG6r8xf/nmtukUEVdujN6Zd8/IW2d71pbuzIUviZ
CaOOhQRLmbhG3uh2Krx42xcszu9+oZPkd1pOvaop9euhYextTl/40Eloc8YVrkMh
/TJ1F+EHWqijJ0KkDuJP3Lk4b5Cpxcn8G+ParirI4113bg/cHHpQMspKDEX9QB28
kemBcO2g1Zq6qc1nMQVKjhuF6tAOGjibTTDD9W6U4OLA0MYrF+9jLuOz2Eog0PMg
LJfHk9lGjBLwuue4qT0t3WxWnoWts00h6cq4VHt5hUOOW8hBVl6zaW03TDxJgSJw
iqLlw1yiUlFYhR6N4FxIdch0siHbysI+MGZRmxzL4uev2dWi7pUJxWyslrjNMISY
TlsYtsynK2HVZm50jOp5zaaYJj+PKfpk3Gqos0rQLRYfctkRAFKVdhwNve3yjXBa
LbX7qdpOLiNLuQfthYBUffwBYeork0PtAXtReX2+CzWjUTpRFCxJQMP8fbrjsNUL
eI52BMfMGcajymyZT+4eTQbUJ/VO/EkmVcnmddqD8AEKfpj2PxU69HdPqHXnpvGP
jfEl8IPkRQJwUEaw0mmEL2cq7G4PXAk0fRb/Pb8THXHOWUqxJcE+9fROw+UvTPor
fQjRsIxWVXABHV2HZfjByXQvlbMSoo00lBc3zMgdSWdHQ4ONdi2fTacsFYF1AOq/
Kl5BhRhK2AHJZC/5FBGYn0JfeE6Kqz7r49VA96/y7TQ104kcyI1eA7VPcjBktm2Y
YAlvkSv4yMVsXof/l5mhwSc5I3HiD1NGYERyTbDR0eWZBK4YfHTnCmQUv2jZpbSq
1vWhDGkFR7ZOtKozlZm1vCsB83oiVaZq9VtOxS5WepPKpGcHkmwk2Y5I895vPmCm
UvVHDXY6lsbgx3ak/vMr7dvPNBmufv3RABsbF6iWERL0CuGur1o5QkomG95YaCSz
Y58+QD+CmTY71Rrr2v/sfHZ4j+nVVXd/Occ3aC2U+ARczn9LCrmvI2eJpgkcASPt
wQxHsDucgrcejI4H76eCZSk8KkT4CqkqKA++AA3ogXdJfdtMXb549UrjPiYKA/zL
4E5tvnD1rE2WE1RfxcX0GSDJ+nsglY3/0LwI1UOtSl+07CLbBcIAmuGzHRft9Ukq
3Pn7tFgDr1CgWBS48vkkBJReqC2k5R48plH+mhi5CrT2DYBH+o78ASdf1Oal3bpa
KTLxCB2erVgRDPfHPGlEVNG8hCbW9uiATpG4G4PLFLziSyGAJpxr8WpufFSOuunK
KFwsQ2xVUNGXSmow2oxQOMnFjnyKevLz+pfE1EKU+cdpLl/tY/8JbtJPwdTItVbn
wX9HqUx25MegiSWdAlzHmAx6mEQcEGrQIGCN6pghbrezDbKUBxTc8fIffnshHm0V
QP8icxTXYM1iuT24oT0MeEGtxdipDFv2odipOFXr0arNwc4IUzSIiSu0u0MCPhAi
D9a9nR8GmhTPBKE67UBedCPETtx3HTFm6VTgzpj3xMGzThTvcQiPFTvAh5K8J5s5
FjIJ9GB6Jv7tEkj4FRzybrIFgOAEhIU5yfEnisXs/jwZyTft54215Jd8/qTr7iQq
DHScPvxKNAk5QB/CAlkJGkWEEMcrnl733jPtqcry9W3kwtWFz687oyzX9Yr4fTcg
VYrTLZPiEmThzgaw4LQ7wDqP+3yYaDjOTFl/jXUqRFu733Fk/RvUTX01EVl9yZc6
QQUoVhrSqeEeRTFbTpiBJpDNary7Z2LQQO96mVmFqJRkGM/kv10zdrAEVzR2stSo
Ynz8xYFtlOWA9vwc1dAMBi747QFg5xWr+e3VZ07iUE62tnAv2qMItFcY2xRtvmbV
nzHqu9N2/R0XV+TIKzUezPTzArKhHWc8qWNhU6lXH1hHculcR5qTrTdCiqX1+/pq
7jqa1Ilj1SU7cgmkFO1DsaWPnx10OCiIvoRiJAMyaqKoGmkIeMVhTB63djGdOWRq
gWvaK9D7Opp+hpPU0rHxAzmm3pDeL3CS5DWPLu6/f6rRl50d/Us8gQFtfE7QXuE4
x/UrmP647h/3sJkFYHUlTlHWVcsY5HqJbEoHD5SOj05aa35ii71QN9+JcyvSBPzg
ygvvppHPA/sd2M/pN/+HLGsMfgAhPXMF3G1nk7V5EQ6Yxrf7NPaWV/GzDcHkt6pi
d81aiILcKfpH9XUG+SqMxs2iRkHcjf91NWqgveAxEOd7tN5gPWjUJYqYXLULVWVb
HRzUJQ3mdl+jFnX5SzPYF/TKcS/+pefuAmjMKClUHGgiv9ZuLH6t4yOU1zY9lNAA
Al0pLU9ISQ/JFxyf+m1DW5YjzDZU+zM5Sn0HcatPc89BqCY+t+mHvX/5CBHVm4KD
U/rPWblyp+Ytdoysc2r+2tbgEhLpI4i3NQRVReuvMThGWA+IE2F6BXqSMOvxh00/
e0oML6OnbfEZxXtoN1QLeGVkwqQLglltACwMpb1Pf1D0c0C5NHKYNFLgnvcQqZ/+
uD/dU/bTgs2ynUnocCsD3cZqvxzqD4mqcamOdGJyLlJLYv3cT1nouP6+F7aKIs9A
7WqRhSe6MyJqKmnVhTbKCJTcuv5F42VnVRUk8pYzei+Sw5LNiO8FiD5cTIQZ7RSB
RFMjrTHI7UxS5yJdvqv8VbUJV0xWkKxtjJE8NX0zGeSIautQ9NVUTuJKh1g+5vwK
gNPBYsh2q4TwyIpIm5Eg8lWUaqgO540s/OlsNYC+7fY6jNWe4XG0z1pulZTFVjKf
LWitoUmHxpGHSmrYlkTOQeczne7qKOgZgQfpaYZPgzQR79cCacuuND1/iKyAyicl
AJLOceLqttnKvp8ZeyrdJJrINtLbn4QNUZgpgWZKF6l5dHAvAXpqpK3W5tsFxAG9
BeQh8SjJbQOu50AfxUaEYWATdF86ATAe0T4S0uhZbJGuWCm8RUc+L6LNdpGs1t0F
JyFymyUsSniZuOIR85Dif7tLu/+OwjAT7xtm0fL0KbFjl3SKE+VTzcsOgy1KzPsQ
HAzZtXR8a4AMlYqOSgQh+vdPq58K55VoUsB1Vw8GBEy+71nnfFK5rZVy+kpzLZBy
o0iCgY3z+mC9GDvzfORVIog0DlFflRqxuI/O3HuLXjJ2pqO8SVc5zeIlvPihiOTF
24L0Bzo6JF8u7xFdSCubg9GM4r0kg/m6jjIcKKLvGnLuFi9G1AMYxPrhmbIvwE7v
kCj573sPu9N92ZqxRtiEw58tzLdqprrtHHQjLmSlhtbrtC0kgc6L8NrT9XGIuyqn
30ZTPojTgRdNDWzmzDlRWuXk+sZIPxEc45Ds7oDLwVU1LU8YObmMgg04Ggh1rt9K
j27ApzlsFSbme+zruEuC1JWxZG97BfKgNnQVCxH/koPEGmK7wegyTAB/3aIeXCWz
NnrSwzRuEKOXzsI+A3gj+QyYldK8p/ESRsYf+h01qXlLjt1kHIMJyZzNsF9zm4d4
L097Brzd/cYD+vnTFucekbdoSlpdQzVqYC4iwf6+3QuPftv8/1utfP+5E8gilvs7
4NepBtokxvuxWmIL8WNJK8EF3ezeMx/alayQbv6YC3L/WuB/ENHUhLGcLPkcHRSk
EUhf4nFqlKLziQLPHO5RUMuKpRqfjqlpOx0+sPYH20O+sEun++yq2jKpklnZ0Cu3
gi3oTuJcONHObIbl4Z+rD4rMkmvopTuFzgMyk0fdqy8I50V0Ch1RzMz59PjT/S39
aGlkkh14SEmiFdrL7Q37epVIVybZBx+mSS+8XEqsTPLDnzPCXHzppH1/ZFB25Wc1
KFcpDpM3uh9wUiOSVwylS3nxZnNvd/tzZn/7Vi6aWasp9Dh0ooGDO+XxwAzhHFM1
GWOg4+5v/xRrU5l64qi9HZONCG/cnUOj6Bn2ZznR4x/GYsLBgOk4x+TTb5/wxs7Z
W3u3HFYKFvAm4zwYtaU1dhllsXkxDX4NoOxMpzwwaxq1lEGNgg1dMW2NWTCNKxji
ak08A+1kwXz9hnkqaXn9mcbPq7VN5KV1PKtaGRAr9EKGTN41ub+dGNxmZEaWw3NB
L1xYrIfRXCpoQkL3iory3pyqbb6b4HIUfBheFNa8jX8Xvu7AGeMaqaF7PpzZMnsM
zYs6uC66QDEvkqxVmiKqalYxJYYUinbidq08cfcIwqWMGhDYacaMuu2FDJtWHuV5
xJCxFZ5qsEOmKVKAMgz3I+8KRxEflsgjl3eYp3LojGzew+lVioexCZmym10yEWGg
uEYYiWtt+HfcsMsmZYtRKDtrk+5Xfh+QXCr/bvGpYQQCsH6YO2WJ+eQLbE4PrG6x
D0isf3eGRkqRRAUPaZJ0nrpaGTnxANqKZ3zTuNOO1tPEzlUfV0hBxHyw/wYGx0+Q
gV+jRCl7NpWCWM9foULNColSi4ma8JD+s1EBQtDKjgA+pWVSPaHf8hbYsRI2onZF
zx55uREspRKRMxBaZJ36vNy5Vklxiu4BHKGlrXm0UHgxJDnNeFldpqtgA1ycUoW7
ToyR4KQ0TFHY1rl/mK0xg8ZVTersfs8IQ9CfcxQ3oms2dFeZzEeR36kKwsh24G5L
wn0ChZVvEbWt8L39UHVRnUQ4bjjogAMJm6M4oSLKaNOksY+tFfSzZA/t8hisum1Z
P64Vs/qTs+2GHIOb+pujHqYXufmHRTBqocBQZmNMw1qsIsaeC/bKKA1fn2jlThC2
BeqCeIdv+xKfT0MrMMkgh1FCyLTrNOTasTcnD8jrkX/mqKvGHxgNdj6Dwn/weJJ6
C+gCn5jogWR7zKtBD8mqFDbpcoYDgclNwyGFTLn9kBt+/3TiYD44tgFF7Y4gu1s0
l1u2Yp9aq5HRYOeWHB0GIuu0PEgkvfoE/S0j1HwfDEb8J+IVZJNI5AWlqebIysmq
MoHV5n+6ExD+H/xwyKlrbdGE7Q0dJZkr0Y2lKhiuudDxqnYi++p6jM57RoMi7Zbq
p0g++4so8GYLV4p0sVhFzbNX5VSOmbiOCL/4mXLdgwssUARnsXFugjFG7sIGHCCz
xnRhkSOLnImy1EXO4Gx32BrY4MOLrlth+gJ1bSkZWs1Zv/i6pHq10a37d9wlPyxA
mpdzAwBeHVSMENDuB/BE5YNj8g1Tv/IPc1k25hn2C9t065ZZiuaZ7AcpG390cBuH
gk57A99dOhDZzrk4b6zkL4kZuRbGep7V3v4uBHTDjWYcj6MtJEYygXGO/yV0w2nB
ZCawIT1zF0qvGXy7RpMdPKDp0nGWF5khIiC6WIdLtxYsvLIKTYPlSZRi0wIq+xkb
+mWlCmKu7nj/uZEwzW610acroDB1YkK9dUYFs+5KzGWeFC2gcPa0si1f/qtdXYi+
+i4+8RSdBJrJpq6xwO9u9SMcNxheWsM8Qiu79bJ7yCkxMKEtwl0gWwaXGo6DPmUc
SR3CH/BZx2BQmpAhoAuYS/wLZ6ox5TzKwo2FDwER+4d5P/hhKTPD0c4fZcAlV9p2
W1dFh1OfLXYghd+7tbsU6IhW7cHgEajyWdY6lfVYygs+D4QHfGbd4DhfYJOF8cIs
nd2SgAv3AJMBE9sILOSKwlSatlJfnwpvbjrM+o0i1j2hpTbxxylwTz9hW9Yib2LZ
uYEGiYRF5sMrMXtWrrd6TxQojMJ/+APb9poQwdNgdi7xmcA9X0PO9OcPV0PZNjU/
yVlfxAYKVV/uuy8l70Yu3Eo+BTNsjtg+gDJ5UpwYWieqAStWxmNONKho2g7YChCd
yULbUqACimvXcCcu4UVlj2HbE/Dpc3kY1QDQQ25Ihv1HcYH3ecBWZRNxiFSo3b5p
kbLftlO75sufj4JVrqFux8H49RC0xRvgJnOEvIRKiBor4Av9rUfzWype5/Syn0j3
ak6nbxxrS1ZDtdQRJGluoQslR686Vz7gEDBuSBIm7twllLZdeQWKmD9LryGOIjtX
glhBiz2Y5+1tf/TpdPOwUU1G633uA8S5TQjWMa04wZKnenXGKY+IeGYrwVg+0jJ4
4ykV2TuIAPPNJW1po84FStxExu8Wf7rR8tvqMXOr+CnsSuZOHwRO7Xb8V+y/aCU5
RfSclZbdFVZGgF4Hugi7Af44mhLiqfN6narQm8Y0Sf+SIZKEvbWdhniK1JJ9Trr3
sou++euTROxd+oFlh3FCIOKGbMcryucZ4bBcN8aU29bicT5xHaXOTADNrc+Z/bEt
OYPjBqypsgFVIxTE2UDexc5dtbvfejdPXFvzwECRX7ZmfIzeIEGwMGMrFLRBe0XG
Z9XRVXs7ujEPf1FIy1oFKKd6IGTAwj+PKLEMUxXRpfvwX1Fdz01uZQfhxppCms/j
44PrGA4ZkogsTAaJJXvaG0qRMVwrJMxhdoMJXiaLaKhOAejMXowKZiUQ2xMUlPgx
KwXLExygmD/rbbkFXVc29kZgDgMgeufCPdYpj/54YPp3jTGyvkfor65Jp6HBv8xL
+R3BvdTJGQXaubqDZFb78ovczWl7SjFc6+rRMwTtX3sc2ycInmp4TdNLNRwZXLiq
TbwMBaRKv7sA1gM++spCF1C2cN5KLc2wTNMrGfCUPjHCIUvq7KmHGH7ecigOL6Fo
HsL/uj2v7ufhP6YKaeDpzWgVugZLYHKErx6IUWXwq3FYZPC5SYmKlMvChEqm2ycD
6mOi239Xetd8uN5l7K4bDtcvbWjuRZE226zxUcCUR9q1io8FNwA7CC9VQbaGuPfY
ZRDZBPwRTpf0sYzRbK7eh+59/VMjoQoE3bTSDjrgLmnq6N+qDlmkRn7Zhojz9n1k
iUs7SSs/du/yKS/7Ab4J8u7OWRuJQybPQMo1dZS/cwh817u5vzPz3sJ3RNq4iUv9
PkmoGQ3dr6/vlyDJ8UwXVJfYNh3yiYYKWsRIgUU7P8ylPB5sCsZLpI0dGLLwgy1B
fiyz0aYwr1z271GfpXRFByuV5SmrFYn5emGlKrB6l4025GO/jncfS598fcHJ3FfB
QOeJl9NzRYdU1KcKj/apF8uf1yDXqKFZqe5suL+bQD3HM1HW27GC3gNirPGXboSk
LHf3Ga1LvhCCNevGL3uMfNdxQL4F3ut1qJnoRPEWcKxw+RBwe1VVR8L/92dJYI9l
99mKGZl05cSe2pcaGU9xBQOwWXDnLBviUb5CboNC6Lj/V2NvfMEa10h+l2HGAoPi
ChrxHnX/3AZO72ora5zGq5rfyfbuJ65W6J8qFQh0qVjlyBzen51pUgTxGZsv05iu
H2DXLFNafIHygOagpvsFPvOutcj4Jn9+9tPL6nur+MS0wL79Mm85xEYe++GMWYhh
4VLI9a2P6YWawPSA9mprKL9pxUvpRY/p3y7DhIu+tmoc2QB+FOzBqj6HzkxhXyVd
zMASU58brJOwPLPAf07yl7zuWWXK4bWRvvGDxLQBPwTo5NkJSqa9IpEqYPRaO6nC
XS9N0MIoJWfQIHdGFeZQ+QYEuOa1zd41SC4PHMAVeLAAXoiJ/708a9L+r8wAm1uU
vteRP25cDrBw0lhFrzksG1rWaeVg/sAoNMzAE1u6hbFSGo9cDbufbHLsEXRHYjk+
27S0SAnYFBeQO13jdIJrUze/ZNTDmFX88K0Y4763C/KFSVhSlUqK+RheDiPKJIZf
fjqvnD8g03+DnCNaD9nY4qGuSGio8vaPlKZkHKHMxmjlqYUYqxw2ogDBA8Rr6zGi
b2fWYfT2aU7ohHpQBKqeVa8oLiTScyCo4YXC4wQIFoX4CQMv/S9Br/q/1pMXNy0j
BJLF6uhP+Og5mJWKJqVWccaWArkHTlKpJyspKGSlGTkh8vXrmjkGqoryak+FQRDq
waNgozAClm7sptEIEcAv4Yo85ldyW1NT4FtgQMh9Gh41Q2sKmEc7/BvWuSSU+K6f
ii0YnBNDjW/NcsW602fTghN6LwYCjtwq01OsQ7DsP7t+56d2ZluPrOB173VO/E5V
QcHFQgK281b5tmuunEGf6nDDUGblSZZ/5aZtTQHE77XacAenctFC/zGDZ84RICAs
irXs2DWF95s2PS9wADL7pBTeov4WEMuKB1ETyTgbtfIEQb5GPPHesBiD/URRWPyW
ncAU26pcl7OGiCDCLtdF6LDDDpJj5/JUHxwau/PTia3BMxKDfDxJYoSRlWwlmC1B
Kdl3+URnJ/4FB+qgNHcDG9yUZ0Xm2ZmlkB9gRGZnUWx8/V8ErVC0Wy2tRIxtfOi+
oVw7ao+ZeWk8g9HnwyIuEYFXNJ7A2ATPG7EjESlgXrTceHqHy0lBobyVEzFm/C2q
6F8pSlloXLiOf6WxZ7wpz9zRAxYJAgkT/WwgDHqpbsZPpbTNqQMDPsD61SzLw6Y7
L7+HEeXwqvT1ECRcMdG7h4vswHSegOpZToDJkwNyQIzr2+aWOeoDBiWy+OJ8oF2a
tyLn2SySciPa9c2A0EU+C/cp5nj6647GsBkiu9kaGO82HrH5yGaBbBqmuIfv4o/M
yOCXvbKh8pnB4FlIEm+OY3bmltQQ2W6WvaCN9Q7DBZmWWTtiH9ZJuc7ljoyg0O3k
oIdkXZnSehJoV8lMWfW3qkxKc6wbz6BWUti7eX17SoBBeqnp1EBL+Zt9Qlv6uCEc
+HaiDDznZpbxthIUMcCD2Paw5pt1GYidJgCkVVlGX+LLAtsa1KncwD0FK18AMFDK
KgG00sL/Vcvuw0Sc2zPiKqgRUXhV9Gu57WjIHNRiBSnISSKOXFDmyvV9nN+OZM+J
77ExnaxBrskebRnAci/enRYghpF2Oy0/WKRwF/zXr4rYSzIULdIJLY7XYAqkctxN
iMWifbUQzmg43dGsmzxLFhF84Gmj64xyvIizP5j04zo7JeYjJF35ETiS0xM5H+cu
eItTdY6sMIq1L7chUlvo9x1pk2GmGM/ab6YaiSOj4vTjV7wNlZ9kKP0V7CQptuG3
K+x7RuKc6RakVwUFT4Aa1C74BiLB7bGYJUGfBsWzLQICTOihLQbIHmyi95IpSAWj
kCb5H3ec+Nqs55A6gFvNo0tK+70efkVs97Ru1xqmtLxsdXKk5y1gSOFGmC4ZR82r
E+Xw0HQQxM+0t7G+ksIYCySFG7zgc2YkcLjLk+GUn5fbCBdlGcmw241zYzgg6R7l
+zJaQS60XpzajSCV6jDcs44ZXkuh8H1BMKalEO10is9pbZxqz2X0KPscs7GAL4EJ
YRsRYBupbM78h/GJ9fsX1ws3YbtjlQFxpq1C4rgk9g+k/Iezg4P3Gz3DWv3At4dT
wajm49G4zrPCTAENDXNXphhl9CQHJSIOfveHAHUaThiiTudJs0odeIaq3M1lWzaK
Z3NA8p1BlI1xr34c7ovkbcMTeiZK9e1Hwn6/j16vNBNme4bTGW9c0qpVfSseX94/
AS1zQbkcJFyQvBOmHW90Lo5uwQkCOR6cHmrWiA0ACJogUBMfgybp3uBiu4FPWl4M
dgoGKNnjOeMlqRVsTbM0Ag9oCd5XyLcQSLxhdEXZyoZCzRJ2sGmFs2R7f/d/DfF1
y3TGS206mGttfbFhSytCIGqZsMqGNP29VUhqIC74cDPQ5OiYBFF/yTi37Dl4kXcf
zs3/llAFtuyoMT/7jcN2Apuc/Cn9TmQSFZbEz9Fpf5LNPMpoaDDMCFDARDhKXZYY
s7DDmp8Pwb/OwA7TWv6oYSW8MLj7DETlJm/uRySHoLnCF4HKUsSpYv4JNTDWERlg
Rd2I9vJY7dSzL9rJu4TGQpOz4NDkdmVIp1FkCPxZe6MIByyrPKLiv+DTKfVUTwHA
tjg3bbra/Yd1uEX5r0ojiC5r7gb0Y2ye8YVIdP5pNicU8UfiVzcF+gwKBonHPsF3
c9pFOedFrN8mGZFk49bW7KjhnCJBHtXVC89hfnb50ozMOxMNbH/Sffs+u9wnwk7z
Uzw10h9dV7Fm+MILkUuBItDZmlHE7Tnvz3TA20DpCOv5KpknWeKrKwmMD2JmyI/l
2IX6YulVAUJvoQx4/l748Qpk85OgxM1idrmfnr5HwEEmgalKCd/WB7qHvdlqrvRy
0rZeJRpOc6f7umURfbdCqFziEV0nW5yVhYWIvU0wzeFjes+p6je5k+wLXlDTJ0D8
E0Mhs0GCRWkFJBhgVRmJ0yxcY1mguh3mW4GIQbV2fnJLOK7DT8DCR03gk9YccifV
ph6k3L5gKucnXoAY+dCIpFUVluT0fo/9zDsf3fJpqsiH3A9TM+1GbLj7OfIzRxLx
sFPB+xymGxhN2JFvmbYE6QLCgi3WsY6yInw05aWUXldH3qnoYsQyA2LDo7tDyHs/
L8nJdq4yaig+s0xjEH+LIVrX4vrwWKo/3ilJ8On1SedovlLlLoMEpIUpIhxoXGMF
ZBz5jyX0WdvcQYLtSTRp4dDOE0Lznt5tNSHroT8hea2O/kTpzt55BJcfZC72jN4i
DGU0p8JDinuO4hwpzn3sne/OF4uIfm+mfu2g0koSaDyuVoow/q69zj5KlKVtEP73
mRkhqmXp6aN/dMPg0LxNx4prsC0Y/fY1gcLtVninRZfJdcS92cfFYrnFMTi5+DOB
eH0eBrTkCSDTei2eFWtSRCoZOAFepV3xjonVdQBVHRtuJtz2oT+mYupvBmIhaqqN
YYq9E9JC/+Pbm9Qfnt8CdPyY81C+Y3xviPV7rPXKsdXWlxq8LlgYgCk9kMbtm/oh
06LROJ7kmSfZ7ZHhEdvl1EW55DnnDd4KK0z7S1g6LBCtIlVC52yfICtAZNnOUz4d
OAh5ADbx1vqyIx3EPBmp8RMONz8HdEk2qIVAO/NCvVceezawYwZbh1OCGGwoK3MX
APNzNmfyEr/CarNHtyvsIeDT1L23lBwIpxHGksfJlumIuz+Pg0DnVGVKZwFz+zyT
Us5MM9YKaa8smBEGw/7k4hvi34nqPPtMCxHd218MqsTYbh8tBlRUVyn4767PHt9w
4rGHWL04t7VTMrp34bjEgsXqth8/izypZNWhdiob7B+WKCcJFoH1e7EXmp5og23M
HjkXAPqEGegf+d8LnItd9RAjQFfk3nF6V/cXUgyMJj+VPxEfjntBI1EuxNjolcIw
ASav84S569yRC51fC8ZkRtW6OCxGZmGNdIJMQ3STkx/ceMr48KS0gEwjAGsWSLEO
r5a9LWRo1y8iTckKC4acIz+FBa5GLIzJhXrYMMckfWcKg6bcNkxn8LJeFRju+M5A
mrohvwTEsioaKR3dAu6F8HaMSlYB0irw6o6h72wCFHnY2SSLjVy0meXi4Ab0cMB9
oxrKh/Jo2S1gWFsy3dCjjPiKlfOLudfMhGmXnglmuOTudWOaLFWKyGDFNc1BLM0i
hSmNtGsvkIYLyRjQR0c9GJgYSeEBlwIPk1kvLksYJmkAZrczNd57mEt7Xv9+Zmf7
hI1WdGaBXEjKPuZ6r9p7M/GSCyduzPEcwKcetcFMZcC5g8YAm0szpZNT1OJaIsoT
cTbubHpckwLvUXOSHw4KI8wn5qb2pO55VRJ6VU5YeDLzOK0fCaQeYjvPuM+44T0e
xZvojB53ZRgN5tNJk51Fl6M1C5J56/ixySyOFTMa+qNqDUkAowu7mM2aBULPF9iC
mT2ZP5ReGvyObyi0Ok4o8+7eD9ri7Faq/sWm/92m7hT1HHsb8safsFvSsnhbpnQz
eYmMQYrHeP79Gd9GDnxjUMkh/NV/ffjvUaniTMR29JINxcSxI2tUjcobwKa5jmT1
h7atXU6AZT1XcsQgvXLogeF9vfWPeqtiQt2k1/rzTEfQdNusnb54DQvMVLB7RCcl
GMdzHQOgN/id0cUPD49Z0Og445hRdgPBw4MK+3egb0xR70j088IgrbCXFvyxElRD
H5d1Nglg4Zz/GwbyvHIH1w9uGBMVoxO2ax3AE3ACQhUpkkJgtMgV9J6r9uxHzLu7
ktTk6bZfYk+6flK4XskfC+yC/3SmXZ3CMhPr5iCUcVA14wWadZICW+HE/LWXMR9B
dB/LR1C5ZQ2l8UBL7Yxa1VYff5lVf+oD3bchheV4ehnC32BtiuwInCslE4EVyd4K
SIPp0bLsaIxiMVWNoKG5eO7Cx21ctvEGbVL/MiqLV0Yu0xBWFvcwPORk8dNKOVDn
JuZatsUbc+cAWIqdrcAgIQUjpysL6sgLIKerBsrhBByEcRo4nCWksb0ZBFxoRTBn
6mE/URfCz5HT/g7CNHrEk0TOMGT2t17vPPxuN+N0/p34b7PEjPI+ZOjlH0UbVfHw
T3Ejiv00Q8AlDfvZRH+jGhDe2Ljchju3rnB3L1VK/drIp57RX0rBxPIyr02+woKr
9GCH9dvZHLvkiVJ6Z6ztpgSbMQlghM1tnjcXKGO8D1LsGaplize8SR8RGb+FjHhl
zebwDhbLS0jBNkuC+bAiYxbBcKbluomoHQ/bX2vOZbhkkEjwadVLC26Ipd0lbYc/
4clUIVhrbMHhLj+3+8E8CUFGNXyyIYxRuSxlj6Wtmt1pA1cVfo+HHJb/CXxlKDTP
4ntm/LowwkIJs9TrtEFlfBhZjyhKcds2J7NPLrly8nF1MRAE2CAPQ+MeHYc75wz+
B7Iy5/lNGgappH46dR4DvE4MgV2qGAxESdrpU16gtWxiT3y9dY907rHmwI4cRZtb
03vsgXHkXGrGn9oqRnOGvenr1Yevb2q0Mt126a6grUvzbVmHHw6vyTFyQQedqYlb
F+KQS7y3l+sKbYul8sVjFp4274RKB7E/XUiGFDJC//JW9PDFCBNx/ujlPBFir1wO
19WdkkySpseh4R+sMJaquI3vuPZLMmzsi6jN+quCXHddfzcQtj4/UygysfimW6X0
sHF5plq/z36zDOYwm9n78RDO9kBvyGKy1p+3/qj/aElerHab8dgN9636nxCuBs+p
vaMBmBrqvVG0LH4H5SZ3SW2ApP0js9JO0ixghvUWQZFaxpyavICp3KWozZktHu5I
5gNdsKtB5uzMWsGct2O5i39euweKH1TqZvoOKz3hbHVpMHgkWbCJnR2CoCgDD3A5
rqpTd+TrqDwqBWUDfAPctfeDQf3fVMw2jgpjkcceKyJGQCEp/CPeAx6fD5W6H71k
R0MdkVsEIm764Ud+exvE3FqhlDqyOy9f4464LdUdC0bDRcZ7O7j0cypRO8T9/2Bl
qxthSNORe15Ku3VziYSRkNtPxcwbsevlNVcekae26uIOqEHB8m0DKxPqrLDKzgBy
OikQAOoRR/KoB6EZ+BH0eNAaBNZmUbhh7VeF4nM3KmwOqelV4lTd4/XcLbuGUQA+
diBCZqmCd/l2iTdXdIpzE0xI2vScRtFfYzplckAZuwHIlv8Rzb+zNYGpWa8ChK0+
VjpvyUmAchyq0ZeFBJK7hKK29klwH13YSdnNO7o3pBi7pHJRJuhsHmwxga5K2jlU
l3Li0S4YJxwLnQBo6dRtTPqFLbZCSh4cFn1QygdJSQyJv3AO/4Omf/+k8p6iglLt
/bPJbcVe9js97SC6a0egHu6KlTy7xgy+4eY31Y+MKRlblZscGGPHPcZ5BkPVzDBj
TABgelccw4uUzcqhhE5tRPLmM87O2Vl53O74IeGKy54wTcr/3izAZAewrUcCEHTg
MXL4AdoNniCj1PWE8uY+rroNGpvVxaFmMeqlW0py6zntYjTPpU8CA1pfiTuQhM5J
W6pkE5p+wsBuRX4GH5oQkRGvXlOlzBhEhbsiCxA2y9515om5jp5PnwpieT1p1JbP
Ax+rv1CUUC7QqaBUF6bcetepnqtPDx24aLztvsRW0LdoqCHk1st3NA42kn3vovwQ
s/7Sy5RWQI8wc3S0VvFtYRRqkbDzCjwrHyTL0ote2jM/r3+Pzs4iJ5l/JOCpdfTX
bsFAhZoEjoZRmnTHhHN/1gPRjXiYpQA3twxqarWlhhue2dAdpxtXau2kmG+v7B6N
5oXPLYus3nQYi8D79R2ZSeMf9zvVgCZYrBliXAk25jDLZ7jWn9ITzAePTJsHP+X2
R0r9jJzVDWwYKvOZ+C8WvqHj8pFs+3N0P3T2cYm0ArfpafUFs+T8UxAoeF7LGXp3
qF9rXb6mf4X9Z6+RSzvFDN+iTbXVHVCZFtWtJPTZ0N0q4POgsGUknhuYVjkmT8FB
B1/0UP9RHH1dmI25VCSmJ+e7Ne+I8j+u5aqMfEFYvOOPXKI66SLS/sFQxOgIwq+k
ZH7tiEgct1XUKw4eeeODWuq53x3eTduPfoG97XCIMgqMLUl2xyLbR4gQHpvPk6Pl
LmTkjtCqZQqLuoz9/td7Wp1mfTzd5xxcCFO5RJHKwr6KXSq2ZTa8NTi09i5NGF9h
+PJNtetByEZp/BAMFlPwJEFbz66NmeYZlmRC7fQZukyvSBcNfISDhkUFqeKpqgNM
tr6+4M65AGzjeG7nLXl4nF+rf9bYigzL8bvKfV3B7iT3rJXjMxjWJHy7FEI6lVve
2ciyVEWSVGwsn83vH88RkXd52RBN6+cHW1H+78PDVwc89+c2VOz3No3naoD1b9yW
uNXML0PXM+V5N5A0XMyAmTBXHfsB0MuxUFPAimWFfBsj+4iYmLmJvGwye9Kct+YW
b10KdeEApz2nu1nYWaOc/yvL5y3i5RKPMEUpn78TIefUQlx5YBiqwZPU1kHXgFtO
8nzl0FLjFQSPb0tYrwClmqpYN6qNnqft3byRsbQ+jF6Kw2ISyP1ouhJcX3dzob1X
2tact84T3OBVLyDyhtw64HtDVdDPsdFcFstM9uDUhpGSOkzOpEhSSrOMIiJcyuXE
G7e3V8Y8nuXUX7aaMJncyi3UZytDj7RYewGCnGAukiuZwrHiX6UwKHh4f53IgQOY
Xqums1RzPNPPhD/PgUlqlEc0YVqxmCHMtPXY9b8+QoO+PBOrdGHHLSM0fuJPikfo
KLJDssCpuXwwtL5+I8hxqVEYnfbj6/sKuzrfwCOXoqwukZteIl9SLncpOH7/GHV0
Q8+LF54BDwaPqDP7c5HFHBXzNcXebEl4eBN6kuiEJtPMPsBhmJN9yOWtT//qRfVR
Imu2sb2rRnsfrWMO9hHkZIDfZRQMqexOYP+gGT53YmmXPe5F8lGa458zn6mlVon1
3Vg3kvxrUnCA2kNJCJrFA2kDRHFsupq4N3HlrAHyUeHg83EKF6LjFvu6tVZUY4OK
L8oy0wDiwHILH/j7CWRX90nTVhfEBPGejPNqwhBR3ClknPiTIQ4wd6fajfGseWrk
gMW+eqJcMa9dut/dtGwmLP3j5PTTaBmlCsBDmaR5mw0+r3c1Pl/fmc6s7KCugAdo
U0pukrZ4Gm+7jIZ8PSxasZWw/Qa3o7wDwVUlWrKHCO3JNCOTX3pJAddn3yPs+Lwh
SlE/D3lrpVObqmnaMjLA8z8X9zsFGpVuqNcP9m8oB7Q0zRSQBBWemuhBZBs+n9VJ
4cn9GahElQOHFVs0dOBZdo6Qab714olQ/mMLGux+F4doUOH8oabfHqOehsIcR0lH
1LiuJrm3f4+qOwxRkUhPp6jdugcTMedVUTNaBhYoGZwm6Evfkojq0Ov+bhc01tfg
Nvvym0jthSFuHwTGk9pe34axQiXEJ/7rzRourBaazYZnOCB1E8pftn1MvoJDaJ8V
DzeghC9MNB2sGkvcveudRMtFLSlq3ukVhnsp+QKbbpdQV4KyFCQsVYRN7yqQRBUI
nqaVuqr2D5lRuLkTopLnMP4obytB3WZsoeLNqO0mzXpLoyqGj8D+mWPd4se3h+p9
kNDPGgFHU8UzWWnEQb3Gyp6RjjJintgw5OlB5olJCNgdJnUhHs9PS+SPyEyEo2dO
osomLz7ODJKYsMxuQ0GwWUaPsfQLo/zXvTejUjAljqvpwoinvWBKWv0oLwSsoxTD
SEIvt9ir6yopxCrWiHQJNbEsK2NdWEj4Yr7Pa0VYD0X2QQPibtOlSHvHTkcN1Ym8
+gG2iutWFy6ZtnB1djnvhZZYXYBx5Cfg12fdSIjw3bj+gRwdpn8oTMznqln8LAds
gNmjXrWVqJShTUPVUP3Ac+vYEoSvWVCK+JWE9am2hlLhrOWduPIPQKENs+l156TS
LMIs9nvV2hfcM3KzGUoBOWayTRRxxjceJwXZxOggQy9r7qNlgtac5+FfN02Ii8G7
dOM+AzHuQwh7XEASs+sVhjJkVnl94li4rXlAWCZTsgtdXm1r/swEmPErZDhPAeSd
o/zriIsmFmaiJmkFcSSSMc8vjTWd0JzWDPZ3R/TBN7XULByGOZ06sHMpTkUw6a0V
dA66DqOfetiEHBpyysHTgnKhtuPaNc85l8oj7BDQeWBHdwUxFQmwiQ0vU4fk/X+f
ysH5ZQrfmcShD1vY4H8I/jSdPsE2llMYT5r7WgJWPx2lFRXRhWTW9uMyxirvgP9n
V1S7U0eqj/+lbt1BL55zNtPvB9ygu6nnkoxa0lMUcgBIxbFoL91aIN4WyX3qouEf
hNz4JnLkDqfAdlcMC5p5MACSpx+GiGvOdptkH3SN+onxTpM/AKr+JrE5E2meT2iI
yomKUkD69n3rG8DWc9Hc9kM2U7y8jiuotMRiN0Sy/4SaJJxppzpp3oDYcfZR4/f2
Q6qcoDr/cn8Fh2lYqX+IknEhBhBAR6T2zep920cf5TiwxrvwXU53wch02IDXGmGY
t3bdKBAIsdxwzKx6plKIMjt8pfwy0jmF6dccuNFwclJf6IIvBLh2dylQ7QIKVOt2
coqOSfrIqKxM+VFlahVjoQZmg31V18MhLlyHGhVlB46COPYPuPdko+az/3Wc9wbv
6gq6ddfV2B8Ikwy3J3y8fDLX3Al3iuGRjek1x3OeIt7Fg1+aQ4qwPGtIHlCDcEJ9
KA7UkQpg5wsPhfmwB/J19npQFOiCtBS75Zv+H80CmKGibGpfVUJu5AcglBbQJm1/
nCiEFX4DvvAfOFF2zLQ66kvyrEfTq9VVlQMVa8nV4JvaQrHrgDIRE9N9E0W7ONOG
y2ZbTFK3kIT1hBE4H+AyMdnQ4L08vch+PKVlDgK+PGxkGz7YgpwsKqcXaazytKFI
YgHdOROwPwPu0fgCyCUvGJJV4Vv1UugPKO13aAVrMAmD/nKlK9r1yCYSPQuiM6ba
rHlGHF/aZymt12wXNq9XkEdUOfjI3mRf3WSEhJQSKHAKL7nnWHw58I/bziGmukuV
2R9CLobmsKJkVFmAXUo+9Oaw9JhpV8isEo8nNAF5bR5bMn76kEInGevTmOoiqheD
8u1YNodye/R4ohFk9o0GbOCNI36cCyYgyyjp6spKiv5xGoKD9FNxa9XEOr/4kelW
Dp2XZ0ZiZR1V+KqBUuvZD4MbAnZ/4cXnM0+ykZxeaLeXaSApdWCw4tpyfCBra7dH
OSFOSTu1sr9qP+8OoRG1Xboa4x7xa7NF6XkTObAsQpvbEnBz+ZQo7478XaqePoQL
rwruiqBHp1/sBMEtKyJvvRip/PfCY+qF1N4ZO8xT8tSMFZ2+X03P0WWfdkavcNcv
8tUbKuAvPDq6IBS1HU0Ez0h3U7hoS56Iy3r4MsrrEiqB4w4WqiACafpt6LQwO2c7
6acdnV5XSKFwCBd6A9q4gkMpH6x8TK3lKSqtIVLNHBbbjzxHgrRXXKvQ7sfGpI1F
nVPrpSvGTYsG9vctF34nz8wrZDBs1vG/VNQWclRD7eMd4tqarhyDXLs6+sDjpDo8
hG1T84VN68yvnMkafjJBBVYdc4inIthM/wsPNyF/CBtYi2oKAGLVpW840Tq4BHMp
cyzRyN2qhCorYWQnYA3cRbx+DOS+tb78ohkAvAElL+YqT/6hIVk2SAXtGFxh9WIS
/SlaEc21+pYXq0D6LpfzRRnxmAk5a/+e0hTU5WszdgCiUMsEe0mn70Ygtnh2/dVd
j/+AvyYqv2Z0moMLbfGMVvC3hYfecbtE4cH74mqmqv9fP3gFOkZQy7SvWXhybeUY
V1qMm0rWfyAlx+dWe5kJJuTMAiVbL8uuD/3GlyMOavZdiQ/7CVLD0h3cJP3zJP1h
iRLDhYYQ15SX14oAEgBE036uso+QWNZ59x1Jey18YvJCTzeVkvXeqnUpfHuEgsy6
wJnpMBWUo5slY2nyZCfRRnIJReZw8NIz8lxblFDQYG5mYK4kJlnh1PqGLXr0+spv
8n7fxlhWG21qvHAcd6lOniwnfdpe2OsYKV8lH++6801XsdXKwhrJWHSOmmoazhoo
EqrvbQ4ttwEgQ66r3KhQD/MIonAf41+87C5UZhjW+vrHSI6pG8LudM2cP3+VMec9
0dIF0ReDdtUb3Zrkx37DtB6hSQ7b/avC9d9+lvFCY2hgcIPqDFjKCvm8mf6p3m65
YuWMucRM5BThjZlNgTghrZK6k2JSzvkZrTglpV4LSg7CADOhbVgxoJLst1JSKFDJ
yXyT4Esf1SFO5nhs0u3WKAMqX1W9z+nMCALvkbYkzskO3bk1NL/ByBZxIzz2JRdF
jE8VHAMAQ2QA/MbJamcEG8gHKZiMPbvUk+KAis2QZrDv1YjxnEOZaaandfeJKksR
jy4kvGCfpWnqUJUJqgk+/LksrbKBDV/01B7vlTIKM4DTorxFBFgEliaUmZT0Veu3
kkJ/L8TbrzPErqOBfl2YWN59YaS1fs+i5KRFJghU6PVQshROZ1AfcbBYN/GMg/Ia
Gj54wuiIe6lkL9WIhipiB24+7/B9g+HRPfBYLM+hSdXmUz6Iwm3aoh/Z0NoIOY/4
Rj3cbFDFNfD0ISRnf7x/+LywbyqYi0GG7wLs/KjiNfFOpQcUYKhTD8KKLVKmweHP
GGiFz/LJHCgf1NQJFS/9gbIKxtImOvt6twwyhLLB84Bksn/zR7ik+SSvXUybCao1
tLMUcPh97TM0Uns6ueEoCeGdp9HKoK6mEeB8Jd2AjP1eja6eJUoOFnHCYkvO7UNe
b5bkA+f2OeA05VHEq0j9fwOsb06m0GUv57r/9v/o1mIxR/7XOaqXdrHCl+4RCU53
xHvdadWhynvT7E9M+TR5/T+LTmwMLqKZybAwQGIYIk6LPfZF51kqh1ueaUAUERRZ
yWDBoBk9CctwbEo98IN0vNpNR/YUam77mX2iIg8QvtDS57KVPnvjmGZCYkAuNWhf
IaJXYeD7BEFFqeH9KqUColGo2PF7cUUhEjGA+FZdiHydqV99fX9Zz3BejLMBWjQg
JeeTao3xDBRil1MNb6NdxPQrthTiNoBYkwpSISY6FsZtCfymKqJVnA+DBBypWFSe
9WmHjmYADGTJrNMO5F8JPWv7uPNYXVr9D58mxHbySsOC0Gyhg0GSi9iUtiap05dz
BF1GSMHI0oogw3VBTBL+mhTP8UFuwoknmysKO6VvMcDvNH9l0pwUOb/8INxjE0Ck
Ily4RNy4oL3MQrGgEAasWsNLpCf1In1gzOMkfrDtykrqGTknQKetO1i2VnNzO1t7
+4iwu2KBnCeAC4fj3pTkj3QKq8NDMQRHeL/LpA8sBL9fce0rk4gwI2LhhBmF+a1E
GWAxJq2xs+IMW4kra/KfMsfd1A3lhfhd3NTlvoFL+CnQtnFKEYIOhu1XL/Zo0/G/
8E9vw2fwZ/zrhLHQkmLfd3Luys6bSbAoy6KzGVH47kU+fAZRMBjyEvTzJvKRCM82
ICiaZFsrKe8b6VYsvagJsLfDZiKc683HfnhGv13OzFHAGhHnAje5tyNANjVA7zCP
EzpDRMDdW2kBxyq2yCMBhbmD4f/NpmN+ahLhJ00wC4wgu8Ke+vIypOQpmXgn8Dnn
YRpDwp9pONQBqUiFybfIvGUzDv7L3dMHXtbCw7YhNQGEF0miKPAonRjUNg7tiwWu
zkkLhAzKxlTbG+VNBrDGoqwUb+Xi/QBaOB3y3YizKokRkqHjedpbexHrm5Qu3JGE
5w1X4w68FHbNtWegDCdfJvBnRqUE/vt8e7WCuhjfEKIPOu4uExeUIafPkM2asLIQ
hhREAuAYdUoGl7GNVgsJ3P59r0ioGCY87yg+AfGiBTc/Hq4L8NR4hx28s1DURacF
wm49KARhmN1XLBOWkHiSSu/ip7gmFUQPJSHGNzb6MKU+GYc+rF1Sw1GDqyzJT3oR
3WKdk1Iw7EOzKTdid/Nd91B1xW/mz7LFg9nF/Ck4gQDm9br3rBVq0gg2dKcJpRgE
R6wiKSuryNJ5EVaaEUWf84BNlF2CxSgrDHafQB7rukO7NRg9TZp1Z24zVHxh4G4z
dlS5wosJwkEv3NtRKoQ0eA9pjaHr1m4yXHET8wRLPzB+REhVHDjUOShlbYDkRCre
l0gehNSEMHjyay036q26qequ/brdBkVSIzFiiXs/GLHX2P6g2QUdgBC7WDbqGtj8
1sDCswW8vUyZj8Kl4/uB3nZ7oEX39CJNGdGUvLlzZt5D78z5XggW71tKKNKEm6s1
0F/vt2pit6nz/GXHY6OeajTwjAuBuTwZpC3KLDjJjwcaZcDW5KSf2Qr2s+B4epSj
JLJ1fsxbNcYb9CDr+B+Abc+4TwBKio7CsNyHk1O6yuF0wG41nQek9h5Lq5Med2Sa
v+xWDPwa6UszeK/YnC8avDt/WFgpWWTtb6n0JsAPDr+NI3srsZhW69uSECp+qwb8
yX+zIPxTGjmnEUjhQVCFpQlEWlIgm9lQz4sIVTz/NSp8lfoe4h9h0vviu+FVrcIF
l5wPeXK2CB+Rzl9Cz2sg7tI6Y2+3XQwNMS+fFduA4iywPykaluwYXW0FAcjrszCx
KrvRcbK56P5gmbvhu1qaPP8gWfD5Fpw2OMkPwmVFEbeqtsHf8urKYTpRwBr94c4l
7TsNIDvSlGXUow0gKGrcpPhg5W1A2pU2ui0UgABamrGwWEmBju1fulqQEBSd0Nek
nRnYMEAZt+5OlMqQUCPMHmgKQ677EMfdHO/pcAXxJz3bVwcX1IWtjN31NQyKedL6
vHM85X28O4QUNqw3wuS5HFLYbJ0Ft9PPExg95i2rXuKuyxYYRotkAmBLboIkZtan
y50Dc+XaWkyvaYgvh+SvBZAQzhkAANqixbfJ9N8F20CvWpQ4YYElrybo6EcdNI2r
FdSYSyQr1/y9ATgdOhoKVlnXHIin1vy+uaZORr1igi2fDaNQHsoagY/KSJYq6qfk
NT7BRQTzpPkO/1cQIBkBigqcljyWsHSmFQ0pL2qzsZoJarSPQ0jaevrkAPIqb45x
DxbKkbbCom0j2TqZWvrABxC3chyCW3viJno3UJkoLgZSU3ehdsMbTZwQK0cT8FSU
xya1PrVNh7Jn2FE4trH3FCVgO+pPyzxClbp8ztvzgckYrTuwLN3arp08xj/qHEC/
vqhZhITpzUAm0bS505Tzx8gS/kBl5qs6VJ+ZCPgkHK6TGscCp4aOTwwFsdEu2Dfn
q4BH+WCHLM4MFqUvw+BvEn6mtroNOK9gMqxufDI6Nj7A+QUR29ey1ZY5LpYI283n
4gsYwQ70vQoKYtXoH61N397WABHL5nXmIkp2LO7mVQkcwYZp50SCvgbBITWCjawr
O/7E5c+8inkQfgjFfSh//focujhnFZTXndsF0zfIbzSXrPKfgBDCcs4he1ci8t/U
o1G5a+QwoLuFBlNdsAUDgbGQxrQluXr45QqQtAXh1GSOAo80rh8yyIwzzkTseu8O
kL/fsRm7gdbC873vE6LRtR+ngfzngLCSb6/HbiLY3oLpAYAGzMC8RNkdeZtVY61S
0pxvybxQ+vNv1pS4Gb7Dwh4zZnHBD9TcIV2YeOaXH0PRaVE6rRKUiJm+4rpxiz9u
R3poZMsjyQ9CUE3YJKSP9xw+pLK8CS8et9oO65L1pUNf4dSZmif7d5egsiUigjYw
MjA+UvX7yLLpG7S//k0muiJ4Lax+Vhnxsn2aoJkJ/VywRq92OdpbdbAOCF2I8vAD
IYGwkQo68nn7Ad3anxBd2enpTP+45U69bXWTz5u8S664VDZKO26Ex+yINuGXRhth
kihD/y++1ACa5HSS8qN6zG59yjrSX2/z1c1SgC0kfOEeIDBhNEvUIroTza7JK3tD
g5Y9OmFOo0fSjaI8Nhw1Q/IKbFbHlnXxqv3Qz/6giH1KYv5/wQrq7GqLkPqBMmpc
QKMpnqzsft6WukdM0tGHTgVrbLW/K5ekeIn7KaYnoFeIf+aLgb3CRlXV4IpTrHUP
n56aE6AmVvySxWygy2HCfYwGV+Ro0W0fFm/CBqarSQX4rS9y5nfPC2dFi8jkGbWm
4ChimwaC3kpPK3O3+RYt6xSbk7KqLkxu//AsUGq5ZZ0RBtU6k4/9NEsZjFWGng72
avhFHHLgVbCTspq1VOLR+CEuklyesMdjHaovtjeIBJsMKQjPvcVYYQBI3J810MZL
wPpYrzRmHcj/soWc3yTddPgigKJ0l12B+SEjiGclRf79dJpgR6KiPUDxudpKwl4G
JAm8lYA4H4PVJJXoZwkaUDq9VIA5vUD440ILkYfqoymyHll6GxQBzrU6+Ft1KFBh
b4kBGMTJqWsbfNqPCC1V4T5+8Ky1KnzEsWj1Jeob2H97l09DiDNN05Yi0SDBjwKK
QEt5iEGX+wwKcSoHtzTungw/wmXaBAphp10hTRxvBPpwNm/fXyA/GtD1ja3EPomp
tdXERJyAlA4oGFsd9ovtPtEsgSQr8ta4EDmmFV2GvvRsE/6BUm6SBELZZ4jC4Pk6
BbEUipNYLy9WYZ3gEH1XgBpJNVDURO0B97T8jRDTnaUlLr20Bo5t29gsk9jAO8Td
LhTVGOReAAF5/52GZOwFWkiM+FT5cbDIoN7ZSPBJl3o8nYDl8qUOaJpS/IQUNN2y
Fbm8IdxTupxB7Fmw8N1yfVSXmqdO1xyhPJ5ZGjJIe0Ei0C+lpm/+ifbVlHnquzwl
0A9yo/4cWRJZL5g57lJ9q2C1nAvptT16TYFBkEd+jG0qQBtlq9xi8L906SHrwx/m
fCY7fa6BS16leimLx+KfHk/4IQoD96tAbl5DoevntVrOl0ofFn5H613fVGm1x2XA
NIJDbzoF4o3w/O5JZrTsV2GTJQvOySPiaCC9PuyOi2lwgmU9Ydqj8qERFaH5EPoY
8gRVT7VyIsKj7pcJhqv8ECKJWWLZexXUgFFbgB+Q9aitTdd6ymKzQ+9yLR3PLrQR
WhxuuwriwDn1U8xl3e+7GXXXTGCKI8QRKkidregtGX8ah/MrT4T/BqwUVX182K8U
/GLbe3W4kfkzeEVjAFs+pVs4+34AuQzntlwmQiPBXScIrycQLhEkx7hSovidwzWP
RM3SLs7ziTDqP8F6M1YKbnfTrFdOLRsA8bl8cCIKoRiNfc9sPNkoSy1l6CF4eZE4
QVm8DEuLkqXApVjvIOSpH/hdqpU+cO4BKLdm0PrKjQPSYRqI/UVYrjdDohUN+fXO
vpyQ/vXgwxpURtzF4ewPAJY2T9s91sDhWDf86bZ63NP4cYmkrlT5EGn2waIII2JZ
aqgFkyMPRZBeO7d/S5XeQhZzFKXD1RBZNX0Wkgd/NpHy8GspK9HDl7yqbz7FQVvJ
1pElMi3I9mz3j6ST8BtVzPM6lc7jG/YYRB1xbHofVNUVbT/+Dc9XBjKeCo6UTErg
+xSjCdm+ByIY6lctvoMRfz7WI6K3edhlaXgaAboQGcZJ6M+ao1agYsBLPogIhFy0
UwbRgcn+P+r0xEzWOHnptv1LH46H6w6kJqoAOnrjhHtwT22tKoQBFxRhq4pOkI4k
VyjhXc0IkNbYcDtoSnR6rndKVCjIkRX6ZRC0oCVdQL6MztZAFCRcoK6paB4vN9SA
zDR40JrVEsJ4E3e7X/0iDGrwNjWJvWHjfsIGzKsvxvjhOtKFY4k/L9VTSS4zXK7F
m3sneJ1zc0PX/twyv5SDKbjd3bPPlo3JfNEjvxi3upQbB23Kao4SmP7DxDav4bxz
4VQ/GwgHmEU/GOkheQE7tHYNEfzyd03tvEcLbSebRTimSh23BHJSIzEpqA/FtqBu
OrXuGVnGQDy2axJKia/plkEcaX3vXV1CTMpBsUKuehr4rG0dg8y9cFk/8oyj8kt+
OrLt/GZeqNCl08D9ZH5XURfRKL1rQ+JcmioTg7npPsJ4e/4NMRz8rDCBDMjOx7kQ
pG4vAzhpkaJucbjgg+982m3URy4/kNyxJvzC/z8CKcA+8+WyYxl+QfMYrWwXHvMj
MjwUyC+Fgw5Nxhb/TsESua63iA0jZKTCjiBddcCIo6pHycPsEF4ovSRvm3j/avgW
+o1GyQUMCjDQvO+6N5+et1IW4nXFOBnzU6mw1YrFQgf9RtVXyPeLbWQ4qFPHe087
6cvBWJrw9HdGgx9bBDLQzUj8nBCY+sgQBWnU1G4b86OeukZTaDjz3NwlsaST2ImS
YpvX7/t8BM7IoKnWQTLd/u/t/t0tLqJ14PMoyuE7TDk4kGD01XWmQENmOjwvKoXu
EReKnpXwe6PciDfT3cKUJFEQhI3SHD7JzfoFeYXDnCFF23eu3fVT7901k+6Y+5Dc
Niaa34ldWjkhs1Agrk2i9mVAjEx3LPXXbbVpVCEBWlBkpeuMN4m0hfkowor+SRyM
nRfqwP8XLUwadzhCMT5Qp0uHWs2oIyK5m8VdD0s1BX2wM2tBDf6OL2kt06XlTfgb
4EatxAPOQiy9eLsbpfBrvxPQAoxskGdtnUiNuIOz1yph7PRkerN1wy6ptctCtvIh
mJq7+AOU4+Uu+R/L5GX1aki6tOZI6v0Jo13gHJVuhXmmKuoNQ8RP/znQfSctZeiI
5SnvpOT+CEuuiaUEV42Mp5KXxvIeTZFJpE2JWdt6Vf5Ug7xfqifS+p9eiW954eOF
SmSUXuY4QB0KqGJT3xsbQwWDOKl0tYtWiO99GKlpfMn1FXKjfE52DhSZoicDHppG
p8ddRJIJ3Rk/kNKXK8BAO3PJePePMWV2tO/osKmZ3GqrPHJ7AWsf6hj0Ys8YOLG6
EX9ZcNoqElmObfpH2woq1XbqRKZ210VySc8+FV/kZsAISZj7drQ4H6ljEtp/TQN3
uITUQ0xTLUoBdvVXTLWZ9x/EZi1cEGNqkkr3E+D6qgyVHEeRX19q1dRpFtqj1oBU
ytDmev4DZUDmoNGi26EdGiRSH4YxzE81KTrb7u1o5JIxSfmyGBxPnfrXFFrZ70dC
3J6HpU5ESsnj95RbyXBgxL7N1k6XK/y55twKQHejdFmVEB9Jjw89FvMQnC++0YuZ
84flN0Tb+ULamG1K9Dlv0mBl4Dd1qhNaZBKVqRevXwt8GGKNz6FN04a7CSHy9vha
YbmkplVR9RnqRmsBeIiTd7AAPc+Y+DxPpV/gNRSmf8uUz+g4/91g7/JnOGc+yAme
F3P1YVuouZ6ZvzI+bE22QqMqylYpbKXJV7rmxQEOac6WAqcRcuhnL3MNIZYpG+ft
tkBvWUDtVH7Sj/sa5pFgS4II73FdnCiq4xrZyN/n44qD1sL8gYbmdKymm/i3dMUI
CoZseH0uAJBqOiyddV7Y3LeUQh+gVzwMCon5LNc+5Wnzw/CdXROLqNTJDLgdux1M
+tfCle1WULCs2sbqII9l6zmRn49KabH7/GZ1qSLohniieaHLAexVfaf4BcHzqKX/
IK8IVOMKfcYpOrmiSjsxLFe9mbdRKsbvELHppnE+MlJ9VaKXurvDASRY/E7+4Xc/
lUheIMB6f7hGZGliutYcvawGq/739rNlg85RFyskmcOOOpKO4+clJSBsvpmCWaWv
Ego7vVHCu24A/mpcsKvmoTeXZJxgLWqyM2qRdX8urT3AMhLmT+fm6OXkfRq1h/Ib
KXo5M5wJ5cUhrIoZGsGak2i5WkWwKhRmnu/XOdYUG111eUpY0G26ElIyFnt3lygP
VERHpKfEOZv98syUqcjDrEiUnV7eTLVd7VQRO19WsMf3bc+zI9ASvi7xldeaFkUR
rSyTTMwa/MGoaRirAPgP7AzXSk6OVDxML/6auQFKN7zzqajIdE/8OnTGVkP/jbfO
tpLUEF3v/DM03h4X/6cydyLtb3y8uy85rGExWvBKo7tlcW7LyVwcLQaB0ySeVutQ
38k/Y8LC7nzxOFErCTWOis4fjjpKAOMvv6LVH6EmddqTdnDaUgqkqI4KUe2/u93v
oKyviDkHXFfgXOIxXQHQgDrM7irPb/trsoPmYJ6ZITu0wzmVs6iCJlUhwUhJvvNn
W3VCuVvMSB0S7vhDv+iskJBV6/D8gVLOdOGA7KVRXPP003BuGyuC8IjtT6PyCmXj
Pmg239z0L8w8wc+q0tXWrUPWOMZGuvPdZqHvPf4OGH8tVOpHSOM46tyY8JsVyOwC
FRVXioyIH1TQxZyhBFIlnufqwPiYijgaPrQauCHluC+oDXgraHaFq+copqBPcDoN
fM7YS1+cNDffCf9UTm+8Zj5Qpce7qPXhYiQAdgp++WHc14fizxFJx1OicBB1Hf5p
sdFI3IXT7BYW3EKsBlPPHy5M8dsMkCw6B/pJVOF/rlILF4xyDGkG8xfdkkDSmOpR
Z0S0aoxjcBvY093PTNJOSvDUWcNIIMhJ7iuV2aVE1o3MXSNBHfWCUDd0A7myT70O
X5fCCDdjwdtNj7uzg+3IMhn5QV3UgFfXEGVn1rtfHxSkQD1t2o2L0uV9hR0GzQ1C
GKkSRs04o8YDB6g1NOer6Y41OFvrebozRx27ht4G1tuJCrSrqORx3EhYKTA5bN5o
oU99fmNltTYnOnozQ8pbdvyOhprR9RndrsFzT2bwZ/HhVyfnf3yn6RxwmWG0htxU
1hWlSiBaP+HVLG4inYhGCvPMAS98wTV+/RHKCkA7aLfpSVs0G4oKZ25N0VPrabw5
TNDVxRWMgN+C+3O2rKPsaQvAFgQyqS9/vZLYkrAw7G5jH8QE8tvizuT/zkhtkxHq
lhuAvhtlKysD0dwz92WVZmSlM37s+lzgkZLql/vfV83tjx4T12AM0NgeO2Jerxdb
PTwVKMCYRy8xwpMl1L8DNXwHBl8fXnB9wiz4TT19EKiXWGtMvoKt0Ly3t+6j57x0
ySklTa+shirQlU0bdyrTV3n0Jx9RBJZos4TJ1B/Md4wLDs24ybKSPZyztH0kY0ke
25SgE6GNCO1BCli7/fXNlcn2MuDqI6ucRjmy1wAZjAU71E9q9ytlNLLzhC66nBY/
4TU/vXDxTrUmRJTel3VqNAWgSte8zAWxAwi3aPAY8QWoKdXJzMd3YuAuBV6osZXZ
n4g0ASCdY+u4vBNiA73NgBXx7m10CYGNXsq6BBgbfd41wBkYNSM8TOeQh85BSPcj
EpsVPxeivqf/I79cEheFAJkJCYJYAt2apJC6fSd9olDtsroCRDnIwnt5c1/tVoJJ
Gj5u5hdfevnVIE4yyG0sqADTxnkeZgFSWD3waqzvU+/7INT4gEDBMbx+kZmj/YMX
3yC3ijYtFcK4/dtJH6AljPEH0JwfgPOlJaoj2IWoukQNgOPGz8zj5M6DKoQ2OVD1
mXfjejXZIucT9WAKwatJbCWE77ksUep8JWveH6MyR0b/yWyvvL3kUVmHkahzH3C+
TOdvFh+0eM2XXGLCFqH5sJLqrdUhmiuQAq77JYIC8bPd9TDP8akwKKxmAb4pwfla
Djw1fq8q3Db+VDXy2RbZXbha5wmxnyWKJj4/lgIBWBQJoLVrCnQ1eztfqqnmgaw1
JiHQo+ggUhMJ9vojEwbS7nN/YwzbGpONJRdoH3+OTT/U+P4XK2D9es+AHsPhW7VC
EUPrnYgHnFk6B1dAzA25nW0ADxMWDifA1nltZxJrvlHfczvzxgEnWcKLv6hDJSpE
lWuS8TdTjfwbwK04Jma9plKJhGx2VpWYPgwGCrXvISbT5zsa+jOzytvQ8EUSy7Q3
vL1457mUBKMY6szklk70OxULD9ZqkZT/gBUHlg27f2uWiZ7syclQaf5xYuRUVQ5R
NicLHyUzb4E+if4g28uRpm1xtzdI58rpOIvywGfOekfDnhRPvm3cfYmB1nGWv91Y
XoIPNg2JFyw/QQ959Pi2EDISdGkl9kJnbuVznrKy0NhBnB5acad6KaVA8h6C/4gN
FXDvS/e2azSmD1skmwXyImQoa3DTIAJo1uf/bNe5roG5GA3cN+FIKIF3kWCAaJdn
J6Da1YbnCE6BpTdLYl1oQNx0VeJwzpzoL5WtgpT+fnSVxkHtF0SJqerLAmw2jzjI
SUn4FUfapvGEFHrZiZxFZqV6VVJnjKmZvautjAKyXqbLU4ExsAs5ni2s4+DW9xAC
1Qb3o9DArutOFIre7hhMSc3k3Av4YQARnCOeeNT2lkAcGGCmU9pxm54Pz3VqVOTl
q9hib/YKFJcztqWdR+erClbjVX4DYT0N5N7ikoW7nRvral6hzO+THTbZg2JpXyeA
brrcJVgEJLdgEyFBhIhBTvyL61zTT80MPzEetRrey94IoXIfpDNkKtrt9fLH4fRT
w8NK/RLQE1301CrrotW4NLlku+e++m4ATWOoZu5npakUgnlvISKtN8s0FPANmYns
/uoWwvs3aFoz9gVbU00I2pvNfKDPJyxa1+cOxYJLrO8UlASZWcl5Q97GnfxBeSWh
QhTHIE07a8uZwGaLz3Vr5fHVMAQ3excGYq4+9X+oMQ+UgZyEBA1F9JxFSvW71Gqo
LPG1W6pm5O5XB2nkB12dH4GXNTwy3G3WbvOdoOftDeeTqDqZ9+94v7WxqRgMoh5O
bjpPx4C9wPoDF7BF0+ICBw7q9Ekfjmp0Fhu8b7g7M0pf3ABoNGHOczRQ5T+J2Ye2
B1+XMrlNGQ9OdBuwQ9TtYSR5qy5wGxcsFWgZHODmPCb55GykboPjnwlOk+6UOKJA
YpwR9SDthbklDbYo/OxNwcOFPfKaP2hQ4SlvCbL5UuG6Wyeek0sEpfe1t3NukTO1
G5F6Fn85iE7Med1LUBICAM4PCj4THRgxoNQtk+4VP+y+wh+3j2nOIjMy0+rNcSi1
dsAOVhwISD+aukxvZFmE/FF9vho7yBG8cwtnlY5vccTmy4dg0pSADRVHr/fDcZit
SZctWFDZjXbiBRVgE4uaDkMYuj/XOZ+9SFLvnWYmwtBH1ZVwwHSw/iclxNqrv6vS
Z9DIS1Eqoad5WnWAjNErf2dmLdL86fTokioVSMoYQS2geJJsnEvfOhqL169V2m/L
xZCYFPJmP7yiI5abcWOyjcydm729tht7r8ppLSGoyp9x9KP8qiGw13syXuP/mn0F
aVLoLtvcnd45YyCsC3wmFjW3zh+3E/59vJmWfmEGKS0/nViWiZZne4Sq+4E8cJDu
aUHgeKScCDuFZl6G1dWRI5CphwrLhFC0sZ4RDaTS+z7yCRVO7nMdmPljmvmQVrRv
INKg0cVLJ0gNyhtsReMb+/aPnmCiCHL4FQwBTAkaQc6EmlweZmdR5JvZIgHmWjO6
ayuL8TvedCOLMU4RvYw5dqnhEC1pfE8lhxqZgfsqvsV8oQrjZYW3yiHsmrVhucGD
20STHATPafcbtpsxhl5tdQlRBkNR9LTeVskh1mnq+RThSb6B6rVO9LmsliwHZtOC
d1v/62kQi7knezw3MpRVT4RS2x8IpU2rpr+JQpcTgtGqazC/kp9J4EyelrQRYXAu
2MVMSJiPKFPFLSJq8bK7yjk6BtrNzCGvqCjKgufrKpc2xtkdfyZy+53g51PIBl0B
NAgDw+gPhhBgscMhvkb9BkhMnmhhoD+M+UJSjfTDb1rRBxDLkpS6Kb45yzYzal3/
VPUNbjz8N5fokxwzSgGAjeGunmdxKY5VjZXgh1LQr4U5SwyM4isfcAWKDon33deV
/wWkhzZDwCFS35IvFFz8G1T6SztBy2c8GNmI9sHigtbU1TFISC1vUG5vC9PFCYJ9
rF59Hp2RG6QNRhV2IYsBZI6vaH/Z74iPjyp10Ak0qMWbaicgzTi2S0WDkjKbCw87
hpX30yhrpGCjdBR9/qvdLWlrEipcfuRCP1wbFVX1cEsMSjbzvCywUQq/fHS4hDRt
84lADswSiC+PLmSvjm1ZZ3JCaicXbx03pZlf6QrUAhUPpXQk2og7xd+jmnvW6tqI
wlv+Umf25rPv5Mdk3ZiOZgxjUEhq5SlBUQ9wmOmtLpM53pOWQfv7wgO9+CmFJS3V
6yUnvxsGn+CDlSOC6snFlrkFc6FPRFbf6SG7oQztDh9Nf1lQAv/XhvKSBt8L3Irz
LobsEAdlY1BG6MltMeyWEzmryzjPzx/z6ihHvMpjsqGpLI577Jrsni/paduOPcBo
GwePv4MlD8X8V+kEb0XEyS2W4ophjUAQl/eEaObGLCnXOSseRgvE7ykeG0dcTiYU
8T9/kmqLUpMUvhOdKzSZ9IdE+DMd0J8o6AhnNEZmfPi6SU3etodvLsvTKBoAPzZD
aVitF8ptYnQ0TuJJd6t+JzAXshcs7EsMkheqDS0fEBj9laVDIXLbzNpo8zLoML2D
zjlpdec0iImICoh1OqzdUnLYQDMO96xGbiA9xekG2kU/V99RKOaWxCkj4ZIeVRlV
uumKs7t4F+0ecbu+2LtAJVVHb8ZlTyfa2vuUcuyzGVGzNeoHgxpFHBuvey6RnoiB
kjsmkQCxWr3fGhbqXRV9m9oopIdBdWe6ClmF48bsFB9oYuysOskxzzSM1lwLgmTm
/U4XgU3g0p1PIJ8nQdjyF1spRAwYbV7POq4FVUGOGSGJhtqte5tWYA1fAGOuMXGO
oDArdsgMh6GezoxXffJobAuWXAS8Z0z2LEMB3GpIjrHgEh2lbwQ0auHy8qpIgnL1
SB9s/pQarCA8HU8Rd6KoMRW9hchvDw4Rk60A5sCv22YvLiN3M+BGSbk/X4viAkVX
70n1TbFhL+EtzMgjfKYJz17FXLCFW8ag2dLwug3Rp2Pv0Unvb3J4K16Ul7jk8VXu
Qvz8WAqONgP32MoqW8Ml9/iYkN1qbH7kQeYKWPDEjqS3EMie5cfFG9HgexobKS2q
luuKjnTc/jlQya0VU2k4RW5frwzGElL5svgLRYgN7ftXpWOGjoCWUOhXXbzTHBRZ
3j/pusqX9Px81Weecy3DGKp4/95mOFoTz//RKL51mrCnmyEGV8NPljHBF1YAzWcq
kyWvQXyxRQFQtErZl8YrY/iyFblRvc5FhPbsBfabvhdwQDhkVvwzwyMg0h+4K0YN
Q0u4P/Zq6r+lg7XjT30LW0sXbvEw0LEw3Hj/GyPghKp60i3OhjW0Ra8rq4qhaEud
wvqkLXtjHfwPOlvB/w4v+os1lVH8KUOfBd9SA6f2Gj335j+u4OKfdKa7/D6ohPdf
WIT8uX2GCww9Q+3KZxyPM3Y7k9wQ/QRzjfwCzF3zlerphdtBdECvep4snlAhl/nC
v1hz5qRmekXxJFE5Y2W0duKRn+oFIsgS7qMes89KpflX3pK7Z+fjm3zJIZMFjF1G
LkR0v2NeoZQYpQ80VwHZiSjBiBdQdi01+0YOt9eKxU5inacUePZ87w8FvZFBDaSz
nnSC2r7hWHDs/kq8z2aLtWcZznfc3CnBGPMwLcuXc2ziSJPVZKurTf8N7J8WxKIW
pt3+Gw+p2455TyK4Hdu7iWn/PCv/fnlgIc/VXA+AHQFqZ0id97ELKIYPzeTurjk7
bq+vKVhl5zJyIG1qohuz+Ws4zbth9iSMvIcoNdnZ3eOJwDDsTySUyLZnGwqP7/iI
9BYZZYpbnVtKmz2qpIKrcmSv27SfbzbPS4TemomL3tTDcRRQMB9h9aJ6z1wVwCQx
7fWsjy3J0AKIsYetYUeAhiOirmVIXj7th8Xx2RAiA7ALENH2LN82h+xKb9eZwVC6
fYhULUeud/jWlgomYpE2HbTNIX3br2/GXrHgD9YfDdewi6ItOrMlmZ5d1kvy5KaM
SeYm4yc4V7/y+B76IUckz84Ik/X47VLzDfESX8icYjgC3td9X9NOD3qi/rA5pit9
aWmoi6+xARaDNRcvZ3L0yGdHNdhfI/W1bMRKdosctyB1t4DIVXiC9uxf0fIGhtos
7QNM75r7wzVBKnhQ8HaGq7Gjl1ez7CvBtT6HSaZTTq0fGXNPUZBIbJRY2x3UdlVm
X2u1iqm5p32O/XFmQypxFzw9msC69XEHXmWpACtLV2Px5XUm3RlFKaMIj5q09tmY
aKqHcM6rtyXony/pgGvR5HdYOIGOrLrgTRCFb7lLSAljibxh5oCCbC//HZ4uoQWJ
Sx4Hn7fby33uVjr3QoVBt9uJHSI+SQU2aNBCPZD+A97T+4UC3TQ13ScDjAx4dCHs
uZp3rmWw34CYcRUFzZdIuc+QM5JQI9h3f2pGMEl6VbJftaP8sXceVx1JFR3QmR16
6EcUmcWnnyXH4poaLQxMPjyziSMF7oSsoYj02yNa5o61WUh0dDGgZgHZOa4guYD0
+7pYguuppZmhAa+FMtfW7TIgITH0/tCENX/Yf4RaDQY2gXh1WYLuIrSysD4wFvu0
L7BtuGNCu6pyBlbg4NK5r+bSlZj5ULqgqKlFNhZVsLPBNxIKbXnNNiR9d+O5GPdQ
1bn42JzPY6xToE9zRbeNUvLFExk4iIYd3ApOhTe/4g8sHk7q/9vETVUKSwzcXH3l
6E21HmU1YTjxaQHwntd/BzSc6bBt1/E6HJ4pZx2mDGJzLhqHKADybYPNHD/yqXDH
DrNJaLaPbR6G1c0cLuL6fAmtMPlPxq06asciR4aJQC94GThu+gzSBMSBhfVzM1Bq
ltGOqo1rn7Q0wrPca5AD84fGLWa5CtOEFODIrS1ZZ6fBKx1wbDDaXPrhghM9aeej
qR9MS6rZm/0bOMbzOwecDEWyeIcdRVPdM3SsDGwD8gFD9tId6S1ayBxJxdHxYZOe
CWQy2dP07zdkOdkdI+GiSnGc4xOwPmU4N+OG/BWO/eK4C31cg7dQ8Yvbz80FGls6
ITF+F2JFevVjt//FjMx7Kf+CO8Q9mlyH9mKyyPKane0RTX/7YPot+OPtBjFovWZ0
ejjDcTMCmD8wOFRJA140aqVI6SCFtflTsSyiv6VTrCTwVxK5WN9FvQd6rnjqqNpZ
6bVcm0lKG8qZezP9LZFCEYrxPegB+G6KXvDtp2Q/TjAGJntqoQbR542bc4kjd8Rz
driaIY2SPuxDG+l79w3ZK+gPS3oGJGOcS2GMvTISz002Xj7SSfw26gSduMAZ9IiB
MeN8Ft0rl5faQNc4b0bPmpoE0QGpPGT1u0RZoQT/XjR+AKFUiwuUzcewTz8EI4a9
Wr7ux8QsTG2N9h+ZuEPfrgVgmykSaQv3mIuNxvpqeQY5uDI/ahjZNnyHtu4ZYdep
jHhHRWvwxnpqIYST1TrQhxtIzSRRIsRhI2YyysS4FEXYDZmKCJ1nevHBYKAMs5cu
BjJqyJ8Wuhm32DiotYYIilm5CFeRpyc/742/NkKKuITR/F/ex1BTCGjDyOph9w2M
F+uKrvgK5QtmFxn+/JDHkpqn4+fFt1LzOIKxRGkk2rorQnLt3CmDN6pF2b/CECgA
LhB059OniDE7XD6kqxFpr8C/l14eCfQ1NZBaHiLFWQBtzHl0JulBkpLWd4Ad2gA1
FLTfip7mUOcMnwwtAcasXSsBr9Vqj3x+qM0TInXKi618ewPSXfPxsNsniRTgSbJj
bCFAXeLgnNeMAuSHURNI/yuoThSsObOHK2Pp5x25TawMFmspQ42xbeKyQK0Rau5+
0wCKXTOrSvkm2PtYf/hyjIYLopboSIAtiWycVtwXSEzENJ6iqtiaXkk4Z2ndigbe
2XT+oGzFMYEznLCQ5pjm+vlN6SyGIWlvPipE/X08c8lwTFkmWctvf6LhlIIrVRGd
ts+naLVcl8UFmnvyjGsWlIatZh+YcihBuMF5iNN4ENE7VEPww9oPlX4aipIRtSQF
2cuvOqDPb+gZ9YGw6oqyia+N2T49Mtgj2mBs3k6YFLlPJGYXfLdQ9X3hFIKGFuB0
fZuePvNfnkGemkPg1ZH6bsCdpehS+L932g4TfvATmvkQrF1JPydHP615spxI/Imi
Ob/RVjk27XtsuiFUso/VfVRT0zR7j5JV7enhdXOwWE8+aIyiqRPkctCt3kJkWHHQ
INiewTI5JGW4Lzg9qeADgjihglBtTi9MWy3kjHCyxC12biMfw2/xq6PUol4Htayq
pzeO43Pdb7898Pj1KW3bzh315ZA2oPFWYHJ2yir3Y2t2zfLpNi+hjr8PUlKXqtW+
UlU8Gnqb51Tdun5rhewWmH10xDMQn7uncgx+u4h+UKmla1G+VP6GbenEfC3+wKJY
HOKHtjXEavdYfRDHt0YPps7u15TuDAE1kIyem+tvw9A4gDjZrFj1MWiqNJ79qDp8
MO0l2vbL2gQJsPB3mJzfG3+pXsiKP0Vrik92Ui803rtp5tW0KXRnWnLYsZaAV+Bu
mEECww8q/iYcjTrui2ZrNFWAjIRnj5aWG7G119x13hUTniBQwICHLsBnAljquU00
hKEkfePcwtwV7nPpxgxbkKTCmcRsmILKdnTqwDU5hVPJ7og+MCQYbe8oHhHGrNeT
enZxumRJhbX4r76RF7nGsGymOu8nNDe1hmRAzQQSLQ0ajvQQbjt+aLjDtmwh06gt
hBSOhvIeAxDXSct2OFFMrcoFuBbTs8U+cggcJDFxy9arCOd9trYoaZ1cd9t9WyFG
EZ5Zu4eybi1rlPciUocRCxLRrHBhA6AD26mfZ43lGK2gXjBWybhrgribBcelQfS3
+rIONRM2CE18TRsnrjnpXimvybwRMObFZafJyKIYei4XdleqDrTOiYELPQJqDjQi
Wa3G0h76bMr/F8rApsXGUdv/6NcRU2zJqaIw4GKLfcEOpK16v6lbffdsU6uKGwqD
qFsc3pJUB2Pgrw/PXT+VWFW8RQyTEWCQR2OpvK15CeOJUZu2yZcFqcYI24O2x75h
zb8yFf2cu1uUCB5nQkEyg3kXArhEjOGxq/wsNIJ2EW89rp0wUPvEdzPJm22tMS+e
lTFMVvpacOiO1XVP645uaVh663MCEGCUChJCkDY8EFgI8n1uaRExhyv9+AXimGn/
CTZ3jSawZwUxLZg1Ne+biQR/qJuxW7psEtzsgdO1W1QRLNs2MfeWwW2Vcw4Zvj+s
s42kbOtD0/xcjjEmLapSPsmiTmri0QqAOK6Ykw3/KMnrsayDFfAnz4Di6bAu5jJl
gAq9dZDbmj36WJYL49PJtV6TZGo2OipjbrV/ZS+jsJXezV0fHxW3yThxZgiYAHiw
/vXXcYmyvev+4Ce8P8U+UtoiTc+J7Y6ugBMcMwBV13bfmDyq+6+muhWValzOTb4R
LEVAfM0VU1uFb887YwkUv6HGd2CZscK8sIeLU13/IhjR9di1QXnalfs/4p43Su5K
99GumKtEDZhAg5bx64hmOkv8XMT+wDqcK2r5d7f2PXTNDe7BVxUvlLpglzpiJSo1
l0o8vTtG2jlQqXeSqDM3Zf9rWd7rc5mhIng08jyWUqbsp6dJI3CRfYCmWNeQ6mK8
21Juxz/vZ3FMoOS7Q1yjBrzvkdfZHRPEosStcsE28gV3LTjhqU2X+vwV+pBg73VF
uUwugwtHBOiQDWcL3eSJdypOhplJD7MuGZApLUQWmG8XlZhy6PD9SuxhoGYP+Wmn
CW5IvGAb5MF8Us070qddJ63J+6TF9dkXmDtDLKseQNxYsTFaT5btbCQT2QT52YJm
OTI3D8Nnohu6u8BGOgcqSaDdtjyan3dFPsbSZyplbbMLYLJVwRqtNb0XwmJ/2LOI
svDdxpIcXHbY/CFmIspSpG15YGYv/dslX9RjGirtKe599QU23hFI3+CdMQrBuSJX
vvLaXB2bG0vVQ/NYJ2tyZ6JQCZwtPQUMFJCLRDwVNBmz1jlJNKZiEBhiUUJSqw8Z
Q/NbGBFmO9hzg2BUdfcAjnDljYJXdGe6w0L/gL/Vbm5M2dGi8z6/rODcZSkFFaYr
VECBDiQZGd3dxYTVozOtVkrZb0i4DN1P6lGgATJVYQjZ4+xUwgAesDazzRXbKxsV
hPgbuz3+IVJzqZXgJ3I51PiJt4b7UflN6Rd1YzKc4GGwSK6ciGr9ZWPp5y/ylqWV
nAVpLUFl8nAFvr7xronH5rdJWakPD3AAlWt3q2+cPrhRtqUmjgE0COErprVcYyCE
S+ueyTv1Zg90FVNXCFGwdC5lxvvQ8xFAJciu+mwPf6LYLKhH2aPGtksXP2Wff27w
GuRWrguUEOADt05IIZTGnC7m9jC2SVNL4PF4T0HiWQZnGxh1nKjlg793tnpCLj4L
RMJ71MowtmCxEccITx+YZRujsBMzukX24HASl+YbTpXsoG2AWCJWajUfGx1+6PV7
NNPPhdFjdIBRizE9v9PfJ+CrzwBt4IXEtbGGxir25fzrUrwVwSdctwBJOxJjEisK
SMkB6wigH/N5OBiLFxvdRqVTl05EKwydXGDsaAojdA+X674qYIL3DQaVri9s/7zG
q2cg2qAdbDnTsnUwWVYOq19ByjYfMxb/PBxT0Yg+6HJeAl0iQvXZn0b0Wi9hP9Kg
tvNNZf4C4vIDfItV3Cp9qRMyUxeB/MCvd4DcVvzZxa9soOZHgWkVF0/Wq4taoSjS
9CHpKgKhx9bJn8C+uC/UX6mHUqarJul5q6YbifV44Mz2NWfDld7r6TTp8AjFRiqd
7/QHXrxcoKSH72lElO6O098Ds/DiHjQ5IpUeBvgQpckFYnYS/YTnbkruGdL/dJqs
k+2fHOfOH9zRuR/r0LCCiFxghmjwVuo/lIKx2pWRtoFs1Eb437whUI3oKhE2y8DM
o2eCjjm6WvGkmD37uVj1J66O+PCVbf/FEzmXIWgrTK7j5U7vGBDB5JSrYRlbygWn
bKJxfow3Zl7S2NGjHEYdH+aVzBbE+HJcu4nhzBRiX9hQsxNDby0le4QD+QJ5ZeoG
BoKk4VmQmMSrGq1cqUcCsrY0VrVkBZ7/HWfuLayUi4Jp9pE8srrtJOGSH+49x0FA
fn1wGrR1FBbdWehI3tlz7iSnbgjsfv4sQexVvDBaHmKbww4VfJpex8MwN1F0l1de
ZQb8vRzyC/Ct/vI/Q7xdwGYpmT7tBY5DnPdpmcj9/ZxQDUq7IfHaDyFfwGDIeKtk
egyJnxRvBFwmRbN6UvTlaHbk55/ZivVC9VSA2EDjFpgMHq3/UtNuVgFr43SQpFD5
0j0XfJl2SzVGNPCzxWRHMQIiA3O4Is5fqNfihqCMFDjv40QNtCL25hALV9x4waVu
kEbWCaD0ZSivPh6lt2pQxf6qvLL4oF+/d0d0Luez6ikLYip0N444s0syvGLzyo3Z
ehR3v9uVi4AYXQ2/F0RJY89QRSlEyCS9jTfsN4V9/mZQGsAqgcWubj2M8SRp9W26
meYXMqJaL1LLwXKlLGMHs/zsIN4+Pu6zRBV088+AleFW/gJwnONfExmVq0YoOeLE
kBowSr9i3VhpcOvqYLtdqo55vBoOK7g1kodgqIwF6nTBoV4SR6EcAYcpBi+0Td7N
UjF9G1/EoCLrxML8uRkqwhY75lbtGsHHOWbSMXQ4AXT2pfF6j4AXv9/IxzaXhgP5
nFIWeTTS/+eDiSOq3AJIjFPqDyULekmmgeEp7VYXEhPJrWrRb94BtuheCQtV9qf7
l/qjO3demSoF8XNbBl98/DOe/3AicaIEZvLEdy3xilKQTsp7y4kQo6ffk3rEhzj6
7wPDfE72xJG3ku28xofSkz+/OuQrlp+vPoXoMq1th+G9gmmCMb37Jqc9DVopzXDE
0N3jmecUOAUK4LUHVJybiBruC1DQ5ZD+be5m4v09MMiKrpJGIhxOpHa0KpuPKVVf
UwDyKnX+KfmjAFeS6FEl09/hSRxVPAiJYoO8XEjBoh6zJRWxFYfp7xK8kU6CsS+T
L+bD8YWbt8mQ5OS3bfL5ExqHk6nnJQFLq1DuMQaq4VQSCaXrUwiAlnT9yb4LCxDj
l4NEW4UQGZIyRnziowzWqSPgn5svnUMRaFOYUtN5CiEn760PGc4gWcL2WxMxNXNq
Ura36QxtrUfcphl8zTVqMkKNP8KGXY/r3Mg9KciP3XnvCKnaDME/ux9tPnOBoYA6
1zjK14Dvv0EKi1gtFdTOIJEAupolALOsqYQhFvIIz8amdXlyodQ1FCUD6K8evPwf
VyMyGxBLLG1qobnUNqcMrmi9BpoZaWz8UK811L5HUWxY75vNIYX87fR++zlCBcYP
eJQJs6tsDYAKzOHIOZXe/vo44x0bN/0T9TxX8Na7w2OHrALrMajlAkALeOW0vkdm
GrVfFjFlgpN737MFRSk4sPqmEI7npKzKO8eAjlKtQ1vZ7KqB+76Nvn9XCye5Bvn1
ljaLG25vVJurNsQ2LbvjDh+dBhkns4wMouKNNx45Iwj1ZIFTc4veCnLtDamb48m1
mn9kvEI/jm7uCcTtGSunrF/Ys3tgR/y8qxS7/wXCENQS9D3XZA1YFpZeRWfptGJC
dtcrdPaXAsTOqpygBbXinZsBtAu76JKqixJmPLupMeRXrtTz83awzCvd0S4X5h86
Med/V1g2oILreb6+rdnphfHIobVVAZHn/QdQgsSaxryyLNUfcxQL326X3PdAqq1e
Y4pIlOYzG56KJHydlFHwzkowRvIbOgpLb50xeGEOdg/uuoDtG/i3D/WfH1/JlrbY
VS2tHH6wGZNCB8KjyNKUX/gGWYGAXnUkrU0SpIk/eR+mT9sIbCcu1yJaR4gtrG1y
9y/O8qbU8tuZmonH6vwfrp2N7L2a1WWG7v7ylQC6OSyWNt5uNjd2USKRRfqAlH6F
el2/lg3L1HBws3g+cEl6dnqCQdrYNPyNK+ai+Bs6dsnS9j8NwqABM5JHCepIcSqi
ilILofeEtpRN/qmLnG1OuU7bSevuYk2r48PpiE0/bq5j5G8r76I5THjKFbcE9OQY
28Hy6LScyJgB0YJ5tT5fUWje4lXHS+mc6PaQ/8s9KlqQAjdpoaK1E3QwWmOzjb83
zTXNeiCbLKILMQhuwgH3vx6prHoiRay+Y/cGtqsByv7NdMmoEfQfVGi45FoIvOtZ
vFMwnLeASpqSof2U3uGAudI30cYDg0zUNFYL09kG6lIkoZ1uvXCq/b9dg3wUUgBt
ZpKSTf51GiiBvHpvIsds0K54xXXPP+5WDae2lRP95HNB1iwYv5qiJvMLHT3SZq7f
iVFP7Y/TmciCEvdEwZiprspWxfIty1GM5g/aGpZvNPPbERrUatmyoRYHiIbmeS3g
3G+19nsmymjT5shqfPRJ42XthuXwLSHJDRK/cSAsOXmLJhgu8M5yWjMBiaqGtPbg
Q4IKfiUEHF7ZYzqgFnpNaE69f3JhBnePt4MTJZafgspq2hVY6W/WtfhqPMHijopS
ORuJmZilV4X3Wy6RID+K7lSSuZ2nscHd5a9piOwckOMI6HKv3IZBRCB6PH0izTOg
cEBiNETBtRTG0syHpw/tRVga3AwGHrNM27NyxUqUYoiTeeaWLikanNupXlWU83hA
ppBDRzjZEZdE9TRpGQBu3lHi+DgG33cO0z8oyea/I2Q/lPYl8Ba0Wv+9Pxqr7zcJ
AQGKwnEC//MxxkeGkoSFekhAzVyo6gbtJq0EZHEGGv+mT2FW/2lyGlld5g6A17S4
SbNqqAn+E4Q7uZkjG0Z59j35XSVX89BrNNzITDtcYjg7xawjwb6YvHBtSpX4GmEL
m90hj7bnutFm7hQdtoaG25iTgjJYxSxnIoBefNOV1fpIdrReZTFi+2Mb34nl02+1
DoSZIHyfzLkybGBzoQr7saCrglQuoLvgk6OO/vCdGWawhh6sQoPaiDXP0ngyE6fa
qMgEW4P3MZg3z7VhTQ8HZQxYfnaMAvIuj7APWXj3VAnrkT056VSp8yzD+FUATWF3
Qb4hAD58/jEHBlhR2s9FeKLRHUdVd6ga0O2+IV9aEPcq6Ehcha17FgpIHXwD5puQ
s4Bn8p2uOtrGOAw/3WCYpuMCrijSzPCFTQQuLP013yz49ZEsY5oQh6VmJhX9pN17
uFGa+HaLdKigUf40vsdQueB1EIbW2V88X2s0nNbEKJSbXLXKFpvxQDTV+YLz7HTR
cHrq+ZKI/LlFNMRx9nIWUS2ur28a6eW0kgKVLsu6Ey/gIONlNHA+ojyDIpOkVCS2
Fo7KdNfqMOyLUCz5/XOxaz1uAIsobxXayAjo6qLScID90sK11CdYPp5zmgtua3ps
njuff3CSW/9g5nF5ZuiQHlZGFdUTxwQYTeeUm6L9RuSOuuFBtPS68Sf0ugyVr5Nw
IW7klCZwWdHyeBFLBZZXbqgbzgXwTWwC2Be/dvWccAh9wYYj+B/X1T7gUaCk7Qnf
iSTFmLtrcKV6c3W4e5Z2CkIj/2gJlgZOXIedAcHJGwFpoNSpE7Igt3aHA1ciLQyp
3BnYo4KCL+63GUpeUIn4RLSSxBP53+tspwHMOhzgKHQo2T3yr3BE7tQk7sQLLWiy
izH4mwpSsyLpx80NUuu5XwurlLi4UxZseGN+wMDDfAWT6nxU8gPF6RJodmRjbdx4
QBN5px/ByHd1q6t2ydv9/hrww8grgfmnGT9NvY/3RsHPWxQscLJExMdKeO8rVLRf
YClEVtAWjOJ4My5f0OjpksC7V4nD+jZizIyJmQOZHtHP0n0g32HBrcGLTFyT46dZ
p1W6ZFe3QgzA/zhvzfx0rlcd5gl7KwbEhywOkzi+SGZYE39AyFazVq9fchakSK7/
J/W6zO4eISDO0ayGLEVbQeubxUHwDV5RiZqMHqWDXYBHuE6LiaGuF1DVd0R55f6Z
yuwIFwUbwqC99mFNELvVbu8S2rJF76HOBAKUZJ4hKlEOchM5J56NS45wrN2mzRz4
6x6m1lpzVf3uwzSQVrQOX3lrJZ4eQ4HB3Rx/zzLMX00eQ4rC42RhVVHGtNtHy1eH
o0Mk/vLLQ+v2kEUbn0bdVYx3MwGuaNB2XU42bCnRCfW2qmKyoVduh6yrzaiqkibZ
t1A96VG1I2mCFd11SQliv7b9oPpnutfbAwYoNbjzym6NeGUc0gjedoioWppZzy0Z
5q4Y3d4bRSFN1v8PYXeZzQk6ZbjMlfdz1kh0fnB/3cZM2g5j5b543tmURJ5Jov66
uVrQBP3IOpnJuFpsrFKnmC9OtZNjwPN3qPm9wJEP73SfQkBrmr7Ex3QZf7vSnfvr
TNbs+CJcUY/jbSaJQSuWH8dRU1uRtrSgmD4OYOmOJUcepdbG59QT54prziuUbmaq
YAa1aJfYkJlutkRDlow1/zXgSqLRPi514kf0ms3LXCrgzaepOmWBlRNq0YYcRU3c
DK9ErS5dl/vRwz9oSKnhGX3DefCRIETOBFqOL8J0Cvi1X1W97sygS3Q6mCe/L1Pm
OHeh01RqmvteD2lX4oVCryvQ7TBkC11PmGmdLG9E5qs/hGu4y5P67xBlcx1bjX4G
39dTyR1NcxTGCIYQlsMVdO65uJZIv5wE2bP+gEgipEOkPHGDpo2rPWSNduF/xYxL
y88BwpIsY0c74TV+IirVc+nT1G8r6mpnxdm4c4QXEBL0oKUay1/DgVkwskn8es7G
KF5Ib+wl5QeTsP+Y9rluCz/2TiJKP5YQs1ISi6oPYmeAhQJar5CKPIf4vtsIrGoC
PXpcDSLzrlIuL+t3O57c3HRgWfz2vVRYTaSHteGUJfPxq5IQPn2s0fEScwgmDIWC
fBWFSBbRUHs0B17Rw5/SjZ/2hSxG+uyQHTniaf8Ix6suSZbQ7eKLJDQTkn4ubdEK
tUmn/s2wlfZ7QSf5CayI2zPwrazb/bwpIdTTwWkRP1irrHs992hFgwcoOLFzTsTb
Pkfq/6n3OdlpYghacPhWRMfjVMWAugEiiyQbTdGkDSgJqcQB+k6qQhb6bA0x7x4L
aKkBAviqtCsbyv4vESTbrf5pM1Br7o8CjLhvK+O6lPHzuP+TJfxkOt7QSUQvABuz
NJSUigC4AItiaWqmAmPwcwxrEvRUHQgYNPZD9nRT5dYgf/vncsPQLBgeHJe04zpu
W/gSEzyQ5AZt/4X71pt7and0CmXGDyNRZ3NPlOK2Fb3bN/bIRf5+qvSfjsbD17Xp
SLjhAU5ViMz9zA3IHeq3QTihTQ+FOk4CjuThzZycIrb9tbPXx3N6v7gQVtoIe1ce
xU7UscAWRNPK/YM+W+OOfyuEe2zsbnTm32oMzl65Sbsz7vCzFDVIizwTJHloM95z
HOWSXGjmcM3VKxF6XhTafAgXDbjx3mkjoBkrdBz16bFP5yck6GNrQ8NGns1VjKBu
QzM1CKV0QggIOlu/Skrzs3gWYYyWncVv/pQ7VUE14peceZvpIsijuccnWcrAViDM
vbR1i+ggjn4++WKz/Lgp+jSpvgAwO/A3/8cYT4eSrin3JKIY/XcSCLe1RB4LGhfZ
TqE24Ar49PQ3zOkGIIwl9g+U/DMOs/7vAC55+xnk67//eMvqMdYdDheLS03s/+mZ
QeqlLI1hQ3rMpBoqEzeK0DP8wgpX3SoQFU2fOlgCJo3KwRG+90kFnGnQEsbDzze2
EJwLSuHmEcFkeV2SKEUUNKa+8N8E+lyFxmfDbApuIcv0aLrTh1k1rMfLXVNHYLGV
WEGUQBiSykNC0Mmb26C3H+Ib2dwS3xfjvD2CsY4Loqz5o5oNZMJ4l5dWH/0aHVpO
zY8OlXR/RIQzcveAU2AnLbt8yQ2iw61DjluXOCrzL7s4tiLmcyysK0jQr80+Kyel
DONy8AboBtzJP9beOIQTlKTkNhBs8S+qlzg3PNSucnIe3/2l7fmQ6yOWfMv0WAEU
MKSnGB29IJuJKxtOFfkR7djs8weO9hl5pdcu6byQLy6vrhDNovrJBYYtFACpor9p
3V7EyUXNOAj3GlGsecHUAaMArgfJHnboKOx2+XSGy2K1S+gPUrrM06L/mfgg5cyL
1myTfIdYdvv17bCmdi4UYLh+rUxTAjwzmd1iFxXpgSvNwTZazmvxdeyr6dFjJ7XF
9FY6IfHP5+AkXP9B01oxgBcrtG9zTa4yuXuJEnIAe9IPgnAzhb2c+QV10WbYoo4O
chLAjpdGad8OXNlmxMJCVvGpVyJi3jhZxxvgBzOdN+cS1/MdxJHoQvpBSp49uI10
9281pCHGWERCMcGDThuME6e0WhmcLMri8dPTXoM99kfePa37SkhLRDIeEEQlER6X
TR8vlAmrceUk2CzWyLeDOIuQLsrDa3phuDjbSwlXEv2XGBHP67gPBEtVzUjE3uaj
JjUL15JeZAZ6SCjWj9vXvCX2tHKjHQuVBTiNVgMj4trzKxdPjfS2nN2hzKNvCL6e
o2yt+lA4JNp38SgBdplo7iAYpqwQk5x6Nq0LrHlZOq7Eg6dAOILASCEjXna7cBCS
+K9bW0SAP58wdWFx7tyj2CfiQYpJUrPN73pnRhhBEFe0/z3G95w7jZQ23NCiykg7
KdW2KOOmIoQ8ocL96/eA8euvvdhCiNj/p0/1rrcnJe4A1cvVIhxbGyiV2E+0ehtP
ih/WjoeCAUrJJqP9M2YkruBHk2xSr44INFEaubGXB7mOWXM4wjNDw+gP+Z44il9w
zGidM8YEX2eoySxq+BY9+29dK5fP51SdLYIyBBbr6nVA3Cu8KquoseSlGqLhGtXw
foccFsImzKkX2UR6Ur02YNzonwEGBCjFes/D4rqmOBncr0FGmWFzczgdnWVj5Op9
Qq5ijSLWfXDut22RApiwUYe/hQtTUzGX7MAsYJ/bCM74gIKA3ir9xGMYp2Xg5tN5
nKVCoLP/lXIRmYjWMe9U4MiJxP8lJZEp2/WrOlZ0Hkvhnfwia/t2fgoaFDaTMXF5
ndmKdOLN4tdOlHriPhTbnUsBOiSLCx7uHKOuiYuFjUma3MqkHYyFxPsqlgibnoxX
CU3E940cTLdLVkzQ+79yNcAb0oS9Zsc2tSrz9tUHEl23K5Q7s5rUo3bwj1v1zxSx
HQf9BMYW+gzOio8UhdhQxNOnTHHLbvWgOikZukt/DPcfPDJYlmBXK04oVWZi9mWC
RPPZkXJAm5uKkMx4fPZjyqT8jEOvUzsROJ7FBWNqHRkKqB/iNd1DAL/P5p0qlOFd
nHYwE0YbJzqiOXisytsLudcOEcoZrm+w3A2gfaLg1O0CAjiplmh00o+hYVS5uFEd
S3wGYFU6udN2uRV3zAHiYVA5IPBkU8/YqYtFHHmjVw7/g1QS7+eXSHJicY0o9anE
wznN3q4KIrYzY7h+NZcTNMvKnJ1XuBA8QiIZonJxMS+ovP9arRiGHnJqq+E/XT7j
85449HRpFY5bPcVNlACYj2KWSktMdfybnVg11iyOa7j0MKFAVBsOJf71Tr3aExZC
5Osx2iJgEIB3aG8kELS/iuh/+1o84rVtPJROoznhbREe0xEqyhWeBb+ras60GCbK
zzLZk1nEpYClLFg1W4ov9EwRbxc1iD8pQQeDl0X4hgDN/8+M3ttsgU2tNb8PM/Bj
BzTCswNO/GLLXtS6MViJuE40HKI9YV03knfGu2NT5+J8BG+LaeoFwQBvPiC7u2Im
EfsXD+EoI6y2gXGhRprTKgSPQX2jeXDkRmAlM8+w1NFXr532AtofazmpxPH7Mrqd
MeV9FFislCOIp4n52/YB091+P2guI+J43nH6O/BNmWIlBTfCYRWIwutaqh/Pl27V
Q616HLZYVfE9hNQy5w5HL8s1suQek8Mvs26OW9TY8O5WSZfdyqNLF1gOcIfpfi3v
raxZvKZzYQVr65m+3xz2iQWXxsG9IJpNxmBkBFrkMJpL3M5JDlxce+ZLrFaXvsnb
bnhW2XKyHS4EBevNv532acvsQQw9aXTUfPHmTUYeqArBn92KUuaV3QKjUsezVyxy
6GBdGP00S+vDEmiii9UD2oe6YeoTwz0aLxBM5y4+U+Q5i504QTvl4NN8mFGL/mQu
27unG3doeM7WppEvUY0dBjW+W/IAiwYotYWnYoE+bLHSlqhH93mNuoGZP0+4oSLW
e8NdKbKE4v2bJX7JLuqRplodwXzAYlTKTWhbvPZmLleBp3i9Ws/aSsPDungyYqqL
nlsGQQwKrMYEaXRq+PVKbfwjzgEWgxsSio9KRw4KhudcJTdg4KpgJ8wm+2op5Ve1
JvTT9vunftJPAmqzLLWyF1QgeGBHo30TvRjBTBE/o9Zft1WTAPQy0dqkF0lj059v
tKuLaHohPOykq+zCClXmMGJLLJPt4HJxOzmsQ7ZWKnY+cPqUoxcqhY7+blyDkUMB
Htl/xBi09Rb4nTkW4KetOaqG3jQMd91dgh81apbXz6JJNVbaxJSd1RELKz5TmyT+
0G095E3ggO8UpD9kvsqLux2SMHIIvpJHHqtiXZFo6KK5TstGQFbjja3q5XwAluUS
VpTu5SvQsV/P2xdWX5MuH1lyJ0QXJuJH1kzUmjiEt34AwzfTCMn8aPaaS4rH5d0K
8EGtuxi7mbZQCOtvclbqOMAwRIM2gvuodQ//xBmv2Dptt6i4ycNDr+s/ECnIQofV
cHU5d+ub3kk/rzcnhJ2dXf8NqL88tU0YgiDy86TVtJdjamg/8JiFMhwQUj0QSWup
biV3M7ZLUky2DcWgTYwvh92j2qrLum24abmWg52d6baCCojQjTSAeD2SHGoVNyOD
OcgGajExU0K8sHR0k6AdJSoX9NcFPhnoWg2FLnNhaTK4jLqrQUXsp0mKqo7Q1fvw
Zop2x6saxAli89EMLTP7aH8FMHNTMevVJvA1B9nsI9iiYPIVS0LkvhSuj1LMitV7
tM/8wHfZGsxh/HS86ydX5VfSzEHwxEMaBnfVKq0Q7pryxyJKo67IFrHvJJGpwKCX
Zn7IKV//TSMBrJBqcWjK6gW8SoGO28cD+aYz625D996HMTXD9AVTg7R0bFZh5zgi
162YonEIl5r3eDzEv6kTt+PAvl0aCm0Wq/8uBu3e+i22hxq/KhtjuSJ2VNyV+FZG
qaY6Gj9K8ChuNw3U6XC+fgMvYnDOAOKmsrsHKUXQum5hw1+j5xVUfFqBipdz8Y0M
6JVq2XIiROP1wro/VsthciQIkN554vOzzukIkihiVVxO/6BQVwWGmad+Rty6WNQH
yMKNEf9bERn1KPntJW/H4AkYdxlad7PMdPzzBttQ0wTUN85TrYi7wPKyrJEQl8nJ
4MNR7454r62yJV99+7+tYMVVK2hd8JJFd5WkZOeWRRpgv6VK8pv0SxuBNNOVuww4
Ac6fGsVfQe+CGgkwQmVR0PRvim7I8pM11xzK9Xx0PPfAmBmQ3eHhDCkxj5yygdhb
5E1JRwXLiDqwYb+SSH1vYYOQF02HLk5d34e9ssIACTbLhsPQs4Oa3910DJiOdmwx
DcFVVGwWDj1dHPr3njFuWMI02Si5t3XxzpGKAPexbX1nEP4THmJ/rk0rpMMeAAZ3
Fgomtum8geyAZ5qtvhHYytvLUp4m8gwjZGa3r6TbRmxOspg2rGXeS6Z6Lhaqy7Th
IjA2Rg6SZjh0aqQTYe6IJ52WBeTjp6zzVdqEOr+QqTa48Lbjd/AYL0ap6nfQ7Ixt
TBdCTUrdjSj1IxRbv1hVXlHCPuvhnTCKnMZmJxkSJXSx6qz9uA4uvc2hnSvs2INi
NFfCrOtcV3M9oaFsu//7y3roTLG6G2FnIBA7lxp2KHTYaOwGyWsEMkXfkVpQZ5jF
KKixNYkp1dfRF4ZzIeTqoyAZHIxB6DwgIjZ6B9ZpUSpZTYntd3MvHlAIA0oZ9OBN
gJN+0aC6a9WLn9dSWfrf3h9Yg2UlqEqTLTlP/A/h5hGD2qg6ZRdnW4o7Kk/JFtzD
/TKJenAXPBgMAgAQkUDfwrzPqhIdo5acBvnDCofb5urL4Ayh2/3swsqkXcvokDxv
6NJGyBmrtJNO0vJwNHg3tTfYQD4qRYMG1szz+mSQD0EIbPIjXtDkxsN6R459rpiL
Phrp+NMpNu5/CVPLlxjrZbMMuiw3jEpxPMhlR/M9fEMM2xchParbA0ppGChVUIg3
zMBptGs7G3jweUgIJvWNmGt3vVFXKITPRrfvmTayEtSTwZ4xvK7zVPlrmF2ag6am
W/5PM0mUEq2S7hg1H/liF3hNp3D19tyWcZ+0Q8P7ONobAXc5kx4V8J2jV4A4dhIs
xwoCBz6DVzEMa5fV7yyrcFAFwa1CofJtVUnsAv4Y1yYlOMROqzhfpdNwWN95s4Sr
sm2Fjy0fZxz/WMxQicOOhkl56wF6DTFEMTwqGctYvwUsCUK2kRfg+t8lheQ4cFND
k021HQUhWca9t5Hk1H9NYjxwpDYkJ9oh3zTclBuV0tHwcCkiiESArg07g1vAhD1L
GEXo3afE86wL8KgYNNg14yzRUyP9zrbV8u+LzEIrHeBJo6X94p6qAoDUARMTN9au
gTHbO0S5wWvLcWieDHamudad+seb4gHsVFF/CmmYZ/DOZMVcc2dxGunvoxTyy0NI
21z8B7Oa11NiuamuWoG5nULqzNE76ddRMtCR0xMQDPRJGWAl3dXPYcBYFDWACMK8
AUguDO08S0VJ2+dDjUcIVQi0PYWUJrFQXvFz11J/d/KliprtqBUBlfnZqfsWF4xd
KgjI+v8qa8gxcEvz1m/2FRJ4nDqgbTIjsz0C6oU7l7p2yGFbtzDTr5gOUeC853iW
2jYMiY4JlwWeKdkFEpxr29BPEHM9rnG9CSilNH5ztQ8pQbJg6nmr6bosP51xG0ak
4mYIqslNDzdNNzUP+bnwHaQzxLbaUpvWj7iaSxs/erX6S8KCuxHx84NbNhu+UKA0
A7b1dv9DVHa5H9JVgzP3mf1mh5TsH8qiitVvyFIHd0E4Rt8jW2It8fbD5IU560OM
QuUOdOZXgWEzr5R0Q9NeXow11N+69pQbw5qF4IDyCrw/3/qGOBaECA84FpM7xy6x
NyhCX0/OLqiUYDuukQOa0Tj6fWmOFWtv+tXn6ggIC3ZInOuiCbcovA+7zqv0iF0a
WEtc8QnDa3G9w04001tRTlR/9OCqxLtv1FJAZRQ5sI2ybp3zr6fa6b2ZAHEKxpyv
IYmRmvpTWGFXE2WKtnA/3daEtCfFWsVsAM4yYh48N5F9UpwkaIn2vmXl0OIb0RWU
mBAlHwCoWFClUsbigsAyTB1NZSSQj5crGvFVrWt0s2ujxahR1nR+/khw0arp8UeC
ZucGL+8sWOTqz+FA4MwRR2urJylkdraknQMiDd36N+ldP4KxXfdcIRiUU26gv7NY
kgAi7WSollOm//OCHa504yE/+KY1ka7LFku4Glss50CNCrd1Daqi7MSF0AfhQ+/o
1KrNIbHZ1rWj0sc9viUQTU2WlQDz4r1j2jEdphSHzHTnMWcvSLSZr/AicSJgIblv
fVtYuGeiUFw+80XR6mjfXsqVnx/gAcV/+A9u0iYKLXlTvo/IOYVCOaTCHXWY+vX1
NMZzOdx7Mdtv+QLMyIppzgV4k4z8+bCM3QVkNoPoS2jt2gyu7fDRNmHxdfnv/z1s
VDC73ZxnFaP0Xjob2UwCIffAhw5ft04D9soCdDIharXRHY0ZNr9THiqYDM7AblwV
mRa6nxFO1jOavGsCYeOvNhTQB+lOXxp67OkrVexwqX2/X6QbVwMloVq9UMiWkdJo
OOYTkrToBkH94hiHploZsMHwVMnXDutgL088sz8r24t1JqFt7AUOHUOPYYZHz2WJ
bBdAPipY/tLVWDWFZtMhGU91F9+md2f8NJnorOAri25Bc1ggTS/O4NnrZaOl9KlQ
3Fs9r4FDSHCMMI+OkpZOvjhUZCGZCP7KAUZChD4ZPOGjYMn1cSoaKbUJNXh3AEzt
wXxa373MMQiKOIg9EfEtiMuqOG3tbvA2c8F29gwoZnPBumPdka+382FpO8E9ddl3
Kg6YEGoAMEuBV6QFeFysFKGombGui7kI1Gs+16YH77Br0cx76sLioZ5QZWCENZUr
o8gpwl9ugxOcJPveN/HHTmbyAxoXdAkggP9U4kf7NH+IUbvwhgxGLH4xow+DPbTm
OwxOnnscDk+vVcH+yEp1ih0M/gcx891TE9NljnM2gB3LJwkloLwO0XPhSK32KJBt
QSbX3FYtKfaViHFPvoZQMga99RUt/2CURcykCHN6alvcliRJB9PfKHzt8L2ZC8p8
CkMX53+X8w2w4UPADi1G6ldHRXDPifzDtIWpmrNzDun9C6nRiZtCI9UUgxxMpjRb
7TsONw6fOSKXtHfLpjJGsMBvY5IVUzyAcjA66m+svfNRZArUXuhJYM7ayvt5bZB/
H/C3X+t7YJdCD0izamHZSY65pqhSrfe5cjCmFxFuNZUVPRpcQsX/oYQalZ7dFaL/
SlJb4maGFiVJH4mQKtc+hqWtPXLr9sFwgt4cPjF/VexTEAKzDmPwS5h/LWaIAVTR
rUpVp+22vhCUK9TnLnQyls1wAFybScQsv19cLtepCtfiAIdKKH8a5bKXpGUO1pbL
2uSD7lPvnFnYisxvpdQzY3sBw2ycTWK0/h1kQ4Y9s9ms+IZGPq3SXhZTytVLOKZ0
rMYbMILokNMVgJ6JInRvBnbrzBIbUN1IMtTaQgjG26nqArAoMzW3ZKTjvz3qHU47
7Jn4evvwtDN7UmTNwUcTdOlk4Adbscv1aDjS3S3fvZPbQ6E0LVd/PpkRAPP2L4kN
uwYxNILBagiW9HKTpUuO0mf0M2npCGD68/aubP1DsFBEio6Im++oPzqAEUOxEcFc
Y8HFSnPBKs9o5sygFKgK/eVnMS+8aoGK+fjOvWn/GpzRt0D2HdLZApJqVyYAwGTz
PLsd9+5XihKqk09XVAWK+DlZDyPNKoncLsF7AaaxRwCXDfOG49mlv0EEYbJMoO8J
sP2jTwPZl7lm6h32ihgYwApifMHlnsB6/6kd+StqDGzclS+al9tzDiTvNeUcRGGt
zK/RoZJjd4UgcDwfuBqO9ksdqvdHJ74CMBA/hKgMwqZP7AjS+XUcPp4nnTb1yCEX
S3gWxnIfHyR+CxMQHlyxASuC0bjiKDpaWiXrS8roZ2UB9UGmDYu9Hkk7v7l4ZAFW
j9vf8cs8xKcbHOjKq6LMZbyDEhBzJhIE6tuXslOOsPKJB6lLaX1/iFMe8uS6N6zP
cvx2/qQ5/Coc438b2xpH+Av0EsWjEpEoXBiQsJ7XGP+YZutk/ztlNcRhhnHbT/w7
Wu1MoCViL1V1Vla6GnqzI/aQ5VGdopmhGv5SuVwlAkI20+BdbHwYqsevQwYsRqBA
FBzcn9iVaSAhJougkoYSLAR4SDXIAoOMPEovqsUQ4RjsDoXSStxH8p1LjBC6MTO2
HO9H5z9QyxCvgRbYmehu7hd2EZ8Lq8fYh0CYck8n8+lc8wYtskgM9KhwRZB2cmxW
Ew+jN3HH6VqcUha/w9QxnsRI8yF2YEcGTbnkS7EHQzWCVAZTCjGjsp4ss26eKViU
ZmVRwkyL95MZFOPlqOzpPJcqmiNVTkuzFuuYFeSEJdb3gTMwOb6j4t/mtZvwX9xv
PmnhZKp/5VIu66iaMpeiDYtOLBWrDpCmHQau9DLAMR0oTGJXyLe8wZMeUQviPOxy
yggxPzC+QUcG4weo0kHYKCfhAxVaPLmBNtK4nv/SHEk3hSDXhYAs5Uvls4sM/mIS
lU0a15A5AWFLIhSXPuajcMgbP4vfVG/1Pk/hl52NKsmxvHOHj4Gkp6zlcAaxQt/O
NXrecThb1XAW72MCVpcGSKDRgWEnLY9K3uugiO+n0di1Y/sOyrTWipDUh7lh3Jx+
f9J35x5MfbX93V1i1jQ5RF3MnR0l+OgC6FWaDto8jytnhGl1r+9cn9/623X2YP39
cTdKFz0fSfVb8VOHvQyfqPiMzAS7JpC1Eof5GvfaXbDbuBZqsImT/6V9LfvM6zjN
Or0u5xmAYw6UCd5PxvS8m7/KAh7SZB4xrmaAoLJZ5NAK7QPGHZUjixBHTrxTm4LZ
j7tadso/yn5QjLA1fKyTvDyHMydZtp/TiBXxnARP0FyDUi7OPltnqSYFJiPWKJcV
aCHixmrXCe3Ea9d5mbwXuycg9SDOOaQIFKRgOsdJTr+Wh2fQJCWLKL0W2Lm1GUBB
zW0FEyFBn89TmIMSshudroUbn7qbqcmLoKlWR5kU3L0b42Q62zqV0+RfG8ViVEVx
3gRrEyHLgSzag3N6DmR/lv+BPX92mFGjOaMCcjvRFs0dD+1iFd3RRXByY8AExX8H
j5soHkqFVBYhVm6SvHVUMurKH05lWHb3foCAmi8QwGpq51k4JCWjYGIntW46nIpB
HMfAoKiMGQnG55ExONn3oJmmAhJ7PNGGeRlSwf6TwCk5VuRz71cc9fYADOwy/o4J
JEXin5h028rxvzLtmOaOgHqsJmm/pzjEO0pg6nBitGTMkspDiE7Xt22SeETtNnlH
yYxs/rasdSa24VFY/x2UzIMalFkgbRPNOlRJr4AqFz0h53mLY10fs2aOX086ecEp
ULTY7uu2wb6t7GzG/MXpM190Puwq1ngJ08Hbau2bTN26us5sjVcx9oR/gx2czw8e
WlLr5rq+dTt/dhYLMMhPoD8WdRFi+FBG+PckXuyTHP3oGSD+eKz7AejKhF4HElkt
QrKCf/76gfm+uTctsvgfh/k+XM2oFwssW2x3v98pEUKIZCvuRJXhIduSaqMGKQ0M
yzmRJuV1XWiyiOIFUJBO7lzx6+0JJ5TSm1xlKv+1c2vB5nQeLC1cGKYEwqNFFRzk
xodZcSQAU9EHWhJZGuJ3QSerGzPBzdRGweVPt7hPEEpD40i7PxpxVh7CGI7MOpk2
P+6W7D5PN92QAfNntxUMdTMBTL+9POt/CuS0GjNZJaK/zKE37D3MUWEdvshHBBMr
4oFCjKBAS5flBDNXFxE9G7c+d9uLpMza7mqhHyFwSUU+6E0AJI3mssAQDJis9SeP
GFLzHB77RssSjr2Jp0xycrqWFfUtcIngnpwHkarVw5gCA7Lw/K7MmVJfpKSTnEih
VzajbbBf0Rw+pCBzH6FgY/U7el2pKHxcNr8RoW+wt/Q7bepNm3ujoDtFeuesOPc+
xOvZ1oZ9OCOchqKD++BeUx9jsqD8bRAgyUY94ve1yyP/ydicU6dVfCegLEFnkpaD
RvJpVwDfSJn3oAcbqxuzB0vM2F5z9yiUVmgRZ586hX1gVzzeSikjlcG60nxqK1Xs
GKEMH/SRjgNXAhCkJJwq6zBqIdL0Rl6sWm7cNuT4oQniri0aQ4I9LNCUulIqnqWN
NEKRriMkH8k9cwRBOjbvp5cemeabLhUkCmNn6J2qQQe+QsO4p9nAGgxGIvFMeo9m
w8N2uQrAOPnSK400iiTyso7T4VAsli95lIJe32rrxr3rUaKB9VaQGea12NniUbyl
jPbuSZRcbTZkYCkaZe3hcvTP193aGV5UyH2ToPNMkAGNqdiNWnLdmd1CqiC1W2qW
hLkuahSy7zfl8YwKliKJpK0cKjOYSWKLXwvK+ymPZJSJ9ycmqBgHoK7oCgDJ/zk1
j/A1aJrP+IB1E9cLTJIh44sAuqkzClLnivPGPVhVt36cHcm2X58ISo3nJKPz4Jsd
nautT9KAAQBRBs55s5MvwdB4JADjdJvZspgejmAjmnZPEfgR/Vk1FV45o3xBdeJT
/PZXthvCRYi3/0h+wkKlmdvsfvbklCCLXnAOjks8Qn/UzY6JP1JYx32T3YRPi/mz
Wui5eDuIWP9Af4W/f2BMppUUhlyciidifs+plZk014JYX/yKCB5Jpe5qtudRjM6A
Fxx0kpv5h+UJGEP5uNNyeVr34Dp3PPsE/5hwXXvuuylSceI2gExatYRIMmp4Rbci
++zEoAfaSBV8rtykakC625SU9IHqZIHn9pOctAEPd9kc0lB8CEshXCMtW5kzNVOE
vdjY164n1UfQyL4MjyiwW8QGzIOrsMgEaTT08SWCmW4gdZbqCtCi+66q7NXB4A2T
7Q+7zdGTEIkuBCZz6vtwAoItMe9MYZOtkMNmSwq6yUbX1KR0POeDP8UqlGqKCcf8
DRNqPo/LF8wVmTggFyHl7cl/Gvec08JynL3cusYY/ciVM12jma3zEfvP5rDIPJ0Q
FqA6Ch6cJpCTJPf9bAOCCVDypnA+oDQnQpkLiw0qXpHWyNW3KqhVSR1w2dNsuGHY
SDjOKrHWR11fbYFPacLY/o5XOiH9W43ySZVhVLuiMwSF5O97Sbafl6BM7V5c9Lp/
ZPeaBb7Al/XYB5L2rMQOtEkaZKCC2VEtmMF9ok+q9gWYWKXdbLX/61n+oQrnPxtx
qulnAYfamMGoC/UBt2PKd1x9C72Q9XQU5zfVHXl1lZ32mEiGHrb+CoRETWzjtTfM
aOVKK5QW4ZBC7L0wn7ekBYiB3K/cIQBEOZWUkCF7k5hh4iSog4B99zkMJLfd5hWd
I2eU/YllrZ7IrtWikbK7h6265r5CIp1NTFAbhlr+EQK9/jOuahts3EO+cs64CJ3k
23wk6fcZrks0IGrAWWqo563c87am1lg0vZH6vOyS1rjI66jF4NfOcAq9KZEF6h08
t8W1V/MlMfT+sMEwzGvRDM9PPXLn8Hb05ThNTrPtHZal//Y7ijNgUwOizzzctgl5
eB6FAHGBmW7VQz9u63XVTOu5XPmOwoRE7IXIqmWVGjd4DQ6Z6fHR9VuToseMEaG5
PsLF5ev1FiknbvzjT+TrrgEuGkwjiYDXrlo0lFLpvKeUqv7/VnfDTuSGJJojc39O
Tihkf0i7MYSesHeujdKmh+KRs2p+PCfOcmm0JTdtmTB075yLIhhqAhGNcmdP/0NQ
OTrypdCQXWv9Bd3RE3dbgx9Tme60MDbfms1kKAGC2ntEIVjndgNQre/g+HF7+YDV
JKbR4BOaV20FX5ECcnETVzbE9/DSwH56fgRxJUDrIvZcfKQukd434xpBOnWzQGJj
EBEDj8QqFpXgAvBw6lFreQywY716//U+pKAM/Djd3TY49WVul78SPpFZ0YdJIvmj
jGEmBK/e3CsWJ+88XLUeLCux9g6WU4EUbLzG0NODagAnhLYcLo8ERGRWCSMeDefq
lLtQLfPgV+Lvy5fUvukJmNbmQM5PsErTiFx4/uZAkKo/ynad9JNQFKIZEjCKdgXa
1VPYe1eaqIq0HkBYab9UQY0gFjbft7INO8oUsIdFHZKU+DeuCwoFiF2OVyqN9mG+
Rc9bur6LFYFPL1dD8+ZWT6sC5AsmPCO5gaW+Dfbrho1xnPJrnj8BgD1Stq5/7cbS
DqiFEmNdH6/fRYi1Zb9OdxviruFYFGqg343uLWgcCIn1zAXS5J5L+5iU+yJQRm+E
jjtISgAgPdtlJBsplEI5UKpTwD5iJ0mvxZo/1mVpHyeJmmw18L5Zb+aEWE2PkQJs
O0K30dr3thWyK3gU88Dpp18m7R1IyJ5YqwJ9ZUbIMtRQftHscF2dw97JlpDxNZ5m
kNGriZFpbp6jXyByVD7ieXvgfj2MpK9tywe8Ad85bywvsNEMsFW+Drm1wkEhqI79
zs7rN8zD+83lQayChv0c/8Ub70IdTYKFfe83l3q4KKpeZsVCejVqYW8baDBywZGv
25lcLJDUQa8p0ZB4YE4GYDZ3fBufU2HFOJr9wEvhbDqlXuv2Ddo9O3fP2tAaV9fM
zwMrIo6DA1SDan6U7LJwxYbEAaclSpTLQYFxPPWuIbJ3iCjV82FOQqMNK59F+Y9a
K/WaG7xG2JbOeVXv9uXk5UAnvnVefIKo0l0B85lt8KYJmstUPLbRTatMcAAs0IrZ
EkEzQe5TgLKCb91tzCrJVSraWFYASCDY9QlVtOb6WzD7rLxt1zFFZw5MUl3/nUt/
z6ZlpgNHuLQwHvMYXxsoy4qu+LTm43OkWjcZrsoicJ4613HpYhB8qT/NojcT090z
BKBW48tPDrsEGmjHVjVqLYHmipdxK2wR8XkPfPByCE2rHvmlxHKc9XBkVs6zUd+q
1N1B0ZV2FkW0R5aAYPgCHDFk6W8wAcwjYYw+GvXowh3bgPKErQaSg1KWNDwa2Qqa
hNMd+jj01/9rK48lDHsa7slGb3280FtqGAZHkzzV4dbgj3CMspntfmaaHuow9eOG
8nGXRtELlIAi6oIwUkm540xR3o2TwpLhNk4ychTXqqokqVbDGi12WXQeOaVa4Gl3
uK+rcQJSoRvUgKtFgdPEtOdW8g0zrJLQMpI1dM9W8UgZPrivI56RXeQ03vj5j/0g
XCWCb8rx3LQ9lpuURhLvS0jm9llbhjiCgkokPcDTx7yW5Om+41Ueg0u9Z4/dkYD1
9WftYE57LNjHX4IfEeB4JAzbqG6ddOG33/eVhx+juycc83sHMC3J+wxFcI7uYnS9
oSk/WtKETQYQUbo9LbIY6MetoFijeKnkvMl0oLNguKMYeWsFPDacTvwj8FkA75nT
nHUgoN8WojqV/eSnRqoQ56+bfomVoa1AoaP8XBByOzc2AtJzkNEhqZEl91c7dU+p
uI3d2T/OM/4LOsMS72m+/d4V3aECJAJE2HW6Mmj/3EYGViFLTmiz5gaJIGLnAAOs
DVaSny9VWQisaSPoGmb5hNZi1swaaD/ZKjbrKGxfzTzF1JvJR+piOzCK5a150KNo
+lcvuOXc6Kll/9rcR5Lu9wmxDqsXeFe5BroHHz/NC4VGL7gzWNyl94jH/VOura0d
3jdebr8zYhY6MNiQBnLdBbaEtxRGptCGl3zylJRhDakFI9ePsrPis8IHBJpLVTwK
1OJ1zc8D+ZmKlrWP1RNffcF7Y2fysrONNU+5PrX1UynEfFDEID4DBlu/p2fDTjvP
bxFgOHal5PZWA4AjIJIICIma3jV4ZFc410WIldzqKgUm+HrbswoWFXqE+//w7ETK
AkHZJwAz1evsMmhAQDoBOMc18aaNulMBhtI5atHsCATQ+1ycMR4nAlBzYbpNbuy3
L5oJLNSp26WVVM+sYc21VfOTsSpcMON5kpKcWhIoQY1AYmyilFCp6lnbJ6qS3WCq
ZzHrDDK0cIeM9TwBAKq/KFM8memFBFi06bH5plk/mZKwJlvqU15CM5eJvNmPWP7R
jMvCG5VVuE4aHgoriAHX1RhZ5hFD0J4S5q7WzXpYCu+Kl+cWfGZskVUvou/uGTvl
EkSGGUdeyRlRuSdGUKhUSMXgQ8h8nFR3WJvLJSwjAe7zjhnN2mgGHgYCViPNrPBx
sL3ZvIqagdvETgPp20oNqNKULi5MO2j5H7U5IiY5D2UAc6edTbTFzjEF68nPKhqo
a5LAVBWptf50sapO3fdpGzCliZJw5Ntd8gNuSjXQXId1YeT4rYN0L9qJWft94hYN
G4YZ9faGVbPAf3aHHDorE+oJC61wKwg2ZTaRfNdcxHQ5iLHi9F7ebT3+0c6hudJa
PUbw5d4RtRREmYpXnPyMX1kbDA0vBZqOLnDdLuYwbkjUw6iQB0R8Id4h8geJvo5C
9UnRI9scgy4m9z1PxlGKv+Fn87pgkM2BIUeLP7QPRXD7IqHE9tL3C4eCHcdXHPhs
CtofaZOITCjZF4zQzvk4SBNv2j3a+NArvNSgDF0+heQ3XU4avg0JCoNEzLvjjsa2
pZfLjXdcxF9yAifAmcCrNm6ibYrQaZdJwcbDlFubV7IntKNZuOPkruhp4NqLpYRT
LNQha+cmhl5CBdr10eVMT+UbbogfA8M1rTs14mrkeOwBGMkjkXnyRD2RYbgvjVKn
5HwcMlLDyn2DMwa5LUiOs8xRrCyJc7tcKNNB6q0lgSCr+5ZKBDooo8fH3TZA3sHk
TUm8NFrs9yHijPUPmrYUp4RJycQmqSM4MSSgd2k8A/zaPaJ9K7RYTul322c0aLRW
3JpZ7Ix9XuEKumaHNJqZatpRx9WjCVjs2cUp3Ajl3UT4kafO/AtukwLDLShGGHLi
7Hik4vsckkY9lYlRXMCKqEGm3YyNgbA9n3E0GMTzqfxQO84x93TbAvJRQ/fxMSiS
BpquoIHyxKFW5VN36a0mesFUjZsworXgBf35XD9Ml9pkH8f4bHJCczjNiv/+n/VH
P9gqkh229GTO3eIt91DmI5tmQtuzORqHNhV/Ktxsc2Hlh8MVozPHpcYU5rnNe5E1
aLlsanJWblGRtU8o8pl+GXNLZkrzF8Fh+yiUAtXfGKmJ9BycF0sDAddxVGbgM8Ng
HnOT2/WLjsfb0b7ckh+Fm9QaTN5G9UEVi9ScWxdeq/NZ3N/f6UKYsEgaTWeWnMCK
lFNK2Whlo2VW1H2u+xDr9Ag8CWp0IXejCAPd7Y09aE3iyf7DBgiut8r9LLVE/YG/
G3NWFUkhh9Iz43/SrvDtsB/Y1/s7xMiw3NOPDqJNd1D7PF8dVUGb9jAjsBuN56l3
OMxRz4O/6EZw5wHD+OSQKPyQdXVsejFjs2THw6KirybLgYHr9cpGrFO7Ok0cMhAo
ePZSAZEm22v4Z/y35ORIjU2PIilH7wacDTQ6zQmLNJWfFGJFiCKeFFSdbUSdfOc9
xEVJXACbyG+6iQS7Ij5ZV8VxG+xmfA3d2Ve/mDg9UNccWa0fntTMJmu6RdPU4tRC
BX+efljHT/D+s5pZd6v+/XBOTyNv037hXp7BN3xUUcRgjMw7mZTJvjl4CZaMRO6W
/2GfZmOxrNqf7peW5pRaGbIH2D2kkexp0vVE1ZPKzot8cxifl+0+C5BOm9yidYF1
yv6TBooZ/DWWrV5dqX+qkkmJ4+KdXZb8jE4c73u16NGPtjc5YE3W9yyGgAYTdrkz
xaNTleyahtuVd6JKY3ODuqpFP3CaNs8k1fUK2cXqq1NA+tM/3umhfLZJFjK2SOsM
apaDrcOEW7cRNMYK3TUPhs39ulvgQP1YCgUNvGl+EilwAaKIKYlrUyTTGd7Oxw+R
cTqg09NHPtrHqZxzpfHZS0P4lZ394MZTeQEk/zlL4HCE25rOle1nuLBtjuPk1zoW
D8Z8EGJhn6IimnPYFrRVNSU1rbCMsYvOdKOFeuNyWpgfNGC5+MT8Sur6AAULXSnl
R0hSN93ewkqhpbhVv1+yHEonBPmLSO8vT2zM6vU4l79KgRckwD3njbAbux7xiIjG
U3Ddu/3pdEgT6QXYfJIU6Je38dEJlIKFKo4S3OIvFPHeHex8AUFnlfvw0aT39mvO
+bIdkwX5pKcb00xfitJymeRig2wDli2sd6d46gZaIvSlw1b3J2xSoqR2TlVNQ/wT
tEnKAtlhHTVUmKj4EGRAPN1B83YTA9freIcrLDPf0K8CqYhT7OqDadDfIRK92a/R
oEof7Rf5rQTdNWY02dz4GugijcvapuYgOZazPye905BHKGYFJHHPKnb7eTOT8CIZ
0ptQHuh7GhH1Yyotr0ZFy9C9mHPBr538g/tc4JgdeKYcP5T5oDngXPq02yEb63Pn
96GgF/wCsmZpNab/a966esfRqeBImWK41Bos8hgaunFoDIE/S+a8kSca6luScZo3
gXgf/6JjNMxmm17P33BmKEgH3a+QIlhGKX9PSd8r6l7xF9rbdBw7yZUbud8iuLeN
RbgXzU+SYudQRcm4Zw8zNfh2rQIH8pM1h7m8yYZ48KZgb+CeDf1Pw1aYHys8Hxvw
4GvYsZF2r7In4PUVKRfeLBKh00DA2xU13f44/1jLeAWjT1gFfbCH+unZtjTpm39n
WXFvDuwcrRpqubWGV2Gy8JThC2G+mHJ3fPKpkeo8lfY+Fee1+2+6oYfSkPZ73TNW
s41IB2BmpAH6uHzWaVwx3GJSwVsIF9FJisSjd12BoIgAKxJueTN2tSHUTSKL3BID
s4OBKa7wSeoTY0muTSw3X/fup87l5eM3f3+sgYDJIkCTObVBt8/62W09czxDl+EX
mVi5xgTo25cxaBVsGQjQ5WfvJjKKxwp3mPr8KmX+6heILZdSYnZ08C1UGR0vajmU
tf4++EWb8riCJLCs2xBRmCneDzKC/SEPElSh91H8VRTJNH/MbYmmju8gCAfBnND9
hwZM/AsZdF06MASJoiH6eJjUB6Uxkpoy8U461l0k1bSGr9+KVorDVf5Zt5lY0yty
2U30PK6BUvityz70M/AfQvYr7To7FagLL4+NqR2463zDiCRfZRXtfPSIHb69kRBJ
bOoI4bx7zREzN7iiu2Weitsl1L49VVMnk0EGHyO+MRxismR4r0epSjup87dkDVrA
Qpc8+y3Ua8BHUc7wAhWtUDSFORETq1naBLd12aScimuU47SgyK6LFo0JjRRYvTDw
yklE8YGQMk89QLqdTEIEpU8k3DTpCrRWelJp37CjdePZ3HlmtqkQ/3vYMrZmdVwe
p5p/PeUIQPymDYpLEboy5gHFrxkAul1xkCOkXBRCiTFG947pLU3HHVyvHx0ACKDE
j2GCebDxMeYFUzq9F6kTuTFYALfyewpqLHfBprDwPKkTUXw+nGcp4p9vK1FURxPD
DDQpxIq4vMkQzQ4Mb6cZf889vxXbrMresTUqVH5nzNuzyI/SZeKNuBOBoD3K2TCb
PMTSX7M3Bw0rP67S/T9RJsV4w860cRILLyhflYOgX2NfZn3g9kuXlW5e6Vl1w79I
S3xBmVA//Xo8V+nBiWYv4WvB6Ed1r5UxOFD6uDZ93FngQXP8q9SV66vG4u/EM/7v
ZzVCGpLl+Nd9pSTy9JvfC9jtVaYfdHjRk8lEQ/oN0rEHf01rmzWJHxhMaVi6wUbZ
MIwa55DfvbS3+WRdOBNHTeqYUxFO6K2ely2+kR9F/EWO2m+nHpjD3lUFJ44uE2ET
WTP6uJOFMzrRWjNtJWk7crDbIZQVBQY6eLTUeN8o0dOpDAMF/PzPQfP8JVxPdHPa
c45LvYwFcMVsdWB+yVWpbBZBnsC+/mExV30u3SWLCiCgWTAixMjA5dbMAacuPfX0
MHYcCgmYPMIIiafFeoFGbw5+0IQhcqmpDTYd6kxL2qiIQap6yzH/Y7DzcZ0vJ0dx
MtpwMPnCyc2EnQwAZY402quFD/RjMNSi8pVMkSzyg99yiUwtsqU6A8SN7ee3GVbg
9SFgJU49J8keNC5YWYbs5w4098/q9d1T360g3ClzEnDsMvtSOKKj9dZiMKW6dqLc
QJrHbiwU4+doDx+Egn8ULL5TbK2jpHlIZtI6mK29cki07cdZb38tLMqLB0VoShrl
NH+X5qZP7k1PqFLlRtn/ZaljypnpsEDLsLJJWyjP+3efSn4uEmE8a8aBLo12TUdh
76RqJCpz39wUhWUv+z2rn+d52weEk43l6sT+PqPrBpY5Aav01iLOjp4X2sZ7BYIY
3RSrsI75cA1bN1R2YH7vdqmmiQMGlYntqCIes0YY3FnbvTLYX0DHqAmKM5ZO55zy
Qiir8SxcmOOHSPnx/0UnLME06cMdpQwnVUTqMUTKKJa9S09tMin9BcC6+GPKvNmA
fZMmDslUwDgoxeEbscOJfZ48F0jIYbBLTYm7mmFuyUsLkIGlaXtmqxsdRYGacWH7
qdhvWhNVr/NxQ+kQ7VrtXT5wl0WhbhNyM2iHTAki9rjewLrS/UKiubwIevUMxlNz
FrVBbfD8hk7yPCmUS+BsZE/hlEfPvIwUWipRaA3+emjdQ1nQ+XxiMeGTbwBLSui4
l3ekzs332vM3k+qGx4VHbtDAdMVWbiTb661h2tdrOfM+/oaAJUREo2KzxLLDQnx+
qSqLODmT7cRoOls7OCSqtFaaL2yPkoovBfjUqmdl2fgpOd4SpaeHRDKtuOys4nLX
FECHdWLvhd0G9vv2mWYW1XksrQAan/Wo7Tx+c7GVOmHg/YtLt6urVS9Y+NskHone
riN9ife76p05/mzCcn8Hy5PxbL3QowrXO0Hs/49J41zx9msdmVYDDRqJiDgGrxyo
DAVTS1Xzc/9XZ4iN4vweMWv3oToBGVf4cI7OMHpwIcrxgkp144HkYkMx5VwW5QxG
git0k2mV3d7A3lknlU9r+0vT06U/RiV4KvwSena2kMMtaqmZMFvyG/L+tIQIdxXG
HQiy1HJp3zjO0iFwhY6I7Jjvp3hSkQME0KuUHyQwTD2mhauoalogw/KeN/eANP1C
KS0IL8FEX2jFHe2cJZWEjOLVSjSLGx36nL+x5a65VPmcbFqbc9CBpF2lCBSX4AIN
kkJ74zIHb+WETNvOHOr27rwc+Mo+ZFR1tGB48r5RHhZC2fljuOuCNu0E5j/ijXEJ
gX0+Pv252+bK3IJlzDuTfUXXKkoIO2M+8qUbYv5TVNyKyKvU+0NKv8MwNiXS3jvA
BXVQe9InfdcNpVLDz0uvn7qhuZ851dsDIlDKJ9BMJONImzUX1Ej5v6h212NusdPa
FtGp1yjEJDHASoPlUpb2LrHIRjwrI4G7o1PM8hcIB7kVn49OTsbLWAkuNmTTIQxU
QpmvfraxAbwk1N9h6j8BIwWrNn61VxughQtdFRkCzg6gGvNp8PxEWLR7/neRNbS4
ft4yQnMjnQqj/NTzdGrlFQj7ej3NQetMIz51l3Xz6YfGLeq1SrXe3krwqExtBqDw
hAn4AaOVvYsB+d1R7xohu1vMm9GwD9s7184KysN5CIN/CbIpIk7VPvnk9/4/oXhx
zUiCpSspM2RH9XlX6jDD6xNJJlnzeHIhHOVwReXQdKG8V3kvD4acYBsuzyyAzvws
Hm1GVyRLxwTlwNxzd9wl1ISZMZRtKH2+sUhQny5RUyJ1+16BCU29JNmiIqbGx2OS
K3AI9MpMw31XjsDrFqlmHGo5lgrf+aVvppjHmPBNTLBknaJ3MYhCSaF8Eqx2cIrD
+P35OZ7Jp7UiqxLiozhHRip4v/9ZJqVwBgyFUrgn6iDjklrh1/vF/H/RqSExxAs3
72RPcEzfweCErfUvTLZP5ocGkHxep3gNbtPzCncL81vsbrBuSzPisLfUdMLbUQzu
c4ejAKUWA9HfAqS596+lKLBQlX01Ku55jJTjsNvVZFZs1OjrCtRx8nixlNhEcLmG
AV+jZte+JhGxxQ6ZEW1eI1jYz1RwH75ssT4oiUqC9cPqMEJytYwj/6VUMc4BOzKk
4H6OPBW534dU3t4bQW5p4Xtdhc54AwoLhQk/vAqJrJXiQAaKzXhXxkZRttjnRnE6
B8O6GWAWqeAd4xmJe6me27n5vJNBsD/qfDIu68Z5t8h+Cew9leb/L25W8fgSOSyU
Wvcouk8b2COFLCaYWE4dEsogUVOlHWVLX/ql+CyYdk9s09LfhPNX8wmh8865UMtb
+/ebW/3UNLxjVbFLH2ygKD3HAYWr6IZmknjxa8Hyao9ykU9iajsLX7rAfsqiQEoW
6OqU3BNYkNf+/GY6HKi1PqI8QeoJOx97Y1F9IAzSs8QECaaxBalWgj4uZJzHtKBa
jB90bkjNcp1TBl2MF8GZ55JbGZ3KUliyw9amhbuO8GdSghmTsbb27YIbBfxj3LdP
3pYHxE0UO7hixSG3dAsed43urzHhDo3nuvSjipcIS2iSI8IpcbAxrzYY5VsBIgRf
hV0H2asFIcVRi6NgkbZ48s0Ksk0+JpFNIsi3lwL+WDZhla8DvKv9qcVdTv9fXgBa
Uk9VrzFh0Ixdnf/AIyfmlQ6ODy1i9i1hF/LEVEyXEC80/WkR9wzSSDBKjZY2UNro
nZoEmV0vTbqOKsOiNm0ayR2CZ3q79niwPX5q/MynhrqgBDCXOfxkDVedPqz3yGK7
6a2xbneZahrin5gpE5795r0N3ZzwEvnZ1S8V2mP5g/G5ejlKoRZ1QcCnL/zOVlcO
QOYHmQJgqhtVRXm4pydnrPyctabH1RTfwVjKPcYOCIctRVTMmEvBJh753ftI+41v
xpEOef7E7CAk9vKmdyGOrvtuBhNPEvEOGZqu3QrFS6vvSL4xHZ5YuYEXhiK981ZX
xk88mbC+qTgbwIGTXsk7fe5sQu9Ydn6A1H9N7RUjtiyT56PpBDXRHw/fidpzeeBy
tCCk2VDMVu+jTAIvhAfdIyovjEa5ZKrgUS/GcuwJXVBf699jyV0oldG6rA6bfPMO
HAC4UfrkVQHzMDEUvL2ctpCLcMqxbGngOdKUtqZulD5Hbrky2ypCIHApiqElIRSX
Y8OEISkT9QFlkkrdIcONxnFPyabxXfrwB+ybiWr+SY+zMZL6c27KwVq4Acwz41js
tiUTJj5oI3PkZFyWUonR+dVu+cEUJqCmXkJozilNr+OFNdjHQA8uHFMVeDWEIzR+
pMzqH/BAponn6MppWtPKwuSBUVW2dsWsajxDpATT6xzd6gLdnlbNsiojyFGhVzq9
8FVM2EPgF7LVgiZT9ckLbY5kyz/N0DEBHfCcjCQfun7VeN9sebfXEWc3RTAJfafn
ya4FmZsixnSp+eqxdHdfeE3869RSS89AA5R8xlKH/3S4UK+88w10jZJUaooeqAkR
eonPjw/gN59S3YFZf5qNsWhY7VypOH1ignM2rLSa+byMPTH2C7c9b1qdgnd/F7Ls
ew+UXBeY9fvZ22Jouj+QdUkqQipDk8GYUOMAEl1Ju8vBQQAMvIdmcycBJcYzCk3n
499rmGDGyaGiMl/dAxxBOe+uXb5e7bG+sfrS+irAXgxD5XWB79ymPG91hLsO2UOt
EZyX6cCGsx1/Ggl/fXA3Q8RAm9GTqLl4YZN4SuDvD82KTk/A9E9CT8atxgN9BGhX
0j4aT9uDLxZ0Mxe+oEBxHX8SrMzVIlFr9DR/a3fjHw934Uj+M3WCnJK/VojiQvET
yZ2RP0Woa3d2ORghsbVQrYzlts6iyDyIfSq00fk4OGQW/KLlKK0XiEznt8nBizZd
xN1HEO/uymjt+gyuO9NrrHV8FjLkU0MxvjvfSFCVlL4=
`pragma protect end_protected
