// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UGV85h4clcgIa7hzE3J6m9WfURN2Gm1OXrZnhtbN/vh1fYKZuECv/GljNe37CO45JTyX6gIdIzoN
V+WWIShfB6tI810Nc/+Ls6GPOvBbxN7pu85RwiahrAetDWu5L1TGP68bZznaQXdq3LC9ThS/+L42
7UivNsT4V3ccXbtBaoCdroyarSiUPSL2nhBVMRtph8r53+qBPWh785HHVXpiwpAR0prm0daTPLTI
iIDkjh7nQf2tEHFbjz+k5/6zUz3acl7ebYhvwIGJNMRasz4J9OFW8iLOlnOLTBJQEQnCPcivgR3D
dVXSTOngF/Zk+aKF1WYlaWG0+1VYwtlF/VdO/A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9392)
Cc2CDEJUYwm0iJyZDpzpLOMMzAWPDwyVeAG37xjqaQGSexdug3sNfcq+yrJi9cAfBTphh+T/Qigj
VlK07shHGgcqLgbyBkAht1l0e3Ise1i6K4TFGZ2ovo/mSFN43Fg1ScsCMWBt8YbgG8SGRPjGAhEt
5dKEZ0U54qTH6J6Bmh4cEFdsi+6lp9JGbSkhzUh73dtXdQ/6eaJAgunpwmLc770aKld1DNhtEg0l
XqxNNmRa3biqtuiawK2iOa5B2ar4idI9vLa3khocYcFJP9dNC7YyOTGugiS2zvu1Io8xE2SaP8dd
psdqKrOpB4s73VRKZsaFgXqWRUKASsIx6Vuop49kMD+Xb9TZgULp0ZUdnXOzwPWHYnDxiTQkMrn/
a6GXgfqn+egtlhwOIJ3DTz2/hLXeVXM/UipqF6RK0aytLPlgF9wVN9NANVb6yn1lPeXm1ZRFfQHo
UIF9bRp0uyVYYvxiXCrisBWMxES7+nXgBmRVQtjxvANgnGbDwQvavpJ/aPaD+4PqL9uAT/wTrw3m
VIfyjwPZbHQ8zDBghBY94h+wJfV3Uq+cfyhhxvbLaEkccbL591rOZ8dK55eSOq1nwwncZIWSLcqo
STo0MUQJyL92Gv60JoIKFDOwTfdwMzr57sQT7UIA0fb3Fxt3cKtYL0hOSRA45BXgGjD0X90fbU7d
Tjb83K4pgRsB/9ZRPt4JtbikOWTESktZQn4QN8wxjPFBNAP+ntEnz26/X+5p9ybIfqZUA5nlaN7Y
xifd/EjidcK32Jcy5Y23bYaBWFdj/ZCYc21jGfZMAE4uHNMMl3G9Fv0M/Rsj8aBs+MGsnDQkOQ7X
ETjRu0tO6E1NMcVEoIJVscpFgK+5DSCRHHO4+wzA3BURrB2LEsne0xr3ANH9FrNTkSJT4HxwhN9A
4yolgr5PibG9+oAmQ3yHZJOXtubpNFZkj4NDVCEyyQ6StjJWf3HmEdqNgCZZTIb/0hLJwYBai8bb
qoV2wixAK+DbyploNqH6IgeMYMIR4/L5h5e4oXrcSdAfslaldNSdFOUAma0P2fxUufHIdYKAjWAD
PphFmiZ1CtNHDPuXNa3yYTi+paupvp7XLUR9sAPOwxR7DjvrG4U9+2xvV3scmrdQs2AKYM0akPlV
Ck7VyxYgK7Y57/lH+57RAWyTZQ48GObtF2rkNYy6hKe/XOA78fIhhf82JowbKptp/4qu4mGHk1CX
+QCjq4CAFGgIo+/CWrVzSKLTRGhTvE3HNVMCpNejotLjLTUsotafT7i2C1wT/R/wFfhorF+zogTP
aQx0tlGml7Ty9XMH3y8Q+qu2k5zH7XIt6HWQoNwZ2iEKrMG2dEukaGK7EpICCSiBckNThiwKMovQ
hMPnQlr8yR3aSK8oNY2HE9WVlCH5pIqPQ+npMLQ3LYfAahIKmTSHlGGte813ZCOOduPDWtDC3iqf
BmyqYUYOZAm0c3A32FZg6RoBnFOTf9VwKdAjDtM8HBNsHYbz45ugg3F0KDLgbqhfYqePhj20xn5m
J0IplHdMpnhJVzIGuxaX7ztFtOAty15yzARX7EuOLHirxk9Ys7t+MAXPVvMkYzRoxKhtfbD4WhxB
U2a/ZYtgGHs9f7VCE/XWidX/T2Cr2wN34Gd4qXQr8ZWGOvdn3SCvgJmJqL32nIKw5h/qkOzC7tRn
lB6KIQeOHy43vywpCGrsui+XoHfmZmxgWm0ZzygFo/dxSawegxS2j9AJJSCck2gqDX3Qy7Z/wGlf
UgXgQgB9fJsXMlsNAsvx6LcRQ9wQlm4i1Kgg12lTw1kJk8HuDEoVxDQRfjFSwoMuhAPppnzMVaih
od2Ng8yz+N6nUMyNF4Xmb5xjgSKIXKidHs+wqRSLzGlaU63qhSjgb16mm2xo2sTPoSAb+y3sLn1R
Q3y8BGFOgONtxaDoysVZ1OqfS8IUJNJ5uQuxb4PealhzMdgmdXEixLGztCTBvgX76pDK8+sgUsIT
3+pEU8HvhJ0qLHEnJv3S595PuIXz8o7HKMPeUGF221MLXpLi9/BXKeglt9vmMqCtRF3cjiQ5UD0g
jE6byW1OOsH3dinlN24349mFaSLoye9Zuzn2dcOQtYO+bo5ANfmpVRaDP1ks40Wp5idv7yBGWvEc
8oKACHrjfGppLLPOEZR2SkexfDq3zzSC9UiRYj70GX+7mIFEkjWok8hh/AWnIHhV/L7CktYjKqLa
DEFAqPAjpKqfHLSI58MmJU9tcTQEHDPvc87+kJ+MNatGdXtbCO+6+Kyd3WEDdWrnE1zEst0+QDJW
vTuv0cyGFSV9f+YZ5QI1sfHY6h4CTfUqERLRyk4CN/m6wT+kxqaXH2y2c5zY2t0nUYi4C3g5FX+R
+HJ4UD6A9ZGQE4VIyWt0gwfMST5cVzboKfdvbxXE2g5ITtoLQLIXBF6hTJD/H3f+6HPG3B0fe+x8
cIwirYDlHLI7GixwM0B10UAuvGZ9urf6MuIVRas7Kg5V9UbsXLOdV9yNljxh6NXCYlNZvL7E7JOg
5EKNR4jCVcELoshgwsvdJDSGtt5mpAR3rvNIFRKDzbkNiOBWnVqbgSi/3iOXy/R/t5GMJkl9PMtj
9d8iNeeHNplWbDxBqd8mDmp1OKB3egtWv+pYf1aQ34jCyTtzU6TydKOHiu//UM2tQn9rmQkbDqPN
9dvgxN3zDx0E8vIrU7aTjbVdT/Pp8wwua4/k39qm/SHO4tKcdbzyPsZVztnHIIjJsYfOYesbz1I4
CJr0fmmwZgKlVoyPLed0fTCNhVPkgdwClfabNrMGiNtXHj8eulTmFGn3eY9aUngPiTOZzHJwndFN
wMaEP2HDw/ult7gC9PPhPr3cGR/qdxZ+yJ+FyqExxZwI1+mKosxo1F8+BnXXLIHyKsDFAjgbd5Ek
w61ehQbwk+pyLAIJBQopY8DaLiEjPLnkXcXRooNnfZSwCo0U9UO+YW6kHUSwFHTaHfhEjlMSqL2C
3jckUVpBBTT8tkBEmqOglfGqSC0jUIdUE8YVfhuewpMhT5DELJ/Ucxhw2fw+Dk9Hji5a2PxTDzl4
SBpFmKXNEn0+5+FOeluDW8CNGhpNH3CYCe35bpu6oHLDP9/G/XpS+w4m4nMFEouGL5NNTIW+qAJu
Ou++IFMbbQdOA4vmsMebvcU1iLf8s5q8MvNciksDKSzqRNDc/fOCDCNi2fp+Jpj9TIPIEfdoRxcL
cJ7PT20Whm+QbfEzDGAOgnbbM4oZRr2U06pyMvxTgwYAAXBCYALUewbr7hSmrGZKVLw7SThJBqjJ
LLZ2FOTjVyAPABZTRmYxmKH9Ut6+5Ofxj5/lgNwo8K4dOF6wj3G8vEP2xEzI1br/ruFmL3GgjZqJ
Ijwde08cD6fzQ9+G32JKEq2elrRsU98Sm8hpJ0j3PRx+NZoP6/EEwaCxd9qHok/4fuXYkvoM54WS
jO3QDb9aOZJe77Za28PvesJpx26KGuRlyc+Q0SQrflCvfJ+2vrg67kvtRD2zktiQUC1k7Z8hcBkd
MS9tiVX/LEUajPcR1FRz6MuqWZX2oyDDcszLPKkAQVkvcLO1IdwVgnapBcyGK0nLL/h6nqAblU/d
9OTeVKt9T7Pz2j3YBjg+bu16NjpIy2+J0mPTZiRPoU/iI2F3GN7GwSGz2DqZr2Rehn40PTA2BriB
5Z7tP1cxgiewG6Bm2QN97OvG70pw9H/waDSYd29I7hM2tCtx6ZI8HjRN1FcVJiTi2zscYVeY2zsZ
FZeyA4mHi2bmzYeinquj1NSoD3B2iLGUVz3JRrTYjKqM8JZWqJwKGYLghik7LF6gIdkg8jF6NyuN
AT93B9GpMUC9VawS0xaZLWe4zStxxUEksAPp8j6sruOFM+Z3lRFsDVHLMjyAHMd5MQCda+QmS/Jx
GmfaB6QoLsHMwtjjBkjnjV3rHqGgFWJb/SwJeyNUrXD3eqGOAuHHRyuQBKG+kcDZWRTnop4TIFpP
o4zgvCkbE+MY8ygmbxLQGsFe6Wb32DPo6vSXntGuviLAfZcF+UDwQ+LNjxCSY3VHS01U0p9TJPQS
som2CuVdtGJrGgO/Z2xkY7puGi9jA5qwo03OuHUn9LKtbl3ZD8Yu8zYS8i8N1bPMz1rrbpYxP4HG
wMr8bUAlreL3PKSeEpq8gjaIncq7h+roDjl3Oh/4DHsc0mfKJ/8sJf1F8tMU2kOn+dvLUr7ec1Oa
J2YM0RuGTkcL3/6W2o/PkZzXRdxryr8zxy5knsiK/BwSNLlNkaemFTzyhFC4/4f0UsEcPe4f97+b
LSU7THDht2X/mc8hqtrRTxzz1F+GpbptD+YuOSzXOMwx7KkclPV4dyYEozaX5gFDw1AkYpCsPprL
U4WYOX1UA9Z2vhw6NQs+UUfKKKVE6LenBruoZePABbkgeVFk8JXNL0bGz8JdCvs+5iwh+mo+CAE3
pRWRCYvKfQoLyjWDd1DgezlCG2gtOHAxDTmZRylhQfSr2aR7U+rWCH22B/PWVVXYsmMh/hv0oWfu
sd0knGVSv0ro6UaxNtnW7eY/4Y6wLfWiRIOSkr29hA2drI23DEVUBbEiHJpC0Gy0dGNPF9ACB2b+
x6m6yGFUJv5MR8ijlF2bn4BRNWfecSYEIMMBKlfP5SrfGIk9jd5GcN54PDRe3cvZedvbJcaRkJge
wU3GjKLQC/72rjjjTvpxVwCnBi6g+P8mAqHG+2rwuuljpPilSglKVx0F8cDqfzRUyxnptlOPo8aQ
+KVaFe1183hUNwhqtekWH57tCARJu9akNxrG+Dk8iU2i2ygCpqtp35aCR+ZSnV7/Bj+OtWK46lY2
rJVHmZUtWEqN1byFw8NiAmqBRI6lpoa97ID4JemS1gFJkQ0YpRbGsOo1UxAhH7st5BGS/xeGn/dW
NxHzWSF2Kb8c95Kl09n4AmN98CEEbfxdP6R0rJBn9wcQk7k4nNhFHsvyK8q9wHA/9fgE3fmHh7Hd
WDSVLzdE1YZ4oaiPP5ZNyhyIeTuNkUfCKDZF5J2erAdg2ibDQmsUwaWeblo0zd1KSLOP+Wh3jOKb
zZe1/jQzhS6LS74WjNMICaw+H1amowAyS9Oe19h2AGIYZg3xOAHYlBuw1/SnyKWn4I6YwgyrQiro
OhTYwfukexN8Aa2XMolXqJke4cqX1iDZF4i+Ck/jAgx9t8TqhnqKuyUrOPrqOYKZvaRoSqijItmi
7KxCHymeFFglVsitfUPfWZludfKmch+4RCKr94iMD/4k92pYn9gglLbUVktfoKcBQccU5+rX4r8i
Gd1sVDxABrxFHQrREisBe1o9XzWAgTnYHcK5m8acPaZsAuJF+ijntOEHTZgCLuuyrCLhYBn5Vcd8
kqYXsp/e4bKZemgit0AjtxuhPCUpOhfny4S7Q86RN53VcNs6COHwl6rSKBSbs+0aSXPLe+TERsNL
6GUHMe2y17WsJGaR9Vf5C6CqtnK4DPfz1aW6a7AfLxCvd6BLjcuz/sPAoA0XiLog6hTw9XkzhyEg
NvI3el5PCdUlZFqGWLw1o6Slvj5ED4JlwFrYTCqicz3XAjZrzlDnVvWo+FOiUrlIBVsVycyz+iRL
8AjE2kkxlw9xtonoBmusCvl4890ygZzabUOzazuE41qSni7YV6S1pVzVUu2x2LVYYQGg9bxc7S4J
3sQgCK89zlEDHYfvVJnxf3ZDyGtt10/h0/d05GGBlmh+jIWqllvwpMCU5b5mp5rrtX9ymnmQNzrh
1aVrdJd9XuTshiwceEObn9vixcb0lJoNr5xCZmWRw4atqWcCKrq7pzqWUTY3GWtbchZVGgSk9M8u
+oLiLp2vHeP8Kb/lcS2b5zeHib2aXtHQHapfaqzFxETYY4pE1UboBdblDeASsrF5g98zgaKiiXBu
hwOPEhfAfG+NcLdi+K6xMxDGmdCriTPasx0phFS/tATQSWNM8tIdtlZ8JuiEvImP915NxDSB42Ba
sw3fdWGZHT/qbwxilrJpV/xHvTwxAvwVQPpEmpwy7pMXmXJqWepYedJ1sKLze+9FPqJdIp668vdy
sW8ySMfCc4heseDEHt9k5JwqSY7Ux3godlcjeaBZ8wGSRsQLdHrZsSqth6Mru1gYJna0l74j5DFs
L1iWRpQm7DmRhiAY4lFqi4cg8jsv0sx1lqzNVhvlOxA43BUdNxE1QDrF6SWPTvN3MLadxnA6Hrrp
j3/bKl0PdYcZ8q9n+BtVC+8HDpBbllR23K6m5/JuOXWu8pdmMNBuuzacviyzhVsUC7yiWKQqsNGd
B1qpZeEGC9O0dPQFATMspjBO/maj+GPKg+lOoke6D0SHqQsOUQSbnfOffA/si+MStiKK4BUl4ORd
qcqdji8bazKNH7XU01+iM1Vk3YBpc1TZe+A4ODA/LfWWjtz0eIYkHT+VkwxPeUvP0Yx2/2NDTvxD
1qu7aRcTzE32cSoZQ0uOY5Sx1+ap63vDgevcxZNNegINot3yrB5HEBSkDSL1ppOY5cac9WPrd4ro
/nfO5aokLK7sOCiXgjD+We44VgqyUT0+8fsebis5S30ReKS/dR6B5Nd3t4aiTlE3HvAg/0sGq3sK
c75JlACdg2YToEkRsdAG8Rg3wbmROq4LsVYbO7Nxm0sRKNHmSs/DWvVtrsC4oMATc/10Onf//FNB
6rySIif0Ad0zE49FFwoxa5Fbr5Xq6nFzuQ6LPuDhZxOUpYrcfjYL39BZ8g5Emm6UIukcQUS7wL9x
jm1ONU8eA9mst1Ms4n2Tzzh2nTnZZ6Nwk3n7IYj136m0U44+wL3BBV2RAyjPs/yZ1rrsFIdXJFV2
zvkrUc4rWPqNh4U+2rrtr80967sSo8PhnFAbCFT71B0+qxmLhc6ABRbg+2xSJqOEsUhJfN7j6PLK
N9iqVmWHBuHEmIDy/wGEE0zdsd2/oEb0otP7W4vrf7k+65xpv4A0xhHE9TqoUo4Xyw+3Qlo5cza2
stmXDADIRDK9cE2/kthg+CWLI9ufnGi9QDmOcAxW0HE3WBWhuaXBphZLKaZYvw95bNIN0o6TElk1
xFOKd8i4wdAf+29vXE1Jrsp7S4YtUBGpkwSnTZ/esOWuHD4xCq+vmh4ES7/AaJLB+aFfxZ5FHGHl
w1/l7J20PKW56EGp7XM57QrRe4BXn7J3PngC7BDs4OjkkpVtVsE3rfBz7AKGB9WzRLq+OcI8z5bq
s/N3YIrZwKjzbFEVMkD9YubkXPDPOHTyZ3PyQo051hdUmWLptOF9Zs2w/+LlZ8oWz0wihMrfOVrT
+5nDheS/uxg1z0BK1sFNmIIwJi/9EocDXqPTTCCcmHCrG3zyQcbGeA3b/y/IZvWDxvlc636rFodd
eLBjHVT7DiO7ejCb7P0b0nOVWzeMn6jVOzxSieFbWqTosXwb4/0dfxqZ76iJAisIna5BZtxHsl7I
WmTdEGy11kV5yDfTPVJqkbVbBZp4Y+TPfkqm3ynZ0gn9LBvKZwtRup+kczMT/2F1TDQbeU6GkqPl
VqPScDEt3+NwpOfgYwP9MfE84gERQjAEtDWTpaeRkOXrB2F7cCErrsSwtSjJ3F+6e6nzNzs+ZKGC
wLF55cKRZQkLYnI1skwETGT1fxz+XKvevmGcCYo6i+zTiy+42PMkE/TPZHmW3DqN9MXnXIp9tnOJ
L5TiRkzEr4UY8J8mzhLYbIykQvpj1YPrkfVMMlBt3FzCNk6gLnTLTfTVcROjSgukUIbplKNqmp3N
hYi1nLQF/752gMZBxaWf/WULIvW+AdcPs46eOXVUISWJH8NC0mdIKAmAVfdIJGIIJkgE/CniGSCo
qs6xNgUDdjr3ksoTWvjEiulk18yQJP1nnoneu5I1bSCItxb+x/h8wrfHmePVwz33RFsW+dRorvhb
RAIsgl5TVpijCIa7Q2m7jSllHeoXtvI5ZmyfaSu+iZRL6mdBn05fbjj1ZHvJkzqxI1sqvCHwLxbl
USAiLORAo/IE0cqf3qvTxO0bDhXZTQ+AXbX9uPKyyRMZvSFQM2ocewaJGL3R2f7aIAeZq3znIjd+
OADdUwBxkfJlgGq8YmBpB04MUzQ8UIYvFy7bmXMyKTi5T1ccp2WSeLixR27c4CslwCkbc9x5q8xt
NeJ/cobibZ+sJa3Uam6ULQmAV1KhXUt4lW7KkghPSZ5o3fnf6yEhKHPc9MmDc+r/LyWPSLoYNdUe
vZTI4r+spcwW+QADR20UG161xySQ6L9x9Y5y8X6MVAXe/tZQTb0+FoGU0c1XgmfJAflJHR65u+J3
JsX/kIMZ0r8h4VqyqTpTN5S+1OsuodEES8OjurVSykK3qmcMgZmgSBK7RAACEQQHWnnk+x0rkloi
NVjOTp8fYNQ93NxPWlSMPJw7UyJtBtsoNnJ5FcfYi8T45xaHmiAvtHI2yQ8Qf2+N3ugcC+ObGqpV
h005TWeAqQHerHR2viXbagSaoyXUR9ods1E/fw0Sg73SzspkGCdkByjxU+PP/lRaglBSBNRvTq3X
z6tQvyFktSliLxmXHMrX6oip2m99Vf/1aG79HMkDn2IupG2ddEztFwlnN3Gvcm4vHtS6r/47osra
BK1Bh81nf2z0Ad8UordpE/a/ZYXAP53XWSHRNAOQTATMnaPgosfrDg13FCcjPTn6VdpvTkx1LTQf
CjYFWafH4wgeBleoIG+vMXzsgiUYlilDkKIaGLKlCJdaIwP0LDJKRVBb/DEYyOuu5ErsSBHCItUO
txS8pesQK9T79zaBc1u+LQxfkXnhUVy5hg+GxLrK0ShmELPXRxIPmAarUpkxVNH71UdGWHb44zQk
EwNcVVtSoGB6dXDym2AlytRIoSKYbrmeTOaUQO40c/Vr88VyZ5rforzpy1HkXnkPHcND1FwcgP/q
1a6xX/eKMCB0gsDWUa4ecd5+aN9J9HILEI2RlR0wTdq78eElqe6XVRipVynDs+kjzmEgd7QIVh+g
+SZYXsZFgv0bP4OuhGfk14xQSoZK7rZi2SFkONY/QskGEzAnrfiudPuT1oXTRBsWMQQ0OtizKGm9
ENxRKzg6locfIvBaNnw66eVvuIM2c02yHYpdk5eYn17pyD7BVIAoWcEBzbBPNai7+YAVHJ3NFVOs
97mKHiynkv2WbO24QruDYdwjUmMj8zeNX2qR+igWZCcsUEkiDeP3CC8HTzCgs0/j4JidcWqJz9D0
oMJcmy3RRrON7hCdMUunQWDJ3/AMk1hN7z04m6SvhkJn8jp/fnNAuC3uaveTuAzy19Al9O5DE4t8
5irBrgkEIemE9rnqYPj2XhTbxvqYWcdKRhLryEEalf/aC6Q72NMGhevLNtApO+bzT7rZr62NMpbT
D/Fp6xuaHcvd0kdRzqR0xFhDM/win3Bm8gBfKnp3MpoxNaJARHcQbJHF54/g7Onm+5MGG9aN99ki
FTuhI4kSDcU0xcU3KVSJsoLFnSj+HWJdPkUcdK5Td6ZkJZ/uEhHRED+KilahRfuhGyHtzTsZl6Xy
6NVCqz0jdtz+j4Ui4C39ow1n9aGrTTl4QSKeJ6gECJbjc3QcTCh6GqP6f6FTHlntkikkDOz3IxMp
o+7Z7y8aWXtZCNlIIaPgENH18k6GemZaNNLBm8b1PxJtn8dyT6e4dI1sOu4GaXc0bj8YWJDLCz1t
MjWE56YnG/UYJsVxTaKDb8rPhU+rePLOVRC6/yX+tObRrSXZFO4cJa2qTv5Iw79fj4u+kHRGuQkz
XdejQpIa8BKdStIBjbyMLiHNWmSKJTBOEwZEiDC+resUmk//bRURLuMzsRgs+CfNrGcEC0k8eDNl
JCumqFl+8vcxEnFl8xgDrZGkeNA0EaUyDwH4jWskAIcPhmIEW+TaBNgpiHXHmePWL98BAIvZXzyK
+o1UFPCMFrsDO1woXI7atKp/qyHUrCacW4sI0nkf2BKcXPrsq3ZHMpTSNK0sp7PFR8rqLVPIqX/5
OKncqzBnAgBN81+w394EgXQ/pNjECVPo657HzdpfiT/810/tioP8wrwcQLRX4DJ39FqybcpEij1o
2XUfCGiuLyFSoNYrKDstHhFf33MZZue/v9Yr8Xpqtk29Kcae1vJw78TU9v+g324q0gUrYH7HMMko
debOogyyiyV3vgyuOT7Q5hDtoy2p1Pfbl7pOAZrI5Mof9NFZM7xJO0Edoe/ZwBnyEgL+FR55R+b1
+xknVln6NdRCFULDQIcowPqb8XKiG0FAau8pRWyez9/v+/gy1AV8ISWz8ja0puXKsosf8/tzRS+U
oAd7dCUz8xIe6FEbYtYlnQsq52zfkrv4ju7PcGrJi/H8zZC/z+wlY4QjcTHZt6fnv5ytBECjy7t9
xPXSchxQRC7McUzirwzT6mKM/p1k5bqgdyN/XyHHjPfXkveysfEvSwe9jmQIucgTnPZhYksqMlie
XzS0FBiTbfMP+eUzZYPKA5zE+mib+FAUJas0HRqrleq6mEHRkZ2tzf/5WEPRD1Vl9FosuJTCLbbG
MTZfCsycDRWQYBWlcM0vgiAUoeuypdP4vO3j+PPF9r4RRp0YAwdYYM+pgH4lDaJH3EU7hh+V/jHB
YHxUdEyrduql0YSK05jc8Ie/HDW18uO3QLtw5T801uB9u2PPFje/+TwtdxDf8bPTp3XZmhngKg80
UmShsJ/QL7xdofVkmTx0PM2fcBG5s74FjhmClyDWakFDRgj0zv94vQr/Ge+au59Hyc9fCkghiWEh
UBlqOYYpZXtFGEmh/jOwPV4PaOqORMQoWQOZ+lvshPKYOoNuMwY5fZp4Hdamx8WzJvGTr7by597y
DcdKS9G8kysCMVAwz+nl68jjiIb8Cxy+1KjfWGgk42SqnbwPZmn9KdxNxwKfZjNo+QnNsFef5piB
057FmFZkgBTD6wdMDGaAeGep1jdRbm6vP4GLqBUNurS0dL1nm12CLDtNJ9zZIlT1KJWEE6i6ZfJW
DLAS5Zs4pisdeqD3Bz1q1pGzN70BJNg6JLv/4EgB/OpV9iCUiU5xH6thF+mu7J+Za38aphGu5vDL
GxMa4Gcu/zBw6gTfLjQTOHyIDwD3SWBX0Y9JK1k85ZHC1icFHT74YMP6KYVhvr7pI/A2Dqwx31JO
MdRI6X46IjbeFeG7+4ZTy/NHrntOZKiSghjpf0XTFfJHcT6ps95MHGY29vk6OEmaYqVL2MJVqI2h
fYWSib20JqwtYuEku/auZsP+2z+uOStBFJ4Y+HTxusZ14qBG44jqqgWUeHa2DAc7gBNPAzabjvdj
7tBZ1JxtGlIy3oTmoJDqg+Jp7qxBZm+PjaygyLIQV3on5BKFUSLi06gGgB9STuDmWUf+vbvrfnW8
weWERnBaRbijbDaNmY/fnxyH20sJa0IVRa5dBKTIHm+L9TNBx7aeWqyQTMballPGzdATjrDmU4fV
XrcuVPcmFmfAoGnAec2d4ARET/jfFpxjAz+ZQP8ZnJ5di63qrLOAlZ7og8AzwTFS51CbelizvbZ7
Zj6xmg0JdN4hmW5MFw038SK71At/0j1uakovzgumQDukBzF2+mexKm203cwdw1ZD4KdbX1/vDAbu
6BwMHAc4yxREGyK8e4IhreMpjT1QHWiPtd2XDYWK/JoiJYkwTvhxaHPllgUVjAfGzVlZ7e1J0zUH
xhr9jHMCM8tB2/ZAL0g9PoOM6GPSLnskGxV+w8sujvXzLKjUiradXdm2Ocj/9bsXUxxSrtNWEEsT
xV2IB13bKPfVMA1cxpUD2gcTg5HRCjQm/Z3sUquVCqeiFHjK5FASf9ZwF8ILIhQ0zWig+nmK15fR
WQLHQjKxHdfouzcQJglCUusNt+FIoJ0gV7VEBQfEsDQeIeKE4zHJXjl8cYYCUM3hjV8Z4FdwkOoz
naF2hjDHo+yz2Yn84usGy14ywqdZrIXYXO7kGR5KZzXmRrC14980LwBsr4OLemdg2u8n58RJx7+d
dcdPC0F4UpdLHDDvPnVl/eKOxX2enoOZV2jkyrujeujWMtE6dgtJOIDlD0d9rehInjuQwCIqz6Wi
t75YyjglN0iZwAV6tjyyQ7HU1WWqMNQDUwy5c9BavktHs4CEPGM9yz/B2K0Eyo/vSVTgHZ8rNU2R
TDr2HfjoguCLUlbcCcjeyU6ab22L1ZNlwh6Pyche2vhyOQjmiTw7aTyZZ2pxudTJ0k4JyIKjJlXh
wWARfEBzqqPGDnXNCgjva6M6JyQdHQKXV9nUo4cIGwUTXxdnh+jUbFeT5WrimP0vXs4A4IPFp6jj
k909TEV+uJxZ4O/pkQNqxsnfM3JMXQM+JMcPnieYkkub0fIlewCcMwW41qwdNDDKYVHH6k4IFF9M
EaFd0SLMxK0RQONMoU3d4/9/qKqafm0YcN0SoVz4Xlqapwmmsge7RjSmKLinwHjs4lpRx9Bao73z
r0JTs4pyb1+bEluzYmidn0hCnPiuivy2SSzeQNw1odRe5Xjo/BWYs1OVxiWwNQw/ibiQd+ky6Ji0
NuQ6WA7wV3BClVsaGPh07xhjocMB1zC3zfj9kiiEB6y6zuN+ZLi9qc7b/Decle7Zg59v4H2jD//7
SsIb3+6hE8OeSNIaG1drzPoesykqRJLOGaiZFdj5DMb47qCfLao/pAqYu7I=
`pragma protect end_protected
