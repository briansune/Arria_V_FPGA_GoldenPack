// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FwO6BXB6ZzazXEj7IBVw7JsrsdC/jV1BrY/Jdp1SK9dm+06pOZ9mAnkHegLetif1
DwfPDFoa1jrjWmgPa8riOHPbRUD/v71GpbWDYdO7sMU+WoM0dy++8inHG0QyW+gt
rXAoYv0w0Sdd2oxKtGWZoNIdbuPSUqWAEgwlN/qjDdA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
XDZgphX5RxV20I03FUSuTk1R+qxjWqpNAQqaMeiYOAFhfeiSRXNesxGKT9OfX9xV
S3KMJqKZImgqlCpyU8VFFj5JxOHmE+BNVnbm9cCp8Vm4L3iNWvjZZeatHJpk0SKo
fefoc6x564B64yLCcyfhwdhfdeHOxYdhsgemf+1KyxuGNjOe1gShF/+o47OejtKh
KLviaOwoNtSjpdKQyJ20fHeWQ9Iam9gWDm09bGGjZeIHX3ALZA2V3I7Y5WcXBBiv
HUySwBpDXqj27mfKNVVUXFqeX6aUUqhhQrA527vH74Z+57kjIML4eesKtKHf01fi
Cv089TuUbXW7AqiAPz4hIDicyNZasqG0kEcPQBGWCOm8YS4EuPZtj8OejaKttnAe
W0S6p39dg5yIMHhm5nriyrOG4fgjf2JrspE8EIWuVrUJ1sXFHB5kvVv/I6aigshF
ElLdPfRkXncA4LjNXHm0LAGOWxMcxCIruR1Db5NB5VI1TfPwULYtjJaotIrkdCpD
hoVprb6Pbm6kugiKeuywTS7EmjqeT0rnGtUkyieymLLziuwbXwpfuFFeFjoOOYEz
T5lSoynpTieOck+3v6b1uU2Jrgyn3GUq4dg9FRnB92yw88HdPJJEKVkEKYMVKgfQ
zKx+nBW/AHFgFf7Piya+Muv1IPBfafaCt3hOhJJVNSFbJStNVY1I7Ry/9aQ5h6j+
D4dn3xVaO7rlnjCh+kEfrULgLBZjBGOURTG2Jjcy7Murx0XGls19NNvQPKOdgXi/
brBINa0D7LOKL0p/TaNSe0QvB2kvHi+d20i8O6WagXYUFbVrX5MF+O1UQAYK51kG
uJYTpzcWahP7ebt6BCnSwDoC/uy4CgjnM51/4qfnwiRgMROL7Kkk+HjO3GHxicvL
M0Nmf5Jf/gtYWFQTonfxqlQVvarP84qYeRpQRgVJagqRHMrSR/tcmUUPmtgqxeKT
K49yLyUxwsjvvn82cwYb9MrLwcltu2yuia9ois0K2hZF8ELEbomk7gJU0scan9u/
IUnt1ond/TAfZCaS1lZTbxySE6ZPytTjgdP2ttg5sybSwOPRRbR+uhfSMLHVLzQW
R0LgHPfM/OAoaY8M7eYLnZk9GuM/IXg+ft2EcgH+mirZIi1uByCus77Mp7eMaY0o
KYc/ZwkZHwjo+6VTP/qhiR1riMdEx6mOgs0Z6zVNnK75ZQajJXrT8u78IBse3esA
/jC9kyoVIxqwvca0EQGMe2RD3sTamCeUVLD80l9FNxEVJDlARwQjJYKtJ7zMbpgT
XmzjdztDCf4IQFYdOPQmDQUdZOxQqhVmdfMc+AkzQ/llzCSXRVR/s5DBp1Bva5ie
LMr0XZ3b3xyM8g/nF0JLsALi5ex0Glh5WpBzsgSldAN3+NQbBmvu3uoG1lLjbFhV
yu+z45t2Fh9pST3WkMzK6RcLR3l7Wj5fvCFBnjtD1jTya4fZrIJosjWGepRtvStH
8HIUSjo8A7oikZgUb0X8gNlqTSMMrfjcjUW3t4PHq+LA50s84/y6bSRcaO2Twl5E
vWdJiIQtjQqEKdbPIlvZoPf6nIRn+LgU4gbUDsXzksJOKg1jlGdyKKfWuVYX2St8
pZWRZiRDwmSyGL97kGRInjY4TgaUV1iDOrNfhuPTc/x8bCustsTsCS2ep50DIIF2
RbkOt//9K/p/dxT2nIJ0vnk9AunafGVhFRaGc2qwyNAOf/est70CL0GE4a6vnQPN
wAN1IcUXUP+N9ntdiDHAMgPviaDrXYTZApYmhRWgA1lfOohhXPlL2b3GSLbSUoV/
WJskutAoMiBu5lFHnK1jwRwemiHtrN1e85OkgPHrNdg4snHOeUn3HI9WErAosnpm
yzKix7qmV2qh+AwOlCgDxh2tle3hTiEWVHDOUccev/1O5QrbaxZNjfkNKg2p/0Ua
S89JgIa5ISMx7MXmHvHJYLRFwubMNdzMMpzip6l2/ICf9WMOY/K2NvI1ueAuu0av
rcQv25qvjD2Cs3RKFu/Mevekcl9uuq10+tHWWYPzQatZfynjTQcymRa5Npa7bTTS
IhuFYA7aQQ6ToEWfLaVhmIy1plsJx38w93QuM0y+3Vrcms60AHcmuEC7jHpOs31z
SogaNYAHjiCDoDeYHNFkh6fjug/FMwUcXZb8dZtGylFX2hqYgU9H0hnzvgxEwYTF
1/IYCzzu9QLOpXos86kutwOShRXejKlxHATS8nvmsyyUNokKK313HyDKmQVLy0ow
LGlhfn+EhNJyDj+g7OkOHV0hlxYJw7ueIEnnfx5CA1FARoPCNf46wVk8M+7EJInZ
XfigrZamJ0HgDUqlNhx0VG/4TKMBXwr5LlBlwa7gkBOcW7posOXF2w65dyG7P37J
lJv7+A9dZeyvre5AiFlxZuQJWQ2Y4YwP4NwTdLjbURgFFCozh6BC56k7rgqWo2Ca
/ddVQ+r6a3R6V7rq72QW7FFydQeYfUijzMN7HF5ht97ZUZxMEYVfSP5cI9V1eIzE
gL/uoN8UcF4Z8oNrmK4QI82yGECw3fjjWooOEfDBMPRjxmEmNygxvHeNOlej1C1P
DpKu0DaKGjCHt+Wi3NEOiv7PJFJd1OK5hvK7Ra4QNt9tldmgSTKfdLGt4Pa+avfi
xwOZRvi7Qdd+fPM+5HWO/HX8Dl3fXkUzXPZeofRqkD+rBJQps7EDknC9C69S0BE3
vmL7tnCNfpQzOFFZ4qypv9qZab+GpdTinefPLrTbL6nfBJRgLF3+h+LmmVytGLLB
3boerxFlN83GcqVrDnrA9GNU910YQMQyzu3PXWe6IZJbnmKF558WPInibb/nLFZg
Qi+rLVy3Z3p/6G3GQ5JciPqJvsDJW78mQV7X8lT/0hAUZ25fCe602xWaMcZML/rj
jtAEhICon/ExXsVuaVAVLCNWV0fUYB24KzX0u7SkJ9dcMZzRS6WKWD3LMZJVNU0v
FMW2tGRx1WjiEbvrEsu4Q/FfqsRRod4DeAX5363M4+uLpE4UZB/Ue3pa992yI4Vu
8kTTv8VjQnscWZH8v/PGkbzYng4mV4Ihas/TnjRixlM3euNdaPWR/0HRNvr54ibp
X8UfHSitWFrLnEVuLDnhqhhQ1q4ae/g74aMogE9Z332xMTPD66IVM80EO9/XlV2g
4AW523dfwaC/c4OUzTzQGZ83FRqM8GgeKa7qQyxtFe+HN0mgjTvZRNqOllJ8WVX0
OMuxQA0FNiVl+IODmQhTu2OH5F2GOGvYCNfW+//wBacQLijYF01ROr/fHe87ZSvG
NKOSvwbd4fl+483fW7DtSpq32Cwu5ZEo8/Bglx4hilTfTVJZlUTxrjstNf3LG9YP
1Bbk+/V7R2khJTKZhMpgIUcw49lZi6jjgppyxn/SY5Htu8ScQjmWTgGNak0GY1yl
tI6McjAQdFqL4Mqxy01ixFf9YTct3cNru92FqwXkYOGMPHcjDfcFM/OWkT96bv/S
tTP7GMCnAe8wxG0RS74rjJSYy3RyCtvR+s41tOibeAEjrg2orOCLWbXvGBYLtjy5
W5+ZoixuvoMxzgSu8Wc92hAKSxG9XqQAyAscwS4PfHo/UeoSNcPsZpX90vYrf1jp
Eg1twET/BQavGb0DvQS40TosvOvueBu9Xgx7bTrsqteSJXFOp/gEZm7+jZY3yV5W
EjGdelnNrvOwuhC1B9qRDfvmPUB4/O1gPL9bRWjhS4lJvjVqMsnQ9RQNvYX52o7l
JtPcW5EXmc88l/yqwYHISlX5GV4Vk87+u55YrY1hW9QmQAq79JtOpMZVLd28PHx8
ZtjKGn8d9LROlYYXldf6BL80Keyhd2QJD8FmAZFq5VBikQCxgfvsfMcYNLNf/BoY
LrLLNJDL49ZkMb8m2b14SWU98WNzmVicJDb5fJGzUS+a95BdXptB8+y3NMYEmc+x
DFCjS+HlPrywLuMvUSD1U8hsZqp0NCw41LYg8SMSfn9orN48wDrEOW/1dmpQzgq+
R25xzC5a82D1wHLatAQCW3Mj680/1ey0eM4WB20SAbqxn2x2YPWWmucYRadwJ9gS
Hb2CtO7HBavwj/3BduOlXBVfwocPt7FJb+ygkRWKW+z8ucUdSAzcWj6B69Ek4m57
QCHDcGTUHnKIAgLpmyyqBQQFPPv4DgJM1di1xA0IytyLGtbXNPyUJ5j1W2FGgcZZ
QukS71520sqsW+78v4Iw3T874Z05zBqmxVrRSqdv+CDZhoxjoJPdKYBbngGHh7qW
Q6mKfz5UuViOqiN0JJrzCVNHp0PH4WLH2YLKhBdwWv4KiF8s0OuDL2Wtgj5mtQug
cC+Ohuo2/lNQ0nDrxhLz/1WlOTH/TPJxtVyU2Xy/TAq3gnwdT4Yeu76ShApGpuck
k3vfD6kE7TJvNUGmrQkI4WUd7OMrmIDPgS8BGw3KKbSNdu9oBnfSokmSOcljNPKY
hY4VE1daM9GhEC0fyrtliKzLNY0PrzRwSOIKVhyhoUd/0SuyyOMDvivnGEmG6meM
jlSc3s7iDxBC/CGbglV+kFVBEJwin3XV92vGwQLAiKfg7NlEimmZaIf5WRcApa3m
EIikkhufQc1utF+/7Ao1/jO7lx04MDPSOa+DHlgiSCMCwYN3JiGcgvseaXA06h0c
IR2+emVh8ZRroX5nPJG/bbgry1/mHyZldJBGrPB6tpPuaSdQ4IlCc+D7VCW1cTqX
zmOlIEy1JaC2/gCeb09FiDDDmr0RgLMGaK1n+CqRZEQfi3zx3nlGfprIEzD22Or5
feOBuH6oxRav04kBKr26YazhiOMc8FFBZonDazxIi9oBiRYLi+91bZ4FcE3uvODT
OOTXyHIBhDpLjeucO2D76bhIY5C3LS5dnoyNf7j2HNiGRcO0wnVn75I0wCycmiOJ
kiqv4RZ/i1VOgVLzVXmS8PpfrHjwNBeHK8RxOd3PjLUF1BEhPMvRUQHQzKNGDcA+
zXYoAWc/wF31TZRYqv9LdRYkwFBruPuZizG/eWapBK/ussEZely7zS4t1XLTHbA3
E47tuM6HEM+vvFPz3mrC5E3n1lNA+cILeqtCaetBaybHlVXBFF3ISx50Kdl6q4XJ
9nhEGRbTXOqI5IgmH1/XZ3bA+B3v36MtzNkYRzmvqJ75qxCdiMjxnLHQbUtE0PAk
j0R7NAXe2QlMpnlXJOdIGGcKdWnkLAt+XlLih7Lzy3iV29X0fm9FFNMpXtxOjFZI
5fVGGP3YMZVl6KsX2qFCStAEL1ObAJ1PGC9G6+IQ47ZQ7QPi7w2OIezpTbWwQ4mz
tLzQdjjYAfKagKYnbwXJl4N31goq3mIHd/QQew3d+IUNyBhsLACeO43ILn2pSDfF
AvnLEofTP82tomR0EqKgtb/l22tnAUNaCLkphTvXPES8fAO7oAvcv+pqm1QNdb6H
Egz0Gb3c7YYAH/jv63p8+h6MGpmic8xJU4b5esp/DPZCOMa+QVhQhRDSXp0qLhLv
AyOXb3/pSu+FpPSEz130hM1lE2Mb1dmrsegdxcFqVMhuccFP8Px3sW9xsf6Dl0+H
3Zg/zsBnAVoh1tii3Bueej2VGrJna0VVO8N5V/Fevpajr6vWncACrqKHmkBWSIqa
Y5dKGj4omWhGXe5bU1TB5yWhdvh7tR8hsfqMhO6dSh7ZHN/i441QmQiJ8BEb4YYf
CnVRBLBPOgbV7Eas881IDiq3kTpuBPgg03ktugFEYCC1TeN0CrPYZYpx3eN/XhUz
lc+Lk7TWpwAyNu6CQcRw7vmAfpT5agqo+XGvlcZNDu7rbqLeomBNwDv2WeV4EBjC
V0MxuX1ukTy/QM9SO+WjBYH7wnG3+34xI9p0NX+pQ811dgMyaO+bxoUnHBrRt51Q
sACGUdVJB8B+427t+69bUFExfvwlMdbJeCxK9t3uI0U2NsLb+0bTN4WVXh8+EWJR
gGbqlDqwI4Da3QSs501oe0exXnfgJwExIkeTl9egy2NpNKTxAflhYVwHHuhkmUWX
m/YRnvuMdxNjmXPdsft8Rut04/1FkKFc8SUv/YTIzFJVGjrgmB4TzH6z27V6KnVu
IF9eobRT5rAPs6WMXApbw+kkqkJLmEfTYACafPIzID3+nilQ7OhQA++gAEb3TeHR
7gWTIZB3rkcHVTHOUE6QzdIHUJ5P/GZEFGxkhrgDpLracTeGB1bB1aPdhE3HmbFN
/xxYjIpNskwcx7TTIuWukF4saJdThhjY7SL8togQmQKnj6yHKbS3ktLTtglK8/Zn
Xty9T+GbZ6qTPxSioyYjLW52J6wl6gp8lhjKquj8tYy8eVH8gZpAaR1e2MP+44E7
/0WMJimtaIS8CnTAnT9fEK8i8WWiXbtPmV5wzqHdLYq3qfWki5abjl78WZOwJv2t
QY+dUfpHomtgk30WPzgHvLGPTsUYpurWWUKcNNiOzTSzGF8JiXNdWW+AcMONTy5U
2hwbALadafbiKE63fgNu7se2uw/SuwxPtdA06rraIB6/dVoB4wX0OVeZPSqHwpNs
YBcDpGpWAwU7OAD0KfJDKwKATPbHoAg4TLWfGnvumo6qM0fFT7ApY/2QHij8np8z
8C+/vovV8z6F8Sxt6IPYMzp6YE/PUkJOjBFdhpj2pIRPc9Ih8buqJgCKhrJFEUs9
L8w7TaVo+nPusDKstZowl0PZOiYovOXrf4mvNYnSkZGyv4pZmh997ceU9xM+1+6M
yXdvFV0bZogd5EYmchq3t78b0gsB65nyy/9MZqikJbt3UwL5Lo8PkOD8gCmp8XuI
3vf/zonyyWE2GyEOm1OqiDzFyIWkvxV2ZGdb8zC3ihjLklc2h6hv0iN9R6R/lbCX
yJ1WSCqexj7FcPG4pPNhnE+OR9hfy+IDWrN21sPY7qxactEWj987TLECUOOe7D5T
WUidt9zJ7xfIuhoi4OqfjDHUZElS3IUWRwx59JfCUAlkd58erpTWyOlLvcJAftCQ
auo90LRrQZizv4z0QhgVDii5Wak9foFD+Bq21nDbxykypB++YDp0366jUBh8lDvc
06gQvOfDGfgmS4NlRhfY7ich9Xufn9fICxHu7Q6zqASp6u1lcqe7tZ2rheyX2MkV
btXx6EYr83su29JN7yJ5exwW5Z14Bx5HHc3o5ENxD3bPRMexfhou3M9y+gpW1RBw
E3srAVekmyWtaEdaxHt12mQiDrwxwr/QQ3B22nVvHE6tPWa0todhbEB0cnAKt1Ki
SGAMilnaSjWDfxStInm0Qlo+NwQSj8ZmQadJPdrGwREoT0+kGiylIlHAoXYt1yMn
7+NX7aJkU3LdyNb5QH6/R/e+AcNx9z3WCcwiDiWPq8r/tpxi1GHIPsY2+DweC+vN
feMQJrW/lR9hyp50ovU0egsU/3fg9aR2SwbUWJ8Lr9YcCSRp2RLhd7LZRfdDOHyn
1MB+K6K2WCpHxTglODPS9Xo0yXkK6WP6CqIEKiIeRTBadGvGTOP+Uiu8Anb8V2hB
TlNIePtAYCa4EnH6yYosqkkXwgwMajLkcgcAHTIzDhGoJmeGC/BW4AAa0NK9kOB2
HoHSRo+XyLZm0LnVR5hj2gaMjKqv2qoK6s3563NWA8vrVPtnFnZAKxEBz9nPVjDz
1rdOaaoYU2y0JD9cRluNg9rHOyqrvxqd1tGtdOuR+uBo1dA1yNIngyIQfDCkknLZ
uycPcNzi7sAn1jmI/LEh1JHjwM70aTtqpU6KmEGedLk6dM5crkaKhBgL6amKRj1k
8RtOY6NnQgxhVE4P1ddhxw==
`pragma protect end_protected
