// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:21 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qVJ0IqCT0XsLqEmznlyg9WN5e9xuRXCBr+ZYgpyECdGSwTe+iisHVEQbPaVA/Wjr
G821Aht0kGaDlp+cVCLT1OLGLf5QtCGHyFM0DKnz7cOwDHhrE/gfQ3AhqOuP3Ti7
aXwsp0EeqlZMIZNxBY7iX8jDmVHS8iKBOX//J6N8onA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104688)
/DYNnVkjxrSYyeqjxgCIXEYXp5vEgFIaShhJO7zRyXnbgXq9DNf0Nd8i7U/2CxIp
T+NqLwQeFi1yCsT5LREdGw0HWEocJLEtptNmyZGO2TAkvb6NdsN3lunXTYVlq/jn
K4wMhR54jJ6EdPvq1x+0X0UnM+6szZOeVEvn1JsBR64fd6ytrjGIiWrQ3EWd9O1j
ALo8rm++Tq9HzyuV8dAXiRE+m/IMGCjhwFcgc5Mho5B7EX37WK38JMyKuBq7jcZp
JFJcfxaiZn9ebvmBWdPMY6pONBdOj1lsjm+3nk/bjj/oMs+rbfmPs23SSilft4CO
e8dLQ8f3Alf00jvxQ9nCuIIOl9Kb5SKWpUKOG0Mg91GmWslogvQu/e6ARfnSfpu1
zBaDaWN/AXEUhfyQFV4LFNWGjdIuSA5F6+U2vo5xRxlFelwRbEKvGXgyIkIFcUn+
npe6V5M+rNH5C52P2VwJ6FIjhLQS1rJP+/lfB+Ubj/oddxQInEF1tMTZKxY3MX5d
YZKEcsRLmluB+fJwZyuMppXfTxRQC8hDgCcDjghGGKnr4GCylCOTYRwFM/b764ZF
BtraSVJUmZQZRK8cK+/YIllZnx4YVRQk+OAd6M8jakrP6nzHXwSq/8Ue59RuYzCi
7QeWEDTR4oUvGqwxT8HeiPUXWYXBDnTwqrSzSA6qUdtkFb/m2OcXKf0MEXj8RRMR
f+KaRV7z8ddfqP+53pMX7pOgw7L3cdd86dlXLwo9vQXdDlmeXiJrR3GwYgHcOcDK
BR1bgu1ARfQlBVWdjN5MmjNRCqEcl4sKRKuAB15zrGiPxYA/1vezx2tbfbjFrEcA
moix+bG1ix3RJLWcNEB9UsFb5hgh4bKu74FSJJCm+d5yXW1fQ34nOGLreXIU9V4p
POxuLs1tNoEpHw1qX1rKhPz2Jui9l/erBJgkwJImF+JOoINPqTPZ6jePqR8qz8Sl
LNAN94vqu9NVI6wP+rQz+//LHVzjmxBSYM80HuAgXUYw/vI4E4I/gsLP/sDYltwm
JgcwRnOv6ZkggfMuOhMXhGGNQssW0akwPLwBP2q/GgsZsfZyrfv5Ymf1dfZUuB2J
umgELjLqT8iTwrGNNkOD2/hhnh4yLLpeN4EkK9o9JAtl9sdtEE7bDBmZpn5HG9GJ
GHcRMtw7OpJhNcBikWSFLSdTSa0P3ByflGxHIREqKjskiNhP6T5wh2dKv4SAyYSn
jKhEFFLYqAOC+uFsdvC7aPf6pF4geKek849IP9oN1poyDzkcdjOK/d5vi/4Uz0An
yGV8IyIUn7wpzB3iVd+nAdlaZmwMtpyS9DnAZhRN6EDc+A3uF69lfAbqj2wQY3SU
pCp41QvxMoSRGYv7KYS7HlToS48mN/WVM0nnH/qoCC62Ic8fJnPdOQhwJQSCAHEw
v+bpTikWWwO/jIkBTuvpDaJji55VjbyWgx/Bw3XIUivkpL6okRBV1F9cVqVvX5/r
mxXyj3sAd0cU2Hs4o7n/iWE14OtXMIQ+ceRBKP4cQKuIjKNPf/56XsYt888cQWFX
FjWwjTZNq6pJH9+4n1pAAZvOCJvQO7W6DefUor9GLizJCf4lrCFecQdmd/lH8Aw3
EHOddyd9CMTnhVFATMUC2C4wAkQJ1lezF6SAgjnE5gRWFdp+urEbtbafHDp4Fu0p
mnacbd4zHx7Xsrn9uxFRQVeDYxrqGXPxt7g9CP57CrEW05tRSlFPSL57tonEtcTe
2ctPQbmYaJNEDGWYa3tJgk91SvPRJdZ+qGs8CflFXvc/V/5zVUm9TDcKZrc2GWo4
IMpQB/M9KyPunz3f0SUdJed08E6OztvuMsIYAjdUJ0iFqE5VW6lC+fyUHQAEl0hY
9Sih+Q0gOcoIrUWOsOW+cfDdfvHyTvPKbc61ar29FRAAP496ndyMrN7K2huk7CLl
7nDY57t7EwW65RBQW7Xw7U2MsKGnY+GPQGCC9UlYD2ICFalvGWSC23BwP4NZ/Okm
LTYauVDAre6QDoXaqvHkD8/CHAKdaxOse7UEa70RyS6z3zjRMxZtXL/tXnksdOjP
FYcNbfWF6cRs10UcE5dT+KDW2IWFVEpCFO5axOF4S8fZQ1RjR/4IDIvuuPR3cfyx
nXRdKes9Mp/ZorqOhPApe3uQgR7z6s50YNm12jzTh53GXhgO6qskrEzq3IUVGB7b
FLj3h6pT4vqt9SEGxxJh242UvvLSKF2zfOGfGaU0O63wpIUlRwFPFhoQZnVWiI6b
hjqrKJRYmfy0XUM3cAsQvqqwEK3zYKnqkuVXTxVGapta4OXzC61LNkrFVqWioq6J
TkJmUDiWfVvE1I4ch09pKx4zPVskKBOLOiJmyTByFcxAZkk5nfF4c0KB3EP0xOhL
xXRxmXaARfdPjwaDgGk/dq4xj5Svl3is+bT91z13qWjxP4YPisnDojR7qV4DpWv6
DQC4hwYQ6niM4leiE8SRdnM3Thh4LJwq9PQwYZaBnQpSpcB7nV2p9EMyT/YKn/7z
hka3QHpq9mYlPsTO8Jmuw8nX49KHz0xZmidAIZ3MTp8kf9NjfKptF3RUL4O5qPam
ndqElwrBcX/BDgwqIUbF6eIzTbi4jKsT6AoBTRA6crK4cl++WIyngeqU6uSKWE6q
5EDGqNZkkSwBAVeCjQJL5vR5p0f2PqmXqN4/eaRO7QQWNbP3Oq83RxH89HCJevPW
emEX/FHOYRXObUctBce6aV5bh47s0QulCFSN0u9FlbCiXXI+ghfILtKsXh1UIPk/
99lUMglBJkUDkWsS1ONG0kHsLNBakFgBjD46vPTN+CNgau2LJD9qaDXT5QTQ/7JO
06dTphjou9+5/FsH3EFsm9jBics2yxJ9JFHpRqs4rbdpZtMJrq3RtiSnwXQDywRj
YsHcuOBajg1T9Xf4STat0fvfTv8e2G2Mt7xMYkZLxHvyVDkdOKxBXazFMQ71iZOJ
WO4THnfVQsPR3z1A0LTpSqqJtzQnBHcgwrszqbnpY1lQvHng11i0RwNjwEzGfzqA
HHkXCtdAEP8+ERfxOhZ725fhzavVSLqFOBu23Mz0W/6agIsevxooePLZYLnC+y1u
qxEBE+eWm0hP3oaXAk+yEd6hgLV8Pe5LNzBYxjZbfJvOFORRL/x9kKuntlia8il7
tTQkBU4wVIYVltBHJ7q2NfKpG29VwcUvmGQblXjzwyynQILQNfDJr+n9Sh3MTyzw
RrtPJRnh22OFt87Pf47HUoR2tM2F6LjPsP4m2y9FCvSgbkhVhV0mDJemnkHcaoWB
ai8mEsTiil6CU9H2WPw7mWHNfG8HncLrzkhUa9zcfr4MSmDbkQyPvdfdAlGM29AW
1l0M9i8/TmgIwYYUww10BTFQwVO26Ojpj8LvK7Byig8bHHhOnNQhLNo8ZjkIJRnC
7+BohZWTWb63aZ6TWPK4W/3f46qnH9Ddg04IT3azksVSKpxi35emeDmpi9rMBKf+
JkFVdxbDVvOn/LAlrKCDz1kdEZR3VQQB7symme5nOYmDpsOq8Ptqko/3HdVAVf2K
vm0j9rmhBMQ9EaU8U4YWuNKwNt3A3aR61BYAm1mbvmqGWEQNAXlAKtCuvGxOLZSG
0H9bIpB1HgYuY56sdIBfpKsKojzrVlgXO7z15h9Y09FOVxwjYaC69diC4Oi3wLsI
Yqre285lJMSaU3+tnfBbHnYGG7KwOuvw6N6Gf0o/cCNNO2rXt4hx/YGHzt76FoZL
f02LBIFyBefQOfbvQZKKSyjLTfpGM/u/VQ897c3JPhxbeoC8GY4uTaCsagvQ3nb1
+H6zzZ8NNMTekOlqB14+/2KvMNhoo7z56exAOG+E5qLL8AER56C4J4Z+g4V6sMjc
QPzQrJzfdsJ6kXnqOyqnV+1stsub5b1Ve7mnKylcya+HPwwUT79hDQBqw1supHu0
GOHVaXMgKsfsDdw2UhD109p0kgHm/OobwJz6QHWE2ATpOv9eSwAKSkIX3TWC9kjg
cuVEEYFqRscEVPSVc0mNSdSaFujZQYPOibsZPLKSnsA0O8r2pslJ4BtI1aB6Jmok
jduEsFa3utnpJcftUK9lqLUwux2adIxG4sGEl5k16yS3jC6KsblAwq9kA+/unj4J
rVLop7kB9Qc07uud04OKhTQ9c3gUC9ROM8TkZrcZLg/BKilA7rANIFtGVbBDcShE
occRtiDAfyhDGTbIIhtAo2EFXabZyY5RrhzUl32erNL+T2NIDIjT5diybLrJH9ya
sVHgkGMriu/Tfo0OJCzU1MpTcjE5bW/qIppUjzogQ5FcSesJm+rAhkh95EfVmZ+K
jWKSRmau3IF36vRq8R9lfwjVFQ69Swi6y90hAXLJh05ncBznDE3Oh8O4BuUyMJvl
UieKhjYc/aUK7cACIetBevXRXT9pZIr7czXoGznnSGXsRw1SIPDrW1BHhiSGs2JQ
lzC+gxUCii2y9zlSzZ9H3BWeGYTh54iuGp4DiEC/tIAhWu7NVkTxsmIYG9AJADie
mNNy+boWGrqOxuM0TmEVZ1t9MvqfiNNdMhc9fjoM4XbHWFbKveoog7ThZQMd6Yzv
3+QnnDCkGO/UgmX+MUCy7dyWFlylDTe7CqClGW6WDc+gckadYXzFOEZ4l0LYUXJx
9VGCPpQnvlWKBTofStA5rxT3Kdvpl98FRbeiji2YUuzV5mb8t7kj1ECbkG1SuqUx
9Z3c+GDvPu33JEOGy18v0RMczXW6GMFG6j3wJU3jVqwICVNIaquCO2BQf8uSTMMg
mNQyIzQrredIDJdtIdimTCXrvvvFZxFmMKbxxsTUn4D7/Ef/YMR8c++bl3AvDW6k
na+iaoalp49+cLj2QJJqnjdCtVWaNyv6/dWr2Jr4/lef6yJcitZMuBVaBQNHGxFm
hbVurb39D3S/g0uCNoSAgdw9CPFAZbOW7IR5qzpvMlft+dJZzbG6BZskNdv6bUTD
3O0E4MO6+KecLLPi1Cel7sORviukiWgSJ15L176d5NHq/kxpXk5CbUpNpGpWS8HZ
pSdcsWNAcIwwg4RI8ZBPAij/2oB/jgd9tnlGC5DOmEW4BGpv1kV2hWEuQeGq18Ve
FOuQHWZphC7zjB/VQNDSjKgn/nD26PfFlfrpS3EUbKKHI/5nvAQm08VjthHbUZLt
7mW5NouizCpkdTLQaG7epDOvyCq8c9RcGspAbxpU1wQzVPijfaN6vr7wCo5YU64E
1YlL7Vv0pGWAKdaq7e4JWoGqgXPy245eLfBmvmzb1wOqOdjqGkqQxMKS3og+EVzH
7wb1WjrM7rqE4cgywaJOg0UMFv3mT480eQ0XQJxc50o419E0SvGqhPur76YP/7KW
GFbdj4qoQPdiODYgjIUmmdW3UVSbBFkG+UbE/zCpplSl2o6KOYU3hGsjUPtpRNyB
9s7Ur5ntkSpN7zZ+Ff0F7XkPGC5jl9d0EzPF4SbfMnFu5r2yVoz0gHs6xjEr6T82
SyygiYdrYm734eRgZve14bN3XuUfyrmHEYBPHUR1Z+7vvp/5u2p7ca16ehXg/Rq1
9URSZSd952qFDyy/H0llGSIOlhOrK7enNnaSBHggbsLGnY7Np3YdC0siGq9uAWM/
1KYybEKvb8CJ5WvSOkdT3FdpwVKE38qIIeKpl11uCU/ICBqUUXOMviA0QjZqOsjy
ytyjH+9aGxaMRs5D3rhacjbyRQcXwurUxpaOVkYGe25soLykc+4Y+mIzaXDGLhsg
fpRluK0PL54BR37SlllW410wG8+PaJDSLXUePO/XcC4n0VsvZKgr/PJCP5nAER27
nt/58s+ERokbMmZEc+a9sylJ+/TI5yNw2hUXuF3LxRc/XkkDfnx0jjV5Hnj30MXO
v04C5HJHjExrOGC5P+qUsAptb1LZP28eCzyb0YwQfXkfS7x7C5QLxaIY/rMlY/P8
JI8E6HIyO6yzTeBLq4bFsdnjQWL/Rl6tkeqbojV7A2YJlnl0pCBh5KRXAX5rY2VD
xY3R36dxvLT2Pg0i5MlJAFwtwit4s9KjI3b7Ncv6VwfMJfqVWCI3Ecumr7IWM9nh
ri/1D4ZyJH9q2I5mElFloL79sxyhqGm2gWC7oa2+KgbcNvBIApt6A+vrmrCt2FNQ
7TCsMW1wITHMwR7wpu8oBdlUlzaUhSsfsP4Uewtc6FAXSqlCNPJF7BXzIf1iOJ7n
3eOi1eXgF4992rRM1LFgmcWYRL4EEtd8oL0Y4AE6jxe1BS5ICFcX+DTSsAuDoJti
OKzCE3gHppKz2caro51IrNIhkpdiHYPGhb+XyKi02HZDuA5IaJ5XSext6++VBkS3
T2k+zYI+olrQfSx/AgNTb/jsPvDlOCj5QIQZ9i5pcrbpiE44tLKtIwHQAsvPTua0
VcgOwcV8PxUwaSKkZrtoVLbRg5AAE/F3hLffudUZ6sqdHnB1FgqYbODMxOybfay/
gD+FyxAdRQxchdI0l+GnXIdBFDLELM6axLMPc1KU4I3i2zsUa3B8PANm578ps1Ft
WstY04CzrJU3aq3veW6hVng3+WuZe4nHjrTy8ssQ2da0B6TOQ13/2FSM6WAyqB9t
N5NB5Fc7Xp9wo9h9zcgrdgVZN3pasp2dQIDXVQVNyaXOviQCk4U9qJjNBk7w0maJ
Tzu0x1rE5h9lUfzroqj1Aw/24mssW3B716xgl7WC94Y2RMAyXn4DrmSQMC3LhoQI
9UjwEFS1UDqM9wcj5muWnnU/j3TpLo7H8b0xbxf0H7hqNpvzNbezQ/nSgEBV7Fm/
9AVdIEpFCq85Yp8du2ZvuydOMX4L0hU/vdJ6Gzs01SaYpTf6IG7nGn2TNfJiwDrW
X5rjLnhQ/i0IHOPYLw9owfodaUd1ynXp1fFs9evTqdIFrBwac4uQnA9KX30NmPpL
+aO6DQ/Bo9LM3h/0HS6pn3VDCOwTRHja1dSFrl1qsN0TiQo9ESvbyr63oqcv16kS
uu4Yf5KsCrhZsXHQ21pA/r1jimZA9iZMie25D8w74yXUruiCG/Z+V2B989N6ec7q
rTCNKh1/zrEMtJJpf+bWZzq5A+Bq40pPSfKOgki0/tJuNqjkl+2v8srlJdAVuGQ6
2G/QbcuFwUdROl9BlrRwZs8QxTrJ3KJXSVUOH5Jk3HEy7EXNA9/A0SxI14X/pn9e
NkL62RyAmDpwFwFGXzWIStCltEVJ+5ys/32/umfTZStufrlU4U3IjY6Iy0xFsG7E
w8HVUiT29NZDeSPVWFy077cU+qXwkJMWGlERMyegoX/LtnY0tHl3hyEoG39h6a0y
SK6V7iWdQ3bkSnFqWk+ZL7+gKrXGHDWApKFzPA4wB4o3RkvBBE2CnDHiVoSrEnow
CqCTmXTLAO2h90Gk98qds3iNboz5EqR1L2tSyFita9khWZu8IArd7K103xvHrbte
g2taRkTiFipQ94hhPKvpplGKaurhUt4YkZXI7h+eK5jDb3Y11U2pzLbceQxQSzlw
Y8jfmiiDMEoSsuraXh7f2hQ8r7uw3ihdZB5orXN5pM/z3Ld7A7i0EyEoIDBczTYb
prs1qefoWIjZZi2L1iBTrY2AbxWu1cdHseTOHdYz4K9xGwRSqJOfAfQEbmq76ATJ
f42hQ1GvogEt/TJ7yGKLEvrd9igS3rotM59/ICq4+jXSSyLAXo0pwfFE0tE6WLAm
4/vAo8B8RIs12EAgRzgH7YtorHImhOWfBtFwAXyvLvfXBBAIA6PSZ+OshbfzHvLc
+cDjGnH4lowskJ2vfe4J4dM/RfqvcHYYECQMY5DlZi8DS22vkIiUPcset5mmH0eS
KesyMCy5cJVtwPuAs7kUBij6B5RV8HWHrLYWEqljnp5RZXYlF9p6a1pSJI7bFSxw
1NL+2UA8trv4vaNud1mFlVdnbajOMrBz2D5t8blgFmkDXDVg8Bydl04djID2hPoD
4Ktknc6pQdnzIvMqD0/sEwPjG5zLlzDfeeH8WUAjowT1Jrvc5XBqQueL8mD/xB3b
PU4N1NFDL4etvi6oe5AIjlR7TWgBQknt7nPSvE7781GKmqia2PsplRIaXHdi1If5
yT//IRobhHkj6psVsVf4/sHjKw7KcOcMfrFgoiLNUzggNrJ2Ixyi8RzAoJzQE1y1
Vm0fQ6ul1yTNtXIDXX5nZ/Oy+LwbNBi0zNFIYM4UFSa5AsjvoONqi8b+7V3THmqQ
RF0FwaJwwYw85KZX2hlihJjZXPzi/x6Ufon4t883gg5JfQtFtCAnmHixnwtjpVDL
KbEhVbnWXGtgvploTRzZRS92namEeAkjv3S+UuFuzX63D/oD3gqYHGxNDaYOb3x4
cVhFZWaIvuKWQPd4CeW5DaEAtFZtg5kO/ceqyFx2NZ6pFdeO2sLxSbgi8SkeSXCz
kL02z8Uioxfd7+RB7pMLPNw58A5lWzoXN6FC4/psGryQNyjMbjplhvjB/eB+Rua9
6jcik5ZV9I3p1xtiJnTFBg4jvvdoGnT/MC2rVuEXoJjyLcxlPsb8+AsHI6l4x6ix
NXvrUNPFndgG1Zqo3kxFc5bBrNS5ogL1A8gd3APEfhhvCxdewIvaXmuelItxxqSB
+l3oCcbuXz4eCzgUwspFxw5rcIGW0aGRcTu512hKULcp5eI0KkxBcXBoW57LNRnj
ZEr53dWh9jLJ95PmvI6reyipaxRxXUyN25p/tWOfR7vOg2jmM8pc64ckFrsH8aMA
SCPu0BqN6izej2wSA3czIpL62TFjMofy64qocz0s7lHewxoJ+XTR+j0FC3eDwAw2
BSKXn90l712/w/jiubuzXIN0+hlclmt2y9zaxGIYOv0jfxBRQN1GYtH8zWGsOeE/
EKz7R6/tF0uXnKoj0+7e9Rui74oZ5I+ED0RKQseZxYMrjplUQNNhoowVIwQP9cUG
KGl7ehJdu9ogpJ+CjAMCXkDsZeyFekciHJIV92Rod4EmaOv2nimOHEdjZdkUGqNE
WqhxH7NuOikhYZQce+td7Eu7RzbUTW3PF3xA87aWBliH0oHQkcF0WSE5YnF421Jj
3m2F9Oiv+pnL07QamAe2rbv9/+VzHBysHNv2CgqVLBQgjSm6iTXOdMrhPOf7SzpA
SNOVwSmh+7lg8sMqwRT/NiZaHNm9jZMfO6zOBXiso+rDw0stp0Lo7+NzlwScIz/F
+zJFY+Wi8dMGU5G3b5/CG2dsH7Etfo4Uejg0xa+P4d2uWVXB40yrfAA8fow6xkG8
RMYtXU5lB2DI567jmHwCkKsqK/prm45TGxulMxLSAvs1d7qF2+b4f8QbTicBSasb
eyq9agtpkYbIK+Fi+xb8Q8r95EVio/dNswfOf91+1ozaajNIwegZPlKTFDsQFdIR
sXB/eAcUVJjF0Cc809ibWlYFiu+QbksZ8yq7EleNWWwgEo+8KKfyNXQpvKcf59EZ
AnyZxAOt+nEvPqllybljo+jK1q18v/2T5DnGpNhM0Bj7+eseHZK5MwGkX7AFzKH8
YfYU7okUUZ8daMIeBv3L4plyNUMSqFgLfufODoNFQ/rhCa5TCxxkLX59FtYzNu9z
PjIB+KNTIoiYyYxgipYpI8e/tUoYLFUCFCEqx3c3FJF6S8p3j58e5/DUXi9GbFTZ
lGN97rIPHODWKclH0gnfNQiQ+c5fFD2JWEbsr/33SrfoA34GoyrByrCeiWn3IwFN
ZpdMs4I2vNyT8jRiWpQ3D/PSiW07BnJHETNeosTqMW+1wtFc+CcCN2t9539dnWjH
XqTmXwyVoejZpebXn2YVs5+OiTj+YAQTs90SP0fZIpqQM7Gj5xthReA4KdZKV7e6
qJCVVwmtklA+v3rD55gHYvrDBzBCN/3o5lpEhBpan/a5qJMEfLmqaf2ZjXe1a9PQ
/9GZEGdc8PnO+MLZ5ua2vMzXspaXopdShn1L0AohdHVDi4Z8KZszKMMYAzui0YA/
i8/TmO9J6sGjKcESDNsVGFTjK42BThcvQdZt/UiouysXrozIYaoVTpdGdH6dWqK5
Dcv/a0SX6f6qV3PgHF60V3PpinzKpGRCydPx4eCe1UjbJEUFWFq2yMiLm80COE9f
lU2AR4wf/xNiU9qZzTpGTwAIal4f0BIKwr08JJyj5Tqbks8pkAcnVOhlHA5jYV6r
Bxbg9p2Z6ZX8d3BDqHF4b8nJ4b6d7h80yTYtwiFm7R69IXYuMf761WyNPRnwZ/NV
GiZBsVkHtzjKV47mNoXYmAXmlaXKu4YZPY8KAgL0IMRWYWnB1JjgoWzs0zv60FTP
PaDDhAoP1JPbCX1GhiIb9kNV0qS8yTWQ8J/gQj/C6D6GMXlm3DtCPwDhnB+BJL/l
5mSx9HNdPN62rHILsCtSODjx78zER6tGV6/Jq2Yc4OObFUEfV5Rom9LQ0dpfjcvq
uKUGVT/WaA+VE1cEkFuDyFsStUTXPbtpSRI/jf+slVuvm1KKDwNHYSX2vwfhe2zL
qvBsrIcgHEyvGpiGXjvP2n5lQ9u5hmMYpnkFHxjsvVtjCVhc1AGRuoZPG3756JJS
QjszcimoUvGRJJ4NHNo6Ds5qWzxnCC8eTa+QvG4XC9Z5pXfqtAKb5rrUgpqsLBZv
ncoiEUOzuyxHaQDs61kSsP/YvYterW0MLXD0BE8OAVv7GG4+hhbu5Kj7vYRnTSt7
0ssDH3lH0CgtAaZshyUETzG+Ao3B6mCWyxj5muhkmb5BoZtsZAdsE5fyHNT1IbX9
T8PRRBHirp+2+q/OMu+ArlnPsLI3M1tA/iNN+7sypSrnwSHE2FBNGhq5Ij9Q2A4Y
O+NshirQUGhL+zbqsnTfvWHCtEufXunl4dr5cPlyMhpQeDIt67/6gVAS89nZbTMW
2ncoX9FbXkC4XgKcfleZiKE2sYzraowRWDTybjQP3VGJ4kyulenOXbI7rBwD1y29
LbDxFE+NpSC7LFOQieWRoASMRgXIq6Dyc7d1OfGKEFweLnLIzguKx6obUE0Pp6Rv
ew4AMV1iw0GfznyUfBQ87fY7V45eGdxk1b/2H5PKHpqzNXNUnr8ytRa8GDAuHend
v8zWxLTvk9fQjbXAsX1v3S1c8Pcf6tMgQkQIAP0/uCX6+mKrw5ALh788EW1D5ncb
SLLQ86TCUFuoiB8LaPUxxXZ+XUiPt4GZ23WSBupPxDuitWYHpnsvIHkz0hddC74w
tOQVy751S0lo7qeaVEUvdxI2+jUtlIWpx74bq90gdSgFVVh8+GvAAFVzC0W0f7yw
Z4Aie50cgmVlyz/OTiz65pmFquawPNkNXxAQ8BuLd2y8SOO6tw0PkvyN5ddbBOtS
7Eder3LmzCNIKBXppuZCeDqsqbKF0FdoLHq55ysR5CtW9TevXoEuf7Zyg6+MRUiU
lDr11lw43YLkKDhRgXnpCJ/YV4hno2Dn7KDJCNJE0YGKV4qFbTcMWMwN+KzcOe1p
SLUXOERRLUias0YkC2CuN7Y7eh2nZRf5g9qon+QZvz1X5kGci1j4rfZHgzCi7PIu
A9jt6vCaFctTEkkL38zN65bQxDPQKfpQm5xXAFVnXOmCgczhMb1YhU+99k2QsSJo
V8GP42SoK3iWD+iqrp00R5Tg3uTwbtsfPE/pDqARW1a4MumuYLH9nIZbCqCb8mvs
nfbZ7B8Dn/JaVcObYyhflrGBErd5e6xfLtMSnkJ0C6bDh+R27Q/Hn2x0DTGcDcIB
YG4ExjtaSkKAkRYnzydNVeT7LFsAQbGJuQhVqMbd/Mcpa2A5xgzZtHfGqTDFrv/f
/I1SS6zN580+E8l6bjPbF7UmF0/2CGavialhbQOcIGpnGRwUq48xTNROmvDIROsI
m25IoE9Bv2hoIvgize4uWoMlZl9bEiWWOcTak6dT4v6TZF/FxrI9Ou0gOHpphR0u
Hd1frQ/6MCSgHVRoMYWzOTMO8+5ZavbzCAaAQ+qqKLo0Hs/MO0hLdX7QjU4+fI2v
J9dxNUfx6Noa9dnUY7g1Tq47rKNK2UEkMhyvR4+lMPvyftSWrTXgK3TIwkM++EWQ
pltmbfEzEse8LUcwhpSxR21iJOrTYPHGW/+u4rZTTl1XlLfztJSrq4oVf3Tf+NYK
dmq4QhuXDuHxZQi0esVvew754kQ7GfwBkVb0dY9LloKrrmXAbJ3DmxxA2j0ay0un
I/lfjSDC10yKT4wkZNOExiIpZIXrw8Mq6uIfCQR111Xu7rjtQZtING3zVUHkv/ce
8VaKCiJQF1lpxunvy5qkKgvBOv8kOP1jTsy/qvtT0PIqZXJboaqArGvDL9/x0GML
aEBuLGcPHUupoLWe27XBsRzyczq+II7Q8sNAduRx7ic2/nu05SKqFz2Hw5sOzf8h
NrTOl5zmRB1EkV3bZ1zIT9CBi8uoH5IYJr2yGKudaHPgZsvj83XqHZ1a+eRjEzhT
wO7MdyKBFhS/mgx/gHACjbvHquDMTabxVKQSqL8YhB4gKtHDIu1tmEm6oCrjZySb
j6x4QTDNwdTi9Hlh6xUewbjZ7Z2TqOBApcVb8HR04bdmmoMAh885hAWZYgiXU+Zn
UwmSik7DNv0eSe8N325GedvoWBqa8ZmLCWQKYaxrVzh3vw4lb9vUV9FJyOYI8wNM
XVLIBg/f+M29nX2OFFdxhDtMlTtNJdcfRkYaRimcwGW+WeU6Zj0QbRN/CClyqfNg
b5Y/f6KXUNiqx08bfPDSV407IyoNQu49BEk5aWRKk9xrCZqo8P1VMXMgG6cgKXDT
2VumWlJjkhg/x9Uzb4Cs90vboUhn52dkVl3BQ/pXq4jYIXVbw0GTIr4mIiCo6mMo
YsC/BEk3lkczkaWgf5XIsaB86x/ryivs7awyXGlUjq0d+K2uM03ztfSwmbJw79fA
BM7DBAy9koUhdljPshcYmgScn6ByX9GWm5LuukQvDzyxbcprIMSW4gfuHOPeGJaa
EMBlfrBTA83+9HtuA9g37ujjSL9sjpy913Gte5aMNG2u9OXl1Ub+IbBMKkBbi/5O
LSvKJPk1ZQNJFIOw/PzPgiPY6GUQtw/+MxgfhrmqZpDaRh5s5/xP/cJDbK/bi5i8
OKazNxjzxVHZI0yRPnCaZyScvn6bfouDA4sjJLtceTcaLDppXIbKwzJyPcLIsfi/
ySf/VYSUthNbjWG1rL/2O2XOcVQF5WSrfs3SbmFewduULbD3KHl+XnkxTjsXJ3fE
zLsC2RK/CLx9p9wMtkTzn2wd3x8Ynf+x6Irt0mAniq09IbOrSAixv62uZ3RjHB/O
KBk2LAGG4+566oh213lRXXMEpA3T7vrP41QCsr+2kww5oIEG7JRLuJl5+3KzN99P
m078h+DVQJXUfk1RXb4R0tk4g/85+OsBZyWDeq6m0BEPEcczkDf/A/FjaSophoWv
c0nZojRhyx4lOpSjf2dNHHgQlNWhQgqbDrT1DgyA6NGSZBa7hznZ+ZdIggJGOqPj
MsRKxo7s/E0rwPtLFvWMdllKBYDJJMWZjX6UY1jzrILup7OoslvXxlifJoRcmxQ7
NQ3OxlRTUxmHexrGC8eh3nlTKlGPlLnRWyoBFjpLL14Qzm9KGS9pPFjfA1/Oocz/
OYY4FEqdJJ0uJTFFnmrr03lRIUz7R85IngIChRDtPUB+f4yslPVUb30S3gaU5MGu
wrtNo6zmZo/OffDZjZGaVSzW0G8+cbzBv36x1qn34N5Q6FotxVgP8JsuoTM32Oqn
/Vkh9EF11yE+/45SUtq+hibCtR5vLczY07EoiGKSquOXfFO9ViCYDHDY90I4l0f1
rHTIZAM1Q8rZZ3b1YMP0qa6sx0CTtNd4Degb5M/QzNfoAfpOyOxHNLJKYuZsXLE3
yQfk+ZKv3T7iJ8Pkhedi31pXjH3FtME3y7bgXAce0sP/vkiP4cEDpFjqupQgIINP
Vux9I636Cm68qIRWZS0SPIM22gleUZNdaEw7K776CI7CTH2rQIlSBqcApWQ3dEzD
48uavGQ1wt1B7hpozKzAl80346f/kK8/XwMB3QLEl/ngxPzti6W5Ns8QmOFxQQt7
Ia5jEkb9/pRePy/ksYrwMg3139XOHLjvsMaUNZBBm/yfpdh+EpeNv3PmDH4o+4+s
4kp9oGKAA/WlJPl22lI0P6MLYcDhDVuG2D1uAfLj0OWTRmDfP0tJHjasSriXObM3
hC/46t5BQQ1zD0wMUtBsfd21/wRRpRFhpvTznHKCUQlhgNJFi00YFwrrPBOZJyEl
rymghbXlcSpXurMM8IHZIfSSJWP0ACa1VHz+7WFzF0g59cx2Qn0xhKRFfyLWv3EJ
XLKsHCHqiRIQVGJA/IJdHdSXXPlMcyt68U4H6USYAnSbF8CldCGFF26dTqPB57Ux
oxNV3OB4Y+yu0FlM01fEbki6ko5LFDHAG4Ffv/UhcWxOnEtt8EcP8ihq5NEsXb7L
Yud0AwIEYHVP5bwrMQl8e9cHh6GCZ2bLpoTwOUtk6AxvidifUq7rxYZBN3VC/Ayi
tx8PUQIrjYlSdbPdGleC565N0HdSZpyXj7gyrhj5OMBq2r4YPndu7Ef3y3ZVY6/A
k1C5E/awpVi0d/SSNZlDfGhSemF4s0k0KUUVDCQYR6rDhfidiQIHI5Dt66OKV76v
iWNHS/508U01l6u9sF52+eMElcbHkmx6UejXD4qXO8PhiRT+ih6jV2DEw13FzLtm
yHbn6sV22eAIz3LfZ99ZaFrFaCW1aZi77o9q/n9xAvfXX3MTMF/HenGOg54XwjRF
uJOudUl15ho6mYELQ+PhNlgeLeUhffiXbC5Unm3/8JS1ikQoSSTDpeI8CDlITj23
h7bBgCUx4dYsLDgfKLHuQAAq+ydlmG1nQzKUGmi74K0ZIlfKU+7JfwxD8EZouayP
7mefP4o9yJWjVRHd01lRvYyA0vVySby/kBln9Kom4FsKEyg4YZ096Ag3Jl35OpZT
7Yo5llxfRp3qWlq1+fVCPqIDwj/7b8Bf+zI1lRLL5JFqhfC9w8yuK8MlfhNy9Vdc
+ulZgH4hWX2J00jc+4ULHhGz0oS19Yo339I3pecQkZfqB3tJCuPYn1WlU6W9EHC4
4fWi7HuDAS098A4DMRU6QFYJ6igNtjW0R+hmchQPACfKPRM3WbnRV2k/wtq20Prp
xOeXw2V/QOdoYGqR8DjfFAXI4qdvVFY2gCHGfognydy+F4+Yz1rxcgsAnFudgyfc
TbWjl+XNySe0O65LXSdLijMR6HxmSMFl4ixEu09m531lvDnfjm5lvcpJa+DFpk3Y
vwKdAbAX+jG37aBRQdTWhHNtClE1ZnCI8jXHESliqmnKz4Mgmk0v59HJkUR+TGt/
0k2OScSgxeN6puCbcDN7oyiyck0Fxd4fmEPYrYHamgTMBV8nZDsGUC7HNbPOw3oM
Bv9ZK7WQElSIvX8zd/ktEDkzGC1i4DGvJgfKlrWQjbA05JVtj1CNspwIdVqTtlCY
WeuorQpJiAt3uGm6upo4hMVOMJCIiPFcFaQAm5r7KzFOvLlVmN1g5zkhrZWVYNl7
ioRYV/4dmoO2FOOtHgEJyI227kHK7o/cdNFWmMYCWCth0lAzu9OcOb4KZjmA+SqD
w3yyfiljcMf32Nmjh/VE+LGnXNlyOr1fTEOQVdE0SyfGU1C5eQXV8B580lsSHrW6
tnozI2fVjHB6WSn6ucaQnwN7UAoK8xGB913OxiTr7MPEhM3Bg42sEXes9e894dW/
Fpb/ykPu44kpR5fJyZ4XPpdhVV1c+dgfX0lDEmvDCmtwW9XpOsdb+2c6OWhYXK+o
7WkLyBJa9AxyQPIh+WfPZM2gXTcXI4c2n2RDFTS8anCudP8u8M7qQTsFxnvxPrw/
KPNbLlxqMTCJMQcrpLqjPoqL8I4GqZ0hDWvPvph1BD1DZkisowtnJofcuTqauYc1
jNn0Va5XyuarkmqJuoRbOVCKdbRusD/rlBLLVfu0zRogoCvHxomeIG5Vq5jn7sDy
YnsQl/huYPIQgm8elA4T5K4YqJTw86N5ux9bMjdroKZHoztzgICraaP2/M6Kn4tB
p9tRQB6JilEhoMK7LIG+CH+sOBzq+5AkODM84/iaiqu7rMVcUAJqDApU8oVpzj+V
qw0pWI+7uzTGUe0MGca3yQvq6wgrOPqeA1HKGbCr5PsJyzYHvFnEMwhZK1lUEJbP
wvnaUOFveToqUqwARu7KWfj24QwcgY97IrC1s+N3HP/oydRqccU+cF9MUOdY1JYa
F1t6yn3vZL5kQfS48+Jkf0jiZO4LModKmj6LwJQ8SjCJ4fVsBC+6i5UPVFMDvIGh
MLLpvi2OYA5J3BMaLD++z/ZSQ0QZmWGzAFARRPY+JczWQq53XaKC5Qub/Z4yOD+c
1LBJ6Q72r996Z8VJeHxLl+VU+Vu4OEWjlwLxUMg32GAtdytcOeEjTgatWyquf6E6
NKS0VBYbCraTy8CQhhbmB92pMYQ/j22TEPZsADQF6Ep/3s3dDLixKQz90u9RAJAc
P+TSZT88QTVR6erha3mONxSKtgeH/c0X0q3/h0LOR5BnEa1icu+qXqRADaaSG1eq
nvZ7M3fzCRmYrOhBrjt2NuCQxbhpt4gLjPxlDE+6LFEQ056K7mppBO84auEy0cC0
+EsMkoHF9SwO6HxRCaf61dpsxbc2COetJMMBKR3gg9rZOjQeXFKZmHIbreCLY+d2
6Mx23kr/3rrNq0SgIPC1hjnbIQ/yTGN9C9YAqdg+wL5EGDvK07+RnYYrkKA1GiBt
gJhZNxH4YLD9jkRnEbU6kYtztwoaQSGWnANu1APA3v4siP2e8ln5f/WGMm1RN+r/
K1T8BoW8cwKJKbsTGimF13ZrE83N8AZOh5+nUK4SCGSt+9l2JKBy2kKxmMFMLLSN
GNgDGM9Q03ym2HRbX0hIR5AmwTSkfg3xUPG9SVIEsF+LQy8eqGI1vpcUXLVITmff
ktpS1m32oYAEpclr3TJxTvQu9fLRk1jxCBPfN1bCQOxrqa/DV6w2YTtA5Yq9ap8L
0Jk80Lit4Pzksfb6hb549/c/7L1CN7ecjE0v9M2AsH3HnDXKLngMzIKons/TCekJ
gfe8fhfDOAtL1j3H62E12OSkSgckn5Qg8wWak41ch4BQeJ2LCsN8VTr8b0Ud9+7F
PeFLOMWwB2XuJkbxUVQl7BCbVBPpzXVzmgBFK4Eg3k8JTTzTfsuBNZViEq46UDqE
lGZEVlH20ABtxOdqXG1CYru5BF7hEqv0QpbgynWUY8ro42ukpiQ17HEr4Bpd7TCi
0nbRMbyoFTKijTX7krBQE1bPbRw/fvOoxHTShsA3gSndiVtaf0FFEqVklDuWypej
SLmIbsPpFfAAudPlYMKTpP6ukqPVjKX+usLTdOj4uVkk3PxyBICapFcu0m4RMtup
PlyAVlYODDQYEBJwn5vVCMYXGqIO9xUc34ttjj3qgHHIw8RZW4vwz4zL3EzpB0VQ
TIFxbGpKnAOUUjZCfjjkrh59E+KVZIL49nxIsMIlGFYcuCPB9Xu0MXopFULODQ7y
9eAf40OjVZavHxN4MO1sNDz1H/Mg/A/iuxat8hQsevlzOh9Qdo3ieUOmHPsJ4bYp
mJGZO/niV6bKb/t59T1zPRChY1C8yAPb4px+JO/UANjnQ/vJwmLBC1TohI028Rqr
BInf6cfuTfTXXoxAW4hOwnuq4MLR80UMxffUxLIgWl+7BjcqdS9cEVOod14Ui6ub
0rJscVOf07osEHHnD8zIB5J3UP4EphMlBnKQN1Dzr24FYD356Pa6PlpMLRQwUWZf
0UttnQgStvMenQX5Ty6J89EqH+WLS7xWfB43ZZLkipwH1j9AHofDGUiNiwb0qah9
0TrCOhesxn6dtxHiubRd9rtFDgn//su63ffmDYPVh159k7LvHvk8Cgbk/VWvGkdG
XEBQU6EdUoaZw8MyU75F3XK620FwewYiOK4L+BPQsbcuF87pg8w9S+OWojb20Nh9
N/vY5QihNUrshwLCIo9tusRH5MQAxvTyFIzM18xp2P+HJwHhwu9UwLj29mYzrRnY
Bxe6meZOghoqxeBV6CLl+sJVANkTAim3pKWZFcQ8OxOxR+6FYvgj6izXo3iat+Vi
kZBnlMtVrAeo8VfyeuM3gyEHuR2aWSulDxMMf9Cr1xze9Gtls5d3lPNNPH9I1/jS
FbjtFT4igtYPc/ICl/BhSmg+wgeJxLDabeesZeKqn6BFsAvLW27HEw56QbXmy5vy
Efhn6eCh6G8UmCdIybd+yKOT+3vfBY9rI16crgCTFXw59tdjya654GsA6FpFeXD3
UgPR5gleZAfFDXdoxOTh5X8vsHwRTv3WRGr64Se+Po6p4zT6mAkXZ+1MiCOrqlKz
3UKmYVeNCXud2C4kpngOSBh0JEvioomoIwMbAiJSu69BbLdiBnTkpxYEzAzDHvYT
pm2fxCXR6JRMnVdOzBIgbhAULDIOdKRTSyNkP64xr6iwDC5+Apr/0AUt13pZSn/7
xzXqmmwTeEyirk7GXsziouBbkYYuDRBej7WzdXYWzxY4haBMUQXPx/1y5T5qjIhK
7ncamfjG3IIYts24hpGvLPI3UdsGy0KknwEHhBRo1Q1Vdwd4kuqCuV1a4JG9HowP
yacPTxGDFBYY0Zccj6N33tjFNYhuV8Cm63BhYMxK6X0vkLlS6WOgDyAYu9w/9N48
QZgK1iRmdqAZuEE44RUTYnbDtrAq/sWojDH3pdhDyD+5y0TnXJeoNfPyjuRbOYJ/
WJ7ZiR2svj3acLHIX5DcxeBv1pqPQD2VuXyfgDP5hOT46L4v5hChGakIJewQD8Ey
JZ4cYqcM0W6FJ8/frP2jBXg1md8hioIHWiLpvuvaYpBRF/rTmanPF0b4JXh1kYrk
8lk4hfBKjcFjDksDP8CJK0iVzfnsxltuQw+qU30Kpz0EmMWOrYAjWLivWjEbAldn
grQSx8KvcBqlnLWMtXQ7VSWY3DIO2SsC0ma8OL8z/5jaE7rQSWFjjF+hfS4kH8ao
lT07nMahf7k7y39VFZmJyw16DKn42Yz/QouiP2SdAp33KtrHKl9k82ZGHeEd9bvU
5Glli/PszfOWGGgg93o/0zYPSr3J+svlpLA0B6JtV5tRdKDoWCXmWYc0zh+ReZDr
xvr1aeRSHtVXZb95HdBNbOSp+9Cm3HUpidUZI0Ktp4ei0l9GRVa++k6LtmCnizuA
vCCtZYYzuUxjbuazvubnzYoVwMkAN1nvIi/KIH2Iys7b/9TzUrzSgugCTdVMKyi4
UeUSytgQzSPkCYt2Ht/qIwW7far34QlF2cTkL2WvXq5LtfKDr0NwQDFeIpZ3sD7n
nBS8htAwy9MfbKSQsFWyz8n7U6pVLIqhylXyrbSx17QclnBGCpKtBNwAX9CQy/rv
o8A/jnEbcEzhN/dcJP3AnY/Vl/GQmg0GUQeZQWytw10J5Gn1ukPC5YCvWtBn4tUn
Ps5f11u/lRvnIkcxAhuXZH3uOJJRrWjcOCGO/JnzvAUQyDRLnEnkW7gMpju/aFkF
R/+SE+/5Ty+3nr8Le5XhV6OG68b8h2x1NgvaCiA5b7T7207f/CvS/ggMaDo8pORK
rTleg9Tf+ohWsJ5TDtR52E1hr9EyIzqzT98JPA7T39mvcCAuxeP/KepIGl6JQoSr
Ouw2kKmqrhStIv4pGwoKtVw4cQWtjJdu/z6h0GONsCSo9AlmRJH3DcVfeJAMU7u1
hOpZRXBpsWJOhny5kDNNCkf+YdOMTAZ2ftRZrqeHQw3DHqdERmlgt18Yp7WOMMoR
gxPugko/tmoFmBxkfgmlb+7evajmABtw2QPBcu4BfFcBC1AxrPsSmL27WBtUxb6q
uVFZxCEvCUetMv9U0FVU+DNX6ZKjwlc/Q4BZR+a9eSdx8C0Sf7xHuAneNNe3aXmk
VCKJp2GRpMpNPYDeqnvOocXZ3+HLjtMmBljEwrENP/xJKvDQDK/5IfHg62QapiBH
VZIrB11ddfTU3hxT3DMQXJYkNA0ow7sBOAbdqHJqFxu+sWbYBRjDIVsMtQLcnVKL
82B7aBTHYtgGMOq/K7TfbmrlcJKglK8RUstMHQKu2IGFnKFT55yOFLfx395Bqe1n
VkFXlRpGG3aZq72BZ0SAFgdbNE2NGRSE7jQ29yd7GmuEUuC13sY/NRhtR+nwDeHu
YPCgY31NraV1pEweUB5ILC4V8mESuWgU+PM6TxydVJQ4l+SXdRyEO/+S/Mds1GBP
Sw6fcYeftcA6QS+3IcUEMUHk7qrzVhh0jXJ3XJWEX+Ai5iKLVK3p/DXLIPlzeRUl
vEZTHF0zA3juM+ZmeL7L3QWvUDbnR6Y+z6SLT3PLmlWo5QTWx3/5sBjIvYI/mtID
B+GQIP4dSyq7+HaGi8xPPoIxMPpTYYbGLfUFw1ybekLY8zlfcYY8owxsVb5OWBMC
n6MtaQoqdXDUxmDBefu+ZGNwTYV8jHOKq36yaFoRqsCxmLlWcXwitUpduDpj/Lrf
gYjhF/P3xgT/S2TcCON7+vjWVQS2JWJ7AeyRRJ3omKajLstppsw9Vf0gIyodcRD9
ptMlWGNAyvqD+3ED4I7wHPz5Clsky7ZG6HE4UaBGza+nYdQGxHs9QvTV/YbqlnVG
zgukXcl46woeeu23x2y5tAsRI/kBQqztPnPEhj4y0iwl3hha3DBZENivXRynAver
KHad++1fLTwU+2qWlxOV2nRsdOacTjo7XPHHvp+Xf9dy5g1GmTd3SjTQshM+RAR1
u13mOfN4nnOn+Z+xxbLnsuTfL0E4Mb4icT+H6bzxXomTZmzxfjApeQLuHw6HUPMZ
dlEraw/l0t8CYO6vnJygBkJD5mI6TXLOf7ude0v5fOu6iKgVAYRwkYqAfrNszyD9
rbXS/kgFi5kP+ytuulzFXWZQ+6q9sBGJHn1wwcQGHFNAzBqmSGIJ0iV8xETEY8+q
+m3JLIbCrsH3tgnk/IZRxh6Az/BMqzo7rYOecuTOpAJcjhih45iEyuio+SzJO32s
Vzeu5Vd+MKgcJApEejFB8kKc+1+H0X6/7uyFfHER+qi8afO7j8/TuwJ9mDH8/fMa
pf+qATuG15BO7mTwoK5Tb3RN3N153lwYhxgZCe1oAbGTOpB3v/pkLJAgSEVzjbxJ
G05I7nmdfOGjZmQ/gPsNMyAGpd/ZU3iXnghOddYockKwPOO0B100n7QhsvUXK/R7
ciHXxOZ+kQ8+xHDz9g9eAMTLIsgqBgQvVmLKyU+y0PsWDjZwYJI/18d50NheTM8I
fpU7y3hd7mdDq03ygeKIeI3KkcsPR85u8EAlzggkY4HS0zoa6uhDhmhJ3Kc2XkIn
cITArbhxAKISrTobBLtmT6IDrjWsw2d/tUPoOxHDQj2Y4yTEKctF+xuZ2GxEJkMb
7PSlPnbGdUGccj2UL9/AsIrSWhLVyO1gTS6JIR/yPAG7Gb62asO6D4MSFUSY41Yz
+hIdqjJRRc7Lmr4n+dzkEDWlgcw8NzXsbqUf5YQJM9FLVYrFcnLwzl4gRVsKD6B3
M/jiVPslkL7E4x3UJ54wyA7rnBIKH2dddLMXWU13uvD7DZyl4iTiXPpDioPFGh3z
uTMDHymKo/zXH3oeczehDaaxyDHy0BqalxVM5XvJurA2KH8oiABWjVM+pX+HoBrW
+8492AEZiRGH+/asx7laizdRD6LoOMp/vAQUkwC4K/xWZvb1lXjp7mDvD1RZMMPb
y8l0INU4sL/zagwwJj7v1Mr0M5bH4RrTOUfVyKXUJkimZ+XnXZdkq3ncviL3uY5B
zUi1hDLfoV4pvNI6zYDF07p+xrFZxQQOmeSDATdeJ89wymyz4Fj/wtmblSIWt0Uw
OBh+T00u9qvT1ll8oT/s5XDl3KkHv/yCjWIPntAoeGsjrhgnACXFUNcKhKPjVtrz
gUIrZ4VrSEgXQCAMuizOcgSKG/wAGA0DR2yp+AvWo2YuZ3yF5Msy/6/M3k6CuYHE
+sbkYZjL6ZxugyxrNRedKbB0lQctFC2IAeO85JzjkCi7qChMrvkaWqXlm3HYyASA
z2wqDoF/ZwUWfkeZKqw8koKLnym5kHM+C8pGRaErj2zYtu+Hq7RiprXqbeE8VGnh
SnHMEUT9cvekwLGiClMDsCygAXZVsYa/XXh6Fm4buI+ndoeMqjE0eogdWGf2af4o
97ZZASso0i+79CRHPuedFDfygLAfhWrbebF24DV7EBMDqZqEnOwp56OetzAATqjY
Hkau1q6o8ZFr6wkbqM2Gs6m1A0NAnn/3v8+XDzbmICA4lZokognIYp5MfI5ax1Rt
mAQZp+/TCNpjthAWz8DHPUn1tt3GgAvBFbGwoEKLPErGDsAL9QGAmrkQS0vMagMj
nu7AFyr81JnOTwKNmTm1fqmVqRA7ergIy22N3V0H3gFPKYCbRkoMi+SVbsPWYeA+
XDe5jZ7R1aWZ5gxxlr/Yw+ZP/vPc2cBCKbLGO62RRfBRx+5p9+whfme2rMbSPtEx
7ofNLIwe8YL77aPXVaLZ5fWlbXoHZ9HHXuEwvV78R5XHaDW8oKkAWYenQXf65lrQ
RCWqzrtfjR/t03eRTE3VlAI7bjq+rLpdoO+5HOkgvZbJCeQNdKo+Ri9Ql6qybyg/
mPmP1MSGQ/j8CwHYm8DeEMtoFG2JqidK7WYwPY8sY4eaR7j8T3JPvVAYIHugTm0N
UFoNceXy/nmyMAunv82jqNyGylQJLHBX4eN8By3rnm53eIjWdQPqAlq3xcRgtvU2
7ZozgeCE0jT4GQGW6s+v3U9kZW5giYnSlg9YVK5GKHNBdOkRP/xAH0CDKfT8UHPV
x5vmah7yIejbJoRMWWr4KKp/Aw4/2be0kJawNHOPq5coB7QhzNO27thjgu6HsZPF
g+paRtHckcrFzzoAwy8S6pntHazPGt92xnQefyo2fYjuN/bVZzp0pazqIemaAGXP
YEh0+9Z651SAvEcEkFCd40thSieY6PnOCOHKlOW/W4fTSF6b7QjuyWaHfyotUY7t
xaBkGdkk4GeqsvMPVwXMZpJERdW/JEToVlLT5xYdjBoAao2OGnmbJmY+9FBersSb
8xYWolmIJih5+qR0rG2Vr5T+rkPEq7fgPG91Iq2pBe9rTPnIKIGKXfhJj1k8SCQe
MP3HCe8YNRZ0gXLvxN8tW8Ai4SClPjPBS4FdMdowIkYuTqCkxwBfsVGIJqoplB4I
UT6dyNyGlZCxBQSKbn8RC+BGCaOhPvtXF6zNxK26Citv/rLG6fAbjVOaLGN/DYCn
cF2DWoL/+crmaeW/qxhq2criKKm0Cm6LIE2Stnhj2Y6MURVSgDkze09hFeA/upiA
ph9PWOP1kkWlG10iW3RLBdrFWPnXWx+eKOlk7ENKZuWDKLiZ1X7iVeQw466vvKYS
zmU1DBZ4WKrJh3NKO4IJ/0U5eUwks+60aH7YUYTTTsufD7krpNJ0KB6GR2BJl7xX
fUEJCsrauwj3a4JMsvYwHsPiCWdhXVBiEWH+6cGbj4oqXpjr81siTUWZn/zCGkvC
gNfMh3/guygwcE9T+qWHt+vtJXCZCToZkiEU8QhoOOX75w893CUyzYESyMCqcA0e
u71k9MfqsbeUSJzG1EfjXyQarsH8BsqnxQGxBZwq6hrqHrKw/fvnjdHzHchZF0aU
PHDKlMVDTDQFQiiPOHA2a3DsWMP56Ok78g++8SXAnxiLE9ra/6X3aAMhDqBqYw4t
dTJyBxnHcHAc1SFtJ69w2whz+imIeZv5HhLzEblKBKY/7i1mN+3ttpil6v8UWjL1
gMykohDm74PqQ1kjWa2tWHYyRGSMnPfhJOTuP80tvTDaIxvRHvis2xbO9dTv6ZQZ
6Qpw0F9nYrKfBKkRPeF2gXVoNtXQXTIHMaE8v7hV4X15eOEY9SHvRf7F/ZrK3yVX
QtX3ZsAu9QQUJUpKPYDItcyGzMN5CujRp8LzegIncDndMm8ENOnihB4rraFj59/E
uwg7lZLHpYo//gGC5wsmwQewMLXl14vuAbq9zaK0jW5Rw4wR/kb5l10K8akq2KcX
R49DOnY0kdCEFl3wfiDgOd9Q1VvptYnh/nIzmeTa8fXs/RB7H/F3Nmhj+DSfA6sa
HLPIm7f/MBKNlXNf2Wu5KEkrizf4pWp3YyqK7puThrBsBdxVWA66Z98Hfj/STYfL
SQAb2TM0iVdfEfwpsI0EyUzL/rbIGAj8/l02mg9DdIWteP9BIgmFwqV166HtsJZM
JFddNcY7+Qj8PIPmbuXTPI62OIq+MQKdt9ktEv4MC/Hjtqm6ck/E+L5fzw+FgKGo
tRsuwgM3YgPGJ3XThuQ12LpPQdz/iOtV2j04FzbNu2ujhIa7pyBYXQU5qHE/FNRK
DrlGaPLObMPOThNYPbT4GlUqKffXnqV4OoATpADgPa47k6x2NMeR8aT9QhnjIzRa
GH8AkaEro05b4+m5HoBg0ZyVTCchKofqSvlvO8TcT4VGcXLwiMSJF/YTOxl9dZce
2nCc8VSSPpa/1+U1ijbjBm6o3JfiVsfTMhkb6KLv35ZZwgm0WRP89SO2Ctw3vPgA
zIVyFWmk4tuabjPx7Wm0+jGnoEBOVJik2gyHlEA1A4IfoTDohJxqiL46jBID4aP3
cY4XiaqleSjCGONO7mkzkSSm9BdYlbVQDsamNGhOXS4R9fs0OcfsC2EeZCYVS8lB
ilrdlQvSLf2iukmv+wJUaMlVi+TlmkcIBceAyy/EYfcHWP2w3JHGUzlumNgIfhmd
uQb28GflzxCm7qjNHcvqQTLB4g1jMeRZp90VjhOBq9QFt7/kcgGxAdG7xy7nHex/
vaoe0zw2GkmE44xZdVNGHB4s2Z1XrDoj4/tiM+AMrc88OZAB1AgWum3bDEbbQIzf
ogysbURSdG0KwOhv+1juZW47eRvGvfhV/WfS3qJDj9pyu1u1G/tlSNGXXZ9FWrrM
MPtN7ChRO24GTYD2PPpmBs09jiFPgQPVJsfv++3yDXLOWLv79AmDhxTr1H8CrgAh
8W3/yWdC7TV7qMGSXuE40h43Oeav5jkr0/VKMszXgjBXCtZV0uBLnglY6DSNZBBv
3QJvHhJ7dG0OzXNOJ4YF+hNQkYzWnnGafIoZDX+/2vXiwqit0JaSZfReEDJYxDI/
MhUwKn+8P7jEK1zyGR2DchJmT0RW9jANQHkBg9opC9xtAFtv+PuBG0rt2+I8dU9A
Op4gNLo9Ld6Gi3eJJkVmccP5v3R3Qdomg4BxQAFputzCwA/MTADo6yM3NbM86ZKj
iXw+8uGk9eD439IBc1hIxAmQW3jXVC3ipGM76AiSRp3tKbyzJajrH0pACh/eLWs/
paDYlIdvuLpIhJDcceMFLTRPrzUPHfng/1K8EZ9rnxOH2CefzVDvj565/vqPszMo
rLWXdKQgGj4loWClRDDwMXQmQO6XRbFWavmW/EwUjrUiCMtEK4xwL49gcucGuzBW
AHFm2yHchgZz+2htmbAgdmLm3F9Mmngs/BpmTuJRGcrERlyabyBkIsawneIU5Y7b
5RtaeYVjqR0iNWChyKlKdLqHnkJKQbUAHiM0PrtvIPp6PZIReHS4e0gu3gj/y9ql
k1uSBhxVTI3y0yOTwDQSFm4oOIUNiybz9fbLd8TACCWDvprzyd+kJovki2HDz8TP
weaU7aM89uXJeANgyNEyPqnw44vjiio2435hC8YsufQpFgNU/lYlTTwMcy8mNYci
rJccy4Dqn9lSF/WOa/hAL7RbylRRc+S8shCivS2QjX7SccSKfW0Kov9n9Zj474h2
a1ybjFsq4f9zqNFUDckjW3X6cHXJXb016ooez6NXZcBRsJ8r1SWhBC5mPtct3J5l
BG6JiR6XDAuFHQ2DrLiMuVFKJTVC8p4M0IoXhqwJCVbFzLMq8PTwUZjIUbRznNAF
hMcWK9IkVhjBe2nJublv4K2/opiTfqXPvEXsOxnjCjCQ4rQ8P8qC/uN3PnqsNIrB
mkBwpLDUnRg8scYF5d7XYru8oGgwKhx8ExEKf7yOXKVbMskbu7qnkq+bcEAglHGw
zonSByVasgWXpvhboJ6YrdSgXfB7pGrA3J7YtyGA64moXydDqDHEyPnTkhDpx2GY
Ex4HZireDk+yxh1mBkq9rHlPXohufyC/0hNKCaqyLTk9tl+QbjhVorLgUiqYVx6t
6D2CkkUQ9LFTOQYMIpRIKfXURUPBCnUOMwvlIaPQjE3+XGqhuxmuUBeqbdzH7BGF
q8kjPHx51ve/qwPjRvxZCREP8ttR5Guo9K7g7Ru1zQVp6E34kLLoDCLc9yFJ/N//
ZACY9hXMw7HWheg17TnVDJ2rgck0aUbe7HqtTwmWYxcaO8SiPtZ0sFEy2Q4QHqlj
An7Eoy3WGSuYRIl+6wm4mmmg/JAydXPFHjKcMH7bZGb7n4zRO3WNKWIKdHD6SXeQ
I+LnmUFWRC5oCSfiLDlwn2ahk5Ttab7zaqOll16j+5d65qrZSCTXk1Pvm65z46c0
uh/IKTuxm3sZJrAYZOI84XRRuGZAXzHfoAsMbcHNGQdnFG40TCTK3KFYIk7fAW1O
hIS9T39Ow3ythAX0vgCwymc6cxel3Fc4sGYmfuhqZlvDUk8UxMG+lX0CVTTMNd30
4Q8pHViV6oLBsJnWufDyNJuOO7Z0SYgc2rDN7AYIrHvlioUkquj+OGSw8nludumn
gVvjiInUZY3P0poSakBbpa5chaFclQlFZ+4M0y3ahOVaz+MvOPHi2I4J62/mKiBm
NXB16SQotRh8PW7YITB5bUZGCNxmJLMCGMrhmZfoNY/zpfeAg7s8oR/tJqIu462z
MH/CcTpV29xNpYun9J5eNfKLnqzdVzG6mUnJgRcuHgEhydN6+ksj1FEMwjJu55zH
VfQbMo5L1ZHPBkcf8V/cbTIII77rTnN/PqxMo0EJnqAvxNQ0rHTkxEouaoKHdvww
GSXFAlMMd598i+02QAU7tQgQNh1uJFrvbavKBDqwpJtGY0buFEtasmhcOFW8bJij
pYevDifP//0450jsAwFJAG9IQcgCk38f2hkIaB+mBYTc8OlfpMwdS8Z92TarOdmf
WfYw9zhejts/Gbucp9p5WxGZlqGdtmK/qU1sENBMf7rqKPjwNCuMglJ7NEmZSaKh
byqJE0yMntRLOaEAerbnuqXmgMIlZa+sCt6ojB5fmwp9jwbzOacS0nTTrQiRrCe/
MnICG4+rMq3PXIYALUIecIYM2dnp1wKLzfMSi795yiiZaDr1eydFlzbtDP6Xij/I
GgGkVE6rLGjWhpO13HIZ8B+lhkPyAvh0g3w3wFQMWsiUnDAuLwQsLP4yWqLeyAkw
EIlgYgCbxKxcienQGDB/+eP0Ermx6vZRZ6/WJlg8K9ElJR4kR+6rRyPNo7omzaXy
FbpI99YA7E0rxsRQhPHy0RtVdfvl6cTFHSnNYbTrVjTgMQSLdCWDrUphstGuCBza
Fps/1NYi1D1yEHghTNkEcKIHIFufX4KxwrXCStlRMSSV/eMKnCCLpkCyrMvOdub3
CjlWf1lSj0UiM9i7JlIu4J4t7E1Re2xn0LOjxd2wbPjJ1F8G22F1fz5nc8KByZ2e
+rRF/S7GLK0UO0asawfgsgOEZ+ZFFwky5+aIj+Til3+tSSlqxN0yltvG/KEnv9D9
6KHZk1Nd+wgujDAPEfvaBGEAoZy0W1ZIBxIU1euACUe/PFNTdVFwpdcL16cN6sbG
RTe1UWFsVk5OwXVABJmhwjq88mp5wvrwrsnS+Q7wvAW7Ke+K2XHyqTxrPGNgWwdP
35ISDF+E7Z+I+gbwRzby9VE8VpikDusbe6e+Wu77uTksNbuIwT5xGD++jrR98AmL
A57G7tYOrh8Td/U8YcfUkkR2ketoxjojyFTPD737bGW/lVm+tBM7OnwJloR4Rdr5
6DA59JVOBUeduz4m1vVmusG6mM0TXyGLkFRxxHtOXJfW7lJcFmAQlSnyIh1SRsjS
1E7eDbE02X+pKbpiBlpHD4m81hxlT/npkgvU4C/5onX5tKYcAtRuJY1+iKRB53B3
ecqqMsLPjoYcq5M1c++Sew6ajQ98ksIDPxHrPBMiXXnv5BMQGrrBLYKBnMPS+4ku
yfKmSec2JvaP8R7hS0UtJwRaCTCe+dRArzvMa7t3X9bh79E7XG3SgALXweD5Wa6B
LRilZAAHz2K5NLiDxFi8nhFWP4UmYByHHt1kipclsVhpFN9H+wDO6jBkC2y/l/tc
LvPKqExFzftTxX3NEN84BQFF9N7kS/b2tOTp2sgRsbbmCGilsSI+ja9pkRsOowQO
pVLDY3POKUKkUrwJ976Oob9WyN33fiQnFj+p4gZ9xidTdGfUtQwSjQlzoEHIXiA8
mzpQWfo/Yebv8GyNrT6HIHN5MF7n4w+ebuS8q9eqRwFcW2Y6TAXwo6BmaDNDn0f9
E/1apxhkTsKJ7gttm0VO0Wv7u19e9gKjN/q/21HyMUESpj0/C5b2qox2ncDt1s42
aybdUjh6WuFhhf3/s1WbVQEVu3qtWwAVjOzDXBXy4vkoQRtt/fQguRcirn/IhPlb
/XiR3iH2bp3cexJx9Ls1/Mvk8S7moEe0rZQ7A63VYsz3qu32fLnMzp4rBn3utOtr
Od/sCnWw+ozTRmlDkx4ZYvnP0yHvX5XspCeA18eozDLfEbBwMhzhWqc0JX9RQaaP
WJjJc0sTkFsmNil2LcJZt9mG0AYnR+pZeS2INtldYQQW16LnGTNnxcGe8IvOOxRU
WMDZ+s5nW3ENrR+YzZw4hbnza74gfsS0GBRkN0UVT66vWE/EojMRGv20S2iUePSi
BypfAYIfDz4YPEs7WlaAXMCUe//1XeLdOdcEFcyU1la/GlUqTWhnnQJaXxUeSxGr
mcxtnKBM42urcxDtQbRKl34JeOFz+NuvpQ7Vgt5jkI+InN6C8wBhPHmeUYvnSK8/
3Vo2+BTbidKXyz5lay0qEDAp0M5pqF+XLud9OjkAbnxCK91kmm6TGTXj1lFOpzfV
Ooysv0c99kUZOuIn+4n0ns05LNzOm85RE7zSVU8yF/Ht1WIcjJVzrCNgWOnwOyUk
rwVSjiwn3F16yGjimf6hW1ts4HF8zsO2JUN5d6inJHM6GAZhVLV863p2r8gqEsU8
MedWE4miKuA9ey8L5e8zvyy+ImlLv9t8AeuQVuDxjZGdrG4ELn0a6iLUB6cH5kA9
4eAifFCY5uhKnOUSxbYQFx+mBS/q3hLcce6jR+OdBiqkMM3gpIApOtb/LOcTUgJA
o9nvE3FkHY6SdOYSuJjriVr0nnQ8aDMRkV+WUTAA4pl3u8vZIg3Qu0MoEWYMrABz
ahk4kop79HyGAGwMhtzzUJtuuhTek1x0vJ6l71y6HW6N6jOYy4iENKxSk/lePFSm
RF1GkgPBeuY8Ad992eDs0MnUClwYb70PKE/JBnaqVXiZxq4fB6jPBhz8Pyelk+3p
r/VowyrRiS1RU/WzrPFChYno0M7by7szgY5dmxm1JLC9V0OW0SItEkseE72inVsC
K/JwBcIEQQvx/uDN7KP2ZiaQcjDYRNqsSz1Y43nQlkcHfzdLynSmNjDY2MRc4eom
84SZCEhcQFHtKlq2R7sXxVuiUhumDSKBGudvagwVmLBK9hQSzD0TcQ/B6jp5T5SP
Z+PvAsVloVpUTwhNlvEAQ6Uz8nlSncF3MCBy/OiKEvF6cdPZDH5IsEl3ax0E3LO5
EaHcjQd6gz9h+c9V6VP5MzNJoTZ1AFWH2yDaeS5TUd85TyMg6LJp9Yo59Fm/1g2S
sstpEvkCzLdUyfHd+KlKrPu9Yo8rx8PVJGdHPe4cwp+DM7eBjhFi3nWdajCDbNQ4
9jAczuCJ0dzBK9SzrmdYebSuVxjNW4eJ2oTnOnyXcHbvmuRVpriGtW6Is0sksrBA
2eOvNOqe4LOUz0DZ87cqRZaX77w7WX3wRSm60NLqvlTGC/wfKwZFmY0s4USZ4cHI
rTekpkdw+Dh36kUK6FiBWJZ0YWsJ9FE4vYltHumxJANWETurfE7MKWs9V4Qiq5r7
f7p+idKI/2VxZvp1DjRt4fHdBg+uPhhrACybmw5ZUGGAzLEscK5gBWbyDxQq4iQ5
rW6NJwbkwTTW+I5NWtLWpqcopzaHf5AowPZDht0Y73QshoCTIrRne5sQMm2BWu1h
Qrv58X3M1ykmTRqHFVuJB/WGDIbmFuHi5cNo8/2rzpEUKN4f1K/+v0XyeyNPK2W9
U/aB4xqbVYXPG1/betQwVYDHRAsUDFclWGLfQQv4yrNj00hu/SEJ4gHXMOyYNYzf
pJYIfvHuL/XU5FYMedLGC5Bo1TUOF0m6lJoF3p4+XiEMTnVP7bc2Tf/tgb61mJfr
fip916l5XYAu5kghmuD+Jy6DeCZJxaFwWqcL4pTOA9o1mHF1U4+LzvG6AEm5ZRIM
D1VgTGFOWuywhI0OJ/dD3hsfjQcfLe0QW2EdZrOOYizHRHXZSR3Rc0dPCCj5VBBx
U7lf5Auvb56FssvzUBPycEJv039UW6ESPGGT+hHT20W1NwlPin5yLVKcbv3U/Jzf
TaU02cD81EIs9k6aBLK1FrknHTkiEUDQI86CQWSFnZ5l6qEibnkCP3wc6Io+LPGy
hs7WXLBjnq5lhLWpLfWWQAOUZOP3y/fROc1zWVBOfLYfcyLAgv7sWAcnynK9NyhB
P5CBNo7CbegAK2rvAFIfxePhnvbk1LLF40xhwcWxvHIGD+zpe4ZhSwnUyb6fD+ps
8uBgZyWwUoUa1GlyzisI8s2/m54u6w+/w9n76Fjvls9XkRiC9N7cmgWDbPYLOaoE
kL6svKPBo93VufrTksu+70kddQXgtMyzPJqvT1hivaXhMdm0QCB1h71b9BpU+Hrj
OjpvQ0OvNmB15BrXUValDZ/xnGiQmtZpHQwgilBrS8iW2BI+Fy8pzGGo4hwn8MuV
DcrIAigRmn6ERnJDKOJ54MUg2602Nj9PuyaPi63pW7cjDDDTFhF6OVP51AFHdBrJ
oMwMSdn5u9ORO2oM8zk1PQS/2pTXWDk2owimtF/M705RsSCZSh0U0GUbMTMbzSq1
GQhM+gnFgy3LvPH1effuU47DHkg3VE8aVTlHmyIyPiT0xX0PbcFPgfnKtpA1J+S+
cLNddqXEcAziZaokJcvjcqEL7bSskOzQ/QNvgzwPpyLH64QxZ0yrOH11AJvUlV4u
9+gE2UTl8tD51a63D4Mj4050gRkp5dlcn3S8ZR/Q+1AHIR98V24vrh1SDhanAOce
wa3FLxUCmtcFV+IiGoV/2IcTifR/Osj40WNOU369WibbvcAWoqeQ5R8mMYh8qwKz
MqciMVjfcX6ilddFnHojdJcFAw9me5t82O30SHRYKPSQPOOC5xsS/pE1cPN+pC+n
Tz9AbwXrJ4D9jcAnvliidIuz2feOYjn4wVCr+df/uwb6i3pvNL5iLq1SxsiWG3Vw
jaP6NlE8sEIqMxKIlHtDSe3Zt5UZHM/nrCRFt+1hvXWXbDN2XuirCjf3BZqfuDdX
qQ/SWYc3xnmtun19IU9yO5D/8nev/Nu8N9B4CTPsiMG3H3DaRO3hRteQkEt1CJJ0
c08w1dSlx+O9SrNdN5yoL2n26QjX6+QMJMf7tXs316FbqE2F/Fap+0vCCKv+Rbfe
h/I2eOFknwB7//azdj3i5hLl1eoFn1Xp5T8jOa2STyphOTmA4a9FbkAc5q6/9O3p
1/vnFvmlRZhb08GD/FpE47iQ6UyzedIvR8PhsEVNolKkWqlE4xWWgDSqedMMyvWf
1mhis1XZlcwIJRbpMUjtMEbvN99Tox5Kd4EJfDUQ4nipbiBj6TxgCDY0nE8CKfvA
g1LADCpRIHB8BQmoqjCLH/iebirD54te/wPQQKl+Zz5lLUTV6P0vpyDjYO0HGIA9
Q29N/R5XcLl4rHLN0A92E+bY1OR2hTrKfsSjJdgpWa8AdAtgyzIvrDQX6RQ9qSsU
KwIjREyDL2gk5LnPZoAsz0sg663laR8ihF7xJchXF1pjrTzGHRuVed1k/WTw5pwj
TwabZwFsQAa+bhVGTjX5XpDdYBLX4pEAn2ghtwOdrpuiOk6Mb4oqhiWNU59lLr8y
EPRJjbT4bXB+Zh0z7LLu+QbcfMTYd+ltgNs71PDFBprGo/Kq9D74zNIenCcPcAF6
Ck0yyT/RjQF3lufrucgjLU3PqqcGizu+57nDMZL3fAOZXcZYUzxsy4tc6BmiziZO
QcQddtsrkFjeehYeQMrpC5Mqn9tNFVeyTl9lI6WJsz7SKTOvaF6Xh5/mlJNORTHX
ureX7+4pDSAEI5PpWUc6bjFP66azzVRrEDYZiOmmZbLYtUPOa0C3+sbEKZtjNtS8
+YKJHEkx3u+G9KloqYySEYH0XkfaZtZZP8y94I8Iq+0+4wpgLogusCNDXTnW6SI2
gbWSmaMsfXPqxhKdxa8kJd3V+JaNVb3tx1z/ZSQ9oW+oXfwVMGYPd062ByDsIShb
GKBswPHyGqSqrwLXWk07BqkfjVGtiMQnbNI3DrLbHOe+MX2BHw6dGLQUjlS1tia7
B1lxT/6l82dvLXY1uWhfT4L/kzvoCwdzuyHSp1O7U4CXOqH7jUECXigwhBc4hUDv
XxOGuU5dCgfGIDCbexYuMsR8yShVGGEADJsiHRCkB5UY+Gnya8RoJZKvg/hs8XYo
2b/NUEzUT4Cz3mtc1jQ+VPnlQrkJZCLH8GUsmr1fbT0u2HeH++mXa4z3csUHx8zp
2ZULfPOyakS2XgMOheJ6v6cfzZIsts2LR7+L5PsMLCWZC3JWomf4jmLSXz9R7Ryd
Eh62LQizbgQHMd4Mq1DGv1jTWAvFsvj8/uK/5EdxHDJbfFKADizVMxm1qwBr+Sap
HLvNCUkEcaC7Q9y6xQY4XSPKWpbDIJfB1j0E687/swjapR43AV8kVRKA/MVTvTeg
fC0cluwP3r5SFpyQmkYPcSL898iEZBkc+r0IxDUpQEv3K7vkCOqKkTz8n5c2QMCy
Pjaj/nEKF/7t7hjVy6iuzcQf63yO+oVQGHxr3B5mXzDz6+rTDCZrMaiqgiK4Tn0A
PTwagsINtimtGgZR60RgP5lyO3QryViaSDkDPC75R5ve3kEke1VdRKqu/YWkkbpW
iSCDo/AePGjlfReqthP+aUnniV2+1wMq6rOYkqvPo3spKKYYFeWg4OC3swydom7Z
vkQ6wZr0C+eBAXaJfWqfo7Yp7ove/fAhkUsRA2xVb/3IiysdLF+xmmn2ukUSrlmK
CX0YJ+vCdxhiItUpnXwfDcpqphm1nTRZr4E9svcDg+L9oUgmc9sJ/hs8/a42KQbw
m2WPw6JprhhJH1m0fj1C9n1dFVSMP1hCFTknbkC/ogd5ZEx10HMkJ952EdUnfm8r
JETxiRa5mArAfVSsQTpZ6uxCM4vxqMhiTxoxT3t7o6Wrkq1mKX2m2FvUkuKPbIqN
skPJG9UJb5w6KN4AMYWn8SbyWszQOzd4FensVDM9answfIUrm8u7yWaip4yWHVkc
gX+Yyb6PlbMvzAAPKf1Ff+D2tU9c0ctSRZ+rpLSwYsFeIMxIIAZJgeLJ82Uc36FL
i5lSiDFCyb7bD/dkH2yRIBPjzFN8VqfOmG+pR6ZzY415vzT1FAbAtHbLOrsBpfoF
O3YuhJj1SAFqCyiOjiEuN9BUVDMHuvDHrp9lMkaAuTwaihRgyryKSfg0eR9WROcV
/NX2faubfZ/oEYv4+G++1ihW+brNqISnw7smcyxCsnO/z+g93IxWRPU/ygh5Yh5+
WXDwDm3KCTGIpkwaM9WjZuiWBSQ4ADA+HvJjzkuZt/4x6SJ64M+hiq0dW1QPgCcw
wbzg7OjL93o9ZbCaPCKsxvnNrgP5byEELwGqs0LDVmWUl55kd9pn7XCaivtmCgIU
EX/OB4cEG21lZJIPBBRaCUNoS4A2PsC2gOz1RjY8KxZSNSfPAKhFr6fJw5IGiGC9
AxLFBdlj32gzr5tObPotoRZGo4WRKOSG4E4/XXvV4C99x/NRn8lAhTWW3P0P82/R
c1wQ50emIf785C5VVZ4gPsegEPrdT9QWQQeOLlt/mwr1fgLSULOrKiGH/Nl4KCi/
b4wXw74uM8LDl+Z3L0a2TVTylLfcJkaeIfnAFoxNDQduzQN0CaZJifEytZ7Taxa9
jZ6Xo3cfmJZuTTflRukcXBDy/lZQVmlknrUM2Pip8cSN8K8YVaKDa99f3sjdiHP/
Ffha0KtJkgbUeONPoH0OnSThudsnmPFjul6qa7yQnMlXRvEt7dDISviJeb+Xv+Oy
+lDGCfj12WWlqDrbwlS01fYH7rR9fhZVwvAPF3hikR0oLRY1USg0L0k1z6YhJG9U
NKBlS4MhNwNWtH22hTI5kbMSNj2lJq0pk3m1WQCakg93JFW3KUSSOqLWLg8IwIfH
Cmh+Gls1zoILVvDg0vDqiPDHESZEkVJkVIP0eA6SZqblV1+7cpNIkjmUs4Qn7PGY
VRG9qRrzlR3xrRmTu1nnfQXYwi+auxJY8FtIjWVRVdhmPi8acBaqOrjst/k5KlaB
m/98ZQt/TbYQTd38XQORfIxiN/86E7Tfp/3eLl3yk/hLowODMiMZeTfs+lAkHPhD
agvU9Ir2kcHaT1E/3frTaYWxyRBO77jJk1KCVdCbgMvxsjXxPiAnCM4mD24JeqDw
DBed3gdnC+0H7B9Cu9SEGjL5ZuhUnDsdaiVC6xWnHnXmikiDlQCBkuAduxuKWsQf
fmPBA1e1DE4RoTRgYAzRU7ItEu6I1yKVJ5WAuy4kb+ayz3uWp6CrNnfOxkp2zM6X
5ki1cTAcChc9lJ9i5elfLDd/9rdZHqrf4gOqc8usKEANDbyJywx9GhYfF+kUtwrB
xItd1ehzWnerzhadUOqKBrnMwopV8KQFN398VKBUUU3Jj3FeS5s/nm6MYjvAPCUw
vE+0+H/b/mNRfd00y2GHyR5QGZK318s5hXYvh/1Dh+tJfq/U6y1f0NGQJ26AzEOe
pc7i14GvqAZOJAv/1x28NywplCzigdjPwTlIz9wTRm7npZQpgHmoD6czj6TSU8Qg
phjazKLejwenTWlX7/bp+R07/jSHsxZYS3YEAX9gMBXhm1Ckndm7MpbgmbD/JCoF
OwjrTRNgXeoHnnYsCLDXG/aOu7YwiTfG7KjnJ5q80lPgUej3M72lg6XDibAVCQAP
PpGt7cQ+A04iiigV9wW0gZYeAwTWGNnMLMWzkAgIHGkWXE8FBBqutxpHRpQfSpTC
GiIsNQJ2ym9HImaD4OCU0Sidp1vjsS3bcMZVdlfH732hx+i12S98xFTp6r2Psf+u
16jFsNLSaMVN6SOJbpLwI4QThH+Gw3ZbP2tFLzqw9Yep/i+mIZUMIMJcYTlmqb8O
7WmK+E3buwBLsigrHDhF/cp0HR5usUMBl4SY2Bs3APud4nY2wZjOvPW0JI/H8CBn
ODlDIgj+ymmIIPCQ9iBxbmf3AhRTUb5M+pi1ksXci8aQk6R0MbfYZF/nCTPLwjXr
mgngbuPdKeNKf3C2tUS7LJuv1YM6ItLIbB6mwpALD1XDQWpac4QBmspQr+xMfLKh
M+ynapdCKIKAK60ASXHL2jD+qLmN0I6gUoACqKAgcJ2fqsDd7K/59L6yfFra/XOv
99Fn7XPUWmwhjlm5+gH9i8+DeGspdqhPyQ18JTgNzCHWBSVWliXuV1QZAG/yPeMn
32hXPCleL0RdIHyOcg6D+0LFD1Ia1EAolmAZ1oPWC2TDP5MEPptrXQcUXIbciRtB
lbgbfwAqaiIPo9PQgBMN9LmV9JdOupITy0ke4Jp0rzZay7G135VbnGHLjfi+eDjY
lRCHO3Ea3Uod3wqYoqJx+V3VpVh+z9ONdS75c3gWhRG/NUMJ/KuDqRcvrIvB7yGS
7vHf577TIINPw1QNG8ORGlRaM/TXY5H75dZSp2aVQ/axR1qmDQBizKs1Pyv6XEtS
Eo+ufe1+k0I1zQZtFbf+qqRfSbppxwOF8kEo3QZyaMeiroIdFZtYRkmRCkXiQZrG
+MLmDckkH+BojZEcQUY9y63qOmqn9Y5Fy3AbFgRO+NrT/5iZTPosIWanQ8V87gVs
5xzJpxSdEs2V1WggAgBEQSco/aMRY9Rh08kwicW8uK2LQjXy26iNyCWlLJslQeX9
N9gT+J2ZWD8lciMVVpWQeO0H2nVaN8PoN0zgD9+393oMMFwbDd8tjKhBVOGsqjPB
9rbBOwX7nHdMBRramE9WMFEAjjf1bTUdbuFj3ZdqFNkT8wxyv2A0+J7gOu2xZxmH
WVG9/KTswPTA0LRuIPCP0Ux+PoAOLf6XqVoeju7fD27gNP3OACoJTsDySHydU/V8
s6jz2cHtDaY9CrGZzftSga2JG67x7ADueuD19l6sMH2/GS+Yr99ANW/IU6JBgjjr
NIrWxBKmNU0MZXVPESW4assGFor/dsSuFVSYhaOCIqs3CHwZb8Ve/mlx//6g7uLE
9I6N+vE21WL6Qp1DDsXNFxkF0O5G5E9iYbACDS69id+xnljQKhRGdKcTJOUcKPoG
fTn1B0Sjf04+jEcq3p6VZUgoz7nAhSkIG7sdxIOGHHMVQhcTjepfoFvGf/RTiAXh
0n6N8APq0Y+PIaptRSDrz7HrYqxXcGnW1NZLvPE8uSYIHTiB8B0eZMUjI8Y8gftS
5IOw289rHLTGJYq5spzq091waxzPCt8fsFFucIlN/lp4qgMGWFxggl8cri+J9IK0
jZVirKAZzmYJXuYcdqWP/5RnUzt54acDWGfTu4ltDuZIwlk3lucgXc3ZaRixGKx6
44J3ROQmWAYdU/cdZ3/Ng4b9owXx/5Kr9S1aVCN+nohvpiFV03POw6zl/CiT/bF7
63Bx5UcWhm47IGwAtZ/F9WHVC8D05XsG8GaWcqoPNdvX04KiCd6xwzb9pi/478XN
8k2v8dj33RvSYQfTChxjUrNoWw/y9HCDYZvusvq4XI9B6z3SuArR3aBCWJYs39Sv
CuU3KekACOh0vdRbQ19hjKujD02w5aTq1aRkRQRVSrkrEF3MmnqG5QKNbrm/SEnq
jRTX4zD7PMGIy+P01y2z6OsyZb3l0WW43wi+04ga1UqHqq2/zwrz2L1WPOSMg3Sc
SLJQ26AhrSJSu8jPShR9hRRohe5dPtwVF82uzbA9IOVTKRpY9drsgrJ7Q2B5LiAV
SLynV4434TABa3akoBRFma3922C1xz3lwUVatsnHosE7i0REyHkFiBuOMilQtRi3
t8T3ahHJCf61whRLAE+hQCgRKjcelQxRpsqbI6XaITmDA2u1TcSCXh41OBDLRH6V
VcEupqJtBImfGWHjcpncmCsoH94pWdDHlNg1eMcQgv26TR7yLVAELH67M1MKEPWd
pmeJxYg+DoL36z0AAaiQHDqbogfOhA6bc3qJ3me7fGwKleq4zv0CZGQCsTYVOE5c
HHhpZGOZm/wokVMJBNvTXFkXxi4LIbn/BfJ/B/oBTSEQKO5h6gANLZvcfKaVMp3h
uGRgv5qrzFuPTcDPT6NDqj6uJCQ0ZjJGAfzimH5dHspwXds1Docz3puTn5aKWga1
T9GnkKk3PKJzkjLHooZ09uqQ69llDqMVEhhYkQWUd8B4ZUD4CA8kUw2vZacSyZ12
BCuzB2vJoc5THX2cB25Jtv9ygNAPgKeSFu5vS6QQAVFbUExAyu/zupdELkclM6rm
WftsZ3vN8HAnUWvhdC1jkZ7Es/IeXTkAKGYXj912HTHtZ/bnaRHgc21Mp4MA+AkY
2p3hD0sNCir+uKGOTATzsCuUSYh94Tme1l6yUMQ6K4lnYegqM0wGVQPPQgtkPPr4
BDNI+J0BhGVCR27dukCSDraTVHK6qwfMVCh0BugmlOaUZPpETbDyaAD2iOW4bye1
OJbZwBjL/AUXMFRXZSpCFlwAw1AQEjY5Vcs2ev7K6w1yR5TWIpp2I1qb4Pe5dTpf
KlO3D+l+rp6TOBcDNoCkz+rHyYoTWxVll8pNvouXWiY9j8TqBqYzuWuWClDfoDPv
WzDiY8w+ZgwLHbZXndtjxaz0wLLdUuMjyR5PC9M9U/SwxcidfVYiHQuG3FIOLmns
Hf71511POkCX7aFXkpL6lcb7qmSnndlwr/lFN2kV6aa6/pAdFWjY7G7cEfdbOszX
LMjJDXTkJDfvvrBJ248ava7BsQRwTLJ7IcSEqzJzeOA1DesOwOD89LuKGo9VCf79
GTP6bL84hggtSLj5tarkIS3JOd48eTGsJgHPvnPh4nGhMWoI7Pg6VpKAxCF3LCQT
uqOFdBWJP9gsntV6+8pFflmi4gAv83A1cp6fX72EbSjxSCUOgpAKjMrB2qEj07Ea
Pnv0a0dhDfH12Mj58GUYM4bM2p2JvHIpkKdlSIp12GdU68c7faMKzWifO5LcEVTJ
+TewFqKVgM9y2BLknzeOoSs5H2xdIAdKlpfVzo5ndAYo93ujkGOYTQFc/hsd4p+I
Z6yJeDfSfPlw32T8dQh+FYJoZJ4K8CPMM4u0Zjlo2A0vYW8VlcG+/5W+Hj35pwiR
ToLwnG+y99kcFxtS1mFrAsi8S6G3Jnw+lBqxzlJYrm0fX3wjI6035ClNp0RreOus
fCu5HUcefCE5/YgwfeP8q2VR4A2+bf8zk+bQhvl2QOwWnahZGsG0XEajwpcmDvdb
9WZjbecDHtLt+YWITk4hw36enBRKM5lzfQDhZnYYip/IwQWJ6D7DC+Zr/a1Txs/+
IUztrExUK3T8grwhsoRwMB/1w4Y3V2oNykxPszpGLfaeBprqW+byT7WaZAInODYe
p0VB9TeTyrnHkw8rVZEfhzNW/jM5NxfPcXWYoriNLqNDSHQjHGuJAPuGkxz4/+6I
BMR5GUsFkxtVtNH82owwwtVDiH6lnwZEJxWaF8JNybHhgWkyZC7A1Ood4do1H/M4
wEIuDFMbY9JrOqEZT3MmbkIT2Sc1qY/YB8S8yjgQTDMMPxqF4ExWrLa4HgdE9c7f
UTXSoG/8vaNPdXvyWFUHnGmHWWLbExcjYRpSBvlZ4HGb30QjzQq8AGWgIhTdtx0T
38U7oL1Ht7L4L4Z0Iu16f09HMIor9E3jjyjWz6AmWxbg0zjsDSZBEeIpEuW+EEBc
Rmq9rbfFtwMCigcjkhX3MzLlPqz2xX1WdRnFDJt/K4N3hahA5cXoO/hbB/GoX3gg
TZ0xFhE0Hfm8pTcozGeTQrutP7bQr/ice38t9VCDgJa6sQCghwVCEK9s22/gYZJS
HW0HJ8qVIx7j2pnihddDM0XVIlubJqz8FZfuzI4oTiEIlQW4XwaEG8ac8A1/LdW0
7mZiUAWO6yIEuQ9bhv0/+RZD0OktYZM2TkXFl8ShJnv7VAcH2yksMnY8cC108A4J
8JyAW2tbFJcBwqvXTQPZX+Be+PINztS3/wXmH+O+6GMd2yMLUMS0nwRdv7GQFWBD
o/R7vNEZ7nasF8tqEu2HYB7Zlon5jK6stzA5jiOxegdY+k9LH+KY0aolKq8YBLRa
mE6jWcNM3efTpwjVE2C/AKm/1jUHj1teAo6SOcipt3J7ViMpKHMi2RuvbB+b0w3O
K4y6T5HhaajsouAExR5Dg4a/DKZD3FZiC+7Snt40MRb2UJ7do+ZmYNdzRQwLuagK
FkFOOKc6nbJonmf2ncBRup+X+iSNUqnY5npQsttopCbgpdFDuXUCJEkVn+YR8T6O
kdQ/AvULRMUWuyS2I4QiWtYTsfF/tNdoozLbrpDZZvrb+hDaChHOTbATjrpNu1xu
CA24kZzXsd61ocT+EReHklg9aW2uVqPrww+aTerjbthPJFMwahNKiilhomann3yk
Pzy4gel6KxaeIYkng4QOXKaq5fY/k4DjCun+zQoaKtdu7wV1dbio8OSDzeUO/Qth
N9umxLQMVRLMLq5u8QIiyIF0ea/B9IH7Kjiyz7lLjAdcknFWxATAkluVwJotyh0C
5HrN6UdwqZJxfM/InaPG/HCoJfneB5mf/sG00FMZ9ovQs3p/HZLU1TkbpgCvoV+t
3UEDWH5fk/FT3HjIXt8Hq2XHZ+NiG9OHOilGR6CrsjDOVccngLyBbckd9+ISl1MN
KH1EAx1BT07oqGnmXxa0mBZGR8+7niNfnWzLWCYL12tPHj9vZVXIpoThtQdnlPQW
uXugTYV38YrJTsATvRKdEJcV7HaSnkOl7kD81U05X4ZFc/rlzybQ5Vy4k7r89aw2
cjtuOTydjj0VzXGa6b1yahAbxD0hVpSyL2KKmzVwQDeXSMgCRIXASzzSQV6dA2zx
McGAJQYKIBoL6Yewtgqo+N7nzywTvC16WQbUt73e7Rbz5SgeGWBo+NqB5/XRnJop
6dRKrDSBSo7r4OjXd2BBCTTHKIcBfrapegiJjktVISQZZOIYKjUAvV90X+YJg3kA
6WOa6zN6yEYn1jArctgj52xyiJDK/2pSo7bBKQLZUxWUxxHq7BJNiyrPLPMseXeL
22I4Bm6nGojroEkYHOUzVSznrFQYKtW9xfDAoYb6CJjM/Uq5ye0BzOzUi60c32YO
8HbhHrWpoSsB2hu+DY2TMSTT180XKm91L0wKVd6iajtoVhmHGpm1nJ4+nQX9OU8E
nqkjrvDv9MsypE5kjRTONzPBE3rF7ivBx9aD9LVnR0JZPvbbOGVCONj84Zaa1ioH
9rhCyVplwbuo8m62O8rcxBogX48Qa1UIz0Occkb9U1CTP+dLQTCjw8j2hXmAYE9X
9bw6lpsh2Y5B5piCEYelQ5tapnuOY1Cduy1ZsATFc6ANpYxrM7o8OPyddbL9f1UA
hh+eVW1OGoW36zeCJD7ExyQR8NUez70Lq5YstGeio41NqegVrbK9+cAjj5jSnPV1
H8HDHhf7lpbjppo7dnnduEJk8nSQSTTp++e6bJlBgQXUFs53GmiGI7eMZOTD+osJ
DqUqxOws8dxsAKIMes9dOHibqRojPof8RfGAHNoF2F1F63Nn2XQhTHmZJVTF5TdW
XXqdvAjt1Vp2n2OJG4IwLhYbxrTc7ExxsCXIFlNU/dWpdX1GncL1z2mNvAV6uHBy
w4WVIJCf1+TuEczCtfNRONYSCBjVe+P5pc72lQmwummQEtSLmPFZd8bZYViEEuDi
4gyBXW6n0RftZxLZHCDQVdlHFkFmA3IuHHaLGMVQ4+OaSQrSQXnmoJL+jjooZXCe
XPothNr+NXRMIDc0VZWGNksOaT3R7LiT3MQ7zDHQWmvf+RgDC9OwC7JMbMlp9UH4
Knq5hHwFSStQakov65dBUgJYQAboOb9farLQUUMHmRcRdSKDHh9nsKpXZG4bUc3t
B6rKLON0K4QdbIKLuR+C4+kGD7uTjleZTqsvjXn+ofjR8tcNmCKMp1r+L9eFP4eh
HF1EjKMVqzK+f3ocDn0/Hx8dbk3vUi17JsF497AVGFBGsSzbVUpOGVS5qzZ/+leM
htdVwkLNpvBlh+3y1WvmKi3MnLVByUZI8rpGOwoa2nKEZP8OAeJV8YKDpTKrcT71
KU03rpq+DdVjdkUpaevFGDVXiixados2BpgjqJly9uOgdDTDYjKo6ukTHOB6v0uR
27pmLKrHRca2+FXCyjSmJiDjBpN7nI/b/txcDCwbXsdfWhn6JArhzIRIlN2tITQS
dELt6XCiHw0bC84lWod9fSiAT5/dxtmiBx9U7tUOcATpckYVD7m+oOyZIHjaPmG8
uCvg21z9HXFTDpJ9JPEpgywaTL/o+2lySmJunmZx05ZhZw1vRj3QwcGU2iN+QzOq
OUj/KSVIwibidw2FEqGJDttiOTuFRUJ799W11t+677l/kAqWS5FO4DwogMmlHFiu
Jttp5P8fbaLVruJMyYhWiwqzODlIt1A6Je+B/BK+khnR86WXAGEYgixs8UcIkcSq
/VnfDZlxHLoBDg2mpXiM2AZBaQ5eUrvYWL3p3ENc39kMtFzgQeiDbQMwSNTgltCQ
h3VjbPkZjITF1pxG8o0d/5omM0NqSwdkjaX5aLUd95NO/JUmhz16scmWNxbZjBlT
7uWayQEq6cbsPGlSbERfmDARZw5aKGBhyTkZxyXLUJvqKdqFswokqDUINENpiHn5
pcZghOTTGq512qJn1nSvkIbr67KtRqr+iB1qNG4ghDDe/xcntgTy4VV99lgzmuwJ
1wSm7d8aI8cLyxhmE7dXyRdFN3nuvN4Dcwh324A5nQqjwpVPU+0priLTMfcXXFwC
sPPcf/Azk0F4xLfT1yBtCzfLhP/kMgwG27NzCLLWRGR3drshMzeQ+ziaLgCatFvF
Y0rAGQqUTNUfSMfGE/AC9w34X2ZjmtSNYGcTU9zsWqG4ylOyMjp304z2H5fn4BYk
CUdMzIe/hytGiYhnuVpMyTS1cXChJtJX1tkUPlJQRjInydl1eLcR+r1ZcTVQRM9Q
wI5OLOB1RBYFpDk8MKHtoRFPggFSGtihUsq3zm4MQGsNSQP0GvZvdlI/03wwh1Vh
+2751+3QPq60fceJPep23SiUVcQcUWZzrXsMUmbvFJHEdhjyoEUlexUlKxcRn6AA
Ntia9EQ+q18IDO7yy/f37X9M8cBGv3qvl73Dv4nPr4EOLlgRYbmZsLLzNvDRYV42
qEBRbqFoNb2cB3O/wEdmwOh0qIlBKW1M+fhF/GoCIhua0n7PLHGagHlRCnmG/1BR
hv4jS247BRZiqLV+P2toF3bBAqenWxnNKlTRXipx64bhMGgdiyybwHa0bDyESyg6
DLx4BGKyHcsCU0gc/GkTAarG78LCe5mMQ7ttCW6JX4XfmRse4gBpy9lbtxIv7M1E
bojIowAFl6B2Vy0/Igkwhr8zvlg22QQKa/sCMc8LLc54xlWKstur2pm/JDniHt74
V2UW8EKzO52ZVL58gC/euO8uM+idP7mutGs+DR8TA5Ky4Pan8nWHPxe66DTLl8QL
52hGNN5ihOx7SYCcbyoA5QmmbmkDmLnAt5PKxj/BDiZVbFR022mQjCTWu0peVRdX
lBvmgZevSK7wBpnq1IQNfjlvSa4Q/WJqelelTh16zfnvtT41LoEfHDTBuVHWcUTJ
VAUcTrp263lsrB2AeYUAlt8IhJgFrdFNVR+/9PgAIzyM/6TZUUAvdyK2lAjvtW+/
adKcOatLNqvXF8EHNOnHQo0boALT1pp2/qld/TgzS7GdjOr2HR8bJrs6K8cQtSnc
cd20OwqB0Y3dOSOdWTnUqODANjAJGtpX8e32T2PNUWF0oarCo8DCr1uzLu1ps0Qb
k0lz8fO6+oEImiaevrunOsw47OqT5GVs+WXfejpBfCyYd1b1W3d/eaPw6+OXc45j
jJehE1rhUAiPAufniQSWWfkFZRxOLxJdIa+YXy5//UuMTmBDS44VmbcCs7dUuhZj
7zyfR3NvCRbtFfwFkiWjW5w5GsO7Krh8V31AwXH1oST8Azj2Q0I16PdMPUQ+1xIr
J/fRHVCNY8G+F0JPS0UzeHZrSdF7YvDX0I1jGnKZ3/YvwLSCkmES5AwR3yix7e4Z
ZklG8emJFGoYqAbFH21abjnCdhKDiKM+b4jwMjeNYBesfu9EWThVp/mSbHs19lU8
HhQ6/nXSCsaOmWdkCGu12KLhCvKEs/L8o3CZhP4FAa4ofkEpG9cLG/lYPByMmhRX
/AOVlv9iVCNG3+ECzo3CSU9PMaFlsfPlJBXAkxgTp5z6nzjEbf+OujgQ6DAwN+9V
6/+paxz/qGiOFYVlt3qtC/nT1Tf76960pql4/95oJ1NZ/we18LfVrNuhY39PI3OS
b9NAwvT64rjNmmcJRrkTeI6Otw+/j9VgNkYWOOQPRdk2M/4/iFrBYurff0NaYDoc
Gr3W/rL0LDR64iQShZOy6r8pBoD/CcrumJ8lzOVeAzECqvId1IMm/rW87Nkroyfe
zxu01Kts5/cGczCj7qrVyW2ehwOPoopqSy8Rw3OATryOuA3sgvMc5POuO4DNuy1P
yjOS+HRX8/CWixt+zRV8tTc/A/xoelL0c7IwEf1kbNbYRusc1GLjm897F2+Hk8Hj
GVK5134x+zs9ew7UwYjNrXd95LA8ldNVOmT9A33T6EdtsSJH71tPwu2mWN03n6aH
haMm8Rg8hITi9azsPpiTqo+PLn7IIACl1X9uUndev0IY8b4qwoAqfP+LTWzDEFsj
EjYzgjqrHJ9NSfLzYSzaswdCRJaWQIyXUSyEYs0ckoN5mTOUB3PRzyJkcLo36YzZ
ZsgV/S/eNuSLmDn/IcRH9WVJ+2zK0Ggkalfe3B0uCJRhlwegZECs+YZrLpbnvmrd
sRWoO8Nsuj6NA1U/qyWNocUXnniKQzD407YB4RzpU2DQ4MwXCi52Ogf6XiwLaSBo
3g8lt57DA079qiyPKb3o9CqYdBv6dUFHWllzL2qyZa+EogHNAr5Og7cehDacMyYB
5r21fQJ7xx3n1RcDGzIkaMAtV5Z8migz9OdonKdOorViMkm8UPrq5VVz8l46tS2M
y/vMZnTojl1d5R5SOrzNA4e2j1rlsKzpC4Sez1r9qOx7lyv186Ib04dD2aoN5kEG
le5o89kTAy0DZIfNwwkRaxQjgvOkTEXPLy/UN8fd8J4cuQ6IpimP54Kr2MnlKz10
XFpqk3cwxONf9kG0vhdNKfhQ8sUcizTEuKNKwB9zYxTLgSlji57BFw0AtoDBrW0J
VT471wSWj73vtc1u/MAz5tYggiAE09k2RpJa0wl/p2Yb/mN1tG/Il+dJFuN+qDZq
AqRy/J2tuofuVb1d8YnRyBDaq7K14GkP/yxYxbIIvkt2yUeWl5Wc538I+PVdMLCM
9WSKIfqI5XTrDzCxoOTfu73/IHoddHiMQF3oRyblhQOHzJ3kDqHyC1g1ux/4ST6D
ZYyCiHyQ4NdrdWvTEw9MXBg5M/9hBYIDKanO4OT/fBJu0cppoInAHrv/w+qkumic
Wxu9WoqfsvQoKeaQ4l3tjzn9NdHpWUjzvlka1JEC37mRRMRKijeoor0TMT2JHqE5
seyCgWQtVXuWd4x0v1oOmiDR73Ft5DWQ+P2ADYrJ8x82uidJ+NhQxe+q/WJMtFaB
q9N5uzSGQaPYxN1wpa/cCWkRRYsXx/TMwEq3NtBgSe4HQurRKdCNaMNlR5630OTO
QNXwsyDShq+muoGKtuLFD31laV5hZwUTTWMuAApr2jUd+CbuyEfylXQWye9tXpWS
xrKPDzWfk8y1/4PyWNlnSudLnvw1w/prt/0zgkQwBZ3WepdzxvrK0PYkA4p0gmSh
A1fUe4lqCFpZLnGbKedx1Q+17Ey/HjTbQKn5xLe8mBvok5g+Ffpgc9rGHqlIDpfm
tWTFxwkgTqRyw4yV998EWUZ8fMVMJjIJw43foqObQTV41+8DXnTGY/CUZfBrUird
H2CCtMtO81x3Da6Eiswt9PMxRIvE4gLzXfTLbcUB4Ayf/vdEBgelq+gRbv8bRun7
dJ+RfiTv4unBY9NA8pcfLQ/uQEIicCOaXB5xfqe2IEKeMPKP3rK7i2WKkqAPLSuj
o7VPdQW/MuDPzLp9VDPvYpueUn4p1cp+xGoIcbJ7af5dlIN6sMgJqAp8+hZCXFvh
o2/9UPInkaRiHv2t2tW/G9c7pzS2uMLmf1FrTKNasCf6nH0hTwXiwks7X+fjjO60
WNUa33bf0b2UAtLgHpELMaVWGm4ojNO24n47xI+wuh4TNr+N68G6UumFaDg8VK7D
pBz+6offW13y9Yu/Vz32DcetuIIog4mJNjmi+Oxo42PW57plaVThLLscYKlIJeK5
KbRZMrWNBdcz8DXjWViUCZUMkjw0ogMZtTlAtimpzEu4zLRQN3ekdOvYXlff0Adz
lIN6/C3oZvHXxWzF7BUbDvU/bEMQuXloEoDSnIERkET4xF9IZ0peo+MCL//yQWeL
Zaj1Fu+nyZ0D39FSxpuR9I48cfVGaGRnV1xyXBxYBUi88WZFiOuWmdR7VwzTOwRF
W8Hn85cSbOyeq//hvcrNUpHdgDQ0Tptpl6+5gr5WYuGhzvnd8c/++oAOnwKqrvDL
9IqVWiDdUs68Y64xVS/nF06RclyKMbH76Bd8OfD0fM/sjcSJNsVCu9K6GhC3uxZP
8YPYzR96uArDgGVQH5uaQ4JWWGD3AIyopzd+9/JnPuCo/RqrI7+xcPU+W73nztxh
k9GUVvsTuiXMq66mRT7k1GngI+KiBUHTQ9C6fSv/TVbf4GL9AQiqKRsmZXXCrNG1
NhfTmx+Bg6og29GRHQGJX3NrLnZu/r54Yq7iqYcRJZ3kPaeXD69jDsDYKql7tQnX
e4ntrXjrVaLi+3WnR2+lv8v4RUcBKxPog9et3BUdQ+nsC83Niv0s5ceoMxItMUBU
IxjDFeX1gwPNcopMYo1aUPAb8rwoh9UyqLObzLK8+kMZO5ZA2AGLMMYi2Ycav64I
x4db1FYapW8J/MYLayWjTpbYEIyZBlE5zaC2c8ElbnvILZ6e0ozzZ3XKFCD7n7IZ
MlFR+NmvG4X0LVriu4E4jaM5tDtWHOQKJ2ziCRM6swN1DovdEn3X/6pc0ujhW5uy
B2L9zHY54YLjrY5qMmhdjGeegStznLuR9CHqNW6hN0dDfk5Lg8uFaygyS8mSmVG1
ltvk5n6R5eFuUL19h0iFLD1zGo+WElZqw1uAeh586SEDzTxO4T3hXi88i7DA258X
79DxcPi7WOwnU3aTTx8Nxyn6RzjDUWlIwzJMjQNEXOdBJcTFI4mIT/tIAX5bCeLe
GQaLw16tNf/t1xBQjBSkqowbAS8APnP7V3Uz48OiUR1C1+Bu5QD01Xo7RewEsGQJ
zeSGoPUh2jeS0lZGnsOZkIdEBRAxRv3JHlUok9NOLsXDiirX9T31qe2mhtmSO8Kk
CYIJd2FA7F75vlOrzO8jRz235VU096R1Izbre1DiniRMqxI4LnPumaSIMYURax7a
+9uoskMC1cHsbq3cnIB/LfOSQ/F7fQdNo1i4WqjTyyiwtUC0raVHr4oGPVCw6W8T
0u84h45p+PRypGTlzi3H6PAn6xqfRJBmYTkCuElqtb6jr2VI6NhZmrOKRtYaNnfP
KOAgr4CqE/LqgYjqvGQL1WeFOuPHyl2bzjzZUdq9J3v1NjIY77UoNpkkB7tpnsyl
au6976Blhb65W4k/85RPkhOnyb1LXpeoy/RLGbX7B0GqAgWWUfXFYoQbKW5Ux7Y2
97AXnUP8s96J7maHOUPXYuau/tzvODy8Fj7UARLunQ62ZPkGFJWJcZLMNPQ5Dq+1
fidJGXD2zbLnHNCF/4ur4jEKBGGquam5Hwa0CX6fnxKIjGHVcqAYiGMxsPHiqkAQ
gk4sFUKm/ruEPgALC21Gaoau105mUttiqUOohoX9KOiSsgNKhvnkRc4ZkWeLfrxN
g6K2j0pC9uA1BuYEYLSVclMFi6zHc6ZTUQQNsWPLYG+z+NAhmQAxdSOny0KJH6GZ
UHwOCQS+ek5Q/uG4OFDFznqNLoQFblxM2poM7JHDwZER+6yO2hNjsuxh+HIMZtjt
DjGr3gpCWK8ZEk+e9PRRrHxbcUheT6JEq0oeAl2WyzdF/ht61GQxlJLOfQvndMNO
7dddotIc5OMxwFMyfVmDKCWLouA8NsC9M6jA0O6zXiIgbviridBkWBxCYQyyWnq0
XrF1ZL+9PIitPFXPJ+3MP+xV8+k1mkR3qWWGTlYaEHAwbTiikgu+mYLkc39tdYAr
MtF8Lk7IVSTZuJoILyAmyuuBUrL00XfY6Oj4btUZzwRUJKEK7KoPjXhDRhmalC7E
OtaiKM2Jy0C42vaiWI2KXkX2Bduf94VcydU4NFH084P4zimbofTO+2HTbFdY1dsn
prexyePlM2Yp2wSE1OmfwZsFchm28ouQtjW6CrZyvWCztWcWE+r0x9ionRDNl4mj
JrfZFSmqwDlZNGtek4xp/PWf5lUKXKXevpMc84vpzqdTLM6Hd248vgrgQgS86pti
yiGZUYmPbv9ynhEphi43xkgHV2qumB0tHG0WVa9C+hL1fwdCp0VoHv5RotgoO7RH
rBaedcwReBNH5AUuEBXLY+DhWmRvhNQZzScaRBIU9yOfSHxiSsAb5oXMlNscGal5
LFLolnl/MV+leq0/3A/Cw46yrrFPQdVTi3hOLd8KD+7mnAmN6Elenas5MmkA2M0G
CjeCbAZHGlFSOx9BMnpr1FlgwMx+zEWVK91CNNF5hsz/Xxu9ANKIEuXXVnukgOpR
ryIquKH98TUuyr7HqD+CCzNImD0nEad8AD5YH2GamQ/Vglh1G0MUdTfUHlkM6vk4
Wv/LARARCaFgWGhEvd/294v9qHo6ixUW8y/PIzZ/ycd5rUHBIzg/4cs9jqzzxktb
x0wXDCXwtA0YdkNyxwryjoWhkehPHHVLFu8Y18BLZ+E1lUj2tvA24tXzI9GVF5rv
pZePAep0FeXATnTuiGd2UXSizfSQ0LkfiwrVdL8koEBkZCI74InfPbBKkR9x2aPu
JVNM9QQr3dY9V7dbpBpqRScWD9+NHd12yMhQBGo4xEQokuf1Zra0LJQHBRLMDvRX
ZucGygoR2PdCUhBvVugiELgq6Xf6DwWxQbHS1fAohGn/ySGfITJrrr2DUPdDga/b
ejDPCJDIRPIF1pMu1QzwI+6GdN/Zr1BjF/3qyTOjzfkGElzFvint2Lp7n0h/jGGN
easO5J5q9eIPXPSaDowlLgINSwiBqVttoxqYN8nRihb4eF2hy+e/JUbw5K5OHwKd
+8XI4MB+5ch22cFOSMTDax8mya3QGFyVv+0RE5f04A5t2RTkV8UMQG8xplPUqdbv
qsehEFpLvIqekl7QYWLb3Gn/9ie1bwpfAfl9x0mGEtccLFmz1cpgjLQ5yE/bBddE
M8jIsb0kgn70vXuyBUVBkxr8yOOQCaPATvEj2W2hR8nVMd1yq993mTyxHq26BL89
6p3KBW18vEGF4GWxieL761PSFWH/HPm2BfTzus+I4/uqO9TX2QZ+9MOWb8PjgDHj
sbm2xM1fwK2le9gQLwIXW5+IAGfCF4XPVDs930zJJKwwMbFAoHLLOJTHB4JCj+bR
l/I/LcL/64w0jvvXbSS1kMj1c8ixuPyY56euN2DmLXJW16XwNCknAxv6ASA5By4T
3z8Fk2xYPAeKeltB4OT7TVhTodL8iBZGS0lrXP6wuqqM/GbSqAVECuxxvGc/uoFt
o7ea/efyaR8Vl4BxVTIzafxFhVMCARMbykwrHTquNONzuiAY4TKlfbr5fn0Tw6HI
unT6jxuSxNGHJLJRKl7mvkfOYCqsTfY8F/M70BtM+7+pik8R2eRGsgBGQC5zsbn0
GPrAs1qgotssgjUuDeiXJgay9CjFnXD2GRycZVphpONSzXo3xNJzImzIruxFTM29
N8M+SIyOwIgXngm29yPcJmOMvv2JysIigP9PrLq77+EBxZur82JGSIrVY37mPML8
OsyDLivIlQGU6xWusfoR/sV2V7iszhTZlwqtIQKX6DDJJtx75qUxess8L58XRj2A
OlyGwa1H07C8O9OlMeTq7Dfl3JfHyYa/WChafnCRPkaX0ab5lyC4wYcF3GViUb41
hWGN/kCFLGMpt604hS4NOQ26KM9gMTnrpqoeSM8DvtkhDve3W0IxsSde9Yo3RrUr
Mn4F4L3rfLHopThx95MVAZ5mINPYyeW6bv4lgDIfXs0fnN6BVQFQ5IKxl72A1Oca
bTvHhyd8IBxuV4x3AmZVHB75gYmEGzBARgjN/6fveQzoLFj3M7kaK7FPgGJzvV5h
1BWzzU1gi/h0gj2esb7pV/J7solEIpOCrQ/fHc8nrEPM46F6tymtT4HiHOYIpVhs
nsK+sN4y8BUJ61d4THGTVL4ajM5l4GzR+6TVmtegW2BCsEqavcy6vFAZjCjH+ocI
jUTf9bujdN7hnzxDeQ2LD+FbUhX6Ad2RymBQysLvl4hK5oyye/NCakjTZJt4iRzU
Ul0P12WKvNGXYpxvEOIVkwFD/YddPUYApmw1ClIi+DShp6urPgZAG98J0u8KuYVb
D9mxq3hg2JXwbebD7hzRZykZo1Fuvuf2hSOo7WgVOqJ8eTupwPp4e6tNX8aFi6dG
JOaUFFQJYh+VMgIPaz+G5LjCTYorNYq/gBZMWgs9SNdPqvKu2+dGU0QDspQDbfHj
PD1R5wbIwak/1rmUqjpEyWZoX5808zo8F/lEm2JTJbR4Zcx5D4zZZF2vjgjwbh8t
T4sz6TJtGv0gXLzKlzdEo0wfiWtbE8D+P4yxB4tYb1z8rjdZcodJ/y7RbGWpLQeo
xPXm0InxSKeqg71dakJpJwJHkVaSmKn+gdQC0ephwf5sb0gmcwxcjk3cRVVLc6mJ
LuxDmJuCUmJ3fyIj7u708BL8yDcruMknYzW207yXMvil2DKbceyKaPINP4BMRkmG
imUowl03xY1fcTD5OEqf7OT9MbyT9uPS3y5ykOJTlK9w/uVIbvcyg5cXptpcdnxk
A3+XqljaEkEzNLwjr69lCCE/qGa92SvzW6d1Sh1xxxUhQaTnoG2VpwXYaxHkX9a/
vbBAakrNpd6vQyRPgTfgTRSjV5dVGhvW7zli1iHRE1c3FbPC2d2vIysF6Z8TDc+A
dY0zgTVzWXleVLXiNsAId2rFBKuwlDYRIzAfwLtBTpzr4m/eT5MYmM1zo6G5yGiz
keyZ4j6Xn5M7J+73IOhi7ePFU3HKiRsjwx2fKKpLUXAS1UDzq4ATFmHbzeOnDYFF
7Lkmxb8tA09IeYm+w2BhztK5oLlnRCnBwNQQWCWbh+1ZmrRfXdOPlspCMsjCk6lk
2fjS2FZVKX7Bc0j0U+kjIkaxCD++mrs+AshvLlCUjZqfIQbuaapiIRXzi5KZLyM2
/cNcR8m+PCgdmksQ+XxXT07PfUsNO2AqSKySXki4dxPDfbF+MiRSe2Qv3uOF2LUw
Her9XqDCNAC37GVEvLn0oCSyFWKBkW10JjXAno1BPiTV4WqFEeiFPSULyiA4NQTq
HR/lL1djI+Sdp2K2ExzPvDFrOmXciT/K3D2DxxxHpN5+A3QrIfTQHAlxEXt58163
DJwioCHHkgKP3VChBEQhOBcSgwZvLkXIpA70SSd4Det/USX1M5Sei/b4IR6+gGqw
kEqCxsTah2yfO0emdDcpFddKNWNb0jcyTWDmExnELNQZEUFiGLZE1cCkqGNrmss9
Tm8dW4+Lg0+RhkYc2qQ9uWJVGI7y4yWjg8mG8INw/FoLn2A72I9/HIA/si6sTZiZ
PJ+G4CjzO2xf1rSQ16jEL5XVNr9YBNxeyWjW54BDTTmpJM5b3ENYMx4JQPOXP2zd
AORNMuBZj4XraZwjW50mdVj/H69dkJfKFZe0yI1FopxPPFWU6bCV3w+Be4r2R/Zd
S+HGF5VdCwaU7TqCseMJ2e4mLrWjLqt+7/yTTs9k0ps93L+HsmdJSWsC+0fn6zwp
CV5qS35DSK66NuguQkOMipSS2nhjwpzoPiG43FM1xMW16NTzmg0UxgqmusdWzu4V
ief81C9Dagor6GxazfqNJQFmQmPcSh2JOO+/fQ3aIXigBzgEUP3tZvt9mIuyqeBN
Fi216nW4YV1Q9hfBeJwM4uLtSBRbayw0g6uvKkN6I/p69/l3ygDQWlo2hofLP2p8
wEnrXJmAp7bxkJAxVS+aYjPEaJfG5bp49DRnkI4E8fEzpfXbzmh5jwo0dpKKdqpr
jtzDg9qZ6MJQo3CPssMbMeYmS57C1LqzCHi5LKgvHVrlN+b+aESVFnkeFhoy1uEg
ebKPHTEgAa9vW6/5y9yWnRd/N8QqxpaSJbkT+Ly0q51O+lmTXtpRUCcif1EiRwzU
tK4jS9XS3u+IEQG8UIVyueIuuv+Vs+SBh0JHuyMQh5VDOqy2LZKaLLQzR6HcZp4l
iSNCUbV1kbHJN3/yaCuM+RbekRwJBAALLQY+Mfa1p1XThQ8q02wCZ6tT5cBiLd2Y
Fg3TBIt4MkktCQWxsEOqD82C2VcRXneqr6qT/rsEzUNOtRAEDtAmFWcoavg8zoKQ
kLk2xexqud1j+AZN5uPJw2bECXXqNr+a+pcxqU3NRnLJX7p6i3vGZvMLyd0QxDed
/3v9yUSlgLR2e6x2uy7dB6qTwLtEE9y8hPtl8N35ZZzDL4AXITBfAjdSy5jbmV4X
1/aOIGuxkERf+NmhL55XCnlRw/mGVM9wExTUUh/yj+kBPkwdU0WswZTZ1Y+jsqyk
74+tjBI3inKaf8t4o8XCANlakVs/5qCdA3oJy0u/t+++lybPv32THpaaq0lz/Srf
gVcSKU3VKwX8v+X+xbq1VcCtMEmkTTEwYQs8hxCVvjYvrMylXsSzM9aQT+drWgXO
vj+B+nQWwx7IMQFw5Bp5eSwOSStqnkZysYNpJvbKqCJG5U0/EkHUm3AoXlX7AS3H
/E48U+dZbpBEwPyCKg383ijFsyUyAFIY+qc7/quNJgSxhm+iopbD5+xVAo6OmD2i
8rAoRxZNadB8r+y08OMXNfaU9x/1pL/mKIuPTMT4uzjQXQWlr8AmEl+b3pV8Mrcm
oEHtG1iSzALilr+qo9odgTXWqYu+Xr0YQTEtr1aiv8tHlOxNds+gX2+XguYJoHPq
kkVL4EYGKNF4+zv9ISbw/0MMdtfFfVa5HE/UDpOIDbOTDKD0bHyNuqooI1m30mNk
XU6xSpq1qxOtJ8D/53QDUOq7rXIrycG4GVe5B+rr+KRH2AOyFYSRSVe81itqLU7b
RGXvb8KHqPFv82gypkSN/LEE0ZOERbhrRKamcfLu8DbaiGggOC9mlSKcgxD//No4
I6PhS21tEHBTqO/+hUh7u/NNwTE3OpziTfg62L0AS6RtD4TmINpVdilBNfaExo7o
F4WvK2+u/bi260la2o4zzNrbminho/N1w7Up8ptVNs2iTiLpbiZFOfTCKXoNKwBD
QzAbvaMEf8ZxVAkcfYCTgzXzHbtHQhEfSxIG8iTj3Wws/W8KWLudkT9aFraF4GvL
9pEb4rNs4Z9d7VNBtV3bFYwy046dULUiKp+xpNC7XqcXVeRE9/VukfPIH4vyAhOT
54l6yhiNcmpE5s/p9I+7SNhA8csZ6GHnJ9pUAfJ1pAajk+E6nKXnrn106BZZWgK6
BPyYM0a6blDnMD/IhDc6woTLjh/V3HLHQLzAOZHMEsml9onkUnNiPEOoUu5nTneS
6+L74s6/GEmU7kFvtrvThn2TMw5+uOjnHhm2xR67wECABpztx3HyP08SZE6zLe9Y
02ZOItsBdPtGkZqZ6ynZrc+64Ixb17+3nV+3Fk9m+gPOsorlaU3nVqDTS0ErLpIA
ZgPCWs1L2T+50/rQU9MR5+BFLV1iv3LbJ4TJoK//TkD3C01nxDBGqix+KDQbKLBP
7JWFeyNQSA2lsEC/HEneEjkfNi7OFOyEAZ9EM8H8LMqkhpINKKKfz0oGiipfiMXg
+LhK9aPUUo1KuONCaPybdyjdvTWP+/2EtjdFSfamT+lb1aaqyf5Jcqxi0LYY5fdu
bMlDwOQ9BETbmMrV1PlhGTNhEN8tuc4gGMLdMcbS/6a6QMZ+ZABNHepc7QQj2nq3
KncYeQ4vMyEf9rNhyapSl1Xf3TEpPxtmEenRAd7SZ1xOhrFvihn65JwVWfADEswY
ElhanayKvtx/aWYIVQ32HIHIl723x5N7h1voq4XdGKT4fRhOTB66Ft8p8QXYaUk5
ZYVHzt0p5uPsgxvlqoJ1JQPxQsIGz9t3jcmEc0scZTIg3Z9KSAWEU+GqDNq4OGUI
Q5wwVqy4XAM2usUQ12B3UQiMgeA+L3pTaKKgVc+/+UC6MxW2S+FbGTHD8+65pjsl
TwIVnBHzBceZKPJ29Vmp5s5bmhfRT/j6wDHPv9R3/R5oRy1GaV6/DGKNXdamhskC
sXEhCmyHMvRN7yXnadLUMP66+Q7PX1rV1RAsOFSC8tL1dSZZjV3o4qSqEERvlTQV
B0bTstR4QBht2cAt1K/MzL2SKuaCPVXWAbn8zu2DKQbcnpq7ctdF9XIvvq5Im1DX
lKd3IYq64ngt/kNN96XqtFvnVEEu5gjXDLCaPFSqldwVMEfheL7rMAjiRRrlYXnN
TxKGxAOBZQAYF+q7bE2ctf9LCbZhicrzCrw627r+IDL2+o0tA+jFk0/3hvz6iWBe
gO0OqnD7Yqp2hVunXQaHu4tFMkOaQ4hRrV6K5a9HqYFxCyWpz81d/4tUaUub4+B7
O/QR/OCSOqtXHbdYNsk0gEVUivNw1vDWIfMXR9U7pE1U+VbqA85/bobTBX9qYstc
dtmfi6l57lT//wF4xAJ2n87REeDImqFvj4PHXOFq9F5OrL8w+0LLwtuFR4vQ5UyI
i0TPDXKnjvxo/THQSoVaHuJpJqDVkCcidUaZpvC/M9TWCvtThhhUKSYxJ6+1kRBr
VqtwL68BmjfQAoqzthkQtc8LM5vEdDd9EIz72SE4pi2SDm83JLCt4xpKJEgFuD+S
2Dj7Rbe+1SdIt/rQ14QJ9R+61047PDRlqv6IT1JGJRe72mpCXwUzm7wtZcgRrz61
6hGktTKOgxzetCCoNKnJ93BG7QdMjgPMxbT5NR4Uj8R9KpR4xhKffPksrPklF9Ka
bveybWh/L8EKqfq6CfCx7mRogpSxjlktIAOs00jwQyCs6dt1Q0dK2XPCwQ9SjarH
NQFQeppv/KMr0iVouHPXtd76ZVSufewX8/mQ25SE5bJ+CE2wx7FXlz3AoqO0f27F
VxwIi6EGGIbBxQOHeMXePalgYYZakwv1kMFR5yZzfXP6NxuYE/DXOdK8WkLz8EPL
gbtcXm1En2I3FgumK4L4LsjCwCvnoywKOxzt62JxQAz9YhydiR1ljL4OEUwAAPpM
UFaVxqy6SmcQNHric9InfxgdrCAEXnCuolfWXjrliIt+cRsr9ZK25bb3Gvy8EnXh
dxcGphNH1O5jZLq282x42XNvKJA1mnU2Kx2C1r47ObaenOVWhNw/P4XljD7QRAIj
eGmXLTsBFueFqmHDcucNUXQvUd+tSjgPmHlzWrt1acvNlXhbFl24F8Eat4ccBsnd
zAhndiCkkC4MPjw0xx3lxALqkP54L/507jDcbU17k2nyXE93uQrKhWfi3RV87o/S
mz6XOVDXWLVAEqONytr2uh8iD5biqoM6hm2RJpfwpOWo3tNRO+82lRSrxQr6AB83
vTXAWpoQrPDYDyytQQYxbn4qiqxOyBqFYiTNuNUwldhQZy9CP+gxIYhfWV2F++9g
oO+qJ5uBJmvyc/gQH4ditshXvuzkaloVSaf+mKfuTx1y812FQDxvSh2JQ++4EtuF
nw4e/yKdhyEYayCNtlWJNhY23TOsv0OBkapWOzdtvUV7lG5rpWufdlhHSWw898xJ
rTIg27uVScltbsdAvK3J6NC6bcMnbH+IaznZDJQzOcOiuNjFY33i2fG0bMgi2I9B
Es7hB8tqSXQ1nsgZK1e4+KeizAyxOZ1eTqooGElEkIWISqu3b2OMJpJBQepH/xuK
iZZ/H8SOeMCj7NinGXwZ9Yg/Ezk7jdNxTslVRNqpanQlt/hqlEez43MDHvE8oXzW
XQjhlSlwHAuoqgKlKjuEYSrKEg1TFCJfsHB2zVE+JquQ0OOFy8MFDynXjukXxwMC
es8E7/76F2yy4z2K2z4SV4ALWUT3+QTIKq/qksdWOIYnWNAb9OMwnQSbSw0yCyla
Z+eB0pXZ8vFSsmalKePvjR9CBC3kd4IxALWB9WDqmi0qQzmHUkV2+AHnzd5xv/cF
XeoCQS6qEnJgAPHUo3Q3pYYnTvO127THJm8seGrzhEjFZo8FtFpbsnyto9lqem5n
GSpPw7Jgj2ybUjGabZxD6z+Wb9tsc/Wv+VhQq1djSrjLHK49F4YrNat399eTOo/g
JhyY8XA+xkWR2k6/z+NKkCBje5EJEqkYfVWeQlFb/O+zmp/O4rhskn8/lfw8NE7X
pM4XRAyGr7AOtJcl8JVOvc+xfYj3vSbJ3dQ17KDoUjFWXqKttEOjuJqLn6xKl/f6
rInYk3/ttMW+2o/LhjOaYpLNQmY9F87WvHd6wXHuRvLYyhAV6SwO6IQDWbigSyR7
LQOd259uB/Xuqq55PgmBp2Ft3u8pezxc/zwRHCTLQ2JdSnM18YsLnyiNsZMJ8Wtv
hA4sFl9a4TUeXlhMuZWVCOrWG9uvr6SnBBIzrGfbmuLHS43GwNcHmRr2SgGruWCK
L36lxypE6UM2jZ1dmN/ELrtqFIDlYjCQUwro4XfSjIP8YEnokOb9oRKml/rRpp7q
tx0HvX4u+uMBSuo36AMEvybjGqShiE1ymKteTfrkWCeLkShArS0Y5Ruaocdm7LFs
0oiL/sqk1Y6/taLqva1n+FzK4suglxZVY2ptJ5Ym9BF2p+Lropn5Gss7g49wtQaL
3BqV0d2//xd/TKr4W8Zj82tSQb4vlDxhl293D8ftDZIWdiWTFuwyeVz5dK6Z+1Ly
0fiAc3kIgYKopmY6D1wdAW8pB4+UAobgk+IaqgXMiu1Bl7B0SaKs9Dmk8yTPIvL7
7+/QtZLKPAh7jVgFzGttLQCL8qeqcGqCIWPTSNlLNeTmuo7QeUK56b9xHfFWtqy+
txQID6h92k5Alnv9XwKwDCQD9EujLGo7f8Eg/rJYghwY3iJcidpNJYXd1yq/PNVI
fSqdKbd7tQxwLEk1/5q12JbdBei+0vWMdPIu41m+eq7HUzlYmZHD4RygyGO86Scr
4cjlrKXGnVVeYDYX2j8ZHEnWbEU7ID2fHEyUrWmBIV2aaqHpE1+SUBtlRQk7BVR2
5ApUbeXg1Qf1GHr1dzo1hu/wWtn4DjDKSD+H9puXML3jcZAwzf8fwckoq2FswG01
qVYQoRn22/Yqr2xZzRhCpPBMN+GG0bp4c4ePVUzq9WPGCE/Gl9U3l1CNHHkx9EjI
n6d1Masm3tSAB+QymqpLUPLe9K0n6AoABmJd6sbRzVf840ajEbe5ZF9Fmha52znp
F4veVNwuqRRJbEDzbLWmwrf3YjWQfXavhY9EzwC2REYKbqE+L9mK22Q078Pm2vqF
227ELZbKb7l7jATS8u/Z1OAn2D/j+B46VQliYTcvErwjG0CiHnM2pJjQOY7VpV9t
IbQ9O5akVfTUAX/P/yS+ovXdEWI3+4Xqv94/mVpsXoVHtn+osm5tI2YZQZjtm/oB
pcSN2gwCr+xy/4y1ECGvjVAIJ44Ninukoj5SkyTBe+Tsyqd4Hx2Mti6Oz2YY7pci
MuwPvre2oguG7M1wT3CqEpzbnlh/m+DTqwUxiryj8U2QY6kUhW/wJi95l9hJrllk
6pL55ToG4RjgBwKZ8d+eDJNLRbAQ5phv6bi+cNO2tpmycY7XRKJleF1OlIUMOPz4
LNV493r9LFHdAgk1DCvaF4mgCnEoe994zpEQ9pS8VSXd9RB2ocxq+Do3fzextE9v
6qvNeruuG24Uylg0Es09BMwpZVDhRMLHXo1ZRlRlWtUIxWDLVea0yTJiuTs5dT/h
bqdnWdLNd+q6LHRQnoi3tkaqoFIctrQYECEP77tLim0w1YF7U7iuQ2lIzDpdJUOb
XENzQRzcmQUurrUuBC/UTDB2paw2Y4ZH69qGg7ecoinO++G2PebpROLPtzpSMJb/
QPw6vW6WK/fC0jDML2j7CB3upUhc4dw4LLALCXJfYKaywiQOuRbORq6YdADAQtfs
FdRXGmaz8dfeLtwNZCDmIcfhvEdOaNoPjNwXbUq55syES9mNXHavfSU9oCsdm0Ls
sxvDax+VKOUn7qXZkJoOLAuj2HnHp/UrkRn2KgpGZmU3pMDb8MgeMo0yGExIsUlT
JotMSGdjGfwBHBPrO0F94HI8bXikRusJ/T06OY1yE82xOX71TStqX06n5uU2UmD8
pZYjTr7Y89zNf5iV7VadaL6lc2rTTbGJ2aVyi8vxRRxe5BBGD/tnUchyJyV0G2IH
ZWhzmqwMjT8ZjVg6o6xojUqhBclpmsQ5nF7+YVJ4Zwqo7fcdsBUgd/UI6kh10wPz
ckXlRF3bfG7QJEEu3oCiSNpEbZEbEC4Bg4vFd+egc/zSOVRYldwm5Icu389N2vvA
kSSnhQAo1mPvPlTTMj8mH01edMlkvhzq9RB13P9SHWB4plkmCI/rHcBZHbe49Y5V
ajOjn7sEDLGcYI9ffXPJnqvAG9CcfgIzXaA2epyK1bQFQrw+lcgqS5lg6dze2sml
N4pWcrSGsJawlEPxID5L9RynAHAEETGKmx4kh3lchxprXPu1WQ8Ktp50N45w8b6C
91+kH6x4aqaaVzAukXTJMYtPGE2odIURqE4Mdpr/RmgKvhENR2AnZqR5V+/sN5qz
FWBnrzUK8Z1kWMRLIfPF8kUhe2w6Uy3FCDuxvZX8qtqac64tH1kfJ5I04uqun6MC
KmNfh/iLzGJ2VbufC0CZ9OnvjKDqY12PbjrpiXMgzl4W89FRbi/3UBRa87s6Hm29
xQQBO8EqSo4OGvmOQXXOjUpyN9SO4OIketHKimmQLUpcfwcsqKIDS+5uLiRoMqar
T5e+JdpywxyiMG95p4D08/8+sDtn1F5AH5lkKL5dDo1KJAyCjFBnzBD+DFRkn/RT
HHqVPSj+FoiXIJe8NIN1/K4cHyCCS9/4goiu7XKIKluEAWep5Auxk3kbYUG0jPV/
Dzl8YNRgtGfDYqwtpLIZHTVW3ZtOSi3NaR7jJ0s93lZGlPZZRFP3H6ShXYDmCLZ/
A2J5b+rLogp3Qp3xNkNJfA7J4kzsm6DE0H547dyhSIgaYgDqKyDUy9kSxaqZkizK
DOZnbB+VQIuFk2eQN71tZmMDf1Zjh7YHhJm08AlvioKSx5mbOWh8IR4zBLSKHZ7T
W61dKrppqNjWGA9DfONwm0AzzOgXnGlqMAZ8JTDaTQyRs9Qou3T6HgM9lY6/1qaa
AqS+xevbHiemLFlSGpd0d5MyoAf4+QugIg3MZov7y7aAd1ugFbLtmosALzc8MjqX
YDN1jPNnw2VSpolOoO9mmJPR9nNbxHvz5gJifrzAI+wq+cKXsfjf4o1O2c59sdu7
DFZKPWMU3g/PrEi4PfcxYKiCKn8L1R7WxRgMusIT3DIGkIrZONbiNRdvp69evLSA
5KVjS/KVIKep4EwlgMud36IxjteH0yI0nXAuoM+KNE/Btz7jKmGGUwcNmazjAKTr
QZN2upKZjrSpHXe/8jCRgSVZUcfeqpmMEiWzFvW1ZhCkfRSeyKAMPyT1cHWmRPBZ
gvRb/jBxGoYQ1JJchJMW6rAXb88rHFi1Pn6fkpG+EL893lOBlMpfq+DsneuHtJy1
LqLYikiF4HI+NqYzIXC3g9pCxqJ0xCJoOWQHB8/osU+f5UNPHv2mrKnHx8SZWgDK
C7wA/g4OfK38uFKemgojyzXEZlCFLk84V7v9XF43HrMGiFsSk/5qCEzJ00pSMTvA
2TXL/dODPFv2z9j1g36iMrHGsgwIZtH03v/oW/oYxnciOjGTQq6Iv3rVvj0r1rfl
Uyxxpzao64J9+4pMElBlCfOnv/PzbGBEABugRZAg5smt3056ZdV44OThVFK+vddR
JgDHoAdGb/4+Zb+p3KqG9fn6mzZM+I4Bq7Tike+VDZpCLs6z9cqQl5gxmsVyWsz0
EaOTW948x9Oie+5bcgxr5zMNMEPKdYUZBLdMWjYjb/FEZj411JD4++VRpoHry56X
8epktQWMjFlz/2TTDUpdiL1qjxML24QxyAN1HER72jL0KeVqL4DCjPvdqrXMyj1D
0oxXVi7kTva+b8UNMsUssGhmPBqJc+mR3IeQwJsaXqcWK5Nw8wgYnAQERBTr2EGm
nJtQIi+/y8vuLDg+tRsf1Ugczy6FIWbd0Ld5gxo35wJIdCNRgs8UOriPw/289KEj
Wyh0YPSyG7cRUuD4DIU21SNDBqMlx/iuIbgQjEUpoY7qvCqDyUUt7MuIjpKYwSzx
dHgduD2cJ89AZxCCNQBe8AlQssMhvpw+t2P/ST7tynNS/28RHNjBvGpPxNToViyr
djdP3kActhVxkwhtqjr8R8cbmYckLacBhKdZMcYzyMMIPsJZgFuUhNqtYa5xfsqQ
gqQMXK/LXwXubwjnvCYAjdbUClU3T4pv9Y8eeMRWLeZHt/i/4NfJ7pNEwdGVEjMz
sQH4EmDmCoXJdDyEufTg64apUMlJFEAGHiE6/hDCV8FNKS+x2E0jo8PrRGvjlQGX
pORJfGj/uxhyFP2CYNu0qcpcpGqfV8TFYE1WDfk0FxHj+E3IdReYX9Eq2/nFqUyp
J8UkausKRpFisUG44I+mOvYqdmKs515fgYQGhaLLlus6ZUyHInuld5OsCtsmlRZ8
Ce3jDlqIG5z64ob3uGykc+SHzJn0aHSGNo//vK+wabpnLcZ15TvE8TbldRoR1yF+
NrbOFhjBXNkqEIFXGYV7YRRnVNe46bJEXD61bGT0W//Z9zUuGXmfmcBN3Q4eY0pf
RAN0Wx9NIhEfx8+t8UqC5zoCuS5tk04sjeP0khPRnIgs3TV+RK4XJL0zya3ZJUlF
Ic5WYuTBTgd3FD4MUaegjoU4SztwhHzzOMbuqUisSnehbMYk/tL0QBNzrMsoizvE
Z/Ewwfvqp3DdOAsVxxmvkrdyDw3db4cZY1gNkSyn6f000JrvxgpZQs6SRpZ7BE8S
O9lOYzqIGe7riReby/Z7zcWcJEI5lhR29z67cjkHcmH2j8rzEuQmuVzOpRj7+Qad
FpdJYRg4uhAWMIvJPmf34+vac7sNnLLuX8JghsPBVksrO2D4MBYq6c9VJbcHTTgT
lJpSO2zVpf0zxt2SYe60UzwCbh9LsNrJb6axJ9Kf/lYp95EW3WnclQqoTdEIJvN/
Uh5/LnFCHDZTob0iPoQM6vZPPDBz5FNqHMevOowKbfQyqoWGCVLNsDNgPZqpUywo
fmUglnYhSsh+cDTfuU/Jj1OwG1E0sPrfIK6AW2jsEXeWxzzI0leeOJe//+E2oOCb
sZ5WmPt0WGP9RTRBvoHXRYognGK6n2u4MEfosO87DC7Ydg6ZZRG3EJNNM5/Ij4OQ
/1GOUzSe4yoZ3Oq2d0tnF4KC4S9nZ4zIvzjifRODENF+8vxB3PvC3ZQk0vTP7Z+q
nelppNXOHDxGEpkLV7Sbqlr5Wz/R5jxSHWdak5nXbzpnQ3yI9YdUhBoYXstAjdZv
dr8HSz14tpMEp6Qv6whljdvcbnYv8uijTHIIYyJcrRzkwJ3Jf3V6zdRM4m1Oh3+c
wSxKwD4tu3f9Mym/IBXhVIVWSHhZrVKEGYMtvke11r/5whs2of7XqXxSXBakjTP1
cX6CIGVHvraMOtEEJ+luQSdLrhDtiAATmnZ4YNSHF40Fxadgd+Y3Oe+pAWfBYmEz
biR8xcRno5so07PVywr/obrtMoxJPl/PV/aYRQ0DC8O6dw9SGSdvEfNSyWx2GGyN
Zw8jy2D08g8QemuMvOD4L8BVs3AMRHJ6pLZBqOe4EG1Wh/DlN1zgfdFy/yJ/kV2u
WUo+L1VDm4LlQHLiI4gPo8Y+MkMnUNz0HP5OgxJjfUmAozj1yb/7oCy7bddNGQjO
E/Lwn1pi2oT24VYIlMIbdFbfRJmEgQTfvWRuHXcvHOXmyOOQM6Car51y0ZBcxAVi
U9tyIJbm5iEaWD7uaw1SDtJXv9NL33HBkGs6tdmqK41lIvOkXyGDT9/LECAv8HwI
cKa9flWNxiT13J/i2cJu8Ju0KNzVrs2t6/guXKJq4uihhibq753xW8e9JU+twvLJ
S6P8UAJFifAryc4xT5Ss3uppw43dFAX3hLfHo8MLN52zxF9o1VaI+OUBEBW1CPxr
N/Df9IXL5DYvhg6Y2fTDomP+Z1qtc5i10FEUmasQXde8E2ti3QFqvZEw1JrSulyt
Uf7tVpKHVQFnCBrGJipSARKnczIcBIbNVzu4vrgyuy2A5J9Wm4RPjkPneR456Sdc
0r0jqbuiNpi+oVBqmRDvM+lduqUrhrR91eN16cP57ES70UmVB/5mJ4mABmrWZZSk
PTu54xq5bLTaPq1MWd66LMEPJ873dMX3RujttyDJWTD0sSqRMxiSlAb1PVDTmWNO
ieKNjV7DaQ3CZMFJeaeLymeLOWKXhjc3HZwaCOz2+FeQvkaW6WGVRXwuxBEORKRW
7wfZGQ2ZeQBZP995pOFB2dfsyXhM1LJGYdWgmTp9z6RIMD+0Fy9pKQ4OophO8E3E
BfnoA1P9bHaSSI8hGdftP49a54OD7W/dQsEZhNvSjgGzX9EcWRmsrs0JDOdtcvxW
hmnbWSUadraWzhql88CL6jxCE+84MLWRFLTRLi0v4jqhigLbvGUkoX91Tmrszn4o
fs7qSu8KjASsCYNJkJBmmZeQaL/myW1mAlkNbMovVrTGM5Gi3kb2/e0xQg7oYUAH
kueE1dviJvPZ3Vb4LeVDyzhd7G0NphD7lo6esG14ibF6QU0IH4EQsDdBRdvfYfhm
lqfHs3qakXewnuJQ1us09lCoO/mpaApsFMIVr81bdluY38jcu75GY+BtoLlxj1bt
XwCoFqc5YeP4RmkbqRX+BzkakUO5Qd3O10Gn5s82J6teG0adJZSE8oHW/BdQ07Gr
v1ock4c79+IFOamdSzRo7ISKEaCi91l94ikn7DiC8LYJKMxxlsXUjAiRLXfwiz8K
x+uplcOvQKJffbVyqssmFZHWkP7zTo+iVIZbZ7pHCgFaYNJDRIV8iPCfvplTJWA1
FjhctcHY3fdvQmvZ7q0AVGb79F5UQ9HGFZ15FT2n8XTt26D59L8pV1qKGfDqlivU
NqMP0zIJoxL6LIllCGYQ1mow+lQGi+di/tN2+5fC1b71od/ZEOO2NMLjC8sg4av8
LzduZNPw/zZxBfUZrZe4lusRiygScaPTQf2TQfwnEO87raN6OkZpfDH4JjTyHfTE
HIKEe1yhlb69ua3TT87QlFuqFZp8PCPxSdmHRgwofRX8s7Jer6ZHNOP3ejgeNeP1
+8V7+19JoV+KouKg6kC17/ob5+lZaO2+bEyusZ52WwfsnRkB8y7Pw+jVdpYfVB/l
sNBfSuZqoCBH+JuuEl5BB3yjQfzN98HakmJcIVhzq+BugZ3P/SOYrlW9vT8sXHv1
OpGJJ+SMJBYtKJ4GdXCLEtOToQdfnOav0nlWOp3yXDHG6qxAFJ5CuRI+SdabjLjj
t74pBMKlZeV9jeEE8EvvvxAtPHU19+CY3oAFh0tftWEdqtdRCs1zgj9pRUUxi3/z
3PN45D6wEXUp6T3rPLohzRVSZiPUq4J9ZbRbhFRWLoA52Gr3AlBk+DhPGU6dSMIe
0HNCkRDOysP5uYtLQIM2m4rnz+hdCMT+cKpgBa3pywsG4x9Qlk01GvS8VCHZUEcf
UkQcYZghvVLJyfGQGEZrJiwz3ulIRD3ZI/kD9Gs32leQ/BIgve0heIhFYygQ9QvJ
kc4ldOaY8MRYx34KwUNPxoKDd3Gu6/HwTxVDqxNtDnNdTow2Xfpo4O3foe7aDYPu
0e/PiWy3bi6r0P0MvAjPhxgB71Ttrdb043BOjB7hE0tlTUuZJEmH74ev4lb+dV9Z
wfUN2tIMPABcrnJHTjKYSw4lhHYQrtlDHkOKRmYAEnx4etgk6xJYMBf9NPQFIY+P
1F6jh0o5vsq2jm5yHPn53V60VZUKIRgOgfXVe/xevUYUEVirP4qzZyo5Bq88hfue
IgzKhAOWCXOtcetRc9+ebGco9NI4mxaolDCDH8/QTVI45T82WkkktLV5ZGSm7oaY
tKXFZLHee7dbOCOjKt5dkCofGYxexmvs5KU63M/jpIndI5PexnYaFfh9gptqmfmA
PlhFI+1hj0VT+yD2sXZL6F07/Ma05C6fNCqBUfGto9Ijyp481KU8BGNX+Ro28Uob
8ehsfB2nOK4oskItIgBMZk5LDlWhU0k4UNMgbC3KM63YbTugkqAE7lT3k0JQnb1u
DuBPwsOLjrSRIfrJrZTKxH3g5bRvYrqPunuBDMjWFACKbyw2XYs7MU7rTKQjqOe9
E/TO90TDGtLaU5JVZIHH4no9lYhZL6wiQxcrhEXQuXaSCZLWTk9VDhb3QjvCocT0
PwMswBVapvbBcafIC6INViMqrLZ9iWJuLMh2iMxuYbevQ9JEHUm6rYvgLsQUiei/
766/UFypfJA4JksFti+PSbjAHcY039ltWYprtNWz7I1vq3oTcWTnUw1aguzgjIST
FEvVeWr6rYxFEp4wx3kTngm5osLEGBtUFnh/1CJiM2vWiONpsnrUdaHOCLIoAdYG
vkic57q3vD1l6MmbkYlgvYcsAWOOEp5tyMakFkolGTHgDF7UIqcLhGZ6kYrCMJdq
tIQEudrfcV+Kb9vZW7wLzwyCpJOMqEuz/OlgyUrSb9n0aXfBfIKdHRW+8dTE6lA0
MG8Y4k0ubp73t/HznRDFZ8DBtJFlYjmDQaQnfGhVnOHfJSBLG4rW50pBdX1F3cxP
JXOcK9OexsW2dWZveHuyQg1n6mOql2p3akVVxLDf3RaaNLxmmdd9YPMs4MXt1bc4
XlLQMH2T+otRAIhgees7axR8CEKVqfVfISrdm1aTtUxoFaHYFsL8YheGwXSGoAVi
l17q9y9vNUYcGHREtzMMhix+AADDR1R2rQPEYHaTZ7dxDQqkRCqDp/zePEp9qyqC
+vEtOoiXiw4PoR65UGDYFKvXzsxRcO8jkAcSyW/9bsqkCl7I1MZyaadaCaqTE7uv
HMU6ZsTibtOgRFbJqsGuOIVkef6P491ZdP+i6FHWgq5S+mN73/ACAd/bcciaxcVX
DzsCcdD7F9qqHoYcQWvnGh3EttVBAOlK2eyVxL75D2nX+BMI+lwonLSd+6ek0yrA
hA9OpR1fZWWr3H/aJFPHAqwgFe1eauNX1QorSrHqwjDNy6feGBi+I7wgLOhxvtGT
grkQ8U3pCqWppe+/+yqMjWPSYDELpG1ebZCs/IKR/hDJtmWOEYtWizU65WpjDXlK
nHdg57hP5fwazYigqJrGVIgdYI9d1lKBEVp33CoUIVl6dXr0FpzNJuAjDYT+T6FO
cT9jRyg2HcNOhooQfUqmoOsgf5xVocXTHKCwMnMY1luaCMvWrp8M43GAPyMu+cml
z1kO1LQGV71g+wQ17QPvzc7IIVIcsB3lt9aR/nLV7ISIXcSb5CBZELHT/+2SnxYZ
g9FW+mXWhZc+YnR5tNfGmBUNsiFSON1HH24bWbUZPYJKH5XuK6jYkiXJsZuo0o/t
vhIsNuQ42zs+fl6vEvXVS1vABS+uB+I0CxuhrRwXT0lqXcUbr/r40MIwbTCV+QM4
vDC223EnQevcAtwqSRNsaUOb9BA3owLV+ixbw17mhVfqOkyWIL1yUxD3g34OzWaz
Bpxxn3F/SZUFdc781HXD6LSflTgU2F9BhY30Oz0nqHvIp87eDeHEC+2QHmIvAaVi
t58waoLKGHIiyFQX/fuuhfj7ztu7RIpwDtZPYmS4ChI/B8t4Ut7nZl/4HBpJjOMT
rgJIHp8Llm9ZNyqZUv5cSCW7tz7kcWnmZ0E7GDxPSq8xh/nyKRjPHhdrETvMKPB8
+RdFKJS917WmVqx+PmmdCYk5woC21jr7il8U7IZ6KIdxxeGWQlnyc6n0SuHXLZck
1S7fkuLaprhUZ1X1fzEBrax9eayLIgyY9wzHRGfw+r8QlOmmw2ri5tkK5KHLnfFj
IXw0nTOQ74mr0W3xnT2hekacvEwPKnemtf3/kZWG4AHtDzm5H7XnzQFZs4hAT841
iLRD8UW875oToyHD+alCtcawIqPIoh6FsFllObAEAxI+cFLTW00IFyekQ3tpKuZK
N7tI9A75DhPbVAJ3mS/Ia8X3gJUcJDl6P6nHir479yWsCfNuYBaLCoyoH5/BxoeP
5M/T3QT5V1t4I+2Yjugx5kFsCfTV0oegc7qOnASdH+KmGVQoqj+/MpnpkBjcfLdH
o8JmaA8YLjAeiCm1N2KIspq5YVdFb8oe2pqwHhiTNpN3x2oFWwpPEuUxm+zTFRuh
Q4TDV7lLgHbSF3tVa1SVe1m3n7ek+m0y7cwOvgnRSWpdKYWLWzEvS0Xgvy9S3p1R
yAHXrsRzasR28ebZlrSHsSmG35/h/8/bt5UtmYo3otvX2F11WG2YGWs7Qmcm50Rb
TmJvKoiGfNUHbreoB6O6QyWPyuARw7Na2eYpxbu8WGYPOzNk+/99tyLQq+Vu2mOx
2iaYRVZpb+ser4yxl947o0jAAK6/ffIETpUciTZW6ZtvmM98r6Iue+k+O8AUbZPA
vTEi3D5oGgXxoH1DPzOW4FHkN7VQbIuvBZBpwG4e0aTNQkOQubVGQxpu2XKRsR2L
ZktqO+GnIeUsyR+jhV0SxT/Z8yZLvYG4QUQ1DzVOSzetmyDJhh/tFhrKHv3HU0Nv
jW9B+QKdK4fdOw4oMrXlmNoYyrcykuSIm5tlPmFn1ta0XAiX/xeMZ4YMrIh25Jp/
BVYihxwayNtwb4ImNwbwHrRGRBtRzwv7XisD2RomP2qF8HBfPSAeDHaC8C0aqyxO
TFXC30c5v5tOv8yhFGrdNMSQ1uPLITglmwPM0m7J7JJCxbGzmsMj6Cv5ehI4eLGX
AvPrGxuX0DuLngJ+dYiAQyw8anZPo9l1TlSi5XhKQyB3lBVtvoCi/2Ql0WTgr+b7
NzYCdJo8o1Cs7VcTQGDjpXNkPaDuEmKboIyNSAtk1A8Vx3PbAZVuQD+E3ZkZRdQO
6BqPHwUg2uELI+x9rZdo95OX4EXg+Q1Rs2rwMkdssKoR9jujZKkfLLKaQxITccEH
XKR8orfRwd1+fbXYhW8H4O/uVcDBbJQra1kFWMTyQ27u0T5Qg/+0ukfpt+rF4Nyz
MPe1H9hg7WWh+HyFtIXhDDG8HA2fGZYh5bf5gCAsh1Zr3eTgviB2Vf8KhYVY3lM7
mcoCSB3KYhjO/T+KKH72IS7L4btGMN5viB1yvL28uQ2WcocYi6OCyXqrnRgP3zEJ
ApOuIDzL059OMAgrLi6+zjGyk2tN+MRpY1bLpIVsC/coEARLJ55Hm4F58VXHcOH0
G/kXLd7URvGB/UJop4kMiLDmugTq/2d3o/AEx8L7KNpnvmEIHhC5y4gPS7q5m+Lp
p3t3N309O7ERoS0oUiKOfK5wIVSEy7SXB83e7jg26q+n5Ks8mP0o6QNdMq9zZig5
Q4XLikq/0szmPV/XhS3ymLRywF0GNJ7lLQ4v6/7Z0BtKp9w5rB3do3uDbCi+JusK
TdAAVJDQFR5dm3DHuJf8f5Enabzr7TfRZvwKbG6NZgK4t8fiDJXkOW96NryDEPw9
89aooqEbtD4XiowSlz63oTp7bXaGVXwz1gqMpvkC7JD7BRRHMVHPIcHU4LaKQZml
ZPGy6ntoHGtNDoZrItuFIAEt3kh0sSwZfO/1w2vQ2d3fBVPzpmiAgNV2qI1aONjL
hRMMA66di4dK11p4PstIwJ7z+XWigOXXYTM8WC1hsKAemUGujlLI5qNr/t+tur9F
fhpgcMYeyE9srx8M1x4bVyvezpQq1zYryqgRSQK2+01ZqrOZOvZKkmuyfNC79ann
Zo9NuvNRJwOJP1dokP30IgqdUzbI6q1uPw7KaVkLn7Vt1+Vnqq58xZjNzxv1W7Wk
yBvgSV73SoDx4T03u8dCismJh/B4BZhkj339QL9JB7d2yeALyHy/Uwbq+Z2ubroy
LE2hjqe8CEAzG5znA1mYDNbRsLLmvTMt7wfN8XxjbXMdSL6F9aAhA1dESuc/tWSo
CUdQ4gwM4agjJp7OikJoTz69rBjHez9rrfVoanhcs0bmuU5R/JF2yZ67UpKCAB/D
6DHHDIM88uVWmH3+iBV0x24+Wm57nTfwxlaJ/Y5+8pRjnkHh1/f5O+4PsXQ0+PL8
e4ohQCv5H6ZXgD/6u9iRqzaO54FgU4OmvkWgS1WHwS+1VupujtBCDhKhmSbofevy
7moi1UlnvB+ES2PtCEeHuGV9clkgdHJBGwkH9qzb8ToB3X8HjEh68ojJ3xJ7R8ZI
voEushHHYqTyv7bNfV+ohg7CWWH5f1r45cuybl54wHTF66JBI98uYijm60MdgRID
QF4o0RkFIMDkYnxGr6bEk8xe/Uze+67+RWAfPWHtk2+dfoCdrt6a/T+zRjs44LNb
6gC0vJgPz2W0kXhk0PKLXgxFXH6KgzNB9jHMLB10uQ9/mWB/JYOiJ6fOwyIEQNtW
e+yG2/RTF1VW/yyemKg/Pw4/kCtLbdu5n7cyvtu5mdjw6v7I+6h2NCsdpFDoulVm
dPYxIs8J18pN2cjSZdlbRIARWKpBK+GwIorGZAWFdjuMAr2hiPq3BqL/J3rcFRJ8
ObWizvugdBrmkE7SDrNALGLgbFgHH5d+Ga73v0XhPWD46vH4CzQyTNlEAgBDkhXT
5FAu13t0v+tdw5Jy8YK5DlEQVOzkt+ONscG3qlYuxgxXDI1n7J1jkz2LTQPGUYSm
jIUBywz+9r7zfRona5Hk184nIx8rlEoY1wpWvVVxzluKpLHU6wikTdzcZF8Y37WT
ve1xjLI4lvx5cf++lhTwDvJpVTrmKx6R6fZtuJ84+gqa56oW0AXWA8ryBpbc1sp3
ExRBaAaAHy5L/yM9wz4axe3IvBdGeUEkYtwx+R3ys/5LtH28xpCkuqhxyIp6HTsW
DAmBcqPtnl8bSoB5jPo5xzN7Z5sKes3yFSvRan4TdeqRPPPG5+RG3HMhU5rpYRoz
Sq3KA6vHjLkl5aiSPN1ObB2HVAQIKKCY/gJjzPeqWCAj+SmYAKRJQg5VekZJunrO
hoZU8JwbAaW53RI44r39Vkgarg9Zh8r/DPxVpefMG8dH4/cmTHpLqs1I60HytJQb
zpEIorSlUm535Sf2yb2mUhteb8RXrYPo4hj9IzqP82C33xa4jductUxgYhF3/Cw7
mwfkp6JVkT0yVFiTeNOUOpvlVGwAqS7jaHmgM+GUrIzuSNPekL8q+T8LO7L+3wIU
U8nlSfbVrA6ef6FeTlfRWu0kBKdEqZ0HWPOVU7Yw5vwMaQeSSdwpT2aiV06Y02Df
0bqkYm7IER9V17v1q58cxlQpvJ3nvpMrXDQGjXqBiH2cxkQzTyYk6wBhstzCjLpn
1bgy9ZTydtwGbb4K0z7GZYYWtkpMtF1h7lKrpbImtLdgfj4QaFSbblvrJK5opQWt
UQ3shE0FF2jnXVTAcds0u1cZBqxNlzDjSKhcFvekN85ZnZ0uLYYYf5DTxG3wRxH7
cKGlhTbtCoC74/WqsOAEB/Rb4cksglFV3YMrLyZhYQrXjnvy1ZDydLPSSQtjrHbO
FNwhoBYGD2b2Xb4IaGbnzoxWIzIhwFYyqdQilVawdlrLSgEF+vZiYdKJQoO0vXiQ
1c/iuEKIS9wpraVtkYE+XUfOiHcRf0ijP1YshoJ5VBKmPkAVR8xkMFlkJafrfnq/
lfCD34JOD3FrsZNyMm/UPDnuR2PnJoRFNjwIx+0QpxOdGmRNKXkNuRBgClD+F4k0
18EnglO0IAli+H71etfPC2UuJhEh/WL+ZTb7MRTGdTVY8qhg8CyBJlrKlsFCAQ07
LJO//jYuKysK8FLBnF6dLDwpmsLg1ZDDryTcAvFOpQgegx8LkIT2C2iQX6tL7l7J
VrrO7QtLHiVvGqHbOWbm/WpCnhs1OdWEG8Nh2VMcvZ3gGeavijQbJxjmamvZnb0w
jNAirz0Vg5NoEJh4kSNxBzwYsm6ZegGUXl8LxD/gV1G4wc8WbgjX2vasXQeJVu4Y
knaHjVG59LoA+P2U28Ll9bY9VvK9xTaFE0HAkL+6n2dMDsR3vd+sFjx2pWcxyjcD
hq2VweSPhbYZxNTSVDs2dkRK+hgSUzAcRGCNHoi7M/b3bbqEdlr59Enub3Mnj3w7
9J8RbHB1JtHOEkb0fF3/11gkFVLxcd7v3VVYk21yokmTW1acibMQHO45NrqO/1bL
GnazafYKW1KrTB2bUzQLAUUJkYxIwAR1wDbkubi8/WZdpxbSH2dJVNpjLTzImXjc
CPLltLvnfXESC4Yok/WXd4R6m6pqGtjdL5a5eFedr6hJIJJqhbN5KlWKlvOmiKGJ
ZaVIrbc4ETdFEWxi6OF8b4RsVAMDkD5FXBplSSyNs+U1y1+CDA+SxzKdkK8AEvFl
OJwQ9aidtoM6+KwGx5npqveB2IxAzdy9FMKeQ9UN8JaY7nhYFixqcaGkrMktTWbA
pUkvODgUeZ91acVsJgKLKD6haG85+Ie+sDRRTgZ3sOzBlpkneTF7RCWOtzhrrEue
lTAneC0LatpryBwHPQUOYQAOFjzhsZKanA302i4NjktOIeQ/9hF/ePf5ugr0LCFp
jVRkstl9+KKxupWYEaiz8WZjQF4SSXD+FUYdB8FD3xTQLZei9KOukNNtf0ggOvXR
wz578DWzB46ahWE0msCFMtTfYs/XeXrJ1Qi+4880Fi+jDOhzFs330oiwujuCCnKq
gHGLeszh43cgJKrz1o8iwfRpvXFC5iMIlUDjO8yozDV3YGFMdBv8tIK0ZvLZAqAV
zsgnoy6DTydGdtezkhyRqGXOk9ZNljr3syFURlvqiLmQpg+Ckldq9HQhtBYV0qI5
FjoaXJht6LKy/50cqP8dHmvv+VDvnR+KzvwoLiVNFwgetv2D8O/5nnAol/Z7vc0G
EAYHzM/qY/J2LFCxr/tcOjGGXuFwa3vPRWcx4gXEr4Rg83N2+h7TJXfeZS2cexV9
MC9boDD6ILyg51Yy4wdDLDDLbM3+jIDPk6DoUj3fjege14z5dV7s9uT3vYZ+jaIP
4kZFNuEkfQ9mD12dH+m4CLG9EJudns5r9xIPYhDLWAUokLYQlFGwpnffZajVTsWu
rGI5ZD7SBPV8ZLv40w0PyQfiirQHRq3sENergGiFOpFmfPvmh05sVbHKXFbxYoOY
8JyQojHneA9s6UB4fyxMOgwlOkUipTrknTKv/+HoHXe+gnGW2A7g/aNPZHdrJkkQ
c3B704yFJSkTC1etJrvngHdSN6xS6mBFi3u2d0kafBTQyn4RKD6u4cV30rSBEk+m
Mlp26WUmeKc7T3qQ1Sb77wNzU2wCAmXB5kVvOvm+Fa5z44A5ceUQwkPiLXTtFAA1
xT31cLOLfKv9lvfqfg6axp6tsS1WMTQ0mZNMY6pA8/tR2vGmZkzpIhVCp5eEaudT
GY9m6aJIPyR28GWvVWSi4vzPsxBbubpAKAsIKDIpTMs3O7Bn28z4Fix8aooEytm1
3MVYA3w0ASayRiVciRmYhh22FsBVqrMIkJA3URacD2eAdj4QJ2wppEUPxwmfZ8Ff
zMnIQikCP2VJnCi+0u/hKr5iCJpM/qLFGRn2pi02U0TKNlCM4dddYlR3ZIePw3vI
3xmXc7urKpePcCaNnNHCutNU+PLzHjcT6q/LMUJxlkrAAplEC7UzmubV5WiCSB+C
DK83bBaW9Ih7xfQQnLfT3VZVoDKOtFyQM9v1NE6Y14xZZVOdRYxvYew4+pvg85dJ
Gzd+ee0Vc1LTEgKmtTGsjvYxA7ZBKvCUMLb+kc2RrHC9J6mv2FQZkFXHkCna8BdY
taJXqqMJLdtgrHdnEj/qCMOXupicImAZDYAGVTEKY9uzUwlYXcvSeM6ZLeT8wyaV
PsWA+dNm28UU6aKFTozLygnemBP0p8cPWqj2xC2e+u9y/MxOdbW4BlMp/Pi8hiZP
QaKzQT8xY8/RNOJcS562IkIfi3mfjRCeEFO7KXIn6RO/HSRLLo2CeWafo8/f3dU+
BSntzw+fdhJ2G74XHeIK1b2U+Hx3yUC2hW8RESMbVubrqkWXjIp4LIc0xacXNorq
5ivkdfm+J148JsazjhXkazJEsr1OzRxWPZjHsDXunCNy7iyEWG2QkfrTtlDOcSAl
CIFT8YwFgXfUSSzzJ60pYHEvF4CttuCA3mcuupjo/6NhEm1hWuxhSXXmpN6ddZd1
iqEkXRLxBhcXwZpDQ4M7DPjfseQ5+jQasGR9LuisJCCf6fgbH5NUnT9tKuGnTDGl
Fq8HOcofKM0uWzKsigNDLB6LMvzAR/YR83ttaDtb4DYFWvv9qHAzPfdGZ9C6A5JN
XRnddQIcZre+9Kt55iLDnHSrvzSJRvchoUrpXoUiJfVyrJs+nreMvO62E0Bz48SW
Y6O4sEe8wBV20lt3J1n6MsK7jFHcNhzS13sK4zZTl1OmQ8aOWXGS9Vr+/AO8BsCt
0zskvesmMLEz/pNRPXUIo/L9lmet5LD2xZVHmOXSu7xqhwpvVUkVa/laCUyc7t0F
/JmM8nj0UTuevKU99wdV9xFVnqPHVNq/cc1kX3GheObf6parn6w8hsbK2azD8aX2
i1TZLBJ8dWLYoNN0MkTgGzA2VdPLu1BVlIVM0vgIrpnjs3dCsfPQCmz4iq6uvc81
FSyKaK6meqthuS4Wg9jSrLtH6C2B96goKfcu9umgZ2hXpC/0ADlK+CDcOESBsF5o
coeHqledSz7JNWb3NgkRtKemafZ58Q2mFiOCV27JrnR6/rx3wP0DuoFJTWe7Cav2
VquWQoiuXyJ6HTHaCEVOGIvakiDHE5hNI3AxuId9Ssgvj9SU81mIpwFqI33bM4Lv
FgACK0crLcRx5IJAOb2kb9rF+wvp09V8800+bK5icl4LfRNMwAPK5yc+Cdv1xj/h
aWul3FKyUN3DUU237AjEc2D6Ifw1YEzEq/lZshbeUjju17A6ar5NtZ+mYtPUB62V
Q7Yvl71qWYktHqAgraA0Vu52jPN2vlA3ssATvm3IEiIgbXr/k9Lgh0vdEhLMzqiF
0PXANSEJvDm066uYbjF44p3z30Tr/gix/t5Jsnyj3JHd70ZUu9VdtiyrLwIwslJD
2CZ3IWXK36WW621Ku+1e9kjoKX1WBbgSHF8InkSZeZ93Fk72e/ZgB9mGYd7+DTKy
hBznlSJTyEP/FgEkruXXyzqFzy8DgOqJ574E8RCYhpv9k4vKRSVU05L46yhy15GH
W/SZIW0rfsA8qjzznd068KTP1nU5VT94E5QnimMPmrsLByPltCRn+gs/4zc3FvtE
nO18GWPerkci9GoUO8wrXVK4JHtWE5d7YvoHN33NeUw7KnpoXEDqjtR8ZlnHeMY5
vOghWdpGvne2rY/UoyiwU5Kak+kVq7QV+mKv5sgo2X16EPCXSLZr95TX1ADhvUeV
Tl5aUnX8DfpEwb8pOVRdd1lGTqpXI1UZBGWOCfsSdd5UYeXIugre0SOZmbtbIGar
baz7iicoK0FQ0u196ickKDgwAM/vI9c+MHnXSbOGIgFcFUG1CXZDd0uKq2BooH3j
An1WgGgepfrr0LlknRoQ65KH28W+JOum1qvQRfnqdn+AuityLXL7AQSoII/rLyyl
INT1V7Yfv+Lz+85yfLryIHc8hmIFPObjju8sU0JYc/Ts7AlbmwknWn8ZrzJ4VN44
MaY0R9Y57FFdj3u26FlPpgU4W0v2350v3mSfsMI3EQSINMigVtc0Nj/L7cDQu9YW
lHRHr02WtMcitD6N/2cwu5Qa7ntQeniFhl20T+ydhoyVevj/AhTAuCm5VJUnyv7U
i2ztSpSOok62mHCLXVQMO7kl/zF6zasO7HrIzzbA/Luu5hayYVN1hu+Bb7sD8h4M
+CvaLPoP512KCACoS2NEYxT0ugyANsrVxywDo6AP6k8e6mYe09nGLvmWKOuLSfIO
Nu3Dyd68tvGPovA94PlAPaj6lsm4t4LljTNP0x/gs3cOKm0UBTlIBjJXlx60oy7z
QuGXgtT8JDFWhtm7wsmgekzA4Zb05LpTgxD9nWSE7pWft3ZrTZxnwbKJoibaht34
15FX4Bf1K5zaxceHMgXcO0abfOI1isF/WK9Ii72E3oOeisQVBkOIcfA2WoDQ/6jR
KpQiKYovewF27/Qm7PnQxGdEHHC4M+6DHp3u1Fi94I1tAsW9BqNs8PqMCR+/425b
gydTb7VWb2C2h9CZ4F9FVX4LPBNGPHYZQKJYAwPnYSzofpjuWvaqDiesBm7qAU7h
6yQk9gv6khJx+0IYzaWLszwWjgAzVcbwgWey5cBhDDK4nrOBrmQh48gFHheCjrw6
aJC3IhOWkpoleLRtItIWeJmExI5yVTH1V8X83So6YekLTU4FyuASRppxSjmV5CP3
QGCYx4IrLITUsXG1I5ofab4C+xfVUfGjArnl++KBhqhP5sWEp/SQ+Ry1gzDiTXWo
YLX8vU5c1J9xDy1qYndqAx0vdwVfkct9mdVs53KyR4eKZHKexb+ipl17tqSoGT77
vqzt30nGT3alFg6m2Ywf+OHd0mDXe+wuT6UO4Q/0J7hrkXRZY3F6yMckrWaTUInq
mPYvmuuVvG2mM8DD6SupR1Sibbaz02cHv6OisrZjvabm4uR0R8rpyQpBO6+exv6L
90PJ+8T9C1VrGkkODFAktdpDsshUbtwPeRTsHyBjAuAQJ+kDS/wbWrahyiK95VVT
uyUtsBvyomwrmCK1Id1F5XkXdX01PiuSliEeieTEL7GnqTGfVCp8fpSnrcfm6pTg
APA3icCE0wZ4iup1xELqEQaK/3fokQRZXtAFonyeajHpOdlHrc1BfN4qpX7h46j4
ChMBa9MHhAVL5UuBrjwlUB+KTFYhUngn0xwytuwU+91O/Kdfmfqo95kNT+85q3GO
/usF67H+PBVdmErhQfQ8HS2OYEBZeQfX9By7321+e403YduqFYUAwiTmANfAOjG5
EA3QQ520KoqJRH2poBpoc8YPiajvpE0iPlp2UufaeBggRQ+XiOphEQnSmJuhivlY
mUO5yqbXApJjnk9mAdoRBlNfmEdMjtq5iT/eybIDaDdB2uMLYFiDNExvYiQCuJW+
6CcFvtx9hiDL5xlh7b72ZuV2/zOKHJo5Zbj8a8LIE7c5Qq4d5LhH1pBdMIBw6ty1
dT9zoh283KqLTIIaCQcQ5T0VA2tT6SgYaoqlsBJXpCNg2RT9JacFSJ/fDBvHInFA
4uTmrRC26y/uZ8q4VfGpe7uJYg0ndNcnC6M67xVBtD0whNmZsfTNHrZJnMM+wnsm
5hHGTeK+lnogwC7nLalCzLj47nd68qCTC+pzrYUaioF5GEtPWfNRcmXSCh6Mly1o
sV99J6XhQgAD+JAmqZQQ2dNWPrVfVgXJC1j4o9P4xGoHsmR9iAMVUQObbIikb4qe
qrY6Z/4Kdn4vJyUtc1z34O7CLBf7yfeQ1NH1gwDESs4wxr2QCbb05niImCKg7XiR
ZeMa9EOwpUFPnHKyOtd3v56gj85eJ8pi8FdWAcLawLprGNz9UXM8w7GXy8Vt6VD9
NgMADBpAIK19vubjdNzwt7HFZnJnBjw52T2YD08Y+fiYie9yISEX/m067E9EYwH8
sp9/aAtkw9pwBBORmaAYBJ1Qh1UyZ03N3NnHLzuUv6fp45Wm4vO149suIZfUY7dD
Dm20c55RqCxbbA4xqwf4vPNHmfMEFNQVGjFbn/J0ENoihC+4NVUhtcFMAap5KRnv
HWVxVvAi5qZ1IaIU6ZuOWxsKLUySfJbV3M2FinerDpDE12qjr7MzmJKUNC289LCk
A9LanTD5kl4c3w5O0KtipmpdQpyf6wlKBcjl/yimWZl4ANTR8l4KA43BmyWU3P02
JprOvLULaaGMVZ3CwuDrqS02gpx3NDKAz1QvfKZgpKMhDZfnXPPWf7UBMG4Il/ns
aT27Hdt2YZqEsnsGuyUFDNRqzhfrUQFydVx0FbtsO+n8k1VyJwaqYErg63XrCbsA
yTZfgFmljy2TOJmiOI4Ge120extZRvjkdJC0oXG1G0nMuOHI6GKQW/aEuGn/zwIr
3rcX4gpzIhTwOz157HUB9UaJ09mrngUe5LGD6rWREF/uQS7452l43cJKGWQOxWSY
o7yoTtj7gc0KxPbK5kQw0ZXOgmeco5Qx8xrmY+Hk1SpJgqGiGudeh815daHH1THb
0gi58hLK/gqaXfey+PW7AGI2c3CJex8twgjSjPCrJp/6Ra8cl2HvvKrPbnn+hRIl
WIchR3Zica4y8lEEacsdf9FkEn/p5pb9YtqBWoTigoNl0+HcTKEHyUUFflDmN0ju
Y2eXWywyjrgzoJuv76nd18kTZWMvEtKkhIbZFMac5/glBLWqi2dZ5IvlDjKkfOqU
mVzUEVv0nkyGhtu6IUIeo4ALVQWo3l3yMqOt4EQHoBrf4sJcgKje0itMu6+FyCrT
qmwPjZlBoQxhkXLo4hP/Am36mXZX+mR6v7FyIVBLWAueGvQzlBgS+eKd+Co7d5pX
3Q26Lu7Eop4e3IOYnzf/BAP9lyvSLyrcxcQgGTM4puLpnxE2yNapJhE6XqN8hpx0
xVqJx6DPlEZ81oyPQ7DcMF5LKNtT4YFAn9RbEb8cjdDXjYOmAvrQ7XydVkYe8xAP
RGa86hVqYBdBU39nOtR1GadmWA8scwkt6Fg42W+9KWR04hC6QwmGjZHE2Pm2jTz6
3jTHE2SqW8WFn9GAsMw2P6bNDGd7Hkm822FuCmndIIrBXziRj+YMLwtfr0hk9DLb
cGAku9JM4Q+sYPMJyTqNo6ytW+5ZGrRxwB0kLbKpt+XQqUu5pp01CKdBOiPBG4iW
ByuzgdbsN6EmbRRCqplspwksw8EMgYANTCq0lq1ipGcCt/TCMMxEdVxFkXz0WXpG
eV/awYUOdgGm5P8KU9xsJ+mnX+hqR7GuCMVly1TEZVXB7IViyBjl2VxBrggN3KuC
b8rvP0u5RObjPeIFi2aClgQiLdJ0TQgNJOjEI2/SafenKNAE5/Z7+x66JvkGW/Gi
/5ObCHeQRO9djjE0k+OX21RRy+GWAuoaal6hEUoXpR6Fuyrt9pW/LjG9zLByHzH1
ROgCIhi/57gIdiG4dvygCVMjLVDhvtGRLKGt4i27UUJgJab4IdF7XV2E3zY1yrc6
Chv7otZL3XQWIaFuAiQxjk+O/D4GfvGJtH3Wt/mC6Vlxs9ncnEaKO/nZhdnIqlik
nTdhPkqzk0FR2raI1RP+MIKQ9bMr+kK2jA1xCwMIpptf+Y12lOyfcB4xy8WcQElq
vaH/NTrNY7ydaFOLOqBxGo5DH3Zs0JCAdUhvKsJTRP5uSUlhZCXB/g39yuzwJm+W
xotGywT7jAlsZnQUbQU1LlkNy6igmTLdOHT5xhzYgCPxORVNTrAYw/cVjHbCl+/d
EizsS8Ierf1EdB4ERujP9Yvlgxe3i+zXmiXpoDofmGhFW28UAmRkrd08ylVfbfJF
DRwFy1W4tYAKJ2d8yD9Db1FRUWweJvhAXHvVcGbLW/kXZmKDX54+BGlbS3a0V91p
uiqE2+T5cscXEArzdMlFPgfQpvjrp50dc/2GUw4aQRvjd707m9YB1CI1zE+zCYyj
p34th5yYc/SPpDQsyyKT1f0O9boKAl2wo1dDQME47/dzEj/WKqJFam/lQQfT+pBc
5AXBxAzV1+tud9T6edYAUPR6vZfXVyPaOzcT4OfBfdZ8Dcd3R3ZYd/6y92T1kmlA
K7bi1yEbv/mYYhb110KIaDO4utbr3K8PQ8mw6GZ1fFcq5SlPDPr5aZVYk0+FBbKN
jjkWFf/YObHVTfTVJYSpMGmum53TQNCQE3lKS3yZ5KlqdDXD0T9K/9Fc2h+Jz5Xd
UnnjpnrORXFkrNdNLCx0TtTtF0GTIoXlE5XR56PcyZD0zC7CdkPHuJfdHCV9oM2X
2XI9BELgZgVaXTXE7RRzy5UUp+fBsA1Iz+AesUDjblRo84WAHAoNh+IMRdUTNC4D
ODS0nc658NrbunMDFKeonDnHBgzg6wKAd3xyyyqaLCa2Nueb7aMqf7M+s8vuqNnE
Rs3VINQK4KSgmdVJTimuC9wBW/OOi00Eyy6IzrD1vn8k2/FWq3HakwDTcBG2McyS
0eJZuLmecVE/ndeZzzKqm9yVFOku4ATWRnKRqka+jjC6pFqLomNAA2p5ZFkGsBQX
TpTgvzyl46U85DE4OPWHWBlCkOcqJlq2gXDTO6ie/Jn3hvc4XMslgQMXNb/NXE04
m/zxlSexBu88UJaHDL0pMafHQaUK1HJdk+0luIOSMRbPZYcVy+PuX4DBqMEqGaHV
4XIL61YIP39SpiPiExI0zmEbWAX5iWHVkagbSXbsgMydmDbagmXXbRB2qr5Xgx9N
2JgAx+3FXXNNB+p6BYGVNvMsaRwGoUOTLqG6nFCBPHfqwlO5pgvX8OfbqdzJ0avI
vB2GNNv/gbS78DCxA5cuCwpds8dbq4rBWmcQPPmR9jB/57EYlDzp6sth8p1w2ujK
+qon2C6n1YKV0WFms//RtRmwpJjfxCLPZ53X6/k1WYdpuIjSu6PveiWS1JJJVo15
up3Ip2bl2FbzbZLx/z/1PS0jnsxrOZuQ8tF2TBaw2K8wgUYFSUCp2zJNpikrsoth
6ilHfyI8EyG/j4cmxu0MJRKSDlLJtl/7M6u2Do/cDBo/RAu24USjJXvToTacQXUG
Jx+BhkE7mMW/X5Zvd87afe7E4NujUGob58PGsU8R9POeprbknTp5vbE1CO9KBzm6
kfjZ1WnOiA1nD06nY6SquqYoT5q/vzayfAkeEsOx/LKbrHKsEeDrGObtQ5TumCU0
kf4dsK16rLFztsHufUVbial7vDavya9BGpd7ckII7/J938zy7MNEaDFr8YkaHqy1
ZjilAtGMT6ygYnHPJkXejjSeOAg4sKgFcnPiT/S1FblbWDx2NXWSqnQ5lEqrvkRB
OSYfLRDFabK6aYanKtCkbm4L8uDpPXuVwx5gY2qOJARd9tDCbaYSTttAxTu5+XNP
UIxShsXrm0J+gZGIROrxWUI1B+O/LDhM+yQMx/8YohghEqzDzGQxa7Sktt50LqjH
xmjXniSrRbxuMLJ9bhEqCZ00resq2FJjXw4MhEQ4rTVCeiEHbcEGLYyyaC/037hS
NYL5XHhKddoH6yc+Ou9zYDU+q9WCLD8hRybTY5hNXbU/f1aF4B1G5j+9cftKFMR3
1Z2eKFKdRbXT0w9t0HGzlCy7s5Vhap1Haem+6Y5s+gBaeZPue/VrZ8WjCaWK1KjQ
xMF7dtXK7WhPEk2vudQDivqFIa073qE8G9AfK16g+7ch9ewgdLzkM9lliuf6ND9O
dZQuKmKMuftUJ9V2A9sLOI2mFcaj8zZvbuBCC6BKojx/wtw6z+KYjQu8rv2zdu8j
TAoj9ZctHX3d5MH+iMUWkyd+EdXU+XqMN2Ia9jSDg/SuyyU4G46zqAzO5WoKaDYy
klKB6Qul4RQphVzdHJLZzVCx/BPgThCD5o5V7asox84Se0PPDiSSYfNzq2VSe9ez
N3irZCp4zdwvh7ORywVyvqdgJvcJKmZCErA7++J9R7xayQfnIZPXEQcSGS+pGoqa
NC4GOlwmYBTjf4Oa7z23PJ1isL37TqqO+P/GVvC0ZZiD1ZWn/94YXj90noWWtLho
s3RlWB1WJXnJD2n4ErNjpROXX7ywR7bFgLRLN5urwkxrz8wj4x+SyyDcTISe6s40
lId64pCK+MdXHr9spqQp90I9In73d04fEZ4762TiEt5OTctxxUweae8yYAtXpPzQ
FgRWJ56hAXtvYUUuJXbYJaqkNoal+z6OS/OyiijHOR9+spAOBFkpEhe68xFoETjh
8qacpfd2nhOoloxA2hDfA2wlstbTGchjutHTYgMdtm2yAmrKJnQwvwr6VGIGl6sv
ggMO7ER+ezf24qQDwCoK8yuXpFVYDnQ+nd/oY7ZhRmdv0i+DIvIh9c0RIrCsx3Vl
OK2YrppKj8k1oYs1v65MlKBg/TpjaO+OvZmSISg1NRtBcSX0pQYSrgPfiotahROB
qmAGuC1iNeLROWkTSJ5i3cFw6drveHtQV5IFGVygVm+iBVvETx+g3UKVRiIq9BxH
jfDRW6mKHRYCTtmE8qeQBm1WNzA4F/T0xwMMuWR52Sx281IjhNi1eEdkcciGtq0F
aStldIZ4YhlUTHNOeb022YYozlNnEw+WVNXfjE6hHSnDo2WV6P637GnzVTd0A2jR
thsQQQsGDCo3CFmUUpGV7HOpGpiVtmh7rl+YVssQtm/ni+rPqPeRd5vsuJy0H6wy
jQoyEwsJaKBfHMT0AnCLtdsYeXqsBN2cUs7+32qec8+I0oWXSTAFwjeIVl2g6IA8
caWEOCraFUjxMO0dTb4WKeHjDvdFJYmJSTNpcKnDph6cdE8BlpTbTiEa4Sbz1kU9
a+ZHpXE2BADbKobbbJ9SX0+mG/cBbL+7Yj3zdDH+2oYCLB14K7sKPIHjzgTANNd7
8mI4w77Nhd6dNYm2wJAPtwvzgVNtQI7O/GivamUk60E2t4mjSNcM1y4d3/qjLcUr
vOhDLF6IIa1XX2MTdtqFw4n0awG9cCWSBlP0glsg/D6UbOzcyTgyifkue2fHhK8H
rQ8fPcOk8sDHJVJTyRCGzd8EEQZ+wXR++U4858OZCin5qxsOpYsunCM/ghow+9cd
tMsIj1d12DaSeiKzcuORMsbtPl+v6iYESnQNByF2chfgsayWgf+t/MXfS6cuXLHv
9xV6rNFlxb3hyZ7P9CBsIMW8XWQiGp5HWk6F0Znapi6OML4MByZ9JGJDfk4z7SUN
DPZ3JVePw1X+8F2A2rvY7kDc/Al9l5zzH7hspWNHP+DMKsamXPk8dWkZCtvHzOXi
Bkno1Qf828Zh7mQW0XG9j5xIuD8WnlgXqppS1NSxVMWkywk5qHqsbIMGiNgdQ8xS
VQXyPVxamOCvmI7Zj7HBED0m2wKzxLJkxNtazjFGZnOZlHF43nmCuBKE3R+CrEce
HOZ0G53qhfbkS+utTaTQ2Uk/Ix2Zam3iSRIsf1VeTeIv3SMHivZ7W0nIrTBPDeDg
xZKVSf5h0L+vbEk0P4NjYI0fx2T0tg+YFFof/EqkJpj5c0UlMgLunWcnwShp4v/l
CqmKEXGPSDuBI36HId6ac5Sg903hyAb3vceqqXwXbGu8glzTkp4Gb5JfyiBT8TA3
1KPct5xwLSWhd2rs7DAEqTqU5Q8ackuAZVDfPUn2PYjtG4Kx5ZENsBf1g20t51sE
OgA3ZI31lfMEYY0vY8fFNLPrQoQOlqmlxzcaUhCXlXLMxwPlS1RU5jQsFzgxeVgf
2lRIuQUbrNIxwdEYER5e5sKhJec7LmCj0VZUM6pZWpAxkq/mp+MWz5mFFyM9XJqI
r2x+qy6UMKkYb0tHltC94crW7R9p7bk7ZdREgR14idV1jAz5jgi6mAusUM620GHe
/jrEO4kqX4cpRWUGO5Z/udanT/ABG3/043+TFPYWW02SWonUcFFLrbYTQJg+DBgy
olPOrd/pi+dh3gTERUkJsRg3p6e6e5D5IDEgGgVjwOKcKepxPcS2/M0G/i9lawTu
NQY9y1uSjPtQhE7935NfnMmTpRJKORIVKDECD29TdEWo7U7jHctjrgzsuGzEX6u+
8Ez6NAYPzVI4LKEcMSi3otCpgnEWnaO6SX9byzk/A7LNG34G5Ba9c1PPjys+wRrP
h9lp1mmIxlmKC4mWfbP8pFXVcnLLKRUx0R98I0G3d0wFCPlNndfvQI9Nfr5ubQt+
C9N0BGD/vNECKB1uEApCqUKjZcD1uF2up5MT8wM0gEKUUNy2k0BDSq+YXaOji9EB
aJiuJ8VzN/49rm3KS3HzpzGX1mwVEKv87zilLpF1jjtglOGREHJxlH6W3pek7+Iu
vNlNf802M4UqbUTbhMuefEsCxFNPd++zbQk5A6Hy3HqGCu5dxPnSqAjuj1y/eTce
e8byeax9XuMcBMUtszR7k2hGPd2psboKwVuyYC3BgHEgtkBoatTe/yc+snPpz5Ni
SXO+rnUiGyGdt6NXp70D/P4K0w4KbS5TZMFK/MdOeR3hgcuOMtUUUdfEW2+aJ2ii
mkuUk5XK2Ve+bcsMG8p8YmlONmOQMSB1jRpIqOw6q9n/1RyMNH6af1RvNYeuJAc1
e7HMdxSXy8smuO/rdRuoX7upJMka2DeepsILOl+QGQpR0AbT1BdJKUWaovIE+dQw
wssUg2kjG/e/RZeU9zczo59l/QzZZTNZhCrbA6OtQqHwm/GEXC77hkBiNWEwJDfP
gtx98AplOfkaQHis2lvNfVFC9uN1xlJdn8+mV9jjckI68ZlK4/sNj8et7WRtihBM
lu2xb87/V9R/z6vWBH2orNy8adHGxlHLLgHzhpM1VjzK+7l2S63ERS9qqGRdnq8T
+v0Ak1+7+dkPANZt06zrtqrivO8xtpiSXPOnlFQgjsPEZ62VszeUpqOQSv8XCLhD
ILV9UjcbmPHiHEQNvyGhQD78FriU9glrBOW7o/30TM7TilZmJCP9CUndk8vSRYc9
jD3jPLLiEwNyLPR1u2NRXUZMXpK77FiQxWmlHs7Tv3BkruA2qMEIqYqhjrMZADMK
Hmjmz47pcX8SRqSw+yrhkY66AbBk+4KZyae8Xu5Uz37HXuEGMphWB3lUJKssfK42
YtU5t17kommuCoi546vVNeKfcbg/qjYIs9Vwl/Msk8GU7YyOCilmNbl8xlgW3Kqk
rqep9ZsURUUuzjQdUcKzoKflKy0XA5qOw4srZbD4U+nTClG+7/VKt489Q+2EkWWX
QNitHJ823J9eiV9zEXmFLwZONR1Ce48s9gjAxlHX0CRYapunuGtLytm5Lxd0hdas
waa2ThF63pZ5S5PURkJVuXsLzPnkWkN6M6/Sf2bmwDWq18BikXRtBUIcHqRbQzq8
cj4jwYi4Hic/ihRZNPSvpn/Ld5FVG5cvnyhAYFtzNuLjZKZLflM4bU3izbaQlpOS
S30blO+5XRknDHqisFdhIirkPMae1K4ajDOXHvutS1FVNLvGThf3shT4Q3nkL3vW
/6frUJDdDHc+bNUfUXXgPkWUqfJRx/m5/bUcnnUoeZwlcAmQAtJZonCT0o4rQpnq
fpNX6XaakpeZVfE1vzyJ9RxIfkFitfDlNd0yD7J0gLbf/tfZGAImzmutlR877p4h
xUdIldxTVITKIV5T+R0cmRE46bE8/CXtotlxjALJmLtZL6ktEaHIu9lowYjNI7Bt
FmfnM5EQt90xco7Z79rKgJaMS2DNzkkPQJGirJjJFUIlaGq72FpPyzIEgW8fbqxq
TjeOUKn/aCRjLg8GGOTW6bJhYBFjm+ilAh8aNf/rmq8g5Mr2wcypQsoX81/boclD
wKcOlR7Mq1X/lnjIX/CAVBBlAkovcBX783oyWvLIlNZn5/M8TNlkCAq+WJIh/lXZ
DE/mBjO+ckbTpPUL12ENd9YidOYlhM90OR5GooRuTBwG54U4ipbUnlrsYlsP2sFD
NIDyL9+MjbpOkW9FDP8XfY0PqWxDzp5U2A7ZUZmGNToUjx22prURvRtMg+QSJaWJ
ViAnb8Gf5QiIMI+iYdhAQaEQNUtWyAAHgIdAFQ/0xIeyB2gV/jb4pu2M7PNb/KJ8
QWXPEzUEKcwXtEqAP8Oe/q8ilsGGcW3i18+j6jR6zWIUhf8ZYyQ6HHfRNZ/SasIi
8JiMz9rNpVX4DW3AwspqKBPXWD5oEMUse39jDx0Z1CIor0ZhGtx/Xj4q7fG/wcfi
48q/6Feb4e/OCW/e+d+aep33+rHZOisDjBmK1cVqxFrIbkZIIHvUfHl69d04stbp
Z6Gee6cHZPJ5w+ry+RluNFc1ohev72COdjlS8XNyb8ZHuf8ok6MMDXap3/lwXtfZ
vi7rMTPQdLaDDdgJySlFCBeoveicNDCcdbt3KfvwQf3l0ruy2svDEV1CJGR0NTbm
Ym1+LAe7fFlIb01rUQXbNoZlFje7n9RtzPnEM868Nb5Y3Jn+ky2puKmuBJV/cFtw
NN6M/PSTdphZ73FsJMR8Gw4DE+fhUnPlnoWhVrN3SWMizW8QOcf3NStsxvIkYz9d
Kk53bO47K6jaSwjkfMjB0/D28mReDqw7gYoQqFEYPq7AEfz9Xxsj4RKapvRAFMzy
gfzjQ2QBEI77lcn0bfB+Jq7BmixJPv1JSQ7pXr990SqnN3KbuTRbFD35zVwJ4F88
q9N+xfVGJGqsMNDhW/ROHKeXd1cbpOu9ycQGcGFJ/H9fYDwaXpr3kz1WTX0cH8WR
U6XelOJNOT41jgkYvYSftPM3N0zoz1ECa5XK8R+wqV+6DLLO/grlw8KeNkORytHN
xMOujpMHHEmB6a4oGCxiDx9yHJpTYaG3vL3n1jZ3qJDkgzcQ4f7MdG+Zh7lQegNB
z+NZRVrgJwc56iwd35e++zmOBmjLrV5h+uFJkgZwB+U3MvMo7praX6jnXBSrlPgB
8tDLGAVc5Bmam/Ih5DT2aK4e0eteyqNPQGbDvZ/hOCKX8zIupvNZixdEzzRv4mWt
zTqDALOXw9VAx5ocW4PFSlhwNrpte099tIZ/lzPquZYRUjESabz8L5OLjlhyOz1N
iu9+03DIsp9iXY8CF9ovhrFfAwcE8IWj8k3smZg63Yo26ZuHq5Zr9DAKzx5Sqnp7
X4t2OGUz1bcgO8H+yDWlWs9m/2IA3CtJG5RMpO9fK1Nzfd3XTTMF6xm0VJbfGFLv
PNy+njvtg21o4vMwH+7Vkwn5VT0jXDFMoYRjPb18F6XjDFSDo1d58JUBsdJdI6sR
Q9CeYMOzrx8UHQGsaeMQQsX4f+jU/Wq+x/Zx+/re/PGHVumSjeNYGRwpOKJqcjJa
K6phvnucP9LwuVI3OfOOHZAZZgAlFmBFZiXO0ONZdp7PZwWgUANWNkBWdkWyxsL/
4QzAwwiBQakhvwxP909EeXfIQO8xDcaZp6X/riXUFQZ4AS6XNbk9HrTlN6YCz4Jk
TXq4g+bFJaf8Z4N4C+bKKqdsqu9s+bjyWpVpzqHiyq+ipXuotMRBA8+BufllrwK6
dqh6xVPqUuEYT4CAhkYFaJyAwWElLplLflfwc+FcPK+CwG2zKXE1DTvw53vI2Zry
fg9z9bvNMtnX76n3HiC6HmU6Wsidy0iYV9Das0kZa9xqM0CfezvBkn/qn9z6xYCa
p3ePXvpxjZtremQTtjH0YJ84/2ICnkpQB1znyZnyqT1FrqvEBR4ga9RnFaqU42DN
X8y+BRNXkyqHTJIlyjtj9t08SxLc0Ans4yR9nnKcvDxh6UuET3UczOW8A2cOOvXL
2BkHRwE4snbKldVz7Nhqkfj0mYhZayKQ9JQ4BSQpjnwa7xRvwcbCZ2X+pyMoglxT
sv2o3QtS+YwDmIXmBdUiD/gs7SmZnCupL/yEJVpo5ex5+GKEHECW9Kvtgn6RbOvH
nQlJRIJayM/N6QYbXV0pi0+IiJU2DsJCDthhBj1Dpk/vgsY0IAIDmgrhOAStkQva
quNzGy+GOmYFvIsFF/vRcljNTw/eBWnwmJKuNPP92ZFEf0JTk48hD+aa60bCO0e1
FQMIGw1hySpv3wUEoHDToe+vxQ7o28Ma2xF59EgxLAN9Mgj7a+b9nT2I0q4L8VGO
bItuFRJenl/YzM6vW5JnNUBaeKbGJ4fa/BNUcYVJ9LsIXivrRKrIZyB4DiULDZcA
v0q6Rd2BSIzJ/jQf7PiS7ptQwpfumCVOm+ldNX8T9iua0ekGFUDz0K4uTWOTnaES
18Wqrn0W1egunH0PPBxYghLExJF/OCiXZZSKdnM2H8POQdO8ZQu5EC4ymSlTa/z2
IaV+OQe99yGOmuJXNYfiDg7H8Y+AWaLHawNbCzMAdlntJGnB9GLN6JbIroZg5+JY
tcblpdC6CcqqOTlaeDyPRZLtH6/s+Q25kc8OkJDrm97QRu4gQUg8G3aKDAoxKMB7
zLuOU+dtPmLu0Pv2I7eZXViR8KTKnnQwvfg+cUoC+R6t6FVF2pw2pgI2m7Whb5d6
jZ7kjWVMJvIQ4wTn5rkq8FTDf0YzjqiXaA8CxAp1M+WIqiX3tmLgV3CX20Q0IbKS
8AoVocxaNxSI/MpTrfU/B72NK8kkeza4cHSeMPkX0R2hOgEr0kGfBotjcOTF4f0g
NNtvkDcny8KCzCCKjsQyNm9pFJLqJTmtovxW7sQKIX2HhAcCrXiXnepqhYsRpYx3
u+lca76T/I9rMy17MWrCopUWmspvBKma6d2pd1+JIsQawXf/Hr7P4ly1AsgqGteA
IaoSAQrcOjHW9N5psrdfWjiit5Kru5RJqa9cesePvwOAvoqUw5QVWNNXYURMiEa/
z5yfzKvtu4Irs7gEIagYSg629CZF/s2fzu00+MDPm9jKyMZryhf1w6tLK6orq9Jn
2CiBbK27IqJRtUKlREbAhswZpkY/dHNUmFDjL9oQI8HULyGTRgJi15u9e1WSJeE2
fZEtnb7HfKRpCRwmH41BDL+VhInqjLbklQyGwenWEfBtgFot4k0/WnWcz6S83mmE
hMIOjyk6m1Etm9rNZiV/8P0fQRhtkhDt8QJ9oq80f5lq/4CzV3rEBeHoGR63e3IY
QJ5UGYxTL7/07Z3361K8xuAPgXBGWZn5npWMK5d2LCpD33s8qSzArMFknuGL1zUO
ixECnax3n1pdqb75diKBeBYwmGGK7ztgFDMLaty+uiciW+XvJPvWGxUbZ7nU1mhV
DWes6pRXIvE4eKLn5QY+A/9bx7TuQ1RcV1EY6DH5EJrq9yAfuNoDUcYKqKqsFkJZ
EUhMF4mHZuuDz4DRdZgdgFTmP3G8+cQ/YxLIM/5YT4nC8IMR1PX9b/cERC1ZkGS8
RP3nHm08gPq5V38DdOw7PLVyLR5nxSzzNQrMX5DnoJXVEqRplI1aTAFgyMgppDL4
wcAvM5qLkouSl+eSji9gwl2pbdlrbwl1nahlX20vQCwN0ziXEluuGHrQ4EQhXjVQ
OZpv2wgNPcOi6F7Mecddr0tm4x3R0CCO6It3303WKRjabAmMtDnpdID89OQ375en
unAj9q545gtqrLucEWIIYrSaN0o+JoOzSfV6b9m54blUc4KEJHdUI7ixnhRKqB5Z
j8TTdWEljgyZ7D9UpGlBeD4S9mkwLEjSaKtYtU/gxs5XvhgfN8KkwB/ME8N2USTA
LLNkuaU0Jsju3KVDeRCAy/qtPGqwetMjSdj0MvFZtR3wkuykvgk/3icul+b716xJ
VcQ2vGUwbGz3MF/vyJ2J4Mw/OjjfFS5lMTqhaLVKleVIyTKG3TUPi3/l2kkYoJ4g
398y+J6+kKJJlN132sSQOSzvLy+FIsmUUIrv4ZPXQzE8h9Awf+AQKqeh5IVu0VTn
rphQn1LEOvDqsB/aa0KHDs7/MFUUuF9O3KB6Zyyx7rFaRN1sh+wanMk/3sy4Lq/D
3irrXqWuV1WKVTTFkf27mp9SvfODshY+NeejJk2yJ4ZnxlHOQ67lf6L6sh1KupW/
OE4RLWDmzgzcA4SoUr45TZe5vpl/hybV6FFHA2E1BaFfZc1mLMggzYHV2fiZzMJm
rJCkhZbUlb09X5TM45EDopDlRtGVLE8nT9dW/n4arUf/aj+LvuVQUfHuAdaW84sN
OpyNq6xKETZ6dSxEJ8B+Sy+o1UcmpQJeURMfobNDeGXepAcLWe8SzH9sFPiNO5AL
bc45MtPfvWgTiKzyoVFUnLyTuNyUQKUTAP3adDWJ++UIYwNP9oroX/Ld58tY8wY8
zLYoNiUKHo8EnpG0QXd0bwfrpGRCqBp1bvQTfEnzDPdbWU0bS8o6mas8JktBF7Gk
r31hgIK39qLu4080ifeZtKW1qhsWHb0tXBBYakEQOk9EoUvCh7HDvzjoxDOV2t+L
KcfLDxU3jZf2uCJVY4o9AkZTRvouLLJwKLgUQAPhLsVyUmz3886mqklom8uwHLf2
rYG8ZpFw1rWBhr1HlUR5PyBJSCBwvIwyZIoDDwaDEEiOvbz9urIcrJevz3JU1OOG
I44z135p9KQfM3VQqAUhoBkbhZkdbSxZDwtn3gDxg0zFacOp0q9/5zRgYx0P0RtI
QKoRW4XwSe6EWg20R9chBTxCW4bdJed4xPg03lXvs+92tMajE38ChN+/x7dHWlVN
IlY5OSykBzq4yVmS6QTIB6sT8Ps8sJzxLiUeW4DSaFvLQH40aVhO9xUlJsBjuhIJ
Z5vFrHeWGfbbIJGD2e5ugskKblSbCzJSDktG+IgOwTdiI0VbnJGaf6EtezQvdw/p
DJx2QfBg2+YoZMK0W0Al4dAFYyz/GudpTn5buHgEf+23DK7ek3WeBm+e74OFrl4u
YipMA6+ngKndfVLg5BZVZgoRXtgH2QyVs9z/nxO2+z52wdPIy1XcKfYW78ij/Tc3
x2Rmi5hclKHCjo2fetk+l6mWThG0B/5OATHBAt0woVTgoF3kVazXXfGJ7g9ZCiTb
bBDBcovCFOaXbZbMRRzEU6Y9YcXEWaer1B3DCrI7e6MhMsd2wI7MyxncqJXEGFgz
SStivEx8qvB3P/8h5zHa7c84C0Yh2UiOwrkQjZzsaBdpfgNSM/IquGo6T5v1Qz4z
HrwRQnQZYhbHcUoEKIVb3yYd/wVYtu3eJyZqZg6o7ALUrJQBwi+ZGwuzI28aIX0t
8EeoEfN1t9+4xd3kNDKa/wWP9BxbtG4arRRovo/6avHaoeGjtqlA7INZ9W0OHcCS
u7CoY1e1+GcLluPRBhPkdMNzNPCr1TWIFXD++Yh02VQcKqbajI5l9tVyvXT1emU0
7eN1/trbheh2KfvZ4TvCaxMKI3AZF50INbP2FHxtQoudJnM5Ql54KqzVdiNggzue
3BkyzMA704MBnOKXJGFb2rtj4X+oXEGrcWGemoNh7E3vT9WgUtYXBc6BcctWA9sN
B4FINhkSyPg4NeUob17NfBbKYlTO90GpwgDlNrX3YjRIa0nhHNZAUEXI4J0a1F24
jCV9ZKvxvqNqsLpI4kUwK2KIdEuyLWKfaGrmpt/DGzV5BZ2zIvL1kB5M4W2Z2+Hr
8/Fac4fhDVIZEmJZQvWyihlIeT/iUPE0+wf7jpafH3np9gvPv0UjILWX/JbzOIW5
2ry5hxwDHVrYHZYgOv+R43ZdXr3fAsc47YZXexn5jswYf6MdomLGsolWPBWv6uLV
ozwNT55h+bkEIYgsWY3pd1uzhdizGZVfPkrbrfzNIojcbUpZ+08hLQFeUCoWiIHJ
/oGwdiTPsPLqaito8kqsjCOFkarwlw3qmxgsin02Izf9hDIxWyUvvzu9CvCt8bsI
n5hpRtSjuNLeAwYRSbmH9A81TbPOcGTiVjgw+onqBDcCm78bgIG1Ob/DS+66/Qxb
8G9dZk+KqTR6iw8xqSwg3wY1jqTfRrCmA2hNH8+Wr3UIjhEfUMndk6nU9IVz7CKO
/9M8OekRllCglsdSq7UhpMaZmQk7G51InTNhn+bnFgGkEA+mle/6WT8y4NTigu+P
fsiuuP6GYVLijX3d0i5BEIzyiAhonWRPod2q6QWxzo2ymcXJ3kn7nCbmKs2QSvyB
pc1NHtfu85VKDRoQTbEq7MtysV8NnRmeX0GIQJHlqS2VdRMFwHAGt97odgma8x/w
5bdvzmtVhSlK+VmxQY884eTHfIycvdDm4gA/NDg4v2tD3WjH/QeL91UWY6fhdqur
c60ilPr5INgVEUMj7NaGF189Ej/HDJxrn5J+uZYWliav6eru90i7uWdseCMmrqLg
YiQu/aTg+biysLtkq4zkMiwdW4nuUvRDo7OdAmo2D4ykTSugf88/BhQQluKw+KbP
TBJW0UBAqHZdYgm2zSURgoh9FZqtxxryCwtnMXr1vUse/S/zHChWSARg9RurldkL
rpVKkP8mEi3MzK8HE7fUFRoCZ+8mp8mT4glfBd19M0hB5VLH1C3x8FJLrV+OYcSq
foibsyTtye3xVahXnBgOWUvN61wdlUcyzB0VVHUVdIduPlTt9grWzPu5y4y+NcVK
JvECfIKUsOxtSaKUEo2CWlG9wBRMeeWufGydbYqxN1t7VrbrtQC0urdWm1q4fupX
AldW58OYHZTczyRX8JvowJe9ODBJOjVG0PVxzgjoq2yPm3in41ctqXbNbexaSYnV
TdpFR+8zgZ9l+pyRRQ7mPhez0mn5CkXCsIxdi7Oq3e19l4n4UdgvPdiqyMe2gk5K
MPsEXqFImDiDlDiU6OCqvylT/9ZZAx4v7yiIFjhHOrMAeg4UK+U39M+jNNVaAA1Y
6ahzHbKjbNUM+u8cm5EDrDAlEwX4jnrxBrCCLO5lqCb3rvyPPh78TaUaxIdcvsFZ
Hz+sySTxnu04OH8vcRJvoQAX95CbgawC+7RgYZhBaYkMT03AtLONYkuWztu+z6t+
bgFxOZUeJyWl1zANVVriRGU5BV/NJ565w0QdI8fTTc1kfPTPMscuXWFvfyVZAE98
qDejEs6oyepqgp5dUEQQjLMqwap4QKRAV4ThI08fRkN+BJN3p4YTTAmfZghCDBlP
lktzeMP5fAdwlEyq/20P00GpOO20v2GK+2TgWc1FbcDrb0rNKC5+vSuef9CRX79h
wert6Cmfv82dhfolKRcBSuGtsVbq0sohPgFpS6FEMHIK5aof/HPcs679b17a9S8G
wip5ai515mraZzVc5FZeLP+zus0+kJkZee+63kTNGBv+ELVcduMocjyYtqHnRVLQ
rPU67ZMUdep5Dk+yF+/TQ6gE3lh3ZPpKL/jP3URhaSTkL7gEeuSo0696quuv3KBS
f6M9iFKY4bM0k896hJlRyRva8pwBuYVI5dT/gzE/z+u/NCn6zJGVELh2Xx22w9Qm
azjg3ulJl51t4hE2L3PNIF5jeiiUxoDTYJ+lMXa2nybKpnXsRZC4Z9w3o00irapX
rvZNeZ6sa4gcGP7osbXqBQOYTv29E+yrlPV0Wdc/TqKCVtxj5GZTrmWvlWaoPqTg
6I1h5GnP8FqKPjVEWPOH+stFpilY1gl7+kdFpW4auywatpb40Li3+xvajuKwunUe
bBAM0d1MFvNJjpt10CzSm1cOWM5bYvln5gAr+ig0poer1PyENs6Csj8JJzAAQpHw
EPIvHRVcGJfarCejhy16EJiwee69a7l+EjetZ/ENFalK4181fTGPrgNq9lf7MpOv
XYrIGRIEt11nEZTQALXHIH42Q50nU+1V9QNAISK9MQ0r07BBkq5gDTSqdX/4e288
yHegVBIw/l3r+r6xpH2vCadqeEBJV0Dqz4PPIYmXHyguG18xDmcJe7cXu90sCnRj
MWVxcFyk+KgL3KAV5ruSJiG6pdfr5TfpYptuXaovyn4Vba2muieBzzNllWe0p2KC
z3w0MZogQTNzVgaaTOrd2inhs+j72TkuHpWvAc+Ek+NnRXsSRlQRj5WXtWL650Zc
uebfiNp9AcfNc0e/75M3Maosb1m3PxVfdT6yHt7pH3XabVPu5TXvM7QnLSTVXFWi
IOn/w+hZvEa68Wa3We+bjhtn2VzCVMlF+RTMfT23xx2zTqQ93X4rwIC6kzIchTpZ
IpFbHa8YjPC5KSrsjeWFfyUYWOKGIb5y1VXCKHZqLeYYIQNFw3Mzyfcd6TwTlz4r
12QHOoCpx1i8Q7DiINP9HrpmpwGzLRdJqQERNTn2c6+px/choVUbmJ0zKpgqw415
Int6NFKTEW0GVo4imhJ1QNwKqJYKJOfQSKA095VRLtm6MasObRFPBOUzhD5vxRbU
8m1W+yeAi8q65YFXkmoKRL2U79ptmpl5aAtScihnL1iafyIzoC3vY+LRlQEpaoGt
mvbl/xN/9cVaMT3gsj7fgGP03dw322yoYYTmMXh771yBVPzEyE7nL+GdSRXW3HyZ
z9oxgLCkOTG/YIctb0pxhwVXjGDsyxtlDYzgdcN1Gwp4ZuQTAB2YU0AL4fPFAMGl
9cK3zfMwwzQ4wBuwvz5pEUjLh6BHkufI9zxz1Znb402Q08tIhUudwcbOvqb9/yBu
MNE5ShEjE42hEXHL+L2TEDU8w29QL3c2hHAaIaNCDbmulyJmkRfOcCrPrgapDoeQ
IoKmaQa/NxSWwOWl5Qt1gZUvsMH0jDAgTviQTkEt0fzgKOJHtmSpUh/lwXdQAjYg
Q1P2A/zE9sjibZQjoR+2+G0kzpZbv+XVnf3oLza77KJj2GWbvjXKcooPYcoT/PGM
VHc2/FYkXy8nlgyhyHJhfwtWFF6zxwLoQaKQ3rCyOqoRHAsrYxcrRBLb+Pvi0C63
gBbQUb5despkfe/jajHTG2oSnEVSyjth5pgvecOSf3i72HhK74N5kWJJjf0jkZ2P
RdwxmN7nknSGyeiujrcKAy/ooCJgLPR+l2MLBgRKd/7STQ3qHfEgDZ7MyFICfNm6
tEyg0rah/6VcFemrn03JY/CJWVPE+J3tUD3ahrFMA8CUXQFt5eoFPWbyY92MZVKc
abv69SECyBOo8ITBn9bUJB0kRR0j0E6HaqjNAqgAsdxgGvWFguIPn2gU2S5GYaXu
8fwuMJBRaNnZQsSl8gkcA1tzUi7UHekSlSsI1AL79JIl5PM82cIzr3WdP/OOdjjM
KO/mJ0RJ3lOs+6tHtB/S8AsOkJoZ4BbZLlAvft2qmWqOGIxxJKgnOxMubbdY6GSJ
nMZxzQlpsRmEMOh9EsCAZbq3MX+nvxIbRO2fzENb0w783Aw4MjpDeXOV3eoWATxe
b2IH/Wt8GIH6po0ugjI7Y6kCbP7/EcuKsZHVGfPS4ZodnLhVgz/X8TBcMrEAFEIt
KSqNAu1UkBK7cwP3q8VAkdavdsKMaGZ5Tdzf9JaxE8qvPA23moe/a0fXzbfCrjU6
Vs2tesAhk7JQWyKQBCBFdpm1rUzavPFldPuPqW+7yeuiOJVctrPi058QwR1/GRNw
hU9fkcgJMGtCaxTRPlWq/LxSqpIYOrknxIybJmqrgeyQl4ZhyWOw2W+rSrdxDMfa
SxZaAFhPDZZYQn+nJyeHo9JcZaoT4avXV16L1X/KYkqBtq2A2E4MYN6UpSQ2/KHL
Hne3a0V/wOLenI9mYjNipvCYQrkoFI9ecbEjx8hBTfUlrirgsD9I9ishlCxF3gFJ
0bgufHL6V3JYTMprEKLSmY8DhGvcvffXgtk3QLblGooxPr6jNMFtcEHogzU+BDKY
NPq9AbPokul3JX1zXyFMeKwdyw4VOwQAR21Hnfyv09/4FF74ddlugsSe3F8zOHJM
NudQzChU8N8AXQKzByozDMs59Xly3biPM6MHV2paZfkqCstIb8B8AiS/qUR/DToh
hqVUOT2gIwD228UxLWbI0Ds0TAVVLk+onthr7ztPClx17VdluGY1ks0HeOP7Tzn1
bE2CewJK+96SMygAZhQk0L/X84XOj1RrTZprwYmKczDZ8+DBGopjuzQctfk6yzlP
Gk0+NH9F3E2Ke5iwfFB7BlelQjOjnrTT2/xSoU8sT7UmgqcKjRiXClrMmIH9H6Fh
bY92tU2ohFCu2KRgu2S49ArP2dkS/OSC7pSG9IhWqgUusiE1WdJ+yrLl+mfLx5YL
4HgcD2lRBK4ttOCrkDedpvk5BVXG4UvuGf5s/vfP0bj1gUTuIZZT1PP8zLPj2ZXK
FDAsbOh2tt4PRqs3kxQus2DyFQQMFgCyj/N8Q5ndt/fwBB9PjZKeToSHFIdw/7gT
0cXb32U6qmL8+Thrg1E+tx83WYuHsq6HRbj420aUN8zwQFhrHsELJ0bg25mhfDM+
9KiO62XLdR3bqlx/3Y75D3H4onCFAtU1Z53hlubMkap2PxtfP6n+Zlpf7aShVs1h
bP8RT9c9sUGJqnD2kecoZ4CcdJ+RN5CmTvh0W6laAXRA670j7INcwTqfQZO3+JX5
qS0C6SMQc5ZrcSDRGc7b0rY2LRbYpNiiuiKZ6DJ6bVeOBH6srmpK+2jRB2Uc2ZlW
L/VJANJth+Y/nTRT3ymQbMN1/OEWFGwB+HrC45jtiQL3+DE6a1KHUcKp0aHmoyI3
+7nuiT5X1Mqc4eH/FzpAP6l5WnWpZzHs8IzkDh10bBBuhKmqloK8JfulVtD2+KBi
AF6+YaE/SXRRe8IoV744PLtxczjNSRDvjPVe97RXYsWFZJR75Qd7tbT7fN2kLhbQ
vY6hwWHG1Bc2JuoWnEM3ZRvSKBuKU1VCHb1cogw/H/G+3AKp04WYgKzwFQMkHoxC
Xl9Enp7oPKYw4sVEok4urt9k55RVI0A0FqD28Mw+JBrUD7kYDPs+QmrdBWm3GDa8
VDkZvQvMVz9lu4kB1RJmfGoA/7iLQbmWZtMR9GY8pF+3uFGoQKe8oG/JQ1K6K/Nk
MG3Agfgd18v8BmVu2yJG0pNDcyIE93rANbcGZt4GpsQnrjBH72N/L748s92w07g+
H23piEmlDHBoTxknQTMCJPEQIOZHG3ep3idrve5cFx7dmNcRatlNSvOSTMtJkINw
0kViDxkKKFU3i6lv9w9zLk6z+23bh+x+lyyzcxDfRkFeXVk3gNtyIDqzbp6AsDS2
7NKybkU+bgVCrXeYpADqmalx+tvxZF+eQbDI6HOkc+CbXIAawyM/DEMklBbfWw7A
JlQs/+K4mmf3Chc94hzTLHYZwhRVw1spY3QrOdbKPQIIaXewF+vDN6wj+rWBM66m
yBSAWqmvq8QIRnQJ/+Xxx/EV4gwv2rHRklunvXGJdXBkO82XGXGEp5qhUCoD2JiX
02d28XZ9I7dOULY+vejcnBYGuadC4f1S4PNJ2gr2586dhqawOjJRBcPw54BjO4mr
jVwuH0sSrsHUFdrvkIKOHJw8RLcOgBILTg99hy4iMB7ERsZ1kSIJJO8eTGIR3wGi
aj4Rnt8EEai3ieXCPmVG7TNm0jhVlO+0k7TgVAPlhGaQsHM5lTBGHSAopAqJ+Eg4
0pY3ZfxBvS96B9lCtaYcCI0AE4ZWEA1Zz1rkL8fQCoRH1vxtonDXfybjSMWYygkn
ipv3Ga9XfX+rVu+mrOh2zw/rlQadqPpwHNuTjcp1NnxTpYldOWz8Opxx03yP1pfd
sjCqoaAUiXshWLkuqrWF40YD3mb4LJrX79iSkV3ocJJB+DPa2fNEmgrDAbLwIhjH
5wb0Hf0B8fCjT8JeftJb6mLeonKkdbOZwFD3zUHu8uZICTmisQBFdkCov7Pjk3vi
5RjFCIe6ixEgdp96yQ/bTCW0cvajQob+l/pJ2bg0ZHkccw+ybLS0bA0lC+IeQfKF
aywHLWwkpDQsLMhcoBb6djZ2IAWSEBrIQoRI5r8pHZOLi8U4qHMMiYnuTDQz1NXn
i0GVdl4rrLz7jG7ISf9HWmdt1vDSWSYy74cFm8SuUer2On58eT924kxzOpLd/J9a
XxUu832rSC0pRjfakvAYvhFyoXAjhOqkJOvLw2w6yRzRUrf7FawkZzyLbGshmtWR
H+nlPpZO+rvu0WA/WoGQ3tENwxJGH5iJL5BPQDC6FLCzhf63b+ZEBflz5IgVEDFY
932MFEqjPcDA2pjd5ciR53Y7jZg0qvH1HEnbkpXdqvMt+mqTXoeT1FOgqJ3eJs0+
gDg6ygggFE/sHmRIlDcWRrqiw2UWz/eMFK9xa5g8Ilhu8pYZV43DkOQOzOHznckk
4VH73kYEhEWcHjwqh46Lh6qo5KHrHtCpsqQ3tgNJY3Z9ZUwcUbBSSberSojWnNoE
ZHLRfAJ+c3dMzlinGIzjj5J/JVSsaD4RyIZlSBeS7TsLIkaiZGggrlFlp1IXD+Nb
XMolw9VVOBbJDDMuuqEO2MOHPNtoStTqCeDFdAYrjMgwBWxbBE52xKH5PBakY81M
tbYHyf+H511z4CTBEbFAWdj7GZLpqaxgQ7VD7MvTVEXysor+TN/dFZAkzNUFYk3y
wbeU1DBAsSa5Tzgxzep+uU/XN7OlSRAH6XVbadHWY6Oa9Bd+y3e678SOtpsqY4cx
eMBj/ON3K+d7XHcFelzOR5yDGA0AcS+fxEgcXMFDF9AHFqLMM3DES9iKPSsK5Zxe
RpchUvm3lsMCcRRB7H77J3jME+I2D1C189ARUQQLgBOkx+bTdhU0ykoCRfZMKOur
SjqYD5D2+4mrGLLinGhH9WJNzaEkZCaxWX8yHdJ28dh9oVrr6KQA8fkw0Rhv2kdW
pc3FVBkpeTzA54RFvip32atMfULzC1KR7ZV0o2bGwrT2ZgJ6gq772aXjQEC32lam
WcN7Xou+Ow4jI1DPEMtAqnpxkJygjIPEiG0zeE26//Q2RYwqQyLCjgrjcG2pDGtt
tvpww/4IQHDxcS9c5HzF0qnU+/xBHnFmDKG4ydZUqzhvmOjBEdoq1zu0ypYuZRkx
3Escekxq+bElgmeE16F1WEm1+TROJY6KxqnBhSicdXZC54epjiPbp2TN9SV+A6X4
1L7hpivO8Cr4HMS1CNZ+ESyVRy4KigZ2NwDxbZmEZhJ6QNGNFKadCRKDKe51tVKu
J58LFImqO+bq43YQNIFT2et7r6vnd1WPyni607QVGwZMfxjgQf4Q2pgvrqWdF5V8
IdlFwkMSU/OGl7OKX03xFztJhiLjrdHG5wmHUe/o+YpTp31Cf65+pv1AP/PDQDpG
H/AW2cT9RUx1t7Q5MUQ53UDt/x2xhPMNFCmoE3KExgSlImx2ppMDEdBwpfYljp4T
3tj5KMAQ44Qrpp445kgkYm/7TetexidjDBFbKI5BVP1HMhXdCTLJdbbCeQJfrU64
2dU0+87vB+iCXLqF6coZPpDigngTi/wh7yEwdLJwiJbzhBbclltRa58d+YKNyvnH
6N1/FaKaAL77yEUTu6/epZCzvYUj1b0nEWy7QX/hFp/S5O1jEtlZM4XRXaAWHtM0
woGZAGI+CfC92OlPFHx9Md13cE5/EGNzkvuqsq6mET3U5F+EEz2Y5tGfg8ZBqSN5
/8eaSLaYcBv4+L2SLpA2VUlmtE585o391m2N6p5aPbSoPn06zCcm+d0palvUR5BU
j2NJyxHnROnfsmlzag0+/pYhpqfhJlGWwegTE4OgJc/e2fR3aGipuyYoLm+7PsYm
Te/pKhR6rWFXHvl0KXVuzLmynyfCvARF9AaUuvcDhJqLYCAUKet1sh7JmLm9sa5k
aTgHnROjlYITEUQYdcteGdchqcTV6bcY5ReBxtW7SwDhc5Eb6rwCiDpRM3AugEyu
cjoo/CBLj0FObwuQofN85QkArkItUWYbbYjeEHxQij6ZLq59iaAfa4pewhdsziHm
fAJH3U4mTZB4QwNXHu5ARkBZV6JgcUIRmq4GKVB9qJegp8eB0i6HOxfiycXYrNFJ
C5MN1p9KUJDP8AEdbtBewHug7k81kkONlj/0g5nJvnRSETIgbsW5wisF0IepLxyI
+7DOhqm+DwiepBhzeZ7PexoZUyWu2i5kGcJuKdwsb790iawyIl0/HNe9NDE+U6Mf
ZM8hE7qPMWzYFr0obWm2W5RXnYgATkDBQQEh4g60KvAW/3diC4QaBV+UABXXduLP
uW9T+fe9PToQZdr4qFRwSzJ9bfTo6UD+TJb6XISFtaFNjCIXwiaAxzn2JEzzVoEM
bwdYVfzvYCpcWidd7cH9lwxyY9V2t/nqgYSf7O1KQWTuD+r88rKqbsv3XD89JDtJ
lnJMqOqIShXF8IbEsLt7Fsb5EeAUFFjdad87vF8gVUj7YW3mTCLjgNJ+6OTAcMaJ
g5PHGQMhOxf1pMyf+x2wb4UJP4cH5nIwu3ivwkYTU0AZLixxbuz/sgDZhkrP9KNy
fqe7qS4TKdRifatcLzMC4W1Gl9cyv2fIdMCk5JzCVIKIa296znZOj4/r2/679Ihe
l9uQgC9SPLQYjXv7BN2EpOAq6zjmQDRMnzLKymAAjkWdK2z9XWEZprVL7aeXdyGZ
LY/0qN+hjfe1CONXlkkCZFIXVB23F8WHP/KpMHFiARoZMoc1rLzBwawAR9hoj3sH
jCCEuAewxYOe+mnA7eXrIuibc0ohI6W72y4bDxWHcyzoLwuS+nEdFdds5H7iuDN5
s96xSRIBFXpJaD9KfQowQ2crF27Y6+XjLzOr6aGmO2z/CsZduJG554xLAL8jJpzS
2KBSgm0T6vpI+BAja8/5kf4S/hucmuhiNiIEZLdYwlj2dNM/pKmAMIur0u9te0Ru
rjadVm/NgEYlBiQ8NWXCmqz+0u12t5rss11zysQEgHcSkBDg6mPM2y616+/wwIlZ
UEGRGG2LndxiqvMMRSHA+uyeqj4F7osVw3cSDlq3zRV3h1iTT84CZ7B9jn4em/aE
SJgFoHD5ozF5fXtEPO+ohokpxwlwwen1KXNZiqN5nmhXRfxOnWo4ikXWAnH0q+MG
Dh8EQ8kGPo3Xlaw1Mr7GYl4D24QxhMpPAjmETBraUlFm/lZOaJh3UEeEPHb3zsNZ
9FhtVznV1qD1l5aj2NrnSO89U/32CtkL9DHtB2AlKyjupaX+eehmBGO3VvcCa1Tm
Xny4I5jtJe10kh2AuVcs0KhQvCMrqfmqoJqlEFyqSXq3KNwICnP7aBgqr3GYO0XC
dGCnjrLPnsZnwb+a7a7TRpU7fETA2WOlHzDT1+otl/jDH2oZNHGaDfyaJId5sv0r
AleSoEpYZn/ivMK0MCqk76rJ/KqI083byHMgTzyAOpKO9gxzmVyZqx+inXanld8c
SZ1Y7z2gJRYhCf6yx6PMvlZkpZLzgN+RmZFqKazbeP9FlgZ5BFmXKRHVHfTWtJGZ
0ZuOcKkeKGIDys+5uA/3UzdN2AQKeWPVGDe+1BSYNUlqW+ZhitYB6gYRGlCmetR4
GhCgCml+3Bw4drrclA5MXaxKvMzl1CjiZVqK0JvA+4BwnynFo8VMnrJ2hTFbSRJT
h/6XFdBA5FsOKFfumLW/Hts9XCnkuzDbzfD6Cv3OKt2y10xXwd98aTz2jzu0XS/+
UyM2zzKbWTKpYSYFE49rN/piTNxOBLWI/UO2ws0tOX5J33CI++6Rl9hzgOdowVd6
8zk2IljpOtCq/1AWV6qIWbo5u7nK7270jp5QI//w9vyQWvcX9BftZ2mIp8MeaHn9
8I6X4y7PUeOnXQqQz4vNEnHkYP+ihINRAJAYnWMTd9BbyII6WyOIQ4Bbs1aBRt+K
c8ji3rpQWH88zud7awGiDsU282Xnw3UmihoprMRDhyPuoSXLsdFa32Ok+F78Qdqf
RZNMwJ/UNdWFp1EcSkhjgfytqa555OC15RriOO/do/vt+auN94/+WJSXnITyAY6N
A4sAzM2zUhPhspBxKnuepVGfcRF3h1FNIHv2EtIoBGepKfihe+e8Or9amyZ2+isY
kDWirbgJWSV7zVZceYsz6xRemA6VpzBHhaukSKeAFHxQbmwSyyk9euVUWKF7AciT
HPkPeGTqKfPj118ctg7S5Uxhlfe+o+uoS2Jzy2lIPbkskJB3Ufy5SZ1w5dxlfAp+
H8wJBYO+LYKBVRZ0tDpuQlwkZB4J5z9UA+QyXMFUd5ePUsFmYvaSxT83TTdhFZfD
ucuDhcm52G3mw1K/zgqPUPDLV6fhk9OmHfgKs/mmRxg3PNPcIlK5D138FXdyA1jI
myCzaaohGqkqUtRViGFf2rvtmcySGw64kcIQMLJ7VnU9vaNLEAnoLO8vJlX7cCbu
ZDrwTa3wlsA2rQGuM9L1Y9q7k50qdZO56tQAwKz1Sdk+fj/1XZGAsXIeWrbV/jMk
Wy5Fjj8J8JOyXrAVLT5TbvlUNuKE7XutH/5ztSh9buBcEM4IZgB/WAetOHAZmntt
BCpUcD4J/NdRbDQBsMFboaiFs3txx/uvip0WsngLtQuoc278SAX7riVhrZcMi/iu
yiuuwPRL9irCdYmB1ZhunevrdsMfhwgirAreZedxws2/iUsC9Me/+VIKYgjW7pVP
LiuYFuQkV+4MBQvaiCBeJaHsZVB650NUx65v8jtCWuTtWcD+2OyTkF5IvumOrhLH
zWQjgTqlubvRW/pZ6PD3X5uF6GarCiY5oNj41Zo9Vm4VFSzAtZUp7CGZpTmVOIyc
qvOyQrQXW87WUCqY5m6BQhqXGs+tABcubeBdB0txj/F5OC6K4/zADz5tHmwtgWQR
YT8fLnCr7y1d0eEQyQdiAzikLHS+/Ek/aDztd9A97dI914J99qCmOSN+YgZRtD5Q
8wuxT3I0hKWNCNgGRzKaK8RTW8CHPPyjW1IPNVNUeYO5JJj/oVxuJZ95bcq6cWQ2
xr3oW3vJwS2/p29GK6dtWVtPXyta1U2BZ6GhmtJyXS9ALlmwu9URMAESm1QX3SDi
6zXMX2nAZCw2I7KtW+Ubks2OzLokevAaQJAsRjvy7dEbUlH6mpYqxGTovNNrMo5T
TozJtv6x3wH3v1Duu6MIHghMhTHxiST5iy0SmEm76Go3wyWkD5IhTWt2pvhXQPql
FZA97e2uTnnpd65cf0MjBeVvWfrAr0/WIbjUFps0+RUdSlMLjJItW3OtiyXuTDIE
kVwIqwWHHO1HvLeao35KSKedq/kR1GaqAMUd0lKVI0KF3UsmZ3JggKtXsf+kuGhH
90pOguOEYEWiS01Y/17mBPwctxUm1ggXp1ewBnPUZg7r2UzIP49OArilv2iSvWTs
dj53h/0Ite+2k7hBB25bWJD0QKIt4cUeGkl68rpjjEKzN0zK8ClxBD5Y2+LpJU6v
BBI12BoE9GTg9Vorix5B3/csO2NLOuJ6aJaNqB0hP6mQB5J4lGXtFuC3Iqdpfpnj
waAt0XTdGa8xYl4ElLGWS/JQezaJ6XNKhyPxDB2kLkBTHwjxtYAUCiS3/QslJyV3
BoVIzfMAMNkIQFRKW7pMUpYIi8xoT6ptm7aSDJIk3APW/f09fWznQiyGgXuMNLRI
DhiGc/DfoReyP1wu4gIRtm1CnMZ75cvnJXH0Qbr2Tx1kCHES+bcn2m4ifVGS6E2U
+CM4M1rnbkxgIUd1gv64dR9zMwVqyzHiXT3u3XVYKmB783rjyZ5chC/5wOnHzd4J
Ac+r0/QLCHkppwW3gUh/IvaUFXy2MZowiNYQpLNiB/vWzlabMnVycpIZ2a3ufgRp
EFghEGa1wNKFDaPA9ncFJTx+lfq8xJuXlq7iqImvUBW8dfC2ktCOH9JpJwsq7m9/
nt6sQw4OuJFH6XBU+j3tnCqFKx2jNZ28s12hri0JJf6f/VqacnQFCow+A9p/rxxR
lhhjixTiDRbqTl2JRM5AxyUp72qcjOBG1F29pKWyWVGu+dP9rlQZdfZO7xDlV5y7
H9nAzYyvI7eSm1e3S3xybxTH7jmGzw1VB/UxgNTTbahenykS0fQOeq1t7VUoxt1v
ZicgnLADGzC2SzVB/3hpoN560xoZKsVynKFr3B4ecz78v5B9+nThK4hfx8djvGQB
nwSJetVAnyyEW13BpZ8xexYER9Azd4ASE4mugVI4PB0RzwM/jepwjaKDlDA3nEMZ
wuqWgHhs71xkwrnuCzBGtRndM/RsTQOnKq/WlN7QksEnxgrwW9+U5PwP2hCoddD9
BGgC/y/0Z5XNQM83ASmNsWAVDDJnEv6NPHsCdiC8APtx4U1JV9lBMTH35tmppL4p
DDLVqFGT4XyVpDNHw0XRtRiBKdrotbF6Ed/fI+GAaGmF4LIHooIb/aUVht6T4ydS
sS0j6wttkrTngbazg24AgvYIlmWbyuuu4tPnBgGUldH/Y+RFzNyykQOFhwnYacoL
j5ZTYu2TlTO4mb6Q26vtAXvfgASKIj2nZBfRMT0GWAJuuR0CkSalIfMrYKkRGW04
+R/LMj028i5jAbQLzIIffU4RmSYk2IticL8SPzRh2jl6f3mkdvCfB6lChgBkc7BV
BZNAttrLWnNx0JX7k+1D9ChCC9brLwrBhxrcjbmOj//0mvshGiSwFrAMpS7o/DTq
yGkej06n3N6DoA+9Ewj6AHhi1t9cgI4znnGMtwUboQC8FaJT79AhXYS/S5On0LUl
7P8pmQJH/nJ54d4sGwrybHAwoP80Pg8AGGVBluEtwAO67TjOI44xRjgghUG2WV91
QSy+rX07FyG/tAUC25mT/r4k4L0M+e8N0VOuJqdwgqqXn2AAU9eCbsj40a0Qrznm
kmBV+3XXSS7lmE11A8iV0HTnHBdV2IKkyra9xtNEspcaFA5kYkGlCUTpraik3fQI
uSicoKWfV4+nxPAQ4JzZtLljcrEeBPykvlf2kYp/xmDbKF0Zo7xmyBnMXNvpaREY
UBi2OK/+YBxZG57Fpcl6j3nTB7QChz69z86o8ixlYbfAk8a2L3vpdZdLwe6XKLU6
yiQtFal6RfVuBxYb5HXbNhb7fNNtwfjOa9WZzbuMtNURSCR1LxqqaNSkDEtDBFxP
Ghd4S1VLGvDYOgbQPrYQ2qR7RLCxBaeKOcp/7SoILvnKpkToLoHB7IqUaAADIxRT
/qNLyDOplXxOCPToig2X9VdhrcCkMb7ZLOuzs9TUsh/mnMpetpMoAfvU+hCkBinl
imgca+ZiysjNRBXQyH2RkJvVS6WwSmrVMTUs1NoSsYI9quO/V0hqeIJiGbYegec7
jaeMQdk5QmgV8xv/MYD4lh8y4Ls4VRsehnCrYWcfbVPyn6NPAZLDZpk0VT+2VGC7
n5HonC+BNxWTpKITRCTkxaW36prCd5c+yYdnklkKLxUCy4bcZ8huG6A/2iICutl9
CkDXo24JDW29buaX6TVfBJTHv+JOuJLQUcrxsBC82gXCbqlbAP+FYOlKrtMmvPXn
933/Rb49+qOAxAfjAQsPYVUtxvkktelW9RT2psEhtqEmOB2pBWm/WdKpaXnDOy0m
AcrfcR/e9RLuIQ8Qsky1RLiCMLMahtsYw4NGEbiGvAj1Vzt2k60GLB49VfmST8zP
bk+LfhuKKJZE/C3X3Ax3qeLlDX76fh3GCho5oZCN2leL+lPgN8mi45TCovaS1z3h
tS1gU4myNy477fvCjfsyVbO2i+Cq9YoiDj0v7QxnXYlC8AFG645gCJEemfa6kVnK
4un/VbvpfqT2Sz20M5g5Cdo7ew8Q09riUPrFzuxgeGUHo/BW7bp9WeYJyT9omN4j
UI6ox8uIFy6r5c6gJ5vxNjQieAzUoviueYtUwtK04+zkvTPHgZWFUctotHEnghMh
6t6GCiFu7qu+XKUyZQ844RN+BqbvuHi59Wmye28ljHpEOMctYmiovDJUPoi7J97M
25RxYjQKNedvR6TjywpxETvml/qbsNhf0B6tWbb4NBEUcqSDUPN+TcnUo6QStZtP
IL0FFCrNO3s4MJh+b9W6bY5xrQMMhT8qrRzJMHbnYg0aQeL8REVm5FZCDNOX8mqy
n2d2myu4Xqmiev9VOFcWl6y7Df3CD9IZK78+H8C3a/PP1iSnRF0pUpjzuxo11i4h
DPc01ENF7j1im6DyN766ywJAkJ2va+ylyF9zBjlK9fYpPz83pTp/RK4SWtxnJo/l
A33vtkCnKD34FoGzxVicY/TznwXj6hn8pQvJZ6PXiOQUG/jaj3YthkgUIoh25MEl
X2tE1morrcxU5BgMidDKu3St04YVk1jgwzRC6IedgvLIYJwl5PlgVA65niYK0JvW
NWsYkC3Dc9zaQxbQn5+Ww8DZDPC2pMgIgJErIm3mAFxT9jB94VfVLtzfIU6y5nf5
3VOUobktyJezIUUqtN6oZPuj8vLf2Hgp9B2PsXZva2uzsZvxAL00FF0qftrMuTyo
tUnHHZ20z+TB02tihL+MOQrmJDVRlK+maBfpkWT57LK3MQjNJpxx/pbDFVfShRU3
koPTMutYCQjlvErfv7BlYVfUP/qJAT9nIFkLPoQ516SmaqxDwos1Tnu7J3z4nGhR
J07CxHPOQU2Ip8bzkApmHmhfvi6otV4zbQvCVN1J8yqkf9oLf2mVzL7WkSjv57f+
CDYLM6tla+aySjjklhpVspg6TVofaj7UwPnHRIaJNJtt0+Nj28etvTuaj9F0j9Rn
GbI6VLeQgM1vhOwDcZ1lGCcSNB5N4wsmTh37Pkj9KDv2B4GBFl2NP3Z+w2StVJKz
vEn0M/Vs0KxF14mKz5UZC7C2Yev8p14BMt5Z+UdB4xXJvbnv/BETvLOp0H+XnVol
l1bDU+gkGV49EdYVYzWYuY1ZJlmMErzT7Buzj/uZn2+xiOjSMyyx4vb+vZnA29M4
HSaSOVJ7CAs0vAkyp85h3SUSaJqcfbbQTZOO39fHs6miHByGodGKhtActSXuJqGz
ija/FYLmPQPtpkUYnAFXKcz7iRvzqBr2YKucEgXJ+noAWD7NK5bX6x064lFHUgdD
WS6JyiGepUzhb6AZvZ3mru05WU7e507R76ApDx+5esEyk5m5c3pEyW3o8JtXtmNu
EFLgJXUcZhP+XrqgK3dq23wNjrbwDbJwjFCwiPRouETGAUJk6T2Z9Q63XGU8npZr
SyKKvzcS+3ve7nWnmJrghLSzW3iOXf1M8zGBZHd2rbcHkPFshwexzbqHPU6jhJhy
HlEn4TcWQJTq7BmMUPivWvSuAK6afMEh0AONa7ZEzOaRhKQfnwHBsUcR4AGZatxK
V2WOFVl+rGNHRTXXFfu2zBzdI+LvhauInLIbvZhXViG9vIIwMuMZJCCm0nz51VQU
Ea1hRIkseC/LotPrt1UkKTh9px9YACG7i7JJvdfEGuUsLrJ9vEFvT/cHb2F/d4DJ
k/CWe8e17C8Tta44ajlGNdAJM7E1ukuVSJCCDx8FvjGH6HAqPU54DVrSAzNTRfyv
i2JXiofVUAoi9lmxvftyw5XT2kmHc7UCv0ax+TGAlzK+o/AP0xOGuUtkyHJ2VUSf
UhbFQbVgRRAYwEcREwLLoGH/9brT4EbzMQyfdXuBvYFBk0yFwLveExJARHhS4HRJ
nXGkyZWPWPrFTYbqRdKud96H2Mfv/PJ9H3A03uPthvbeVMuNYMCvqTISpO4h1HEX
rg32vQH+Tq+aVpvSVoHjZhMoyL0CV7E2UPFwFFC4OSjVNJLw3JOffGYXcekgQWEj
+5Bte003ndy2H6o+/t3/Jh2aPuzBJEYvwSBr3CPooPsZt6SpT+j812YmQFxRZ/NZ
69mr5Op75zPYWnHAdo0RiWVSPOTapfKdHhfvSedEy+NedDFfaVzRsurImpEwMvhu
1s5tCM9gV6N+xXH37Bez1eqYwGiarNHK5gdTT7EDCYRwGH7T+0fzMTSb+3EltNEm
irh6BkE0mSAvFb1HEegGKM5crK0uhKTH+cwpk7IZTZng6BqcDp3xRGL8uFRelyNE
Au/8SEtXV0ul3IdG9Yf5Kyxa+PUyEBViovmjGXKwW1CTcqD/wAJJQWJ01kt30rpf
I9i0voeuXJG4i3PTIyHhL+WIuSGee/OBroz7BJ6lacNAMA6yLXzDkAmdSHKmMO22
3EKNt3pALv6OOe8xRto+HXd9b+e3CwnUtDo9Bj38cCUA+K2H8IRKqKkxBK8gVFHs
ncUF5JEfsEDB8qQL+kpOi0jx9gcTidt+fEOxD8t5UJx6Bd4+LbXhBX/IVgEK+L1C
bW3XKKsKGY0KgiV2Gn5/uU07IxhDypMy3F7iboxyZzSf7Xs8Ke3eN2/mvdLAGA/N
ydXn0PQ/PQZ8AQ6voAaa/1gO+3ZuRELikr82SdkB2nI6NZ2VLVYnUMHMDRriPhP7
cEyWtheW9tInBRSq2SWLi1s20O9PLIIm91pnb9QKzpH7hCdXWmb+I9ucjYL1MiAp
fiYZAo96Z8ub9WLSHUtRwPs0myNRZO4ePWvjBXxVPouOJStHLDwzaxfN6/wnwlmH
EkFUMsQ73mVhtf8hhfGSevrL3S0/UumP2ngB1/F/x0IfSHRYkvkBWVzscDqK7zyW
pGB6Epuj5qJJgPPt5eVgxEH42TafMd7qcojePI060ifTrEsPBiPiD8fJYNRG7eR0
GPB504f7LsYHgpM1H4M2QQuy1h8a4di11KyLYaQIQ2k8ckvVCvKnm/v1rGYi15kD
zWyAYPxFRRImnOW5YqorzF0tcMrcS90QxBmAj2n8hLr6NCwwkbV9JmgnKB+KKswu
xOWcwVMUThe31P6VI0jt+99RN74EMMrN9KfD8KFW6mw1mBvnOIHAORJBgom9DOIF
T7ItL7camt7Qf/qSobM47jXzGqM5Q2r+geb9ZXyTWF/VhLNfA9ilE3l5CkUFl/EC
cGBpt563X7vfx3s3GEQjehXeyrO4IIvGbMwdraVScGTjr+N2HkKYj1AAnFGSFohu
L+y2TcQx4rW+albbUljn8OVx1P9jL5lRLE3/0ZlgF5tvy/bePStNQyDOdC1mejoj
uA8DtM53m2n0MqbBujJHGFdxWsb7SEWyn9vHGMEt211+PFG0dA7C+9m+Ea+zcQPb
sGWHivNDPDwWV5AhVYKR+HMtGh1twLqbs0ECeYN+4iYBzssym86LLrJKXAnVH5ng
tJawXh91NOrlkyWv2e2FPtsnW0x3f9XaGhMxWnHtMYYl8RnLJJjxINXjiZS4/uUp
RNkhM+VuZpcLYv4AxkBgx6hIgHmSbFNCFmYcHZIbvrHst5kmi4ObWBj9UK0aPedS
MU+g3qvi3zCgmhoZ5uOO/uDW5QTrvbZ0kTwHIXQfN2bzGAC8TS/46tPKpN/L0DJ7
cBgePMAtC83wFaoHKT100wXWGg19qSUrYnHX/MnRvZtX3CG8k5zmt+6Zto8sYE+5
R7hucNuVjCVx9Ev3dUijwv9v2ePYOSMbNo6MByDn6baUa1QQ4wS7643kFB/ZOp5o
FSEPKKneiTPnLLkYpPcdMSz1D9uuBjurQoPw23DjwnHu7AIW0yh+trvGYEOzcCtz
jVB+qhJS9e+fSMiVEbUTuIxYYHUKoTcU0sCPrvpuDGhr8FFyHfgdHLEo7H9Ukhto
4Ihpn1DtaIo45k50d9dcKOpGkFPelzEkTqEJgqLFo7CzXcNh/Vq9GpxeAvkyRWwB
7MfDTPY8s5XldeBNe+xdgY3iygXMZlkiJnpvcQQb3KjnvxAnci8gLVyRRxYBcn0b
PWHQEVR3QRArrXQdGA6JDs5UqXq+h1mk10iKd1DQLn98Z1ogeK8z6fc1kPfTIXPt
q8vD5uAK7Asr18xj7Yj/DObhC8rJV75m/+WBFOL+6xxoijxXXSSz/1QkxS308ghv
YJpoydoOVt9Qw6TMMWlx4PqDq23PkNFEZlwxCA/YkHt2kte7nUOiT/cXouTwdcVZ
3nRla51fegagPzaejWiJm8mElTPKdm+JqyBmFj5yymgnF/WrZNXlCisSlmhb1ttH
RmYNpnj8+e3h3tYvZNhp99o46WiTWy18hUeXnF4o57w96dS/tw9o1CcHQ3h4SfAK
ZIAIOU5GhIsDw2Z4xiLd7yCLbkqDY0paPQJHF8rqMkgiBC3EcbxvrrWvXUEKeS4o
jFE3b0vguIKBaHA1grrwus1s77nCzqHZbrrlD9eQj5UMKZbfNa9SOhb1vHePxjYb
HznsFdBmXyU1FpzwAGzF3XLRAeUMV3QUBBZF6TAIZXXJNAIbVfrHMwi2IMBazVOz
C6UpMGaRUdK+ZBLRbtwH/gOLsU7DvW4Fy/tPH63mmvh7cax+gQhQtruzbgWzAU2O
0bIkllCv1Z8etkhXeSLfS2a2Nxeg3aKfIecdYu3h2kAxaeLjliNrZx7mnPiMHrcE
Zt+dxhvSOMZPoJ3nsvB/udFbY7b6rOC9UFEjfE/6tnXowcAuXhWSU1EOhff0gPqj
BdK2nFo7JjL7JLCqF22rS6sZHNwsjwhqqM+5G0TPvJBfd3Z9Es7V89+Rypr+oML2
vknUZVqh4fZa2YyBzxf7kHQxjjPfG42yHv8gyALUjEXewNDEsvrK31Fv8nghnvHq
UaQbPlaRawKuktmq55Gu/+39QBaSaADiJiccH0e3KUztw1ChsMAGUEXkFWbkHV9H
SuzSG8M5EmM5xicmiCJqgepqnFH/QXi2z5K7z24NUl6kyagJ/GxZa2cIa8gt+1Je
bBB2hbNf+vfFnMGqSssyXWwT+4nCiPasbU/Jl+1wCe12aIAvJtVzumdqOrQ+Hzcq
ty1KXeeFO8qDmUeMOW28ZHLIviMSiORSMq32jC5AP2/CHnkP5AP+hf/6APS+vStm
QW3BPnlPkWX1jyUWETEE2vOnxsMkI9XUO1Qzk9/pHfMFyCqeQctzOmcxShLSS4QI
g7JqhLKUY0I9zTcBlltUD+hDkrTQxGhvM3+2cqmBfElLMywqeXDI+vj5iXstMtBJ
9HnnoPOZhlh4SwA8xqaO5vDX5f2yh/4wFr187RaVL09Ub/4RjhG1+ydGRTzp716M
6DatRwj8IwZwWxJCSbQflhr+6KOvHtV7AfigsRuZVpO5ccCe8sm0T2hVkFI1NTL3
kd2ANE0xWv26L06O2WeAgfI1s5hsz9k/unkpYvj1cy/6clCSDxEhqIvnayuEk9lW
NC1v2sk9L8pR/MmSGbyo1qs3rOZ2l3+PE/6bImnNh+/LSUEMRMDmGtQVWYQ5Kjs7
I4LSEFaWgzcjCvdNkQ5kjaAGEgGY5ykmEGGV72jtpeifiWGr7Gyr/TLymMdK6B54
pDmkMDKo59aWFYkEcXKfhwbbJqvxIVq/z4O3+Z2iIF0E/p+YNEfsFvSb0zjpsJjL
T2lY5tNk5sY7EB2eCDnbXFCKgu74s7wPaZP8NtnYNknXB8Qbo1RNfS5Nn/j8t2JX
XCYUKpTs0La4BRSg74FEf8G6naDdGZk73wNdkhWj+1VKy6yWqAOz1RuDMrJdnSsy
fsPmoXBMLqdJaUTGryErrtUCXqTIz5AI8azvs7ye8n0DkoHP1ZXE08J57hcooZxy
PzqG1eavXZvnGBwHrG1LqT24tvkbRHnTnSx1ydp8Z/aiShkpRJtOwi35xYjXORo1
ivUCV6IHUVziNV0Jfx08k1uAUJrjbnI0s3213OeYPAZdQihM3nvzHVPUTLyomV2P
nZit3LROuuk4t53idLEU8flolgHeICesKA8UiLI2eYb1uyaKTxVXxCoraM/B7mwn
6qmxj0uBugJ3FMBHUrH3mzT6i22D0Mhotfj/Y1Fk57GvyX0x+rEFRL1KXj2jTnCm
QVKNy8pJbg+ML9uRJTybZBBpe1gzaHJaqIGztD5TN+lC51KSfyMwG6xtFFjRdhjx
sMCTuF+LfvgDcFQynz/CfKdbyiiMnGgZnB3dwAXJurWG6r5KRoHzqRf+xkazO7O3
PSkrGIKpHw/MG0gTD64onBWCfY7N/pq4YjqAyhaVjmSlG50fncmpih3xLo1SVqyC
5pl5CCC1iu9rgh1XLrGqeodK6ePwgzuRMEtOinGO5QmIm7cutu07NZcfh06vZNL+
5Ap5dUdbu5M4FO7JcTiBJwqQvByBqpWmrQvB8g3y+3IJS+4D48U0/3+7duJbXJRF
uXfIRTVJQzzawq2kOFVYRw+OZpUa/k+qOMlb00wugjjHhNHNwQpf+pS7/q57Yy9C
SgZKyNK4tD8kjv4tW8c0d2LreEB+ifbsfUu6AlWLmAmEzWTryRlUB4XBpfs5PB7+
4fyJ1/AUD8kMjQ61cf+i+Ijbhqud/6vcuNn7MbRSK/bV5zUxcQG/kD2kx4rV69Sd
GPgj3cL4Q/BCcvCmAzWwbxESwktsLa1shTvqksPGu/cNPCnCaNjDjCR4QHMVquxn
GkepGgg7M5nyn09sNvCEiNU6mKEfsB6sAsO7513ktPBPV4NoYc9l1dda2kzraIMT
MxuTNppGriSwGM/Nz415TVLQ05pmxZd5uuCpofdAPOHwQNafCmJEqdLjTEWsshfB
93EHOlVBXXXvrR68XhJCnULAAnQmN4NKWpNxOXIzb108O+eI4dWsCf+/KtsTj7+m
JeFRyaQOdeMsazNS8k8HQkozdepGhWbsjs5+64qcfAwwzODrJN9uILKj0KXzk2kO
RKXaGK1KKSe4Lb6ddo0lxH0LZUG3Jtea8suz7OGBulwxBx518Vmp5eQVAiAMPSAU
Z3aaDcVWg7rvKSqp/csxBrHgjjoVbIi5f2cCjxYfAr+STlWi21lAuDC9Z1AOIFfm
GSuTqObpGsrs40nNiSOCzUKP1A9xKxrce25lZJHGPQgJj669BDCyd+lSb0UAIAob
/aRdTSJJWMNKWaauoAyn7V/mdUVvIxtd339NEzCpKKl7+ea8i8AzbAjLEadvg54P
mYNECnUPRZ1V/RYe1LpwJSAZR2o9B0BltW0JDqDW5JMt14p+2xSRjzJPw9D3fkK7
JB2dVyUg1YdCsmlejm+mwzVnXSJVwWrcVldQ3sm72TPDnXlbeIVse34x/8j/NzYR
EedzEIjsD7ruPMrhV4xavX6VSlUuEBe0GQSy7IrXJRnQmbcMkwJdE/vi47vJSwKp
SAIFq69xkgUG4G4swm/ZMRamQdG/44cbSgmiyahz9ITgRKlwOyD5iloYNA6i6FKv
ELeMF1uCEXPNv+756SN+/3ggshed2GlucA01tL0gUwCLuH5Y1oafDezvRwLrUkr4
Ccm3IUWlAmx3AaDTcPyIamF0pL5R9p8zgJh/W2jJrKZZZ0OhnvtH3dQPiYuZNzJ9
pegD0urL33j9fbIXiDsv8PmGU3QHizj6ULLyYbsQYt+aRkgNhglWxFibL3TBf/EU
b8FV3LVaMVhHrWH9tjgFPpvKkXW7LRBvUzF1dnl/UJV6N4Sh2qfCt+wivWFLDWgd
t6mZSQtFIiLfnh0pDtO9NfXvdbMmQEIoKzJVzFroQaolvS7LeSsXUUp7smqq3OSw
l1/cVB0L7X4TssOWfhhGL7AAt9qlFfsxdXLhVYsYin64lKikwYHa2nI0vX8l0K2E
SoP8eHx1yH4JQJhG5/kt/rqtfZD2py+1yFZkjcNaav8t/Y1oBH7rH+xJKHvArmio
RdQKzruzqyS/6DT9Wkut2Tppu9PKBtFi7upd1aDMakd4M8rP6MbkeZfzqXwvpf14
syOeseDHh+qq8NP+vk6BycDHganYI9jxBLXtYIymfXWAUkqct7K98GjFFiHEEO0i
j6sXdmB00McEI5D5YtSM5/z+nKUmtCGLyP1kW50xTNy6m7jc026OH3xX/xeLmcm3
oG6Jnuwd5B37rhKrx0ppebuQLrHtkjwUEalu1Xt78W6QDcpa0/AAUY1J80FD1HXA
QDGu33AzjHedHPvWUW7t++L85JI2Y0p0gI8ZwYWsU7V0y/VpqGm3GaB0SEMMdWI1
kaez9xquqPu18cDKU12jTB5+4GNZ0dDi6eBtSjw+UucJKZcHNAoT/ifgOlgZ2l0e
ZYguJ+Q11PpEuE95ChvGONuShrvRLN6xvK3FKmgU9ilKdRhrB7clx+GH3sjJkPlF
5xIWGvPNuOWuBv6BKUmg98N1Ke/BFcuh7VHZuWReYWO0do29waanmJc7cvBCZ2RN
hvfI7rIZbDQwVOkmW+W3s2pDMU7MjBe9XCT3hpuBJ0RfjI/15HRt+ZJfZAX9+Ev1
gGIMEyEZkwLOW6gRPYA0EN/wE1k0LMHBE8YemJDJgokPIRYqbEzb2HBQ9qcXJ2nP
3Td/g2Vowoog9iKuWDK61KUzCkYuWicpRsxb1wo+t8mts+l85SV3z179F43Ner4V
A1PKSYqXSDmczg8NzCGUCn4GYitF1oef/msdugpeUfyzG0xsXe06lKCHC3bUURWN
AXMhh6lw0ZKrfA7Cqdpp6D/EiIHfbggarJtwEkzP/+CElva7QXcSE7ygeG0vM9L4
qftr3Bs9PEBN/N49av2077ADuH8bNsG2QpuX55psm6K9qndSr6EzfAzFhlnOvTwU
qp4mREqAke8GSvfO4BcejW7DBi0L4RIXuumaGtDjkM6QaUfdWuE7MkSw0otRWM11
odsXPgUWL6Vx9JQlJz0coxOtfQwJvzrLDkh6gVl/dPLgivOZ9oJGOLmAcg79dwZH
FHy0aFh6tYosL4btPmIMGHhycCxjvoFZmFe11TgZEKuc0kKbdpBNXi3kCkrh8bkF
Nn9jAr7Zpoef0tevM4A6EtEnP0NlvOiVxh+O3nHnwCfjrPs4sE36uP5oMakJ1QHs
bNxsG+QtQ+72ttXXJK1ZklzOXNnEp/cZfi/C5z6xkVEKQ/bOhEm6ouiW6IglKzhO
+MgfkoO0iGQB5NfoJY5XGUyFsOTXbx1FktJSJ+ktwEeOxXhOFt0L5st4J/TWUGpT
8Ut6VhengiJNS33gyv/6xCeheHylFIEABbGe1dPaxjc+BvxAQKWJ60p4RK562VqE
pqAxnKgqIAoI+k+vOBn8JDc0qoOJB9gYscMrOBqggVWniQ+/8tiWimlyfsaKhoW2
zlDI0fC2bp3u/skA9pU+qTIlsm0OsVAD/nqAl2jGW3hbrOGpzGspfkmqQu591bb0
sDia9GP7vVjThj5DhbXLQppGjKmVYb2RVmB2ddU8hz6a5PkIMYaE8malkcr8PGEW
CLrmF9WEQKgo0Bn7x/Z4LZvQ+juwpEHxkZE1V4ksI20X+G/Hf+uTjIJBFtVj0vvB
VrLiLVoAsEbJwBo7qHDYktudAE9Qs+Fk3hEbxJau6avbS1hcQRH7L4PCl5kQ90y1
UdqeGFd8sOSmdY66DQ7vdgluZNXU2XqRB7pLuUuH7BgZQMMjwSBGbNU7JrWNyDTL
9nSsk3GOeDzBLurgTwxZ6m0jWxGPNPVs4VCkxQgkAPv35DvOeFEawGwVtxkMAX6o
JxjRMfQMNw3ghhQB0YuYVyIcuRKnNIjIpAlFOT/huaF8CLIxczb5t8dCR7ucpGTC
8Rjy+sZHdCBKyg/4q+vo3X2vU8Vj7O3BBDEP4VMx5PfLKMqnue0LfttPNK4ritTM
1fx6JkU3DjIOg637zG44waoMoXbH5nT2Crpu0knBl92LC8Nhz+ZUxWaeBJQchtFu
eI9Q+yzItoBlxyJ+m/KitAv+XRgdUPAVNBw6Qe08HQM8F1ke1Lan79lH+LJFzsCq
U1FyHt4HvKe9UM+Tp+uuJa+pLJQeafWKsJ/GUy3iVDb2nGcWujELngOig7hwSBoo
KG3sXBH5lTTzxgnDjTv8hLvVYdhjKGPn9hiA2ujJ6pPfuWwBtlZuRdN9VHOOIo5E
ekz7lHH1VgAHHKwhKVJsvisL8LSXtasrgqUpcduEaEUn6YM0Srh1D2LoJ2BaPiOb
w4YSYVPiV++Lk2kmVm2DhcaxQLCccIPzJ3yw3TlpLeeeJv5Ppv6FUqLbxZqkje49
p4fOATdffpORlZ/IMwTwwOWgm+/mjcxE+08Us8i7KIrxX8gNMRaDmTthg46CtkX6
4mwq8Ylp5u9XB3z4jmbHxBhW5rFTwibKfkUbliCAY8iBT7ZdA5tBCBS6NIl+1+0c
xghdKMhFwRuWRikr4Z5UhvXVUi3AlQo5GTqfzosuZFrrUrudWUhYvB0ziglciwOw
ibtNiAQg6IGvMH6cAOCgLkeZ9Ckshx8w1JpnLnFPk5ILAIC25TCvgJ4ZNlrv1ELG
fYJmuyTjEvdpEiEzQ16+E57dMjW8mAMlNoXWZbLpti/bkrqJnOnEcqpy4ZYJMHLh
9hB6v0svIdZKyzXa9dwpyIVm9ogPih4Xyg7Kv8V4nS/OvcWZBdQCoH0EniB+rHBo
sd9vxYoMyh9Vfa4eKpZyxPJwnDPZblWKBKy3ocBN/XEBEa5EnoAUwBXONO2iW6wb
22agdJyXHqXKSMufBSABH3GCdPn7G1r0lrhCgsywjFbrTVp6YZq8MGGfpR+SfGez
eLwP4wGQ0Ddx5jN1FTFhzWVRa7BW+GPdnQ1tAKd++YPVWlSDFjL+X4gPC3lHJTJM
fFdPFu3SrHdn+hGH4DNRyUgAuVGlr7Dzw7qxAb9PL1Bg4hgGTaceei05Id4Nt1vA
KvDPhrGqGxvR62A6sYpfEMhu+xIO6+XMqW0dc2AyCCxFwHOqlzHtdLQmCLt2hFYM
NxzaLjZ7EEvA8JdEwBFrtO0yHwahIiTxBN+o9LAGJDVkFkBuD/TVbEzob9RWu/AI
OLY7Gjl0NrGkf9/5YwVuug1sj6T4hRQSjRMcpXgDedEFvLeEphg5gw2IdSgC9Gyn
xyCt/DW5hia1wlTDlQhQenAy4Ati3wZJtqtQfz6rZyekZiorxHIMEB3Gbw66Hpz7
bu+cynUONxvPRO5uWHlGxlG6toQPnG1cZ8oX1oKRoOS0+f57ISlUFsxPpydhdiRY
sp3UMZKvBNz07fT1KILiM5WLhkWuSiXyAYuf/zgFC+3xjSOc7ENqhEhfYBq+m+Ew
Zcl/1WF/CGXoDmxK6POvfxFkR6AYVSBYJWOOpE4DUQnpGIhJYYtEssUM4q2dFbVg
FtCVd9VYi1TK7X3SENc1PBu58Vpq/h966NllSaFAF4p+qzcRiWFKgAVc+L9gagsM
AK31ZNYQjSnsbzWD/ekWWInrEPV0R1yPh3MCuVQwsjfFd+WM5FICV6gCcHk6cokQ
wU8umiyZECF/fVgJ1e7Y8CpjYrJG7ogp9vYI7kv4PC4XF8ZVzM6xDezKi+FPkR59
iBmT4OytluqXWZyNLAr9mmF2hmjMJ2yWslRbWCeGbS0Le/oiD0QZvDXcIp4BU3hG
zA8ckycycgpcTP/VvE+qvg9dA9GsAwSOi7sRHYll0XBAPayFnCk5sqko/igwe/ix
TH3urwTX29xX+UN5JI9wfJq3jXwr8xOSVSgDH7wnW1gzacVa05anwFAHHKygGuB8
XfHjKrTjE4VzH5YCHTxt5GxTOrrQZkkBI65aigj0oN+ys66J4rLPGMbxOwQ2Q8c1
OS6+etmE5nUO41iIXzjshzk98sWe+7271K9hZtZsQ1yvLRmiLNH4QPygA9zKu0ZB
l2C01GPmykZEzbc4J/bN9cVmTCpdYYOhFptvd4xHtmBrUBoler/kblCWmELRTTkC
+pLYr63hHIMvf0b/q2iGq1Ebe3KXDRa5GEC683o9+1FmOHbHXfsFr4VKC7ZxrsLZ
0Z87kMmWRy765dHHatyx9iYi1wakdVTWl5afFjKW1yHPX0kQfRqNh/w6pnLj/XZ0
SaCD4HkhI2gb+k0V6yKTF/V/mrsMVxkYOtzXSsVpKHQ2JpnUqssPELrudhclIJls
8GvFDntxhM2GC5X/kq5q4WSsa0ykiVzoxwe5wsFxbN434lQuqAUXuEgPJ9IhcrFh
8LH3yqcy4kO8din7p5mNA78e9z5oS9WM9xllwBwRuVD142y0INiDGRiYTe+J1Z2h
cXoGWiWaICRS1rPjb4DabQr2eFQRiLdBCUQn2JXP/ERGJOp1aAZSFOoIlRXIEloL
G3P9bkz5BU8haOSM97dtXaP8ryFErg27aDX7imNdCcbWH0E5bn2XOz6gqZGmJIhG
BxbYeVEBt1Ho7ssQU0c9jf3J4I1Zaw9Gi8ViREwvAWbvBA1/ylD7vW/hCGDy8m0j
ZJpsxdu7jaYBtVyA0qNKvvrmsfJOMWQnhQ7urZTPOks8fRSxj8nlMaFo3Ji0nMZJ
N8jotBZS3HxOGBr8z0du1wrw4ZgWkJmv1MgItPewG5bFaxgCW1kJbfdxHpbF33Sd
Oz8qaC6iJjPioDgqag9s4+3Dp/NIY0bOYMVru7UGUZFMMOEEnYhrXaAqo/KHLSAA
zEHhMOjSGKT2WBiKG/0LF5KPnvssSsWIwEa5ZIIL3FzBH37jBpvswZAEtFGQzony
OCkIlJC3k1+003tTyZ0240XOVwlHfTca/O6rmw833NUTLz2DMJsead3GnDcaV/BV
DfdPhYK1wXdgypkgNi/eWHYY8p9DQYH7SoECRoZ+77tzrLbEq7ph4UkEmkLo7rj5
ZN9+ODRyYmym3lq7sOjmY4b8PXCYyrFTUhuaTpDgAwsrFYJW6gCZ8IWo8PFP0v+F
1ny2GqBB4mFOlrvhXyFo4xKNadtnNKf25FjUtImVgPBkSM6O1SX4D/fnqtS20fmN
34S53MtlX5ZLe3l2Dt7ZJZcbVHv0m7jRjHyCHevzZ1HP5EB8mmLny+Y0jXyhFpJv
wyMbVWgn3fi6xw632tg/KZBjmKV8AUVdLSWJ19uQ+CVcNgy+6Ew9CZGug0VyMzak
QRFZ7DLfHqR8vezeFZZq/jnGxbrPma0791SJaVM3IsCpZmyjvp+gk65C4a2m3ogz
E0aWIXF/4dXvMuGVwBYNTWc8beYYgTS8VRoZzb1r+f5PU7q8zlfLnc/I8hY/aNmu
FF30iOqnLRGFpVsaPYk+F/YtHp/jZe3fFOZ8mPME7kCJKRzJnDjLg8PXfMmXfPOL
78Gbl0m67BKLFxdzkYFX6hzG+elxzxHHMj2Xv8pxPnIAaoEer2TJ4EdYY8Qco7WN
Sf95FykWhCjtTdk2fzIeeFFElYVvpRvInlFT7Dq7eUGxoUqCbdhY7kmwe4KpTwEY
wb6iDOyhB6M05i5FW24fm/3WzFDdWI/FWJhUw4Fm/w5e+vNb3+d0n7Mh3kwz5Pxc
K7FtAaI9vkKg5cA72DrTQJZWmwmoxXd0ezQ3ga/x6HqKdzN7NeGInKsEFW8+PqY7
3J2OSXgOeS+1imYXUY5iX66DIzPVbTdo7OSVBA1SJKHa0DNB5eU9UVhPotY1eD56
0BlPVx1b2uMR+5Kb4Vyiy2S99PRJw80d7bN6JrQhT01u7VjSIm3EESm5XO6Zp90w
BRIGm7/n1IM1AnZPRylOg7dAmeSQBDXUGzD9RbQ0gHmuQN+eswp/dHNnBO2DDmhj
/KknWbyW6wZPDZCA6I1H7HLlBxblkR112Cyn3z4ewz0B/5+kRyUpXrVlWjuBsL3D
BxebmGnRR8Yc3WrDKcUA6x6eXo6wSSgdTa8gUuH9S6qjpEToK6z2T8b6d9y9xoNw
RFsapVeW7rSjGpGlacW1vfyz9k+/ViXDJ+qYe8PSZPVLyrKGQhae7igimxwWbk+4
IaoZAk2yyqXIlMjMooz6/Bl+5ieRYSlEal2foNDikwe3uBTNgCjh7mQFhWuG2w3t
h+CBxp1prQMXwN3U53ff7FYHNBn0QPJLtZZlnZ9sKK8/xHw/1BaJJzD6SJMCBJ2T
4uxqlsyFQUVKq6RYDOF9hu6LCbuDKsUi8qMcGWsYEGhCBz173Ry6xztsXHwiTVYf
iPWTVASUQImthd2SPscJORrnyli0ziwPoloWHpVX2/XyCIcfCfsACZrNI/yAMcAp
/8ar/kv6hDQzCAZz+3ni7yF9OdhNCDnBRLGG+CLchPNAidK1x65FH3sRZ2rJU2ry
idjy2vCnnuSBOB7eIFLiV6JwRqNJ3BhrQJmlwUoXfMkjn5tVVxM5OY0OjxkE3LWq
D6NpOExgvJ/ArDQpzgmPwcWspMw4fOOPeSQyiIv6PntE9svmMs6EsAuwMQs6dNw6
if9L76ZiUe2t0XPVR0fHa/gbmvOFdmGCSJsetLULlJoA9kBLPP80+wfanWrW51Xw
8cfoG/IMfU676TSRzJPBKFrEVOjraZYjVuxkDrXSrmfFJOsr+UCCK+dSY3Hp+2xF
ocKYShg6Ss1OhIPBfVU4wH0pBq1WoxX1HTadIlpIDd1LcQ3OMgL8WcJdaa7jawe6
I75bN45/FZQKwDQ0CGtRuhBLi5LW37H6UNCT2JjHf5Iu7MSe0nho+WtTFem2TeWY
GnN5lHR+Cn5Ky/GYjFZwJgwA2yMN5Oo/CtPcLNQMok35SK/+4HW6eBMDguiJ0x9M
7EmjmCvxAcF/PGtJfXqWp1QYo3uW7AlHNmPfrOMtwPWXtOpfoyDuJwCtpwvQ4SOE
qPAKP+PTLmriHck533z+4VLX3iBuu0nfyGLTTsxkmtLf6LhQT8hglp1ZYZ0a9RL7
SSLaAZYfTER0H7yITEE4bM2ZL+u2j7RGLIDssHqNyS2oFOUqzalv0sukVjIPzT2u
f6gfMrxiKBG+Yyox/BLkFmZI8VTLKmxMACAoaRBEdd2Z0A+6HB+i3XeudChSnsbS
muW7M8rJ8XaqEf7UNPXPvsmZqvc5FP+8V1CZayHjfytXbXYYBiluC36qKycwpOww
jPmyMzOhGjvCWCQ8lNHYW1Z4DbQAVGvMy0GZxmkzoU5n6BwpEN9zgWhOZVy/JWJe
9Zno5qpraH9n5ja/ZdS8X7NeJqoPL1Hp8x83urnREmhYGMgpzFur4RG2N7w+Ss+P
dHx1PcW2KLn4ETmfpSjS7wOhnSpFSDS8uqLBJQJXiL5FvfuZxzSRPeU4K9gl4BeQ
PFaVEuf2cEX7h/tX622vYkwOvNPyHb23qnUfOCNVVUp+bHxqREC9em5g0VqKQIQc
VfkOCaVwJp9zLNolUjaRhuuROqUOXPb0OZsAcMBHqqF4xw8JlHbYfYuI9KopH8+j
6FzcyPKUvvvlGSawgDZNn8DyZslmKgEG6+MjEyNmChln+0DIflkwetFGEeD1eoI7
ocg/BB1UncgrSFUThNohGArjlfO7P3rNNfvzIr2KwdRqRMcpGuTOiOqzcFON8c0r
U6VS+S/QEdS+Za1vqwYL/PEwuf8mk5eI/ISKmSmT3WlnjgpaiA4xW2dA0ybBB/z6
cEBdOzFyuAjlLW5sIiwtbW3kMf/nbhCftCiJU7NJMnQ7AmW+nW8y5Kk8YlDFNlXO
nrvBW9kCUzYtuvftPzn2zQ52DsngJ8y83rKFWeYL/jVAJY8pP9yuhS1QGdcLpy9k
40obtqvg53PXJE9iH8txR7NwGw1+LGe8gNktBLfOJ4RnYciz/+Tl26Nv2cuZ+Fll
Cz+sCQu1kJRdtSDYfjgHv62NTZAu1ib8rQ815w0kRR7w4u55e00/LTIIr/aSSoVH
13jxHMvovBBrC0lNuWEcNmpfASKrCuyC2DXNHqJxWhMf9EbODB/EupCftxmxIqoF
CLoh2MvBMp0G/HZRY7XJ4oImivNasyHOlWxpHs6q2cRmn/Lu278WO0VFxnb8veTb
Yc5Gm08VA60SmeSn8LknCgH/LrUH+9P/Kjo1PC8fGlPWUMlFXSGPMoU4jd1XYILk
NTN/EVr+B7XJX0xWohXr4JW58KLLVZwFT67m1E2pkHuSBP18QugmH8oncf6uiITb
KTA4/MDwOVLogBL/OyvIePthZ2kxZIom285jANC9EPjB8B6mUMNg7+wX9kSSPQ/w
XJ33gJRnq0uJE2XkCm+5EIDpKkJ3qV38d55fLJEG+D4iq6v05JFVo8DhEzuCYABu
UIAhY4ABsrkAWcnt7fpBF1qMTvKr2nvhITTPzXsAu8n9pMLHpPaHeazWV+mxYmED
1EsNLfihKs3i2W8x2XyG+AXWbQeucCCN+6NWBH4xrUftA0aucefpiKxKXgNbmXcU
FWBSFVqaoWfWlq6E/Vbl9fvDPTc9Jp/NCaC/Rx5T4ELX5EqSV5HRhnKtnZvsHrp4
nKxU2v8eJ/eAd+/TiBRydspGdUdolbebzIabgklbf02lxl4+36EP9yoeyg7cGLqV
vys5IAPvwYRGBjFwzRENyNQbfQHyqhviQDm9MR83L/jSKZWNZFwyAP3BZk9WAWIp
6dFmzuFWH+dDR8PTJsrZpqhAGK/hnM971A0nFsXxBUDyVwZJs5ivJpKVUTPuw42L
R6XNojgb93cI8wuVq5sadvtPLkS+INa5YWUWt9qqSF7CZwDKJ09kY6Z0HVYIBrcL
sk4QAkV+/U4p07zjgLbOqWr1qNYUFQlpWZN6nFduJdvfs2lzFHeIhPxMyGv7TmWs
ye56yV2V0gPNaYHYOO3ckYbUkKwD9hwF7hBpEZKnQX1AnswkF2aBdnUXUgww+M6z
lHora6TmAonFUvH3KxGjKcjweEB2/26APdAXjRMgsx3XmYjKVFo7P9F2cKWfLMt1
gRdSBOQubqk6vaxr311zefzusTWQZF60id2VXkKsiElazPUwJUVU4fTcX4M2qXPV
TaqjOswv0UrGpkcpHgDCRRVTa/t++j0zZBJyWcErYRvrgEunFF9i9u85qee4OEkZ
36gmDkpKr/NY0+GIKGnRfNObaNih5FbQC+pBfcLL6jKKuC+GrAJ9L/gxIo0M3qPh
MiqK+0QoGCGx3HjW5TgaFTGIv4rkS0xOVqOjdCTWpNhU+I/IB2uh7GLgt0BeRwEQ
BenShSDSa4UoAzt0RHrSB8htJ4K6fzupu1L0lKuJO8Jpd8aIoItsO8if7C1P4OGm
lv5+xZ9oXTxfbJ9tVDR1V9hIiav8y2yUxVONxPhVt9WNessZKyoVq6ZMNNYHyU4j
ChwgkEFqwdSanDaPW2APOIA7UoWIdawmV4jYhTVT2r2TbY42O9hsBKx6+01GJzSf
rqLFQzaj/X7/o8+m0GqygyET7vSGzEjrO294PVCCm80arIXdc3AHhWdbsoDS8prC
1A8OD17x2BoS6xIKewXPGAf5bqe5eex//zep10u+v06jBmEB0rcjb9Rq4pXc2EXc
5ypNZ1KivcqqlD9/wu0uAG3uP1Z39hYuEFFmpmuby7GmJ1eIt/o7H2YB2dg6Npg3
quCq9Ky4xK0yjOjC5bzujsBuYL2wG3aFmgBXQKo5Bx10gfe40qJHt7+sKqbfI8qh
JNbeTIbQh2hhIpa0RelTednWi7KyxTS3uATPDw7lZMaWPggVMVAtZux4whL/FV/W
50JTTUkqMA348PDHq3FUqqesHDTm4QyBIo8IbO7P9dl+JOg/PlgR7x5zG+KzqHuB
dlUKTkfsj2uE1J9Cb1wJfkFWJzCqxHwF+K9xzAiitOnFdKqJpMuDmudjKryjyjUw
OHtzKePuFnP6B4ouQolXJtWAhq8kttsXNaowXqWXdntD5KHjos0E1u+4zfbTfMFv
O4dd+CMALNmdQ/t2f1/lF7yBbEVY/uLFh3sbobWSZkfsg+wH8RCmFfyzisRfrcT8
2+JEOijV1KP1azDbazyJ/2WAjtFiKe1HOXVQmJLTECuFMXBRgKD8FQQoWk08P6fh
ycdAVVDRl9a2Grkv1HO1nJ8k9+jdaA90yO079UN6Nk6+ojB2B1ZDYnfpOhvkJ6DC
H8WpEodBe3uOAQn24L3/72nMqqklgPkg2pEXqi2DsGeBK+I77eITIJUTQOoynrdZ
7pkvRrC3xKpyYN4cynnokoy5EjrU9FPr3+aHEA2krZ1aju0NdJRps9WgZ5M3W0yl
i2QRsfiJfawZyc2ms/e8aOAI2iSwpV9HX9UDG2H0hiyWwu7lBrLm++WraNrPItqB
PpVN5o0XS3Ev6u4xYBU96wthT0wTzI59yGBMoP2N4zqQPC1UREdkuPCaquWSNSe5
EhtKMJw3Z3wjviavKbNgPEpIAEFGfFIoVDmwM+K/6A+hX8ox2pcc8zxBOQ/YZ/Qa
u9REd6H9hT5SSMxW9eGf1B6o264UlfM2yiw6cGo/nhL2WgADbkHoXUyPEgL4S29Y
vU1lcY4o0HAc+nTfAqKcYsCWdNmbC25DmWNI/eZrr+Ke0EwJIK+Hn2TtvcoVRtun
63Tf5BINHBcjzFDFaR6r5EKzN+GBZV9gYHySTsVU32JLKzdJC0Lisa4nqYkBhlqG
VwyfG6lVD2dBLckPluPjZTnK5GeWPTGryAexd+GEq3tSCcLSf6mNeLP1VBQTNgYt
TSqxjvFwAjHkSJSU9xGTmsjqQfzadoVSf9LT/oEX7rkmvoiU3FmS+AvImO76GpsB
8H2njnp7ITVwemhJ2ItjY4i0yj/NmW8AELuz+BsdRS4/Dr3nCld9IcwB1BlBEkYi
nYVKNHM5MRar+9yrcnNPhSflZ8KxbyzvDcd3O2hboFid3+HLy6Shqv7nkmf+qrKc
5ZcfEM9o7+fvOS7i9br68BOk3tGQgHeXFXHCSbjPbZzslxlA/KP850uh0X2tdvjW
IdUu4w1qIctiJELOZB4AtnHSQ0XM3yeSrnbyuCHosaRCo3oZpZeZrp6Gt8z+dW3i
Zrfp54UJRCe6nAxZ5nXumLS3JQJ+cx+3ZmYyaVncmMBevmWUCsi2SMEsMyelh6El
2uZDFtzVH5Oq3pRzhR/Un39GV8jgs7hQqwAL1DUTyRnAzjArB6109hy1eGsQNv9Y
qbb6UbHgfvpQ9taWZvpDJwcqm6q2+WwOBe4ah81q+xs7ORr2OoW3gtG/2hAmSrsB
ltZpNFZDc5Qsls+P7942B4NDZXLQ63nbd3129f262Obu9+iK4Be/I3RLaaNb2l6S
j/XFZDfqcIpaARQb2avyxKT9oUHSKBKe923Vtc8zuNUyq4eR2gtrsU/5+LoPPuBh
5xdrgJXpt+8rJIb4zXmlzQTRh1gUKXAnxhANiBVX4ekLzZirXf14Gh2qVOUD0+jM
BtELEVB11+IN8yQlTvgdZ3ElYnCL1GHQpQXO/cxa0oPQrGpLRPv57AbMlTDoCTQd
wcaJUdzFLiF46MmGmRxYEA5wWT0aG0AErSKy8YOgRblFlN2FbV87Dle6dAfr+2AX
W9kcztr4gmOWNxdCqXtslQ2XChDcVU+dSVbdEoYneKt0nLFQEiiAJpgYx2ISt6s+
5MNOFJdG023VDLjHxkBxlEXKmuFGL1fIfp56RUJbcp4upyFjgg+0WEDloLHdgeG0
CRVlDZmmJSHzN5sYD+CT5ITJDhi8rV3iQIJQo/P6BCixPtStGfFtie7MUi47t9HA
b3MGCNQ2NfYlc94cj/cZ80fmAxl1+sx+LRrSlMWjZdimk6voH0LLrye5EOHS5KiL
QlaLBYQVhhpbcWOUJTwgf5OGLPeOaqUVF1voeC1GkH3XHixGDzDKdBFAxU7t+9Rc
UrN7TkLx+Vu3EcIxRVPmv95DtYr2h4tFeeCT3PUTHnwlF85sQ/eQbuIk4S6YIfn9
iaQKrtJMRqM3wvIjKZtGajd8ITzRhacUbJifbLA4iP3WulL3OktDuLi1sA8Af9O5
Bpi6UPg0Z0kXtjtVatWfwsjPQX4XRrOmbXxzQJuoA28p3pHFCF0PG0VbS7QhwyJd
TjTN1unqBnsarKHtSjLWbfRinbejI5P8e6Irw1x0/mJY2IRBD1kjSYWWrh/i3Xtm
jHgNOVctzOd//NRlBC9Bnp0T+7Dh10eJTX0G45wFclW1SxZYXo+E0OyCo7CYDSsq
n2lpwsnUNX3yyJG2rEhAktGiMg6+kLzpTr0NK1nY/qh4ZqRVe6d/D7mI7LPeSnyQ
l8PHMafsAswynUDM9+a/9bFgYFMSW7ug6ZNG0i3hUs3Qgl8O13Cid5CqgS2rfJcH
5Edz9rRzO7IC8gSwIVDbxB1E8YRybz9XVwh6k0YsWYh6btb49R49nLbHUySHINn8
XrHKWky95CRtgsMLftGKyeiZ6Or9gUWo7H6jaBZMZdup8oe9KqORKUcXy6rN7s9F
XJccLE4ldWNhtqTmForB82CRr3Qfh/ZE08TvXt+JGXOLTbEI3GuCubTJb6nbDX7q
l4QASA4yT2JihAXvfhiBwk2gBU3rPGXHszGoRNvFFACjwsNDzlY+lX7pMkffNctZ
uSD3u1I7mgrvbAngGOQZGDVMBpFrUSW7zEDl7IxwOMhT1oCJpRIpVS5xQRDy+Buz
rPCpSANszOLWhWD39HCnl6GGnDG0DSJJi+42PpTJhowFwu0GJom9aB7ri2G8PjxK
4AYj2vf5OaVycPATDv/2K4a8sKdBusz4mColw/PGDogQ3b6UiEMlcx56J5UT3goQ
OTf3aer5ax54dxv/Qav1zstUg69+N7VVzNbcMhKyYm+n3asq6qujf7a6R9CE+gHo
28Vy71XtNk7+RE2yfeiF2Y3hIclBJSoFr42sUbeKcewuwxMAN85SY4cf12z7DLqp
gDWjM1dYae/6+tw4mbL0fTWvpeciU1VrK4oNkqL7/niirTlFkrYZcMGwQUbT1frI
9LeqPRa+TPqG3KuphINjUPQ1Jpt2PoduCcb99At/XQ3bbzC9Slj7D2anGC/yVnJW
9Nst7O7dnq5vHcrOK8EySKPYa3Yn9AYMcOSUIkyz67j2mdHq7EZ5PaKmo45GkpRb
Rv8u8G1bYzH/YI8xY9gsN15DJjgGMvHh6kB6sGcA5ODNE7WfT5sO9F3vO61P18b/
2BuquTGZLmYwIKtQmTyDNSdWtS69hmy/6utawB2HuI3Gtj7eD3PNNiSgui3Jh9b2
s1ZAAVJL9r1FiM1/2Td+gMhr1iNgipTNazZWYaq8IYEhD4xHAdP6fY8/WpRUl1lH
eGkN9//wntsqczThcmenbHMgFa8Z65CoKqsrxdVgqOT8KW3j2LGLtNgR+YR7Eode
cdEQJ+urH6wvoTjynS+YSSoRVU/3L+N1sWzw/+70B0HhpmfYnLVGxZhc3+1VF9wU
992XIzwLwWQYMR70fntvFivN3iciSBYZsxcYwZxESvFcQHJUxy+gY2WUD7QMrc0G
o2l/0x4tS7zhA55TgYM8YoPEHqL7wlSSFohiPEJQQ1MPeyx9uu7etXShhNX0gRtV
D3C1iawPFrxQ48ydn2p7ShA493CFgWD5b+hxfGjPDu5TXj03p3zWjmLrJkaDaQl1
h0Yg6d9/LhSduQFoqYygKbvmbSN8LHfok8Gbq5YZGf5YniyMxKldl5uZaEjbijKo
7LXNoNlazb5fV+dFRK/yfk8cQLyte1wnPITAS4nVslSShzmsum0JRIJYpaxtnwUK
gT05sorL1AXA3wcp+SDLP+MN6MVyMif5sYdyCr0F80hU0MhebvYfEjXI6V80zJ0H
cUc2MaeY7tnxAuC8O4VhncsSl1lT9LBw6x1N8ubCqDaAz5ZIqWjweq/18TYdxmpF
f2mZ+oCJp2PTmzqaTrC2rrClIY6/KBIPoRQ/NnzGZRSQ1AP4RDqZmt4BlwCvSQ7w
TfaHpqi1utwuTXGlSeQUafgvC83OO32Pw33IiqV0bOOPLD3J2mhV/IAQGV5lNM+d
RY8uHwwxopP2xUqvOd9fPlZKp4k7BY5qef5Ie4JCGNuib8FKswHVnq8pRtuKBHoY
QGYOH4xIruRGr7MdUbxUnPycRvsFsQpaiBPOw6J26SdohCql0jd+etZYb9/lkcag
fkaNCbeOGd6qAi5NLQ0HREddUZRd7d1h22+UW6kJe1AMMWatnutGzX5aqrCZQXSS
iiNHPyBDP0EVQtyrzkXRdluj/8NzlC9kmSVSe6I0E9bw503y4YSnsmUowvihp9N7
gjkTVtG1dxvY9c3D5Rf9s5+htfKnp7ReLFawi0bPeH3d3rmk/Q3DxFHRSw15dNin
tR06aNsHI1tWbQ+xqsiqruboMRcYOYLBwCHqkwLFYxA6Oic1vqqsNZZ5Q6Ni7gnN
mf/CcJI8maTO+kmCYO1WAz0Qb3n0SZnv360fqhYNgJ2vVw8pFHppgWREOaWDD65f
P6n8IBRWMJAhIwr0NXz4NU64vbMtejv42d+YzaDB0YRD72ESD1leYHC4rfiGqNWA
aJ/RBmIdnmB1/eCxworDC4vCimW41CKBD/XFiXIZSjJKvPhuwD/NkYF3+9whS+o/
L3dEGBTVzbWjvGRP0M3mB7cwryN2OFVrD1Bcqk+lzYNqkvJEBLvFD1YqIUwJVvu0
Uf7I/VCsg0wGxvL2F5hY+9qbqtQJ4lWTau6yQe3v7bsP+MsFRFcnd8G3m+dadfgb
aU/FupBk4KNN/jsVUAE1ivfm8VOrmdHM0wYpjHgv0PeXBTq/g2OmjXnUTXNBLSOq
ID1fMX+j6J58m7iWnIqSEJZm/s471y3mAINul4NW1tjej/r210EXoIJ/hFcuHG0S
/SQZUSbwwyfTVrsR5A7ZiTuCm2SNfjioVt7z46DSJ6DGBxrM9at4QvHnAaXaXUDQ
IvzgZ4x+e4pHDQs0eIi/Yt9MUmqW5r5xqYGjTgmaLJQGlfBpugPv9ESRKW9mFq6q
T2MoLa2/ZxcfkchuOnlDm5/OTnF321aGn/RVCAQ2Jy3Tf+KBAj7TbJbY3/p7hN/N
zCdwueSpuLdu73k1KK9b+y/tauIsvxThh6yim1Ld7wFi90F6RNYxgLL+DMfu6dTr
npJK2k4rzTnm8ir7tLBl+OCRxCPYuRu0g00j6vrWL/9aejI778QabmS8VOMopQji
lRwoz+oQBj1YaDC/qDtlE7qB1JNUn06U99nIKI3bLUk8BKpxLtju5KG5zT6f3WbW
mVsmHHTrLx1UVQrh0jVEPYDT4F7KYWM99TpwIH/Dm9sPTTT6DpnCNNxgXPy9RGdH
peD+jYs8x9M67T6PMkM3TuT4qpHOtRM8Fm0Jtl0i6EtVb1jtWLvKRIunvwrRooAJ
KPiQhpVe76BHCmBYAVdyTQ4wsTzkWvH2vXpmqY4+L21fR8DgklkEwlFhPAhYNbtF
ygkhMHuj8eOMmTrwPpkCrK8E6YrLeW4dumI7JklGsyYnj2m3/MO9Z/YTEfxg4JO+
4qo0ncs1yzo5+4Ps4UizM653Vx/H3yIwL8NVpDOVCaeuitosLQLYr87bKb789kU1
4OMJ73S04JmbIqxi2/DeZMw0JVJm4FMdyieSmRbFPeXyNcjpZcCt+v7Bl8sOUhgu
WbUJbtNiVIsyT9STjuahryFaaxlT+/6vVrY2KFYrEcyu1JuGGYVjadrFneuZntQw
NkDZCfyILYEdH0MyokJSXJrnMndo6LNGpGMD20okvt0cenCIApT4zLhHoX+myXA3
8Vld5G8F0UCBCjnn/aGPOyQrvTtAArBgGB8jExIbAv+wpfa6h4CKlEXfELF1Qe5h
2XPkYY10IN3Z1aL9B9bqBAlmU0iqn2Er8Lbj+GXxUFdZ/jn1o2ZGub99WDXLyWHA
g/QAJ4nwqLQVnkqRgEY2cGRPOJ15jKnK2D9yputFogGA46r7kTSlGUiYE+9xqmMu
3ueu3D7Uos/lFXXBNOreVxZbpoMqI1rYih98ExSvcrFuQSpSi8aKbkqeC9KOMQH2
N8eBP6DXTpKFBO73MxEwHLQv9uQisFD3sfpr253Jxv1tq4FWHSRa0yh0qM0lEkYX
8G9Y4Pa9Ay1705gFoQUeO1mlvjwht2I7aIzf3Z0cq24beKJXyrM4gJUxW857/m0w
QmkH5vqcQERCM6l+82Tglo5nclky5IAUVzhDTa52xgiEEGGbJ/00b5s/wDTxJFuf
vVXUAqNM6ehkOIjiBKeaV0BZJBVOuwrEDMiKN1hZ9eSqZmF5l+Vg+C8awgNDpii4
3/reRtm37JeOLLCy9e5ND9NAHJYKE00JdIeEnBGumQcspZf1RLgnUwsRduXOMOo2
+I8WW7BisMstZy+ZlnDL+e7ZBOrqzfhfMcU1hJLkcQeqm/1gifDJqrowyNijvo1s
wI66G+ObMwZuU6a3no/zzY5fEzT8OvbIEStrS+Nx00vRVXBOPvJ5LNwFY6sDMPke
+IwTgGRNKzlwWV1g9/NqRA9mSDo54pGy5Q598icDIuYKrH3bm01Ctao3el5lgyiO
LN/W8yLkp8atbC5XVR3U33aPFlkvmU2O/3IAIJUPe+MZnE52uCI8BtWFUo6vQe/z
4+/dcJv1/aZ4teRNojb7HkhkcccaCqnNTOYWXuLQa22K+9kPD1eg4y4lMCjFW5ww
9SvLyXMaNBfJWVERDa+xbWJ+lpyAnHPAk8h8hD9H4NI1ZpBTH3Shs30s3XGL2CX+
LIRRzAJOdDsx6ku2mJ+vYFW7nvFrOEQrdd9jNbCsh1/1e4t2t26wosknjxaZYO6Z
KdDe//D6x0Uy5VU54qel0qZlI38Z5HnhzYp5xsG8yDZRzpyS7Bb1+8FvCTLtpdd+
wblyPNUu/c/5gowQGbeuz6C+BKQLRllOHmPFCOC3ARqgQ34j68pLb77PJtNLtSuR
rXFoQd/NStyIxwFcnQsApJ0F2Wq60ZgK7w0QLvSSofkJt0ZDk3NlVW/UvsJU3spF
36DyekNtiZbeW4q9OKWAP8M5fmTY0tzbCWiLqCtop3d6dSl0NQ3wXglndZ2brN1/
mgcd51HCgbOxhoTP9ieZWeiIMvpzKw6wTkRGgMh8ZehLMgKKhZeKgTRKod+rtKx6
MJOaG9ikxypWpPoQlYb/gICxWb8XSTB26nHmCRESvSOBq85G9GpNZ6sIAsRRzMWD
S00u9hIln198POLzWK4OL6841YMriBL8Gkpz3SoUk5oKq8o9Vc6poevl96XXR/5Y
XhqgiDO+mqyEp6yY5+xI+ktZ3JCuKGv+EiWOfUp7jMT7RdBAxf6M7+BnIYC85e9d
+3KRFrXtEXN/vwxUw2m9t/ffwtgyUj2UParo5A9eJnB5rg9SOsmYN1knJYSc+DgX
8UdJDH4SVamCjqRQaGxn/FboIiXaBiVflwxJFluDJBI80EvQIag1bH83GB/qPuUc
ilwLDRVNlUrV911LmXVyRdmVXBd8ink5+kuHXxjMigQbdT6VH2cs0jzWbQCfE/jv
Ax+zrvJz+SvPQ2NRCcFKOIhD2zGwEw4IYDSlBJx+buwmtSvz3QInLKeGtnJFF3aG
64DSXBIz3x1E2wSC4iSiQQDXD9CIGnxUED9zul6gHTrYqLTrGZaB4p+T2LZVDTxp
zWnP8qjK3+uzhXF+j2ea/a0+XzeWSPRsl0S1UVgW+NNDz3p77r8s2rA79VQ8rVHY
IT2WPFXVwXqWwT5bVYPa3iY00Qd9QfF4TaAWhmcdM6epVlA6tg6wY4BJMdfKzDPu
ncwAwRuFuEDXyzTYPPJ/LRPLYj496TtVWESDcoblbYzmkIJUwhY6dbBBr6Lg1BlG
UqO6isjwnSKDyf0+qpdu1nZwxLtmrq7wUNOKIHpP07TC0nHxw4hY73ABeSTZQNo1
7jl+SlHH2hyt/q4ptU9ghw1DqoI9XA2w035qKokL8UgVpDCTwdzVXEmFi/n6cw5O
UxxXE6YMbzBrytOwFoz4ZGWH6gwNUg787VEd1LXMPL2BFox3ZwiIyaHphsft1FdO
vOYYRfQdcnHrdTK4vtq2Mh1PWC2oHCEu3n7bZT9zh5VqPKR4XIPUdTZ6TdOUtKwc
+UaJuuG7KiaPfn8BPiu53nF25X0XyzUuD9LoiUL/Q0Z76FmbTf6UjX4+6fsFnpLJ
9a8G75Onl3QFUALwHyMjtWEu+baj11yVy062uO26WtJL3Dcy7QIIOK71ar1dBKZ0
3L7J1kUC8SSn52V7DpAfyZBAJwlOnkSGCiSbl+tlgu2jpT3iYg/0kC1InpRmFArI
jmz+kGn9kF1egTh+ygeW20XqwBsdrhV9Mi5ylUR62xVVFTtpBI1aTKMfhPTKE1PJ
KcC2RtAHBMwlhlbMMqWbMISLAFxhx9gGUP3b6DBWX0ccXANivT+ycm7CsfRW1hXa
5fi3OZQpa3KELuc1BTCnpI8wnBmWBUxojvYFat/dht+3/TXihHCf+hlnLByofRaR
juOCSATtSbq37quLZD9vFKBTbDlSMvPLH6AgTrLOCEcyo8s87rDdT+mpb2F0YRJf
LxV126yofhaNwUu8ZgEy0DExjEsiWaVBrpG6DQ5FKzu34qxvGB0zjc7yM8yROr3L
I43QOiPVD6b1m+XYgM625l8ksOMbQtXBEDPEx0ymoPltGTJvu4sOkcsnhkZwlxMc
3khq+MW3DXyrNjpBwO6AJMeljYimdZZfv/U/xU3niSehNwRdFs8wfpz2s6Cw6x6B
LgVpRTJVqls9AO1MWAyOmNfpgMO3M5dDcy3n5IorS+0cKbFprSpx25IQ3CnfL7Wg
yh4pePyt04WUK8l6+2aJ4H+xPiooPrBKQN0R9nIhHqP3/Jg21pQgC5LwAu5zS0SQ
Ijqvd0xRfRXHUlcYP60zOcTZVFJ4w75fKiVvfxWtweAyNOWOhegF57IgayZgK+lD
3OJS17q1d8CeecwXGdIH8LR1Wwsmwp3n93TApLpjBZJ+Kzigi7BhmMjN2rKayYAJ
+gjAc3LwpkS+OgAzTS9UtwLuV8izQxj4s8h7eXsE0qkoVL93dBdxVthi/Lt7R2p+
FHgyQ1c+CctP1yYI0aYEkZlcXTzQrwA3kRCocfQjfo5/P6NKr8rvoFEHh7gyrZUy
uEoFzm4Y0iS6ouL+e9M4rnNqS9GI/rEvXQv0a90GBHA99dAz+ShS3QyhjKrmqToW
l6Zp8HDsK+0z57qRwvDXVbkIfOIpL2WgUJ231GPoWKFqQkhCp7T8AFR2UTkb0ZXC
UgyhZcFv8rhZiVAFn2lxdobmoOxoF/QDc6hjvX6fHpi+aWhSr81ibVVlmJh7h28h
qFuQ6Pjn41Leh07xfsnXjLIpBL0FLG22Cms89aA6G9V/l5wu5oKOGeeQ91iZO7k4
XZ/CEcRed1hLDkKHy6KEg9OvnAjs7sfWbkVBKNpA00GclRhxlSm+zJtUScreNqKV
w8yIQjF51m8h+0IJRiWDsIYDZw4668+DMla7Tm2/2zqyaCxOHQ0BuQKii/ssnMAF
o7RustSbWUU7iZ8icBdeB8VENgS+6HgPtEH/O7fiNGWN7ce/HEPgaGF52MrPXj7H
w435etKeQHjLcFBJSRXMoDSkVNUgRInYWWZZlYnRkorP83Fc9Tf/Dj9qN02GnE2x
f6WDdmRzFWoZ9kqXWHPKvzuT+smOZEDOpmSN15W/xn6OHpnQsZN/+voZlP64SB0D
blxuGODCS8s8i+g4OhyWItQvVpy9r/NQ12lSB5fJOIsYi2Rnoi/yo6G9m555TBeG
jCliJD8RFuaBaxC6jixE+n4t+50L4CwV+JqkK/KcAxIYls3/ZgVkFf/DsECpB1ng
dTzLcQzJY4PJwsWfg+cIf8NptDbT/XW8rUnfsHAqUSEtMcTRKtl2Q7XP+C+AQOHm
O+X8NFF9JQszRFaCLM1MKPLBtHHcyKisvoEjyTipXWNSOtFxhaGOxYlfzvbuZJvW
AhOen7uXgAWL/K9BFPDiiKI4PyyBzVkrmMy5Ui8qZ8H05JsdYIE055pUIzhK26H8
8BoN6U13aHNJFcNjQglKEXR0zC5qd4TzgYOqCo90AsIbvFk4wsxGZe32Z5YL3EDf
YirLNMMX++fBqQkJLjjqy4M22CfNGATEpuzXgjgOBgJ/KvamrrLMiWk72aPlAkfX
qHdtGA4gyKdtRwjxHZec5d28eP3BDdzo09SARGrISxsO4FP7FE7ur+h6mM4l5uI/
7ng83H8862a8ID7t8XL7Lovhzwp3bbhwLhpmuf/ZmeL/3uJvlcC7c7IYztA+Q9h0
bj0C0nfCfHsE5h30l64HBh9RFUsGqtNlUGu1+LiAlTJ21oIbOi9mIFfa9HK54NbI
i4T98VrB7KjTKHBtu0Ul5iUJ9jc0sb+Kjydg0RqN4whsJqAbWgrFIEsM/Ic1GYCE
3hKl0LVOTj1h2jWXViZZQghAQyPIxnr9i6zmLRt3NPZh1xvS0DtDNybYlnPjUkjU
i3j6SiNfCLubsVngQDBB1n8teV/Z0tL+6Fr8oCesn6AK7PCe4SSbWZuC4LaoG2Lc
QTzfgfiiyReD5FjOPNSAs8HXNHAkk2w9FAAZkVCwjS5adsbUhj2ShoX8c+qCtwAk
mfoTfJxgkuXJJYPPolUdNCOmGdLGNf5J9BlJ3v/kKglJYZ3oUKja6z3X+509o1EG
fF4C8lwhG23SQxKVr+shnyJBdyqKuQHab204mnXT1hXl36v1aqokmvpKHBan3z73
zOsd49vjb7HCo+YroYvU8Y7jctrL30+QrkdHSnSGyhKczly4lapTczeN5nMZpgHz
fXfgZVsCG2Zuk7QbSCgr0jr6+adtSlK8iXRv6DenrCXIPDdPvyBySucsTgCTP0vD
M/r9mZ5wZUxG7C4gGMYIQd6jOOIEEe+S8G6kYgm52nGc5flbhHDQPaL++0tvEn7k
6SrJN201ycUAiBg4J9n7IZOqFjqUZ0PwSgZUtW5tZjav7QRf7zA5x6q2HyKr7vAR
j0fRPUc9Za1omvV/v8OUxvEJWFTAlpG0qgHSVsJ0uiquAGaVO/pAaNWBCmBGXmF6
pYR2aHy3C2I6yr44yvieSyDF4bRiRnNudm2wdeu1T/2q0trI72OVoytPRRO4pb/s
JK6nOVWBTnKqcR4wKEc5L5KWoNfVIjI5YelhLRZzk3EB4NI1TOY9dUlKS6F5SRWm
pYkrY2feMcxxhr1TQpCaqDClckdjF9MEHi6Tbxp60KU938k/+7K1EmD/SlOIC3g+
gBg0v754oJfhORIRs3Zu+2jdl1E18yuELOveNLVE9oc8osk+AGcZ3xSAqXF741bo
4WMshF2tnpUc9ZAFrJhdURIXVbeExFb9Iy4wGszcf09P0f4xChBeuz7AO1U/Wcum
Byv3/iopihJuU2dlQh8Ejec1iGMUpzq1GuRGAT2MeOCbBTTRXbqb38uQ5D4RA/Vw
Nfs+4z9Qi6Zg9uhq45lL0BdvLTVFHvjMeCBtKdlbdJgokniGWmQw0YniJCRjyXqF
b/cOqeBpI/FflsXHp7YkWgsZlO1bF9v6ai3YvA8LAQKvS3nZftO19DJLn6QQkUtN
bQvR7xnuiF3x/UYA15kqKAszE6S+1iDXfQQyY3BhU7yglK1fgN0k2kPGEUZTUHrH
vulPHP1e1tcV0ld4dR8/V2Qdv0qSnxz25mgE6S5NCnNAXSBGKCavQojVIoTBlRTa
PZLGnpw9etwG3C3JE95PiHtp9AZ73L2onOVTCvWe0HhaRdv6A6HfGmIz5RwdVNvT
BsW7+q/RokkDoPITgWL9gz3YGEfg8vbgjuG0aNRziebPGeXis6VHQCp47TNTTlYl
Re33MvYLM9hu961O3fHYcxoCK+m8h21QROnQp4D0zdSYz/7wJqdbh8wIxc3XDhts
DWt66iEOTxX87ZNtny8ikjhiNdlwyoz6I9kBOnrsKx+FNKOy2oX+D287JsUKyE5T
iQTx+f5lYEfH9+tq5of7ULdEHJnP7yJ4PbH6mKzFaLqQ4vZp5G0/4/myMDUko9Q0
MbTw7y9sLQ1ZloBkwjMgWtMJxzOc5ULqENCYp3t3lW7EcqkG4bgijK7zx/K6jHEA
B0VbyDP9gj/QojRB89nFD0t87o9QMJj8ti1O8dD9eJmNhK3PW73DOh4nKMrjA85M
36/chRO6yvpPV21T+MEnB1nv1HMaUwYUj3UkoZL4RB41Le0EKib64JOTxw/ZfLnF
9MS3QgNgfhOHcBTvKZm84OdVW5KZLb7kW1hzFurnVCcTSbIXe9yQlLAL3UwsoEA9
UWnEOV2+SU27v3qDEID62VfaSnHlhx5lhJuTc2DXX3TEM5y+bXKgCdjT22BNyAKj
rGVtMc6n0tApKrzA4wdn/Ykuwm90Cyvw73KZNjbRu0hEJmL/DbcDLfSq0VTv02iL
bGSsoXRbfKYpn5MQjb/4upXnktMqDIjbjbGAyY5ObhaJEayPtAYPcjAQaYpTjhRs
a0dyQeNjjsMw5vPOUzxDTnx8x+S/WpiK3BO2pdeQhRNNYkdkV/IyBKAa/SBJmLdJ
reTdiurqpooDx+VDEuCMFdgEbNC3SNngJ/cYPoLb+HjQvCo2+MaFw1R93EAe//Vx
PfZdl8DL9pNwnHrokpvk1PubT/KlH9y3zZgv56O5JO6k7jJ9p0aj6uuMDTL6QZ9Y
I0/dctSeXVL1x1Z8NZ0WOJCjXn4sHDOitxLVsa0IlldBSsgBTbM2RXEiJMFO2ioD
rSjrOz2X0zy3IU7KTWtz66hAxjiSKS8PncbQwxuDxac0YdhmBYfj3Y4lU+RhYYw3
gV0mL1Kmmk5jDBvVzP3B5wtC+TJX7V1kgWsru14BjDwuCFGTtmIXs/u8gwlHjucQ
OiEyFa1MBHfkj5hpbwfqrd7DFR2msDsikEH1UhcjU2xwvfCouGenuIWzUv4E4rH7
9yDFfSSVTlbrwWESBqwoy3ivllzVoiUgI+5QJ7SH8dcQoMnT24BFpFExkkZxrJrl
QqvSbOGOR40PKyyl4OMi/+X8clvnu4DPWzQM3DFKyuaocrklax3aMr3dNtKYdE8N
pfUGJEgywJQMHNn6hh2xkNDEGMbTij0ehw4sdru0JeThAu27LbiJfT7a8YJAtDDs
JsTjIy208FxBuH4GT4Fo1O4/Eb7KlUrzmgGuPVmgyHUAe7azVRXcvWkvlgeKrJ7b
efKICmoa9QJSB9vWzqUE45enVHnk3aXkVW37gdigSbELVUQtYD1JWjtxMyRqtQj2
0kJ4dZVWivwGL5+btPMxCasIazrYbfQ0bzVB+QVB7SSxrgOXG9dyzO/0FkHanQ/u
etVrPJ1V/0fJZ0dQX0/zbL0Gk8nNceFp/QQ9j/gtm2XzO91zNENYVvD7JY6oCtVa
E0c1EEzLFeE0Lc6O/GFYHica2BZRJEztzUGNLKqjbFGqsQ12mjZBs672630/TjFv
fnd2ybsk/tpMaQ0iVXQIrugCXCd3+1UabZxXqRwDovZSg/E+EWaIw2KARbcOaTQ2
ZzK4MYBxfwKzXCYnzudLEiBe0i3e/AmmZZf+5YafkJDAR+k+pCmgzgmHNZHxAcie
2yUUY2IYFwEQyL80DVCgyVVUOa5FFNfTPMv//H87+v/rT9DTgZeJigv7jdLS7mSb
9XhIMjkGNoThLgYwqcSqU9eG50sIWS3I/xo2hSDP/OtRdraZLwNJ3z2GnCw26G1e
YCF+DUtdS8HwjgbTSSUarXESoFAKZKVz26SBoF2+q3Vb2dQtM4ZLTgS/ILyUTDQI
vim79Lu49GECI9fmtgqKoLBziCWwuC41sJxdntvQWzS7eYxqdLEkgq/9WMFsVEyD
JQ8yWA+cAqrhdILS9mkqYrvUw9DdwOIV/jX/eRFcuX0QIX6+HIk4X6+c+pQF0UVS
bnyagV0My9XldyIsDQJLLfw1SPKNvTdypeP9UkDoDps1kR37HY/YgYbLrAm3IkLe
bPn7wMke/JDYlC8/29J/V40vSYmDhqwFNC32GQFOEqGtHGuLAy1c1cLUsOz+YCiY
m6l0c314bQNCzHMwDClnuvkjRPxoHlIopelhngfpQ3/f9fVcjHihiZYKlCZ3Mfkc
Fs6Exs/Jyn2aFmOmI7NeFi/vydfKyYoNs2S/qw4LZCnsPKD07n2nqFKLg4XjOmJ6
+2yyAO4mmGAUyFrZVVozquPx8PCHkxoEXbWppcfZY80pV1kp3oJRyFNW6BbPMNq7
sO0KDUrXin88wqq0/Vw08bN/xldCDcb6kThvUE9yGlNJ1aDZOgcM5NqoZ5Upx7lC
5985m/GIScyVN/2UT9MPLk0FTPWL+5vF5WRvZ/+6jNVMYmTiwBKB4HE0G+1ZfB3M
HLjaGUNGT9kz/c0NS1eXcntrZem4kJeOa0DzXnynbjP7lZ7ATtA9pYBU2dQmrOgC
AZNwNThjyNxWkB29QZy+NntfO5sI+JY4ypr6rSScLpTXISzxqv79vKgGL7vwkv4M
Qp9ohOJ4KkFPLHv+OlL/OmJVf+/RbDFWT0LMJtjoMdFDI7QWJiP8JGY0LmUk5Qv5
qatCrrM5PA0sCt6asyiHaOQJdNl7K/HhwXTqZroF+Db7gR8nX/Dx06nEx5rW47P3
u7UBl/Vav5GzwWHKEDpD9S8k24XG8osZCka+Ec+EvYuXHb2E10MZ8+Ai8/BIAodQ
mDrE7al60ZVpnksTbj0Pws9BeR9LPcM2EhlGWZ/VA+TMd1AvgrWH+okMAp0LWR6V
VVUKkly8t9zujEJHzwzSXifWHrrn8CXCmQBYXgOJ+RbA4xiyUAyomdA5pok2NcOF
yi3euCkbH1M7VehQX0WL3p+bMuP3MNprZgEoiv+PChHE7l16eI7dooYb4tv9or5s
Nw/MwWXuyjquE4uoIZhw9ZMyiQjqK1Gq+iEONQGyi9iR/sXB1PBxEriZ6xNrNOvX
jESBaQmSe+qW4GtlQtMs9BV6K45e12NGCxzRxF8qISUhJqjkpjD493Se3dsvVVkJ
YtqV5a2FVdbWp9LtA7QRaqU+nxSF16tPKovS92kxmYXx5R9I+nddtk0zoOxH+Px0
nhjCCPnQ3JAiV26qqVimGPbhdRH7fDaP/MFGOieAXaSNuvDZX0nQphIGHcXvNfHS
9jgcx+aAp5jum/UkClD8vfYxZDH7Unl9pN4CzbfKohrgHSy7q4M7bP0155XYMrZO
x5KlNRkmXdTtovcyPjcdwjAmJKHmLj6Y7+YgicfootKNESMLTQFYHhVrt1aPiuUd
PUUoUHlXPgkmMlKp/XGPhjdvLKtGVWFC6w8ixMxR947r2TpVvPGW42ZMuWwLy31M
62T5mybSktpFxvmu0TubWO/XUpg1spsytyAchwVomNtMFUsi4ED+zPlV00U/I6TD
BOg+34mn6GVP159/xgbOda3tcn0xbLfj9YFaJUp8i2bpa8yJvuJK8qVtypwnd4l8
vq68FftR7F2QMRJ1JC61Y9LiU6TSWYnNWVWnFaOLNlnY3g4Yn08TD9BrDHbHFr1m
vuj3LqYfuIXldcoOnzCPRQvpoPlVabzrqK2M1SnBqoJBWpLppqUz0V3TIO2B08xr
25tVFSGaPJLYtCurGmtJh5aVe+CH527nfZOZZrfLDOzCuUpji046e/AiI3n/WcOv
qD7F2MZ3exjaLM0i64JPBXBfMEKiMH3b8dggQCzkzbm5zN+Xrs44zZ9XbqofJyrt
u3Y0Tj+jXQuO9Yo43w8M7GENwe5xZ+tXaQfSI+7BDbkKUfVaDJMKwX+lnjyT5jIr
/gAaZnmWzaUO2n3s1emOze+FjddfByo6tZbsJhO2NqqTLsMg5FUPoEAVys005jzR
M0tJKAdqjiCgje6l5ka8C9VFKPqx2FW0LlaJPfn7cINmAeGGsjHtLX6LM4bdsIiZ
K3GBdK96goHvHq78OGyYdpYGqdPBCUORkVgsgkfqAyHiQ+vfW7AK5c/l2AShNwEf
/7eseyZbYsKcxco/8LzrfXLAImGtlhE8hTFyBPS/4oN+fOmG4YV8kRoE7nzsysU1
5Hx3r50uaxTBefa9/LVPUee7fIobzrODJ4BIRbzC1UjOfBGClPj0Qk1OW2KWeSfh
tPzlndH5kbSZ88ICROwb9c53XB5YrPfOpNAs73GuZaAY1Di85nsqrO+49nc/ufNa
msPwZqxxlmtGU41lMShWfOyVrRedM6LZ/iEFh8dd0e5mQSgGltptdS3pQNARm428
il6rRFbAQ7nLh/hMqoWKyas1CxSHW70S/5gvTNX45MTBuue+0gKkQ7/bBdVredO9
/y8C0wwa8nTCbFl/9MT411SAuntKQiP7mY+aPw1u3VmMvstyYfxTyvT+bIXHOmER
kfMkcBiXiM7NJg9anOTZ9vWYYFieFUfVUovejArQo+gSzvKQ3uPS4BwCIzduY1GF
zLigTvZQ1O5nza/eVeKk0FprxTVw9hrV4cySJ9eqrZPdRO809UW4tpuYHjO5ZYvY
KGEPTToLFApbYla60wXcM5+WsZGaCdfRm9KaHQMmXEtU7UY4vlQFMS8njGJfeCrX
8e9vpJrtldLaMBQadxEMHwdDsBBtOBzPdwO1eaYSRccI4q1Q6vIkOhIwcCVyvWil
E2dNujqUqxD7rGB1TKlpGlWJrOU2eTJZjom3Pv4dC8DwqbZEI9UJVo0nRY3jJHm8
NZJ+GrCX/OxasWpA4yJnD1mt0++A0U3qgGtAZ7QdumFk2oziSpza3N9ldn/huA6U
wIztk4izoRRJC+YvvZ+eVEua5FEd5YGVA36UFgPYAmSqioYOdOw2tj4lG1LOj7xV
LRBcQ+ZQTwqZXbtbfqZ72CA9uiauLgxVjPl1crMzw+Ak6oryPQHAlLBQnfpx8PjW
qsBSOfdCvSdJsKA5kYBjhsmT7XsCLlBbe8AU23uSF3Uvc3KU0/cP4kI1E1AX7r9M
nkaYiqqoXyeBNwhIPFFjXf91o/2T4sbPcglFEt8fDIRu9aD3p1trTfNuf36Y2fJT
gQeq/QU7jgACKLtcEV9kDCsUmlaau3WFseaObudJ0Y9pjQX9LeMIQnenv4VmGFjx
+ORADaGMXj4CZYrOx6yoccjmaBvgVApheEYsd05JETuHi/4/ZjZJNvdGGEZxOjSa
LO4rfJ5bN0c/3fygzO0MG/kf7yPnAoZS793J9e8rR1l0tJL67yX6iVRhV3QHLuro
Q1MWB0VBXJEI17cYRDeFhR9gkxQqv8H4MWyJWKfwkkbVgwk3C+HKVm5WZZpBZI6j
yR13QlhuCFDWCGLjxUlyv6anTJaxb1upHAcCH/Gx/WN8QRfYsaPtm5zNhDOdJ+dn
icaOTDzzsp0kOFSLXubV9YPzjADQxiWqPZTQaZ+vIQKa/YjnQn8T9sx5PSsPM74q
z1gQaGIy07VE3ioq8crsxCt6mySwIBTo2n2Hx9icdWIki0b5Adi6jri92xnL4NjS
E4lAvKeYjO6zgDx7qzbSJ0tnBM6bOGenOP4M0F1FXPh7ccdEoYYezibIzpx/SEeL
TqUAcpx/lwz9vBHbE4HlUbg28pyJCkGwlsZedmVWIR5BySjpUoVtrfTr6pYz+Pma
Rrp5DZpJyZAN64Mu3tf0YuSlYJVw330DD3uH5Vzr2lCz85gDNB8WCRv2WuigiZB+
5gySPewTWU3toMK/ZabPG/nheeSHp5MYEvOt2Hx7rNbhp/K5I7KIviFEU4EK0huy
OdFgimOfjvEvjNrYM+hTy1IAWkGg2owRVeNz6RojvzFOIhebEQEYACLl2hCP7SB/
BNKF47NGuJFbRTMpz1UfvdFrC363Bq/zokHxB1bdja/sbljCjVyp3VCwrOQJogbk
qyYSr2FPlU1gjydYYz809CCYlWS5GTxjmfPqsqw0JrajWI1+MtzAYVDG5APLPB7A
0gtMHX5/mPrHkEiH7XEwXHCpzahqJyG3MohVuXoXpXDu5Bg8z4WAuBtNZcSK8zZF
5t+aOIoAiOrXAjKhk/W37HC45330aOpPaAcRWO1rzZewJRF8jXznB9t31l5Z+uou
sYKcL8YDkddRry0q6Vb4TE25yT4m/3DTd0i4wtz4xVHNV+daCZP7U7A3HKbg39xH
ASxMtJ0OyAboH9DQi38cIlEMulEukCyYC40eOo0Gzr/wiMs6tFmeqie6D0Ehq9gO
cN/UT8irIDyC3tUot98FA1bcdZvoJuMVSNNTikrZr4o2UAPVTkmKIoy/lSZ6eLh8
wd9LVVWFzPHQt8ptbRMyJSnb6BwY+W1jxuud/J9LTb7NtHw/e7w0aNdBachX8dPy
fo5hIFkRGGoYezlavxtiHQMqyN4LhPbFoWUNOaWhNR++AkegfVRk3Bi9cEwSP8zx
Pv7eNic9iXS7e3WZjphGX8Wi2nQ29i/+41YUWupOai72JCxQLHxyrmE2TbuRjQtJ
h9YTyvf3BTVsPkg+GMt8RQ03hZb06ItJaz2NKSlicZjl+nm3b4RRGH6XLCabC0Ha
O02XvipWuEWI46jEabhdeLdUg+uB17awu/NqY+08ZfWS7F6YwPMCc6bJG76MuHXJ
RJvFnys2/zwmofP8YUdXDxASY7XfPIkQqOvdlbLzqcw5dHqgiB4RoEwZmn+vD8dc
K73Q1XxBJWI1WioCoZUSBbIbiYkS6ZmcywelHgnKeP3JQicOcvYwsTJOLtATPQMp
w8vKWef4XoMSv6B5GdmQgATqDeDW20Hukh5SQQJwIzAnod5cXvSDlTpwbG2yr4nx
RbzXHNo2EzNVUs2JbVVnftnPT+85nnye3Tqgum8pCCreq3AleuNur5fHq2Zw29E7
+4C/nnO+VUZwYJM3YKFq6VFWvK6eyUzVigcNB4mEMZSkV4AlCqMr6PIeMU5Cxs9+
YsDKAfIPq4Evfcn1VDq8Q1sJnDwsXLCSP0ATImAqCVc07MtG/xN89iZ3rK0kDdj/
+wyGT9/UzI5O21mmlEe7+QWh63r86hhj1I7Razhy6G6T9kLHOJa5oBmQIahIuyXd
/tITdrLJiuAULKNIkLCATOZcoTqTdahBzFsICpp+7Iy/q2rLN5PeTFuw+CjZX1ab
5r+mFBl5GTxCE+iLpbo9dtd323yK7xioJEi1TiHU5EORb+jY+nziobS+9DRczCUh
zWJndjVyPZoPKkGil+XtbUAbQTispod2E/tlvYAX1jaZIdmBzghAYVwIIToypzpN
ghxlCotZOgo+QfNd79/RVi4UTRBIc1LRQbE+cbfIzzvJ3+bb1wh2cPZ8yBMlpLPM
Xqe6jdUH6+Xl6KGzRSBZyXuY+BaZFkeSw3QXc77MPrwiQJdgqmZbYSqNnK1xMpRt
lQixK7JjP6uToZP2EhrfZXUjEPTtTM88Gycl0bOBV99myBgeMIveEAKzRpJWqBOl
jItxKVoPpo/Ea32/3FDsNQqfQmAVQJpMcg5eeVvCOZlninBWFMX25yawTFuzocqp
sBZfU1IK2ADXOAkCN8MKKMFfKJrqGNOzuUBRe7Ujs5IEw2OLcNKKfdleWLzmIuvf
ILNWTAaATGejGXsAuGtrVTxHScBR33TAFro+T/V6R4A0bS50GCzkUQCuidWd2ng/
JAiAg3fmh53FNe3AwXYp+0AUUu31cbdrt4oOmkYc2LMkdsr6sZnUfZIfdI4PnO6q
VvNiA1u7e07zRWerrHLhAfR70FQ9MYke8GC9PBElZN4v5nt334H+yVZ/W7NX66nn
UlHFaEMtqTc59LwlpUiYaR1GhYvCjiSX658YsSF1lp0sieNig3k61NFwO80zuKmD
KUezlhX7VNIhcyeQe67oGp+6TcLCP71msOyNOS1VqH51LKEEBeg3qWCx1MiMxBWG
4rlYqFVHqVxog+dtB32w9P4KX8+0tOXpmNdE6Hm04WXwCTVhnX/qmSwhHYVYp+Vn
GpXn3/Z16TXl8f2tVv2MCyo2jlU0bGyhdaRWg45ahQ8+8TzIIw6FHWIM3m4QX/Pq
q8sm5X+BNspAqjG+xcMIo+mrN66wPzEdvOAtn/yCmAVRua47rVfBq6cZk3ApBA1s
PFLv1tJohSXqxhSepbfqmz/4wwShLdBy4lxoxGBMpeJankDNv1MYEcjkgdj5q4oX
2rhoC4GgaTtucNtTRoudzbLIFQKhmCWm/+QyHNcUtyuA/tMNexrAK09h0crJD4Z1
`pragma protect end_protected
