// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:42 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H56rvo+YczWhlkBh/Tc6N1/KJwB59aFsOq8J9AsY2UmkL6vDHap+0Vm3Ha1xr/CQ
NgJe8E2PVaWtLRaTgZ1K64AuvMgWd0wxeNzzVGzJeIgkHljj05sEYIwFaNQB8VGx
JSoo34/Za49loRqsL5UZP+JsraPau7l0mfjnhElP9uk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22448)
yZsePSiTPzI6R3pvgRAhfYuHaEbHuS+3g2W7n8O1syP5UegslBqt70IHEUZtCTCO
PX4lEqkHXDyxb2bS/rLy7X2hXubPMi7YLKtr8NWG621PCW2YWdUuxp7UGLAW1kKU
Fl/Ay3xCTCAUTWCMb4Q/OXWr/h0w6nI4OmjT0ch10ZSo1fU7pXZol6srOFbbnO8B
674XBkeicdzN7AV8ackQ43NLKC4WCmLfzv0QsOex+MWHmirgb41QUmmfb2tekyGY
0zbPS+vIhhKlOFMMji7E4eT70IiEMoENlQqvWkvoIayGUm98fmofjPHzrIjXbWxZ
5oB1Q5DuZrlwzo8AP7OadRKR3v7NYSfxORG2MstSK64s9W4yBJE0WpGFno4cpJ0U
9Sb4zbMgzgez951xCaXZBOYVVCpNxlLacpKaGoLpyuGY/7BadiuHZ2/WPA1fEE1x
SN13ofr/yZ/GS74iwmqBcL1rD0MV2N2D7UPkxL/ql2ccXrPUMI9ld7TJOHhBZRWt
mKp1vpkUrxxRaESFz4dQnr2zppTt3EK3AK7RPiQM85qrQUj0pA4j4Bo2p87UEFl/
sHPMSyU0rng4Uz/iAOyc2JWb0EVi+c7n1L2QyGy/vp2LBP2QeH+OC5AcHhFfUmDn
N4AGp1FhHKhc/u3CVochysnGWsccWfKaxWz9tr672I54jUL7YtyAk47/Kcyy/gV8
ewmriNRY6Df5x+nkux7QmL73nxQn/s8fR7byFmLB88Beu6LOVIgk6k3W74qshS4H
lCHrMWjSDn2LHAztkTDC4ly2Y6LiPfaUSe524U8o2l1Drg4SAth56ksJ9gksF0QF
eWyctNSIhdTrM232rhxwjggC6NFNtoBg/3QOTtR0pOTcgfPBBxPMLqx7QoQrtbdK
JLgpuec5X6QTtqtFZ7kyocwD6/7o2UzA/jCSZds/vM5gcPp7u57c9NUE1XKwIw+/
ZaZnJMJsKShwSt9DeoEbaR9L3TjQpV7IMbH3Z3xLhyL8lM7RK5LUzIZ/xJlD1WWJ
rWUxyVEU44HkaPA/PZZeaF+Ir/SE3+d6krag1PX4k8T0Z0abCbXq6gzEVNeF8O3I
0DUKPBIw8muUEtQrtWLRQe4QuYOPqvucr32za+7gwyOC8ra9k+eVoJBS1WmKz1MO
aJo9RnXMuQhJMrMxPWpbbt2G6x4OBG4f5pK6N/mt7fH74MpkutCzsyGCfnJcR0uT
SVJ3UxBSvZQ6zs5PD5uDKsGJn3j5jiwbuiloXU4RDk+NNfdNjdHj3kmMGrCgdDmm
hQSaHkyztDhFnEeDzMuvWXUtUT7HI6k1xzfFH834tL+YFH5Aaetwzy6GCWrLR2Js
Bm57aJEaIffHChOt07ZF8Gsc0jlOl7bv+V7mjmcWA6hEGU7Jt80lYu5cx9UYV4Uv
X3ZF8hvQO+YaaFHlExJ3UjsWepaomBiR6EI/uZHi4SIq1dBy2q3x/XvIf4c4pLoo
U3qaD4FampeMW5qf4/ntBNzMpjwH38/v1n2On2EEF1atQUKMWvByLXt0EmE/qRZE
NbyXq/tl2au1cCqkelpObF0QzYCxzE0WtsFZmxvGYyc4g8lRF7XSyp0uBa1AngHR
nhw3CPtF/2ihHKBJ3njVvE8yhg9cld+QJ0iVV+mNWLKTrOEqn/qtZFaC5AONGhGy
S7+uZ37j7//c4Yt086AFiqbYYV/tCSKJHhAQmlkS/+/8ZDgj4T6a41PCiPxwqMFy
9zysH32OsQwomRbzwO5QgrC55sx5KzL1BeMCPg0NHyrQJj3Qb3+T59L2F1ER7d9+
jWF3GkyrwloWm/JoN/KgjQ60FKT9uq1tnwhzYLtc7OsZjc3GAu1iJqxt5Q5+vaAb
R+adOV0+WXIzRhKk3WcDc76WrhnIEzvKwqB+Xc1DERh0mTvk7p5LF9AezK6/zTXo
HX1Acr7to/WNJBLVbmL7YSjg1GqTbH654LfuNMI7r71NF/ADT/H+LEX8+tJrpwlz
31x9YCTgT1uCXaQgjzM/JE1kw8ti6JNpnCyzCwjuRVnI0M1+I2VJlHyWs0vvYeGn
Jw9yc+MTzV0XNztAWjnXSiqmU3Oe8Pf0on7xjGCstVhTb97R2cBkuMX7YsJV5fsi
WXjQrBsB8Y0SeaScfr9Uyd0WmuPk80sKDVonfeoCL0z2fq0c6L6Aqgr2TykrWhzU
nPSary4oweVJRzWogSDYuy2FTQLxIvsNDxJFFMuWEqc2vMcVyf4RuSNVi2Aaf9SG
XemtTa3pT4xg20VdFU9aCQsAR1g6dXJBOoIGyXqRYLA0JYOcd68T0e0i0JExmG7X
B8CUmBKTsHBAxqYIgXKOU0ycc5VPZ0CITCtBqSbGeWHuhK3unq1105SEmd6R7QwR
dOC+aWcBSypyArxLFRKY5GB4lQL88gdcp1wqIXr7M4ch4yWO3GTvpfsG2Uh+01Q2
x52ja6HvJi32WYBvPwi+FpElRcmIzebjmDb26sUOyr7YL8mTxxEeI0bwNzwSXAf/
8QZUcoaUMNiaaVOWCHiyH9GevkDRq6c83ZIheTtd00m6//DNMOni7CuYq0rYvomB
V42lxQFIwrnsacO7Pt3+UJQ5TCDmMfQQisOwSmPZdsNcywitJN01wV4Cfwh7w7Zh
g/fO0eZdp2vh6ckcS57gfTbJpWeFmOFqgnCfATqm37+kw4fvk9fxSTcDh/2jbMu/
ciXFr64UnGi+Xg5D6JBzKN6XN+ZMaPfbtSPaTbKea2cQ0+NbkV6qzIGiwiib64QB
2rY34S2qBOeV1fQ97O7KVCDgRVAyv2BzRytNkkf2bU4taafw54s1CZZpFizrMOHM
MJ9RGva4LN4btCiE9wQXR7kXGhMGheTWNdQ2ZbDUs094BZCy0jo454zxqymX+nxz
QuQH56mCbLUxhREo7kNfbzVCz05OzbXdpR8MYjM2cMQ7ETKbB3rGOrkzEgs2hCzo
vjaMtKRFh4qZ96AXSooOA8ick0B4Ge3/ANTP7p5u6toz4V5hK5D89C/rS1/HxbeB
BiFujRayAgKYUz/36ENdPtIIUSApk+pzhAvTLH+UUXqfoGoEnpf6C3VhOR+r2BN8
zhxfEAAYJiJDaWgymHbbBA9Bvngj6VdbYfNGQPCyMO8nXCcAhvciyHFL7RNhb7iZ
RAqvdd0STGAqdsgqEOImIV0Wmf7EaltrDEMwb1IrJPJYAXA50mhNBAIfpebGosfa
npU8bRoA0apr3XTtssVwGojl5tKtzyd7F5PqfBhT948bQuVw5dPtK/UjAg8RjMHv
Lzk5GU3QRbDH9P+u8L7R2QU3QIOh6pGgC21PQKLou3CHZTwe2QGlnH66eMC8hCCa
D3b96RvR865fpkReC5errlvyfMFeoQ1hGf3jlZzJSKA5UVHpm1/6o4mz/NMxfcG1
iLWo4dsrKREyWcJFFVmct5dZzXfDPD4HcuAQMFSyHzK/G6LAWHG/eioXMj6P3gmw
V4Gb6Zk9UTiruaHnu29zy8BPUzN+Yl3DAU46Vp6iJyxHqjbxu5RWYBYKIprzRJRH
aTTmP+RSH3F0OZHy3FsHvPLQd2wNFqKGfJPywxQ9XR35iZWLKAFh+IF+LBl+8PLe
0EfYWviEr0mguLM/VhlUbGZDK0YeZBV2Hnhtu1MD9kdTxGnzlUH2NmMAt4xWGV+x
F1BRXOQ0rP85RJpD3NELkEHyDJOJDBhtvMIorFk9XRJe4vjpvq2gI/k10+mKCIpZ
CYNYCIy6COZyYVyyQAy9aKa8CBgYiPvgdwciTUQBFXPY2I3fqMce95c0BaFBt3l5
EmSglUvnIHSXSkI8EmAXcNwL2R7wkMmbfbBet5OwkfW5uGysLe/noTW8VLOKXjUJ
16wLcOFLFtafYF3QH8g01b/kGmBNtBr6TkYF7gZtgRowloYLKwXp0eNJSXnv8tQF
sokpFniK7BqC8gi9mxishQScdMF2siAMYPQTXRU1YbAA+ReIac73cH6Q1JstE4Oj
Kd7QD+3f/AS2RgXJHzHNpQ8jG30r1mzcwdJdPmzZv9dxwwI/iQ7Tq8+gliDZfHSs
wRcHcFjDBlBaYQeyFV+K79/XkMVoE0OfAHcdbkyGcMyFr5JmVhB/5XwgNrNN7n83
GVKM5kT2B1U5mgQLfoeCAgY+40+XMjjEeKjNutOjAwuwbym02fHtneB1KAu5bfmm
5opcZ4dozfSQkk/9rvwpoW8TgXfXNxJlDbQYl8uuy6ZHGIVE9jXMRTjbS7C1Ze+M
cOa4F+8v8lTOsP0/Z+53pi+THSLq+Ck9dKRMehfo3n0PR7cwA/Q2TbDZivyLVK4v
m2qKcYqGsVEVXbdxHEdtQHXtaH9QoX75KnJIx5ezbJ9nyWBrfhtijB+22+OIhYQF
29uQlM2ntE0aagy26th0FZV66nl5FgMWqqI+H7XChGXJN/6MSHMn531/Ytb+aJYZ
pqA4jPskkQR2Jh18c9l4vKWDXQLI2Rr65vF4q4FRw3ATQlODj8uFnjthWt4jthmx
uwxfsyXHvbsT1jpHb4UIRgwIbxcq2hrm1ECNZOrwFRtar6hp6AvrkLIs3GVHtWKj
4rxTDZh/hccqqRf3vgMuo7D73JFBnuhOFp5S582WC9Db/TGv1lMqK97Hc8Qq2f/j
igPo+JYB4PQb3IuUmMROV+I0XohFHmuZt0gTi+IZdhzfS1QPmPTEDMMXcITRwgLM
eW/iimAPFAYVUyLzJ77Fv1aXLFEjw0taDO7NH35XCIESvUMv3AFh9Z80P+gZl7M/
N7BMGUdvfq1wTeBVxTAdvxCDnhwHdG+wyxsvILGKWCrzrTS/rn7rx9xixpDLKyuv
U15uJNKngeUVqfieKJzYum7buA6PGRg7JJWrGoV0iBmZQjxBxmgtH6354efhgiw5
JPp+z38Iqq1gX82k5mWyxI1yF4K/wXOgdbohbj4X/6fI6CrytP15/nOisxogW+Ak
io/YED9Z/XtOnsbWoWj0+gvYeskyu6Qey2gygHHSdL0KWprJc60o7vXFnBU9NwDo
pXB6gItzwGqBWx14KhPzCJ2YWlj3aN6b/h/el3FTiQaEGaGlpvO0Id9nX4//rVEY
AfJpuZ+Fym+ul/Bb+B6WHt6xUB42De1ShnbEnFTd3j8szRcz8B/fpbz8a+H9VWUM
VfuSuDEEG4y+SCfz5OLVxXF69O7W96SuWMPKEk0GKzXrE/GHnW4xzN3jzyaZNz67
ZRGZh9fAfiaUcQEzPDrSnaYkQGx5loBfuNe/Asdfr88LjrnDPYFZu8e25FPKGulj
2yu6JkVnIkInzgndbiE4ZCewAVq5hfuZPXiy9axrQliuBRA/7KK67KHmd7RDHuen
nv4Z2d3oqubKMqhArCmjbNqp4dkVmy1sAjkWzzgkwrPRCZeqt649LwHOf+O4mOCe
wjYsA9HOzkCoBdn1ZyFFs4ETYEiniHSoKvK7cGuBDUgtvWeZTSIsHpDTOQ0eAAzq
U8a+XK4nPBrVcZdAgvmmEyyqlljjZLHEb5iZB8BIVVtTDJsQS6l0rBXGcLPydrMb
ghnnS/3IZqD5yyDsvdnATG6ySAV4ZVX7qNw8qMT/oYjyCInKdW8k4eXvc/RJGNMP
02bXLqRC0s+ojYEcAXrcFs/XpVdRX/uo2GpkWOTVXPMeH6qwDwLMfsXqBtZQMP0H
lraQY42B7WEBXqg99HxDpE0bSBYzHSww3ZqdAtgknUy6Zg2wV8cLZVKLza9swvPg
LgCS669Vf1V6CkFVRjQSR9sprajwA+CBN5ciIa64cuYxMZFck9EL1EjFqUT+yP34
DYDoyG6peii5QiDkMTeHNko9e9NgoHNabF5yk69wR3u+P77A2epEnAtsrtO8NVMJ
nuONQDv97WlzPnettQ+JYwuj5B0g7Jk4zTmf8GHdX6IW6hOifJ51vsFRaMvlreCH
6tdPn0keCE1Ie2OthzfpJQaXrYQ6ovXAFpd86CWO/fqJxDb5bCVbZYS4IqwdkTy1
QwKFJXv2Rg/caf8DF8ibffhditR/jRS+fHuIDKovVhiv8/FDt+3M5tf+aLEyhv7d
4lpj36CqNT2G35BkFiNS/bQLZt6FRmTNsRqeZSkc6QAc0w1OrGw8jJA+oqpcdtgz
lK99+Z202ZtuT2yBt7fnbKpKPnO+81f7pE6tVhE10t80UEPPtl4ZRbYPtAOBZtek
lyUVm4RrqXyIX9NRtOeydZW1fT6+yYbhO8IBSTWDPtTzN3gcLJVrFf8/pAnkN2BS
5mrEZRW4PrXGzB8c2r+sNDh/sooR93/Fzs4mPbBIb6u4QQEsasU/s92w28kUSVJC
CbPES+3aE2CM5P/BuAnhEqBCSmvjxbBPcVDTmWg/R2yXbboHGoEwxCWAWa1sZ/+z
gg8dRDgGesXFiATYuZ3O4bLmQwpA/49Pjp4deNKMF74PFpYcQHdgl2csGZyBWkp9
7IZQFoHQYE/z9KnZ5or8j8XCg4Mz3TPcHpYpw6OpQ5lruXjU1Y8AJ95RNqjfzdq/
K5FKrxl88NA4sDU3MOigLM6nnzYURs+Bq1VWsnJFvs/3tCSlEAzbSY6fvbxx7/oG
Ey4TXp0oRjGr7JYPXydXvsb/qhT4DzWZl8reFQ8BxKiFejW9O8Gbl039WCPwO00q
5G8Um/R/YI0OXo83eF0L8/7GFj0wTV2Ssz55EyZXudSyI45SWqCAjDSm0PT66BJ3
ZARchqm2NodF27UAqWinagYAsCxql2tIkEz5VRq3qRgS/FCic7iVVG/ZHXr1BWUQ
zj9oJDWo9sIoknRwQ44R+pLCu0SnvXCHHVWCdoGMGewJdOfEmQuzRtXiUFzpHl/U
fBcHLvX0b1CZKJfqE4LZtcerNwyYRO4x/zNCypLti5Lywehvi089DGNWmA3mFUwN
LLyMuBCmXPfUYaSdmSZCZLjmxeHumKIyaqR1lprphpo4SC1TH0PUbluwC+XAtCTF
CMimJ+De6qiol6+/TeGqLYNFLLHqw4gMQMv+T5kzcNGY+YpJg9CwlIQN20IHLmJn
65sY2XQ/5nxplBTOl89KE5w8JYt0VX05utHWUZAiqJ3uLImPLCSRiQIzBhpEeT0I
fCqkUJL6K+kGIkzTORipyDoW30AQB/USganC2Kfey6G4GqjuQefx7AKXP0aBt6ix
C/fKzZiSOldqchsmCp3jmhtbNzIHvSc6Z1qGrwrprnG3dTOuGoQen3anCtWmSH5U
+DZcr5F5i4JBS8LX9eCKeEGMD4vB7M36OSB9N6tn5n64VHRBj3BCHRrH9RF1vF7T
8QQ5Vx9Fmho6rs9OU/T6TlhThhp9bc4rpUuCNeOr0aY7Wm9q6Nb39WjOs8mg4uRy
8P4/wPuXU4H5TL1iFWwD3anHtGeGAt+ZxZ10Pox6SNhtFFz3H6SZ2GR6dv5xHoFd
XwMgnMEa9IbqaMgCFRs5fPjhTi6/96Wg5/a35MTwpVkf1b8YxQ0FBf+1vcSKN0vO
X5u5Cz63vRlK5pVdgBghGu4thw8H7UZIfpAIMYI4xxk+76Et9jDQ0LvrWmF2K7zy
4W12euwrSiC3t8yZiTqUYSaH9WXrDu9PWuseIiUYtU5SBza16oYAU5iotf631xOV
3RJ0mlL5guDjdumcqttyg/2YDv1sA7jic6EEp7+qR889TWTLIjcNCWIYLWJddMOK
GfnZZ6S7N4YswV6z+JRxqQTlphSbBAv11OvfA5rzo8BuOzKYS/XYTM/NbjB/8JA/
38NNDG00ZhL0BSackmTxabz5AruveKC4sgTDxRv/Cb6mX+H0FE3rs5smDkhMo0Rn
Bs/8r/+Ryk2elCkE2tp8R2lx9zZ0T0IenzPjILYZQxaEApbztKiDIX4L3WrBXV1C
n7kVJvX22tFt5+TJkBksBYXilwvERHPbPg+PbhkkmnAf4MFhR0k5ZG1yg+aa9Qeo
XEc8Vlc5Z527T/Cj8ar9w0NxYYPKz1AG11VpOotIdpIw3yUW+69C7qcDU02qb2HY
ramoih7nMFcpckNPeyY4so9g8h62XA+qXGwTRAPlHgBesa0zMraXUGpt+dP3/acy
2NnhAvKxHFsffnjs/x257ABtP3W/COb3TbLyvWZ0+/bosRrltvcAwQw5C85RtWqr
tYTKMx/kESTJpxZUFQ0ij/6n/5t3o3hPLbvokQ4jqHXyX3QacUa0R8VJcQNmWMIG
2GyIdxToaBPCcAkxv5KqsAmB4aGZabr4PjmkV9wu+FPDlCgV+6rsGoX+Z93nW63e
GWMmdmrX2iT6rCvs3h/szZMNQslVwDgJJlVPXj0O122cP4CqUkrBs1A3C81URBkj
oqydeNjtOkDNooSfUZHtmQyBSuC6tGKeI/CjEgdaqHGAQL0mhflaTMKSDVDMQmrE
/O+IFSGiLPyg4to1PBw44UOZVfoAaYAvgZMXbibh69HL/gsle46SJeqMw+Op6bmq
gYPV1Kvkl3FoRhjgpC76Ix6htYz6FCC63oqxPZ80rZIwCLUWclIRkO1SFiE1Lu23
i3N5/QWaBxsKrI6XGA44cDrbu9LsG4cy2p/f5V29aPEpiZXqmvN4N8Wri85zAIW/
mun2GHjECGhHX9LeX7xLKDNxxgAAP9/zDj5mhJiJqeAe0tc2AA5EF9rKrtO7wiD2
FF1iw5QB+hh4FUVOVpvMVxL976jYviQyhs/7yqHimTFjlnLg6c5Jod1VBOrWGdVE
pi4adg2QTLKTuM+3YFWwC79omjc8GZM9QKPTyjdYVUVzAS76tpYGf2tKfghG9+lD
3iY3xYE0XehxzG73zGs2zXXYnZzqyjqXvcisM8xSdVfzvYHVvfejRmdcVRTqwAyG
z+HuAThRrLWHx4BzEIg4Z4n6SH+sq3hhicoh9y8LcjhS9XKt+nsxgW3US/n6oF9y
CTBXhJgtMCSbXYltFNpRqL5fvlYNWb3DuAIN6SPIMwKE/N4Hc7k+ZY6Ot33io3fB
ST8gl1wYXlT3mkAmF/4L7nRl7JhwbuThdzzuqUS9GruajEWwsQHEcc4NKaZIJyR3
8xrGv70f859HhSeuDh/N/sbfwtcHxF5eLRt4h8eK5yQlp5cN+JsQqR75c3RgXTVV
G/ArbybRCIMrS9Ngc3Ju9AmsW+ibQhnC/pesAiMvG/usAyCDU8Hn3AS78oS/VnCr
/okW9W610UorpwHyGSkcF/rDN7Ov9dJPcZPmkYcGduV8vTdSN+JL1Rn8qVYqgeZi
QkuWWKXPvQeL46vrPZOLm4LhiW4OTcTfOC5mO1zlVxD0gt0gueBA3FDFnnHwVxSu
PgDttkWFbj8WvWYi3pg/U5bIHYhNIq9yyGT0CM3NYFpxkr8HBE5uJyhkQ2J0B0sq
DX1hJMF0c1MBc6KX17OYcur1n+bcezp7pHlOkojDKApLlr04JbYgaW+lfLqkbJ5w
XW+GskeCO8HNtzvJcZd08dAbTV0ihAS7N2p1g4/iqSMkCeRZd7l9tSLEAMn/aAP5
uUw4zECmxbOxXn5vz/A3fTsel/BVoEIbp28Sx7lo7eyojVJH/HiEUEFwbOabeu44
S+FT8GXbYmyaQPK4ZuAqriYCDcH9+9gH7jucsf/SjMyZ775jfklTjrAO7LOtCBsD
aSWW8yjD3XjYZE8qLAWsmNHIoFXl+xjacsF0Q8w0CEO4pzx6TKPlK60iRtCv4urK
3Fz6D8ph2bY2z5eWu69sJuBtgZ2npmUuNEvFtrsEFxhAws9002vl75+ZeOY7E0qy
XaXMYoO19kwpckneuKYV/T7l3h6ZT9awT7nqPWxfwHl9Dns14pS7qLPPL7OHPOeI
Cki3/JjpniMRcSsPQBRrPZWS112C1h0fW8H3KWREMvQYjmA0piRG3FDKg/YciPn7
S52dontZ0pL/emCOrqRy4BkFUe/M31VJDS/eW/AsZHf4AC1EutAW22lWr7WM6jkX
dtz6xWtNgHwmrV7YNbuBbHo7yRcRdfK+VfFFJZ5P7ZNN9IuU09UIqSZmsbkATzOu
LsHCVsYBJaYNlKlIEfDOEnNXddfFtILs0hIfuohbOXbVtNC9Laico0pZGU+oP9vr
gilm+7uYb4iOZU7xNDswuyH3uVC1M/aCgYRP7JiTOsti9hhj6ZadzHNE7tRa4MZ/
pUJBOdYKp4BWxn0PyubQd5CICGnSPH3+60+wXHKyXcx0wgjIzKJXWbLbyx3hO1Sd
n5mNxNz3P1A4TNeq+inrcT9zvCkWZURhSixYlaOghJyOFEEkwIPzI080nu/Mkoxi
lQEYyLLo3uAwn527nDgIl2drwMXAUiXat58aFz5sfc8vD/ODug22R9GM9F4IThHQ
jRvjcw7e6S7BVRP3P4a8ir490vCHkJBUCcVx/OyXrlAli0DfYzFPacHXgjtotEJg
/AOTNLwuUMcaM6pT0z5gtBMdn8A0gO/yrRiBsiKhfuSbwgnIy7kzDUmGmYraB98Q
MoaLiLCCnPCvy34z4oMoF2lzvizu34JSiVRd4KwQcnamFaCp5QsXfourKx2D5e8A
yKqsC7uUmodzF9LWUztcruVPl2d0jkLZ350J+3oBMGnpAx1B0hFixiUSuNfvB5VT
sTiNNpLvst+o5gI+TkwAoIsBMy1SVJ4i/mHAI/Tj6S7Cd7tyL0a7OHzrlgzQgUJR
Bh5m6E7rZ5FQFlf2QJbAaiH0WU6fyJAE2/KbDdeG83FKVaAiiKVwNA+ZEl2Ilw6e
eMH6qAbvEkYpI1h9WqA73CcyBTMoXgieAdqQOBDxI1uE4wtetLD7Up+eeOrgrz+u
Em5xg3j7q7fjbn2flhQVXlT0aB5J6juEOEoQBBGjRbsPVHYY8WtYpmvdCQbWT9AL
evtlq5xLjHj5kd2JzsIa69hpA2BW6QGnLL1RVB8ClmtIOUeY370UsDjHI0q83bRv
byPPGyO5KM46Z/6L4bRJoqXzelg1t0xB8TQGVsfkEmzDNqO/E1xSyZBOZYNoi6c8
LIRaDmdHIJY/XHdq4ORgF9jC/AEofc9gxPMoI7coSin3Skp1p8dNnpyXyfWqMn7Z
z5/eJ3ajm6NQj+oCp4NyJUkhIRzVCwLBeoNYIbqqa8LIT2ChjMwwA03uJcOEJRD2
eDseCQpLbRsiyQML5+NfotM20zdm1Zi1Sb83CYx6rzSn0LhBDSfd4RMop0JdN2UH
GKlki584QkI6nybR4UY1WJhthSxI5VMcyzM03RRYgT5rpS4kSEqVYR6Q1Ao9tpe6
wGJydeJTl0KC3Xh8i8aEhoeCw4y90ANO1plsZ+LD04ivv0g9UW2cjkAnlUA+97OC
l6Zo2pq+SHcTvITpFql1M/LA1miZ49pWtrnBjlcHtb00DDoaOX8R1ia/K5qiJzAW
4qwGCftbM/Y2SQXk6I/pXKhcZDMEYx062uUzUB5l71SytgMLAcLTu+08pcH3w0mk
0FjyhITWghyyXXyEdvVLTlvewCjKgGqL4558lipBDUeVjVYWu40e9ZSCPTXHWSDW
luUkKWEsmzTZRM/yqdxPuU5oBXZQrr1tLHuUMgpTYe1nQZguA29kz8u4j1fFZqxk
D5g/nSqtd4lTUTobcigQtN4I2s+2Xo06WEgrDBie3SLKlINYqOOJZIKeH5NzYtAn
72PuLst74+LpysLmlnKQXiK5Nxq53bbayO8rqG9ps/N8Zm/PTQu29x7vMWnmu9t/
H1Ze1J62G0iEkUmXVz2w1yv4FSJ/hpVltHVJ0AaKUhOA341bDFu6OPN7fcfAhAIS
kI6zLrAzBOSMnyrbCTydjq1JlxiwBeNcvkYtcu/He01lZnDPq74rgbco0i5Es6di
yYAiqWiXIeL9s5F7z/DQJs2MC8vuc6S6Ncl0hJPdWWvPqjh6Oj5/Xp2kxPkFNMZv
7WT0ZD26vAij23PZ+9nURocfWiu4uBD/BRFfJGz96ZozyYfY5+g553bQoWUwtOmA
cNfClAWHo4GDuW0QNwnuNurKMUW3ht3l823D5FNgHkIAtTTNXJ88nmb3aQElX6nO
l7/5QESNTkkmJ83czN1M15ez/REq/3E5nf03NQmHuszBPD2t5tFhqmk1tRXw/2ps
4U+NeUlKEo2k17uMPDUZWyaKaNT/yyxEiyq62RMC+uDSoyiDuzC/LIat4X+Sq9mC
MinYTwnd1HF7vzWUZbzGiHs1aopzVS67uylqC/Pwe1Qz48UlSv7V85qHAq2Xfcu7
vKXHKNddU8C5LSKhjrFZb/4gTPwUV9kw5bE8Po12h8rdGILDvECiyNXgXOhAt2KK
IQL5rhE1Q67zQCyowvbaROoyd8NybErZm7l6iAvW+zK1y86Rb/m1yX6ZlbkFmPPx
uaIXk0KPEUPuKX3uKW0VcMgHHq3EhAOSqNFG3qraiEhFiM+XM5cnhAVCxtQOVm6C
kpU+H431pKZVhQvdgFtXuW6E4ieS68+TYIkz4iMziP8pNH6Pk4TROU1oPhIJyqF9
vcsZoI/UoJcx4FXswU0ETZOnLgpu5g7hfAveayUJlqPCFAF0zBZY+yU6R4v3yOQA
5XnRNz1GvjvMUeSBFL4S971iPkKRADfPotb2wt9oWX55h2ljQ5bYnKb+a/tc7ImG
eClTZjCkWHucNBjHzf5rWqAG4johEUyePhLmoMJEb+p+duw0OI01S0Gpnc0XMkmW
jVvOS149mhhrz8eSPhYHx44v6chIWqJRfTbm2TSOxSETgYfBYOT0VD8WoIcqBATJ
mEJPLMmP0FWx/fedn8hqP8w0lE/JXO4qSqv8TdI2DcGX0htqMszx05HMlXODZoZD
kCaJa28Yi3Idh3uv79/Y0jpjr735QThxEta7d20g/125jcEa4yftbdbywBKBeZxh
HgWWt4bdlm89KpGATqQTdXGU5qby20LsdiOKD+s1r1ZeMIx3aUbfriGD6u9iipJT
hiV557+ybL+LPFzUntUJVPxbhn/McB7XsdbKK8pbty2Pl9NMZxHtMDZ/fSv13EPY
LHc7J3fchHoZ4NUdBq9UL913vpaDkKT1x4dJ0Bq9m7mXCLcCzx1XHr7nwEGIrT5/
u/xzvpPlsg8jovv9xwztmCsmCXKh42toqZvEUU8AaiHMaVxdZOtkSyzt7wALA+tb
Vo9ODZ9Scwff7+0yqbAqIYH1YKYZNqcPjENS4W6JNsCAFMm3Ieg/dHC8qTG5AfQb
61gN4AEHjhUGY/+9qy7GV8Wylu4vlURz+S17IvRygHp5B+hUk0yWOXqjgsQ+lc1n
QXHrjYEL0b+WeebifH7oSn9jAUtUcOJr8vIpS1e3XLVk96p8q9f97vrdLyQM83XZ
7ddt0O3R7OvZYKakh2g967WMbgAimft+QvIEQrD8zLbjFI5OebEg7OJVxa07D+7K
xU+qjTd9QLDxfei0PyM5/Fm6g8xNQdYg4eIJSbqNDMak4FcfCB55NASNAYZHsF+T
E0CYMH+9qi7MiYlJmSKCYcP0rbl2rrKxkEKfjEbfM8PZq5M+jrx0ExyC9nlkq1KA
eP4kx2q/YtvmF83xRS2Qj1juA2FO92MhjlSkMuvoeCYwb9PYpvMEG5Nrzc+be2Dz
CgiyDBSX9y6tC8XvWaH5OMmEQpb6A/6VNmAyALNZ67Vd6Mifwn82jPoRJweZNzCh
TJhoOQCXQHlftrUwuLiv9yFGHt6mjpr1L74MGa1kDs9kNwK//xkh8IoeAtsyiGzJ
5PBwEnQZFPkp/+oDfBkkO3/s4C996N56bIAUZjQnXkEkZnF+jMZ8LptK6tOkVcRE
xXVm4F/i2CBCXp98BO1NJNsb+SehlWg930zR+aKKJm4u5Ljfzc/ErG98jUPkxBuL
ikC+in5O86AbRnCs3EJtklMojpPFUyiP69OuoszWYF43WlPU4i3T9B1b5nntISo1
wxKDuu0xtU3HJC1s1E1oDAJ+6qOCp0tR1CwG+0QGBBgFBMsDZgCD8rcE8VDzdy9W
xbMUwfQXF2UaP4mN+Zdnqk8v8YjYefVSauvsiKilz87i4aCpBlnX8Pk5/0CkhO0B
dFCeotqy7n6VIwu6IXYI0d8QRC+o8kr3lQgU9fN0QiGF0xHpjFlMCdZMgjQUKfd6
TOK8A1gpGw04HsizmkvO/QVX9pIta1CKiRTWt5KCl8DVTxpUHC/GcNHC6KBqfGKl
0vktnZ7tYbF8+cmAq3m7Raefbg+6n6wOoypGAP5JrCMuQBZinK6bUoNl/BAcOoPM
6Ns2p5xsHDKI952XVJFwbc6d8W3eJ6lPtbHFjj2tok7e2pvvX7PxMh5wT5qKF27R
YNvF8dNJ2zTLgq1pQTe+mfGX1MI1M/gmSaExgtHKHwpgLU7E2+8q/KoILzFFp2DM
v00wyhlQWWUAvSJlJHHuKHuKl1em8KeKLWDi4e6ePDEGrR5gQok9kvDKCtc3t95A
z7svKuKINfZXhZ7AIicIM9Kb3wmqsmYja56A9/JeXvBhN3nTrTFHTz2y2udnsC7D
QDgnadzEYeRTgSJlQ+vVOBzaympAqahGE4Du+93dQDILG+/ri9ZaFU5ajb0Z8D+P
sWXZ3S8eLlE3BmuZV9f0G6+YwBzaT15jvOG0qlqeH9k+O+Yh8LaTVWFXCan8nfaM
rkDbLmx/V//9qqYsqJuf6/NQtKeVB88xIzJUmjDYxy14/cIZ5BkzvyCJWaCBtlmA
qhzHKsho2Ndtw83FS4mQ5aVjXy0U8ge5E0ZbjcwegwT3t3IiFckZe6m6QFysnd5A
tIjQiZheEp9yw+2XGjSfRpNdyQEiiXHahgLmbOQvfRp8AIkDQw1y7m6OKJNiFRMS
sjNJsozyGp+dhhBMPMMDSQvAKB47r9PYsIyzfov9tpJyKWD1AJwDgAWVU+eRN/tN
a1cDuZmaor1IfseVWFKaCh2USHAREy2wGJ/nWShJmWzRh8RUgy4B/nfnSvkoefBR
GIA+7b6iW8ErnqK0mVFUG2JqKStnnzzUatAHlt+Jr8SX+SAfNTfEB4KXwOpgaWnW
HThnHJOLM5u3r7LgZMBiNWD2eFBhgN6FMANJIygnOe8CvKlXgvftuEjS8BlpSNGk
CglXP3SdsahjjNFQo8v1FnDE7NUAbZsW4PiY7KRdM9A1oBGhXM3Irm1ErdYq8cYO
PLGqoScqr1BNQ9fNbPtmA540zEjNe7iRpLteLyTqtrxlgF3sN/gJ4I+RgkKSCB7K
hl/Q6FbymJaUgjCSEFDaDKRPFX/OORknB5G/p2b7fWLlWjfwMpXNdon6qoSfreMe
LlHDjy0T7Qfd4FPi24VRPOOypl2VLGMfzWHBesDzapzO5XjESKc5iHtStyXlvkUX
cXyGbCE6V5GvJJPKBNc/RZfYNfSB2lIzYnpmb93FcpcHbi8fBAX9AUAyHSxw9S6u
cEJB/na0rwE26XMDHMf3zWUG1FNBXVQ6xkWDyeb3tJ3Pcm6PVlt3LqqZ5J+vQEDX
4jS++XJiSmupUIC8UK3Xcu7BMvMnqkzIoBLLWEsLMZHuviNIUAHoZ1SmniClKmjX
VKsMLIYww3DxzC0Fld1cankPxv8N+khqffP/0rtbSrtPv1wckk7hRUboLJClZPya
DAIsPohy3U/HcprJ0o+TyGMsqgDaw2LHlgBO0pkO0UdwGan4mVTUwALRX1ghia27
nDbMRQuWh8Hu4IE5rpAeIRXuMJ8iurmiQzc57wRyUFMTYOloUxX+SDUB6OIUR1k5
+9SlSTwXmcxOPryf5e26U1iFFoyZgSH5ezcah4bQL6VvnGPaerlMG/jLSkVxiMfx
oewlmmXkZxdKDXZMkcgWxKq8Fgf7cAtGXfu1szOPvNDX7REW1XPTR0msVlEXk0I+
72rAWsX3P0B7EZMJEvaihaU4GlbffRNiUV5rzOs7XulwJzSVW4gGgg3s1CAY4LPE
MLYrgEUi6azbrxFlQY3ZvJ0DIiFRRsxL6OMAKXNmAVSYjtnXtU9EQLpQ7HAAwWE3
VTlG0qIfUWuVGY28fq77L16PqxfBT6YK3jvuDt4sMrEZtDpQLH8OUaiuV4I5xLRc
uRssnwNdwwSfKIm9QkkBHnWrPRzo9gRvhJbppnqX3gQtiIFcgR/xLZNplopXBT+d
3Jmz1iDRseLoyrlNUahgiBiI43trFpwJR0KKgG2Jx4taVFlJqqdqsqNzaz5I/nWn
BvavMBMgjQgsYMcwzqj/F8OcQU19Z2cmwvj/hXT156ZR14fsuMAO8N+A66tRsHv3
K8teESw/HgeIcEcEoRDZZhSoaxdcKnKnFQUBkF23WOJjw4jy5Q+nxgy4TZjwVFXM
9xpjcP8G2FC40mHasS6yOM8LdeBmQvXOwc8KktkrIhhkZNuzKhaPiFUKUMztckQH
jvieq4iIWVzAm1KD+oahx0H/x/ZpcTgfs9kJpnVzjYUNAN3c+vPVE2hYbPbz0A98
4Ggih1EfaKlSlVoAe/P/WWmoDyGswyvyM7V5YmOS+inU6Fh/crD83nMyjB+77dG7
FaF7sAGBVVxX5//Ubmc2zojR898y+KiOL0yTxhbXo9Yz4tQV7ZB3Eq2hS0Kobsq+
W3QRuVLCKAyajWNASyKDevUlSxcyQRkhYcHnEB2xCsX812hIlMhMrHPd0IqSn/se
VmQ3DFFdDx6kvI73R8eKfwK0abTXgwjH+F7M1iWrb4VDLuiuzBCnL2sEKzve+GTH
tI64T8JPkCMgYTS1Nvb+k2wQ6mZuA74S7UiQiBDbUJ6zfPN6JA6XyGWh9SHL/26W
62+Dy08Zetw6b8D9rTPdrdwv6YRgO6hPsI9kfBxIjXbfBy3MtDwMV1B1/4XIHqXQ
hjqkZcHiVLS+tkcpgI1tTSwIYq9IDykBJQlxpxl/7VKkTtXPvcj0GDyIk7thLUPk
jCsX08cxp5UrmLQwCo307LVs3X9e3l7pFc7Hplqh/SThnnD2JJQw/WfsMLUCBMuS
zD8mbuvhNUP/iIlkoijSGW8glbQwLJaMiBGAuXpj23LquW02T91f1/Usne0u/yKQ
tNobQOAOSoF1CS0jl+IjTtOv0/tjRB2sHPNQ8YjiOXmUDlHFLP1pAJGtObtlzHjW
kgmba8+mkNfEo7GQDW7NP11Ful1hLxZnOZq7jSc7z4faAjZAA0AtZvEUty/yce3k
uW6eunxsWU4h8EMj9cJrbwjAxWFt8GkGqUaIv0TwXqvuiYRapKrlpe1tb7nMK0b8
0fp/w3WjDDsdOtUiEvSQVzd2C1zWeC243TxK6saQyNNjtV0oO7sge/XmEnkzZrke
pTU1WaWzNrSiqNMCwx/Wa0yfgf5lPCidvbqTnVX+Uo7KH+IL/PzEbpdHomv6JT9A
lt5ifIWrPQfvlt+1i7XPJJAnfaMiNXSOm/s9HeQmWDfV+mMGZ6ss4EsuJkUNPodG
xDzbniqUxBK+dx8OB9rNP02z1iIvE7/Z+hFJ+L8NQ8YZHwxL9ZNOYpPP8Td5alNN
/loc5Hi2xHB+i475SEmGriphrEEc8Jgmp0PUra9G/URiVsYcXuJg4fqOrHK+Mz2c
PAs/4KrxLdaxtd2g7N68Hm200oAy28iL9Gh4uJKxNiAUSSmfn6tgBfGtjkKMKX8+
OEgIwfi8D3vLIowpaT7m/TtCHeNRNyRQ4BQtKsxLsMez/RfMYCxEemRxMH7X41G7
dnA9YimzVWLeupsuTSW5rmiiBUqETUBgK7uezvnR0T8Vwq8Zl71lmyEqMjI1hEN/
UFXVvEXTA4yJEkyFZr54QyVbGujTMJgPUI23wMN1jPEbPZR4IiT+OflnwPK6mBPf
x17pvYe/jszdfMkFVeihjV1lVtMaZ7hhlVmaKMhEl+FsHpPs1qEZs6z0BaERnc/8
706lJ08pBxiGhMzBWekHqY9bl9Bj1yHxpqxthwPEtskfPcGrbcVLUEJw/uR6ipYG
dpT/rFGIAnhwlU8iRR5dkiTXETQPAEoZ5Yp+FPVQyAcTvroPibm9mzWoRSN1BHZA
DoYfM9K4rI3qk/9MK5O9ONw1rvmVM7M5lqirvrV3xSWlNCEjLQmBCSG528up+UKH
/dPC9tisrp0DJzkzy3IzuC14PjL5f478PTHd/SRdagsrpH0/LcUmI/trrfpvvf4R
AsOLq3Uh9H3Mj5GIM4kc1mfALbuf4Bvc0u55LFhOsb94Vo/C4Fe9Ykg4BfjwY6w1
GYA1VlEizskGauw4ZTCSiGsr5LH8PafRO1DmjRNWIPPzwiviP11GzJLr/hIi19v3
WRHys8wYPFob1lhka4qkKPbaXAbQZrqlSdKWpAFGC+BiMKTWDoYXnrBu2ZTWmMNW
dLUVzRxqNdE3MqA+pXcYPv3lYqeTGv/aEMujmDYdrV2szdMZjFPiP2LiSF3W1kBK
3dlQzGjhjrL49lWPdylJqgasX21n5u3kYFPUFGKidQrnX0rOcYg7Vu/mIOvg8wVx
mJPIjgQ9rGbAbG/zaBmJaqABHq0C8DH+jfg9rzcF5hjYxOfTDiLy6ZgJ1QXsHCDn
lyeMFhCKAzxAHIKu6qHDufdXSpQ/DArNIQEq0N8PtK/dZOCw4C04p0msjumcnptX
w+N4vRKHCAxp8qWNAxgRSLSDdBgqY+2NogPTIw6UFTDz+jr9c0Ursklp0OEMDWhu
fKY/Ry4XsezADoo0cZ7yNMam6ImlhmJePmkHsmSM+ZGGVzYzS6iNWqnRS+/BjLkK
KkMhuwwlxU2t1IQ6TKELGEWGlj6kYoRG0D+iCaglFCkRgbrToNUhrhBbwZfZgifP
xWuRMEIedLVguqI/mXCH/i0vgH2KVCV8aQCKjogBYmfuLTAfNOj2yqZ/O7+oGTLF
2aMmoUAUT5Bdy40qyss46OyShxkoQsk27CpbZcVuUTpNxZOlOMrdmvr5DsXGMtzw
oyljDMDHDQrXtHyiMMkzL5y1A245lOuFhk6wzF6kbhdPuVOkURCdGnrxNG+ji1+J
kDEfh/4zTh/gM/7XPlgk0OyanqY+eYlfv7tyIspazhIi46zkTK8qGwF4Qg+6lsfN
GAx6rQTpcpkXPt5fsg06LEYBGbYBEBYBR/U1F+Rggg5MJDctCAkEuxyBpOBNup0Y
SKAv8Zz1ERyy++qFEMb2jhT6dCBJtcvGYaXL5vyYgcRGNnsbyNuNwxHENqeTIU15
nl9qZ9xAO/nMVICKn+UI0M4qcHkiX/ReG1wsePDXTBME5rUEVxZv3zuGQugOh8V9
m8mDt+yUE19Y0BnFaiVCe5Eij7xiwQUlIc0TjWiDib2MkcCXwcHx7xfp+Ztwqo3t
iKIHdWQoKdAyXWcBmUhRDO4cLOifzl/undtBQFoXt5oXzaA1dlsRSacgVX/TZOw6
JxBwAmf4+7x3ZIMwG2GM+lrW/+chEthZaAUcNys4lFVy2t3Jze0U3wA7lwb73+f4
27nUt800v0kwYA84FObw9CZP+1YYPlwe5nEhT3kz+y+OsZFz+H7PYSXF0V0eu7Ny
eyvmQv4OP+BKzj8jso24SSw8ms01C68SVRCsSuRTPxolSFZw5jAPc6beHSmcTHdJ
kWcYfU1f6vBZwCzP0AbLlatLOUs5bRYx62lWOhseepm77znGsldQPWT+RwRigma9
17ynPbXwDSwTDHYPB9/IyrD9XY7q0fAayPmwpXiMQzxU3Gywmltz/i8RwEBWWZFu
Q+sV933RXbNMbhl9x8cQB6B6Zt1zuElr7tkAD1glHMp6Ih2ASUVfZzFy2clLi6um
vaEhMSODktKf2f3mMOUWLe2/AkaQzCS9HAx1v7WbsspB6JJHCHZbMvvlFrIlUFRt
Zej8UhkUNbE0vNkrk/zFfKHFEN76be8GAnIT7dUtpq29vq3zvHfVZejkyZppNe5z
3xGuso/njk78dtOkdIhYkSEq8M0JN7PEi8AtAfDrn3OlqHYIEYqi2EmIkjq8ukzP
uc6zIzZGStG5VE9BzMNJgDpON47Is2bVu5I4ll0jfzKilY/m7ypzJfVpo9pPHyrc
O4/OJLD5IIgNHzS8mnoBITQGMnRyf+ouGBgtt+BAxvE2rv9GIaUgfN28QBMVzePc
9UTrK96nceDoiCtbXPoYSZz5sLHlhwU1siLAm591kRhy1IyDfaqJ7k7N5TJDmKeJ
dkEOIQROwGaiylvo4WxYANOWfGu3o8C0U2rUS/fYHxpY3kCfTVk2Q7IQ9xyi5cYQ
dDRe8l4/xvpzVBitYgLzaVUji/UVvTWZkdEcys1hFHGu2eI/r/F9BI67P5msxygU
7KJdx6yZ1WxCfW+ibK5nrGIGnLs63xypOlNaUXXbc0jqLfcWRwFx9v8FJf3W2shG
iUqEi/tWRxc14J8dv6bgXqIsIMrRjreqINuF1mouIAi+YSnJLLhk6JrvhAq31GWA
R2HsPjTDl2qOqDCk9q2XbdXlKqPOWaPVyINnuRQ6VGMj0xZhl7u40ohKd7bDEjfK
1OFPEDiQjHwCbOd59/LDYfWXdGgmZtIIHsoSbvURnG3lKoASPtWjSGvszv7JJZ7q
V84Ofm/HVtD3HnEXlPrtm/eOBVERlPRjWAVy6Bkz3ULhgqlqGnOf5SPVSTepXVOy
RhxCIhE4g93rKQZ1cQGoRodO4Yh33BhHnbtDzm5xjmLNIlb1aooXwNh1NGOm+Bqm
+OvdfWWmNnKjrE4Ki6iYrG11lTM395RZrzQ7NgNElDrrWwu3vIXsNw3Q4uxdaonc
Z30d7bJ0muwqjPqv1OE3XkJbGz8q6kLJbZ1dwMt1xHEtJpEaTdXLMRJyJnMbO1mx
00nhPdfKeckrta2lMpU7ut9o5au0zyAvQ+a5i7KQlDK8kenBaNLIOVkDu3vTc6M+
ZLv1cHtztzvoFTMCg7WYHzfPQJOW0Ixspw+zWPNOPFd9AaW0HprW6EbeAL6jQeIt
y8LhJI7jhawOlfvkAKDcap34Ve7XRqUIQwiK1SpjjfzBiKAGS8ruiqjQYTFTwmcw
41gqvR/87c5jOrprz72tnxJ8HW27uz+9N4REIEP/almN0d655U9ygFQ0/PMxfXMP
xuRBJ8ozhFYWGxv0PW6AdPJ8gX9PzFOl2G+v/f/UNBsGLpZWEmpwdGq7IiuApnMI
6eNdBdllLaAbUZ3NyCKnCIinJaAkqU3h0ZE5/d/H6cQXk/GZB1Vv7f3vsLbcXOIH
7ehL/X+jJWUjAjV+2yD8znrDf1Aqhcblt1c7fbnwQWrjID6RbJe4wK1DAecSSptZ
f2GpSmyNDF3PG5pqY8uMQ1pR+40D2gXBz2MD8lstSt4ibDNde9DsqpAGWrsZL8EE
FaJb1p1qrtSd7P/jdvchX7WyPuFLsWz1bE28JYupgiM3oMN5SxAy1NmrMik6dSap
hpA10LrXbsg1O2egYN6fNzRnc6kqAUAw7PwWOdLDG7s7eMF9YO2NHI5tuWAxmfZE
egHhNWWgIbWarFkbJfaayS5qP1OJt+9nzeupHPbxZIhkQhmPOw4OXP9BHJ8pU5T6
tw9dKWz+L0lc14+B/xZXbInneqQ0DVz8AFkaXaHawHkwe5mb1IyA50CMweDiNlly
keqoarsed/rjBds7Cx4NpuDR9TiuL4B0DeJ9CZuxX23T6AkJR171dsGAfIYp9tpV
9QfkQiuXIt0+NF4Tr6P3QZ8mnZxsjWrSTs6x3pAXVtAFSz8sfFOi1wMAWTz12KKI
9qU/k/GOxBB9s2bq61dYRTNIncON8uMp04GHSNfboKn84sJyhXUYdomdBjWmkRzM
ncruHVw32LSBe0LlT1+x8L/LGXoG7ZPkT+/HbxikaTQYOEtcoge5GU+1v8LyDh4u
umlRHaSxNbQ0yW13SElxZt8ZOT+nKxwGdCss+fXy/G06EaXeUKmQnU+ey5jOYcvh
p1HDMhuLKUFrys6v+KgQyYtO06JPFNxiz77tKZy+VfaILGhLiCxs/9RHkMCtIHq5
VFEi2irpzOhae3l487Mv/lkSEp34CelgNIw/xZ8PA9u0RzE0SuiMujN+2Hpj5gx/
eVRYwRwHNV5WZoWkMAmbFDadmwW+MUqnBrN8xd+ZNtT8MeqivosVKCYWgqWuA01K
8y4Tw9QojXNDLLHoRfmrkwbkAFFYbqyjbLIKCIh+2MvrIXpR6zzeTU1tOh39rmZk
tLds7w7a9xoLTgrtmOxjLZnJOT1rqXEHG1UgvXFcMhC7CL/YHKGu5/2bQIv5Tgo+
eN01oQlUb/m1aegymkRI8IYDteEjCGMK9gxPdmgXs1nwdLV0BXZRc0xngVKgqolu
MMfbYsMAPvAJYspJkxlaSo6bD0EUh+wkxC0fQSqCTdIzWRVqNmanFoh2AZCIao1w
bg+TilAzFpPeRNANN4x98fDafRnL8y7xvUOCjv2RuOyh/EiyXXcRWo9CDnOzFUJ4
jLR/cyKlR2q98lxnOFAwJPvlrgf8wWk8j8lFtIrXHhGCm1ON5KVd0yCtzZDF+LJB
oGyOwVGv5dfSxSNXw2oR7f3/qIZ81uiFXIp2cZbaFnTIBu+vU5WervDM3veSvx/e
ReW6WCg3kQwfmycR72QMkgl2kGJKia4qfvPi3ttIPiIsgXHzXHNJSpse+zR9pmX7
+3CLYUk8SpJwGN2RnXPmwGvrfeHlzgvyBeEwPLMO07mGdmooqjYiPVDyQCW5ngKk
wMI2ayH8+Lo1i+kEzxusypLk8LioNU0cExRR+dLSfnFIL+dULeueP3SJSscKvAnl
hlUWmuzCNkOcro3GbfsGO3ZK+WvZwk5oOvheKBSLwWs4DXvLLMvnm88CwgPgMb8d
bX2VYfIXIk2R/84x51i1z6UAm1h6NUuVoNRf8Si4C0f3BpfgFRdlu8w8Rhi4W5Rb
C2kQny2yW+i1r3zPxMW/i9Z/Auh6r29ihD6vkwpK7T+1mN5znBQL25IyScG7zq0T
LCmZ52HlmFVIsPSpqg5r1xl0auUQx2PO/drikobg3d5Lf4yo0PzsYiBPDTCIeKsk
VfgT03BbAo3Ebg0VDBPj4KIBb/TDwI74u2GtNfsTrn2miMdeH79wJI1OfgVYVTGy
xoqU3pITjao6VpgyCZ7oBzW+Xri5oGnmVGE6cjkXac/n55rd/XtKYpWjKQqvJsM7
e0Ka4zVE8pCYL/5ZY+jlaYUkqw2Ho3ShLLuOgwqv5JauSsE1p8cIJD5BiXIPHr1w
6dU/cXMvS0aw9CngW0mdGGc42Y63PcYGifWX9T7kx9hCBWtiQ7Xs7WD/XpS3MhSY
MEKYNhocAF+Kmt2nlMNpBwrkLhtsv5wV0HjbOdVFIpU23o5DEn3uybfqnOLLUpUG
e4ozCllBqmqu5TfQ+sQ1j7B5u9gnUOETu9W8LGLlDNoCWkPhyF+OVue9zLzLJPV2
Qz9nFX+5WPWbFT8kC6khfyBvT3UpGknoOvyvlktwaS43P6cfJhtE8LojAWe2iBT8
Opyy2hnv6UBFP1Aws1hw/FxuX2kWTxf1AkTR0d5TkgBnOEV3GFopitzot6K3FUJB
9uofd3NgYDLmj6+rI+AzyZspx2BEw3z0+H1XI95EUmQSy6tOtjlOtl4wFaFutlsN
6inKgpciZIwnnzqQNdvGleh+krxg+GHyxEmgVCG+mss3edtZ9ew//Fieqses3WxB
mZO0w8ndxlZBmYBgGCNBPNGBFU3eabZ+UQ6+5a+bg6bb3Bww2XwkiHwAAUI+RxXE
FtXZf4K5pzagkdq4s7L3Bux00HfqtEncJYDTxPf/AuYNzEKL2Ee5Q+AQ7czh47gz
XfzETEo+SKYl3oik8KHhDz3Beu1s8lxWkrl7X0H6UjccfncgdGOL9i68yxI27nE/
muxwlJDcX0+Lup4QVekXLetU//mXYMkSPW7G9zt04lIbi5+TYEYQMc10M7V2yav1
cDCpqnVhuoxnw35bETER9FN1mg6QKHYUSMTHXO2bk1L7ivFF4DHR7dY+xeiY6Xkv
gppdbPIJM8sXXIBrnljblZ/HoJETEJy8c2iQClq5hp2Qr0sVetLEs9KKzEsgdkGK
8RiDQvF5lOphQ0upXPJU25QE+BUlNz4jezOG5f+dBbT0Q5xJLo15ffcHEDR27Nel
Db8wRxBN1N2BKZJ4GEeSoQlhccYfKeCaIcYu7gQEk/Z6JLh2nShFY/EFlupdRsVy
ypNSfdLjIbn5rtuvKd52jXyU+5R8YgVaeRAhJfOt5lADuKblAUMArBIjTK+8JvU1
UC+bWq2eyeLAiHbrVJBT1kTEf8TAKnMzF18UeysCdWOMd1WuGjZkCnD5Fpv+tjTP
TBs0gR4EqEnDh2vTiVRsquLwWMwH+WgiT3xbDDN73e0Sw1mf8DdMdXS520x/PpR6
qt190tTcFYaW2bmkU1nY+44jwwi78iBuZHckI4NBz2Qu4vf4/p+jomWj/b/zr63b
Uri6OW91pogCT1noqpiBaOJnaTt/xl4Z6tPOZcH/O1fb6w3+BJDjRKh320Me5g4v
jn6JUKgPOlP9I6VZi8BwTA7kskTic30zeV0Ynh43ALoxB+JJ5irRxcsawAp+PSPC
MxcxHYOpW/nA9VAD4swd5kqPOZykk3gvYSakRkq5y2puXOZeTh3IO+C9p7lUO2Dw
y32zvH0QcIHIhVqo6rYerhHyZJXkGNkAAW+YvmHKoz6AGa9/x/zJ6KM4/BAtznr5
wt3WUq2ueOVs46R4eeiWv7cjKly9IGPjOWNSvKXm9dK4ngr2amHM1v3mS5ggfUV3
PAtli0BoiAg9PUX3HEQ03ZfaLPnCa1Ds1pgM8dsQYPwG/nM1O8H0r/KywZfoqUxM
vMgZVkd3DdQl8YMbqQw54k7sOLxF1eIHtuDSbiTCwWef5ibV5Yy1bnejDEpHq9Dw
krCiweac7aWqg5GJCS/CnQAo9SRrY0/wmTUs/IurUwFDoTmxBmTqvbX4RIUwcfGP
Cz0ApaV3aums4oXz2xCLhV60lahk5/6WSh/Y4WyvIeLrhH0qKdxk6YgQVTKTTlhh
wl1Csu5ZWMXBecRGgLHsOQmQhh1G2Q/kZbLf7XyOqZWJZe3u9ArOP+6FxKhfXc9n
bdgpsf6QnhOmrhS/2XAu40wmOfwvWL3hHM0cLxxbV/Atzf2DGHxNZaNB3zR+UXmd
4YePYRgAp+ebjrueRrbeg8V7K9NQ0ZSt4VTf1PK7faLOJSbflKLuohSQHMISDQ/5
yIxQ1mVIfFBQDhkyEARt0nqepFIO767MOwmo4sLrcoiYdgKi5fTjL9FIArDCNi4A
aIWreLY76Z0t7cp+LIu66ODplKQPHHHbytghtk7n/31W6TAIwPUUa2fNgp5M1ejE
MT5d+6NXOnjcE1ucX+k0WoHFCqYxOoqP6EHOAoJGta5YNa7PGgsIgtLBa0do/Ljm
xIqadtJ+LPncDvDCYIcIAMhzpKAtbaT/C8uBLPR8JHRv5pvMdKtOmbdJM+hVlnuw
HOWneWaAk+UfFbt0SV5NoFl3MkFdlTPDm7Qfuor4MUsj6qgVEa5LK0hm6xMotnZT
iVfZn6fWcy4ZOiyVbKXbmWk/EARtU+DMCn/bIqoNH28mHznzl/CZDHtgeq+XFYAQ
ce/Mc2k82PSzcdpmBk186gwMuqOE8vjFhHUsULYiauLWMCq/JQ8R5MrrbpML8ujg
kB4VhwWva7ZHrQ+25/CLyHCkVTwRQ/7QFUMx1+TdNJTVC7yDJ04K7/TRoipqTAa3
Mj5M1Qxg8qSP63cN1UAElvAZPnISTGTh9SVS+ky+zU7Cqd8+MYzGW1cB8W/JYTur
OAIlDCrS8Kx8Jv+Tj46Pj7bZIDnG9aREXSndg9xM9czoF6fFqjbHEKSgsia0Vvd1
bK1BdfYDgP5UD4LdBIJqoU4EzXsNfy3txAUgTBjgkUBrMJIZLLTeFsWwEE+wVm5N
HLXnkGRWRA26emLKiLj0MknL+TOkXR4d67l/d/DLO0ZlWJQyj1skqAqMQhEmG0oF
fXDTgcshhEqaqhDBZMO9r4hY0RS6Fovxujp/IxlnkxjRMhmGSKIUaaLX7ZSOq3b6
xMG1uI1aBQskwo3+DkOfBvGA++EPxh1tp7aVxgYDPrIOma3Yvr8CMOYgBfaMKTnj
8dGD07Ozm7OPCNRtJ7lw1TigIti1KDeK5VmHVCfIpSzBgp8RQvS18sZZzvmnXRUT
vmZU4nXtEO2BPHLxJXkpkqsMPueO0R4ey3xozfOTxrzeaI2iWlK1wYKY+PySbHaW
3BhjTI8obFmPg2mFPRNqLVYvYUeGI46kDVbV7mJYGAUHi5HoCK8fV+eKvPmL1zZu
F78iTHvDmHk5fSKMotqrRc+6hIn7dx67CurNER4QBF0+kuIdsumaL1xtSxEghmx+
np9v8CSJecnpgGtfbDkpuAFjiIFoRlfVSs0CjU9Fxfus2VhAiUzLRX8P43aqpXb8
0dQ+kM5+n9rDZ64QmzMZb1pwB7qH7BuDgb34X/LxrK6mVINiTXNtDdAw6kV/JA6D
CsPprgzZrVC9A7dzbyiVMz8DvJu++NhqjUhFdc5RU4yPLIbt43wO9iF4cBa0P9aa
WmR/5YLDGB5QxSFqbl1u2rmjb1sH81VuREf51kwOfiWwGGC/rY2Yz83/wLdd2w7B
EqM33N0qh1o8RAEkPjjbu+Ghz0HNDLM0A7Z4vceewc5hAa9XzKybLsZJYi75b6di
eltD7E94zqR91QlGY3edGdWinRyBnn9sdftCP0xzPtq8OD+71FYPRfgu2IgUWWJu
DF+6cxd1wQ9m0KT5kkx4Ih9wKRse9TT0QsiefKSX3c5XSHP6SvnzI6eOf1p0EuBf
k4A6rPJpk8qNQROjDWWwp15qc+ILVtBlNo2sdf2q/UFLjHvbvB0fbnL1a0dwTQ6G
i0fjqeRLoTF5RP9RBExUCz1voD/UkU2/dnxydSwYEp/igLELqnEn5SIqejfCx525
vnrnHO6wIL4EUDm3xCDsgEu6VFUK9vHzjmi2KeeAZ41x66nCcJK/m2LL6rkE1KIW
XLwtvEpTS0d91Ns4q80aWVLmVieWwrWepVK9ceWiiiic89nuVzf8cAqHhUvmagVM
5cW4yh9Q19d7JXMimCVkZ5VInc2PH0uUtHv+by/i359rKnC8M38Q1M5VAryw8WXR
V0xqVcMbkLdZbdbykDODBnDrlvr0TI+/AfrW79O+TNQDIycp5U18ZcrW+Rmrlh/B
PfAvxNHpkNg7xsWItfqgyzXYe3zxC4Rpavni0bdB45QB1pZjcaFhxrS5Js+qfmEo
FaoouRWZL1BAFc5SIakTIXhoFZEDu8UnV38FxV3fClqjPubqCNSOEnUtjYolrcQG
NHhUuQQfIZuQdyN5Ah3CanPPI9XSmqVYmGT0uR0BITtgqlHSYt/5W9XWTFdfDz89
pGjUTD+KBBDdXSxK3ogQ/8qBH0kX1f5SstoezqX1QiZqs7lTc7oBnAjA/4YxEri/
LZW6TtU0GB/00WWmBbWNSJjhAYsanDCHSCX6QWRC9nQnMzNuc8lHpinz2mAJmUEI
8Qf1yy0CuKCq/rNP8/bqTbRBYT4ODOSTs2Lvc095bXrwVlrF6Pk9QcwXwy+DD9mN
E0q5N4y+OQWOcuOzaMZagiAe/DWoxe+KFAJZ58pm1vI8GunZDo4cSo5DKYGsxCIT
bTXZi2CarOgKf8ZLx6En2FLSlVwix8weoqBmE2idZAHBvd7okmKyjiKpfCc2p+wk
oTWqH7xbKo+Wmoa094laYG8XSSFDdpG9YRmZV+pBIV0UvOnHMufBkrICanA+4hwM
gfOY0xdJL29U8khMsLVecYfdAYos82Pz/RQWw5GawqnlRXazSBwfwlDBKvfNIwlZ
oRG4MzTY0Io30Pvj76kDz1MMHg5fRWhXDRIZMK0kTZzxsKINNqWKqaTJVgXgyjZ0
/l2Kft+ioUnH6eUH3kglRiducvQtOVbMjjtTYZyvJ2+HXmpAc9xTNnHF9jd9TT8S
DLt9QP+7HzPzUYbB7lT7pmlcMGMH0199priIpyQjdwCrKg7VjRPVVdV1EW8fKIZX
9rDd3eiRYaR0pWZGjf//LCFsS5VejD8AmMiiPqoZdpWUmxNiExBD6vxgZagNe5RQ
glgVNLB8oD1WEzgpGg0Ma4k1B0cYBEONg2ezUqRxfMTXoJBC3DxzsWW0MdLnRwJ6
ZJPVaYuRdTtGbg514TVlZSYNCQJxxlgsCw+g+98Bd27Slw8I0d+13hr1zJl/hILX
28LSCvNrggJmElp1NsajUQYoLooZbsxANBkJx/WWyROMPp6bDl4TPo//30GH8tXh
D7iV3SWfI0/R44SFT729t+0rMeIpKFyZQMStVczhA5f9FnEeTw34W7HRmhd+IRhI
4YOJ9Id1ccxgzS+Q+hdiSkDH/qtcJfYxH/AwjEzavt9TgpR36ijoXyMIRU88fkI2
9ldEA5w3LsOmrUJiyHamZzZTbeCgxwobzmBNykQaACNLGDQ+vFzfTmmVKBPG5G3g
3kH0gCLKTXK6TYDi47sJiZJ0nW2uVfeyrbVEIcuLp3x5TxwQLm0L7IJJiRNpR1cR
6YXb+RLmGKvdFFBN8BQURKeJcWvuRaZJRn5yWiajc68dpCh6/II9/w06HQW25/BT
B18B3cRH/pJ8bsNdIp67+osmoQr9SGo6bfSUZgKflRl2p0Xlx/Mb3iyF4YfapkWr
QZ2WQReWp9jcPhMr9lTTHE/aOOT5tZBejnauWu52XTi2XDfbe6eI4bxeRDsQk1un
o86N2Py2JomWg13ZleIS+uY48L/bgUxIp9fKyaVDPVcMjEvWhxFIbyr1mRswuqML
cN9mX8+v0GRbactKjxOvx8Dp+S71bdr2UqLswYhD6n5iev6N2idfDOVCNLI+twww
qw6ukNo04oO3SMBWEdDbvnAMKQCTHEqzW5n7LWOCrPcGlQldj5sjd5H0nf28c+Ii
A1K2/M482VtCIm3AbD68jEsVg80s1udXMQEXfQcToEawjF8xfpEcUXccaNuZjpLi
Q5JwS1++H/niJv41lm9LlQk9Lm8fHhBJwFhmYnpTbwciHBDaZTmroHjsTCyalMea
Xv0rrvqP8NP52YTEcI2U1Ec0NIYs0ZmtwhUzmPFAvncZ/wpD0x/wxIwGRpboH977
E4eKHIDo60ydpO6wHOccRwefbQZNKlZu47C6XH+XDADYeqzSFuBsZs5iLTCUw6U0
0sRkPNw4OWSo+qmf/TRx6kmFvawd8aZ/CkVt5bgb+yG8DHHtiAKgLq9GoFFZA+Lw
qoHkiBjBSV397ljVIPi3RCoRzsNGDwxAEdN/DXw7BYFIXVoNfavgNh31ByJLYuz4
MRQpD+wq00zfZAWSHDZtUQuAgZdlGmJR8v0KsCWHVPhe/UJ9aavh/Y4tisCanfaT
toGn/0hlixzvWkif/rxgIPuKbtJHL44U3VWiuIcBJERc26VhbicPrGUDQJbaF31F
Utbxm7ljM7Nlpt85pxVBgqMpOQbaj/7vkg+6Mjf7xcDjxyG8siSavJ79HP0/LsFp
RbJwABL98U0qgXR0I5e6/bDg8+zkubPvoSNl3gRY8joO2y210pn+xzIEN5+o6Gd8
J0FCqZ3Lr/sVmgQrTxB2vlFYaICxUud8KIbiNda5xzFlDoN0EPF2jxq0wqG7+i+R
HcXurIjzGV03NhrgMQc4Xn20vVD1Rflbu2xwfTXYCXNh9cpK6HLc9Ping5xZkQgc
evV2DDQrkzjsOSIoWgA2HN2pFmoGtZYVSZRR5pAtPQrJtFrQU+cBhT8xZ/XVY45y
XWnM5lVh2973up2XpJrJXGWUcIL1K0v1xKn4PznbEsnmIzW4MMefXSzwYoAae+JK
DdVBIMnx/uQ9bJ8SHhN0ZO2RyWhHqD3hJnFhb213A3FVd2cPzY1SVvf2kNry2ht/
M0ATgQsHMKQfPXyJsj1kTWBGBW6h+LMWPGLEyGLhpuNcl6CAHzcHdcTb/7JQiu8c
bbnsxvGfwY9xaxk1QIwsstejd5VSYyn+IsNbDvYB2mZVFuzd6iX2kvqej/xoPOFE
doOlW0QpdryONt8YTYp7CGWZFSHjWN3WhtWMFq3BC18kZ47e+pdp5qmtPS/6uXPn
zXwc8/eOnUo3nUExmZNyez/THFs7yChEBeVuuuNq3HXIHsWooZQpsvNvWcr2wuXZ
yPLlmYIaCWm8ywqiypZDS6vFBt86r7KLBu6qJtQRER1FlQjVRLJaHqDpKvPhptIo
n9YRDYze6C6ZS3fD22BV/h4VVSQsgskjlzz+wtv/+Mo=
`pragma protect end_protected
