// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:28 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
I373wBX22giiOrM5NokKnZcMH6tl7xVzrCe2fYwtrKM8BjU8iCQgamJR406poZjv
xNNhocCd55b4e71hYdum44kVZPYj4TASbk7rDmWSoN2WoLblqxe93vRUmspMLNuV
f2Xb/UIplI48z8xbCiQIsnu7BlSv+jK5kfg+KyNAGA0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
QwZdBjpWDe8bPPHGYzkt4LnHPiIws8/UwoGroO98ZWoOLQZSGPBbEY/IrzqOgPUR
q3352qvBmxfhC1k94su3mjBn0uERr8EDQiqgofYivzNOrpoZlbp2t9BfbRpDxOL0
qxWK7j5oVDmO32bY8sSlzV+wvsAUwxuJaC0n3r7hMEJ5/fUtF0+Q7Y0WLUrKi+B1
/tlMqXV07EJin28R5f0KdkJsN66psSC3fJCaXJg0QsyUVSpxnrz6rPoBpIPGblDg
06W0mRRiT+RYRy7dk2q2KwSJdTnIsjBI4krA/lGfHaLlaDVGV23i0M9lRk4WREl6
3+HTCuj4rD2h45ncPaKT5cKtFg+S2sAeP+assiZU3+pLZC2EcVCjCPpK08n5Fv8U
xXK9mjl8JTGeyqmS0nLpndz1S3DLtrMzHQUZGcAA+StOp0fJ7Ei/dugY1M/zK36H
AdfPajoBH5YMB4NWzfqh4TE/K7/gZxWH8EpX1A1ygztZh+LkoNPHV2F5DA++xw0A
RsApkgXPWwfL+TpxL4Rp1u8/2vVTCl6ezhk8/j4r8X5tuSfVKHR/Y6emjjknT1aZ
sidAx01OqUcGICyT8BWhXR4kmxRtd2z+AcUKdZIj+2SNaqCRez+h3cgA52vKKeEv
NhiLs6woMemTxchCKjgEGdnO6e4YAoxHZh+nYDUF0+HpuKH5wpEXlHwt0eP2J5oU
GPrgVcvu2lFDcPJiUSD2MS2RJEsn9+r7vX1Dm9OUWSbzI+kLsBjFAWdfRuczHeG5
vfFNEyKxgtBOrfamXkh7CWUmpP3Rt7zplFccSyokqSy7BdCMrTz5Ye3BBEoRl46T
ZUP/JR67GsCsykDS1CjYaEoagTOh7su8zB6U7bxQqK85dekfb+vf7dAh3GmQoPbj
XTznR7cfvOpj6lV/OkI90g2ZMb/3IHRZu2e4aSlcIpMS9SgyAOLt+N7OHt80V7Ht
Lu63AU1iRrI6hFInJ1U3i2/n6WfOpEpFh9oD4IC5xpKZPTiSUns0uLdpArevbENP
JVoBGd1ma1bz427n+Ro5ZaeABtuga9cDziFR2maj5NXKQVitNOtjkjiE8zwKpygQ
RyBDraTyNDA36nh2ZulICMbNBckqsGH7ImgwvXDivrzDC7XNELEz7DVrsygfHgsI
v5qgFaxR5F9W9DobTCkfJNTAfVtJqTziyz/HThlTDOnXVF/SWXUNmwH3JOpjwrz5
oOAeolOyFd7QLzy/Iu5Bgv/A7o3shBD7HMFvwDjoFkAAzZZvS8GGAG4fLjchRgpN
sAQ+Fk7Ovc905xM7NuWYDrrj4ty+aqpyc9WmHKa6yeqzs1LYgEMP2x/bs6dU4Hn6
AAJpKWcFuba7rlmKCbAuIkt/rnCA+qaAW8upqKE25yaZL/pBYhwT50J/OgJ9tyjb
Gad2HDVL6w7fDfJD/xHkmbtYI2cMC5CEfO9YYyhKYNGaztu1h57GIJHRQpTWyc51
1w0gqR8nKf4drEVZSg33DaEo3pVEozWz2+Z02hT4lPyGJLH6V18CHI5ueEK8RuaA
M+4Z3fp1KIs4SWtpv1mrNcFAMS+I3SxRw3PSO7BFN+4Yytp/m9o4mPMVUeEKfwId
+dI1zQQ7ZUiiuVL4rwsoDLNeUcpg4u42Do70Zk+CaEec67L8oofAvX2S1OL/mXEl
Xk97h5dUorY0IoafqnVWh7mYYwuA75R/iHQmOjXwvAfEFEhzCyjxEalYSh0TKIf6
pOUbVC3YDph8a0ffcCJ5pelWLigVfG8EDiH/fYG30Pksc7dFWn9kKH+Q7bzBWevF
n87LQmJUY2bZ0ewxWzIRfvkTtoQXSzhKxwZG8wptAS50e7vuvakn5KSjUPIknTjN
vbb6Bnnb5rpvQ9/VbSua3BuygxCLxwWAtjv6zB4swEvn+ED60js4/eIX4RA3qTcZ
Tu/1WoCLm1jkXuqWJZV+RVD/RmPbyGv1Ob5G+EaC4e8IVchYQ0j/jP9LB6cUTyWf
XgmJk39KAdaJQGd7zVtLObkBm4Vzsfgp++gCCf8GtQz4r3Qyk0HDYXJjgKyEIB44
PIScnJlx36FTQbVt1vuyDG3A2GlfNzwGjl0Oj05J1c5Sw8OoOQBM9/CL/q2GXCDU
yItMZjF8NMX4jWL/5qLnewy92qUh+Ll1Nh1rMktj170asHH2ZW6SzzYVoz5DDDMc
zzILtp5TX12Am4mIItnYC2106CRqzPAikE11rJggVFfT/bbhFfLQPjeauso09KJX
zswoiu4VJZhrRnSke97bdsvuvsSi9leOlHd9aFEYb/QuLzWafEaESwmeRd4nLOAV
Dmtvb/XoCL0nPb/m5VezCkvoi38afGECG0/1FfHHx77Mtkpl4R7GmFRl0v7IjIAs
g0Qox7vrA47J+Im2sDtozJRfIJTOiRUW6lEvPhyYyiS9zf2SdbGuPCG3DwnllroH
g0EBDPNZ530XntVukY9q3tUCMsTTCO1mXM3uEWMuEKeCyi4rguPWb/sWFh1hs5Cs
/oTG31ws89P4gkl1Pbcd96m7ftPDEnQjWEGQ40vCjwRQ0sgWDUuwM87gn/nsFYZh
QZmHSpnqziaQPV5ZTenRHIoEKHoeSQcl/36xAbYrLvjXH1JPHm9XE/hmW+9RXZWc
G+8yI4bgbIMvti3TOE7nCTpwYA6/Tm4a5nG+hoY0z7HT1sj86e2TcKOiDFp8W9B6
q9owrIt+KBb2SE6IMLywwz7Uo+EXogWfvYk2kHuNdSft5LWVvpo0Cm7bXCW9Hycm
q8pYe+M++UCUEUbLyPhrC1rxYEbL8F9zhp1hZ6kfF5UcoIdhhBQ+2/3lMGIzGEIR
csTW8+/Q87PUD5HmsQOUvO1TYW17qkwwlXsmM8h0fNo2ayz2/DDEaHz77YNQ2dH8
4zoaI+rZvI8pZWybAdhVWOp2h20IHA0NvC21vDZw67/g5X1kn9IJRFVmILg4z15X
b/maWDzPWyC3CFkKpNEkduONamNuDHWgpLRCWe/7ZliQdbMkuleK62h9FE5C5eFY
e+6Ir/6kiMB8MgbOvHajC5SrnsuFhDYqo261o4zQLDMAAek4wRo0Y5WMQIOXiecY
1kPPFgHa7J5ftDnptu2WoVr2JbUQIre/CpbYFJ46CgaBnRmX0baeN+9mJin7nC4o
xxk5IxiJHu79UwzYrkO0tNh+MO4/1MW4KcEC2t+MxgXaY4WHSKierLCa3W7ywG4Z
82FA+ce59R4jcPCQ0KeMgiie6Wtd98qGLFRsAmmzPm0Z43RT/gJPx2Y3VkTyYzGd
WqSqqV0X1V3X0KO6wA7kERmDoFPmJ6G7ENiHTn5k8DQC9qeNiut0C59+zAyJKob7
fafRFBMBBBPr1zrPhF32w9srG/l9ypo7tuvYP5Q9VAFYcgKcMj98sc4JnEkbOl6K
4kQ9CfAI/aOCWsqyHfm6Kqa1RUPp7s2USceBjcUCpQSTzLY9zuj12Peyf+kwXWaX
qB4OKtaWPobDBrl84Yft5REcxa1UEd4F8H7Vp/dqSCLHlA4YQUsyPK2PWekk8O/W
M3cv4oB3DBC2R6La3ETXby16t4dyPfT3eTqBGOwyK78z/13sMNQ3UgsbelgJywEb
dYLqD8ReybzZdtZPMjxQ+fVJEeCGapEc8p9wCBnxqDrOlfxwAdfCBR4x5X4Bw9i5
p0JjhmkiHpMBkfedsvK/8+3Jnqylbpyus69KNeNtkLH17Lvt+GzwEkVRciBISx2T
6tS77gaXR+0wzhwzlzQKNTbnPggTg7iH5rrEsHWTfwjrE6rj+jdrWWLIRUJu9Rn5
ySR7wFW6r6x015fEDZYCAVZooQhcqbLOAXNmod0cLofaR4zXcLvreCFHRs7pFpNz
SW2BJV8WtjUstlE8Nf1kMyc/du9rLKiikNoS13mXxrp31iSuhl9neIgp5UJBqndZ
1PH3w9Q9+4EwRE+VKWBIddrQDQk0OCwcCcmybIqS8Bp9kgsZeA92x09tsBUyPAHU
FkudQrgshhFaGEPBO5lk57zK9WNVVqaINvL+PY8EmxjUArD4+VOZGihLRNABn/CO
Hd12VZ1gk7BV5vsJdGZltQ==
`pragma protect end_protected
