��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)���vG4��NB*v�^%��_�rG�v�2�H!�W��m�e��
q�˖��������7��8^�G߶��;9q����M��q��Jh^lq�cp%��#�Y&�9*d^w�8��Mrb�/�9�'yU}�/���5Ps��7.���	D���7<e�.�γqBBq>߭8�g�z�LBL4�bRn���bޔ�a��xX�3�y����qa�e8V��o�@��kUw��U|;
��p"��g4B�K�b��P�������6,�̿���U�<!�2Yt�R�$'B̫�g�!�U���:�уj����A؏�V��.���7�%U\
z���r?��e�����M��Q+d�	�&�Xȏm��.T�Y�g7X�#�h��x�V�U��:ǉ|O}gB�_�c }P�6��-�;E��<;sD�*�)O��3
ưr��
�p�6�'H�&�U�`���@��y������z@,��E����1�{f�8����D��8ۼ�� f_���.4�qj�T���E�F��}��A7v�f��
�vv����޾]�+B���[�l�'�B�W�x���7R���'���0����&��vWޖ���N��}�;�k� Y��P�Hg�m��4V��,�	���a��oj\�,H���&�3`������3/�i���ź�_��3��C0p>���צo��O�2B� z�Ru���}��h)K�v�h��>�dӆ⋋Z������,V�1`ep�S4Tpy�~)�7���ޤy?��w5�w[^}����+<���Xp]s����9x�|�R�H)�"�1���[u�Σ���Er�0�9{�Xq�I*U�f�.ώ`����]U���Ʋ�R=�6v���3��n@�^���KxGQ�]���Gm��g��=R�"Ē6o+p�_�{ D���2�j���M&�`�qJ�ߕE�Q�H���4�ٞ`�jNeg��>ut,�7S|���3�,c���j��Nx/.c��FX�t��tEa�̳�^�7|���������A	�#�|ԫu�{�؍H~�a,�L2�wt���bQz[6�/Y�@����P"��Y3h�4��X�(�.��91R�,!�aG�O�H=6��u!����b���(%8�6��U��؅�@�5��������W�,	j+V���U�D 9I19#Ϩ(�d,#eT�?>9B:e��M˭7��f�cl��6~d�k����s{5=Y�4*��G.�����>��N#��|e�j
�Ike� ̑F!Q�:�?���ɒ(�k]x:�r�`�{��	zf�2�	���J�����7�9�<9�l�H��qW�hu�r�ż֏�����G}�*Ħ����+a�Er�eU��}�I	����T����$а�^�a1��������7��_���Q�zo3��d|���O�g�H ody,Ƅ�H� �^���BNN�J���:����F�}(%�1�{�=�B_� g\���9���~�����<a�m�F�u��O��d����,X��K��_��qɜ��St�IyM� S�gMȄg��74����Q[Mo���M�G0�J5^z�9��}�[�X��K�g]y]�Z���!����ۀ����-eL��L�!�3͛��U��M7���_�S�;6	�)�'����e\�!~�\lJ'��G)��7/�.��$s4W����uf�(|��b�e,�gˍkqׄ�)�U���*af��A2��	�D݂BndH� ��Cu��R��<Ń���S���1.�+4T�6xXrIK7���^[���)_mT�3�����N����٦=�q�A�ǭ`�&]�v�`��L
�s��	�D$Y�㞴*O��]�!k�&�ċ��ߨP���ǈBx&�W���'y�n��z�'�!��5��W����C�<�j�������j���꧔�Yhl@�F������`a?F(�|h��	�.��>4�Sg_j򤝺Ԑ����1��ğS���w��̦�Ր�+�+��b�&nhKo�ao�Ǳ(���8@H�3,{Խ�̔�K������`ul\Oid��2��Va�Վ�p4�;-ސ���'�y���j���)�#��nW#�33Y��d���9R!�[`:��YLge,f|
�������/t�Ǝ'ؠ�A>��#Ԃ�*X�h��H�O�6b��H�w�n4��^�}���ZK$oD&���a��<Jw*X��/},/�)�1'���~#>�{wN@���Rę��V�����rmT���0��G�&�h�~W��6�n��I@I.yE�]�Ԟ� �C���Bf��Pfu{����2Tz�?�GN�g68��I,hL�x�6y�>d����ZF�#�fV m�P����0t��`r��[�3�����3q�U� "'��[������q �Կ I�j{<q	'��������?Þ �no��Ã�����h~� �Q�ڍG�gu�pk��3ڕ.��D���{�[C�G[�'�h2e�sJ�hp���o�M����,:f��I��;~�O�W.����[ry�ºV�+/���p�T����{��|��uy��aժ<����s>��6(�n���2���x������#oۘ�8�bܲv�i�$�I=�%�IW�!,k�}�G¯j�:Jg�rH~���]Ƈ���!I�}9��2�prF�>U)��}B���Ac�ԫ���3�$Xi�+��u���.B|*V음/z��ĵ1�̰�=��C&7���;�Y? �Ö9V�{d%�=�}؞,�a���L��s���iҵ�����ԑ������u�7����m��o���D�N[b�u�O�7Q'%�UZ�l���*�#3�	Er�c�ʈ�7�ic!x����vML>�\L��d�4�Z���O<���+*��Jʷ�c��>�h|��#��4�2���'�d�g�8_ ��)B��H�K�<)s�h���3�_��Q���6���*�#&�nwV�)��#��
6�ݗ���ؑ.��:ӎ=~W��5R9^Vwh�z0>��L�ǈ/8��B@ ��0�
��D���)'M)��	U�t5n�7c�*���pw���8$&��[�<���ӼUg`<x�.����9��A'�/�*m��i�aj[�:J����a�2|-��"Vȗd�w�����2���J��3�q��A�k��O>k��jw��}��Y�LϨ(Wa�:�N{�U����b�[����B��4d&��S,����T��ye���yԀɠ[�ܵۤ�E��\>��(���Ԇ���j�޷�_�'�i�@�Ģ�w!#������A���^�D֡��dG{F�RJ�A�+�Z�=��u�����}!�;cZ���!��aw�>dT���^Q��ɑ�ԭ4=��(�ڬ2�I P��Ph���P�¨#��o���`�4\~��wuZ�W Q����qq�[6��3p),���?0�`.;	n�+K�\���k��^g�/�,d��(�A�h��E�`�1���n}���y��J���#�B@^կ����_?} [�]P���kI�̋ɇ���/�b����(jv<�
_@�������A���O�b|�RT��F��W�]��bS�q��O���%�x�w�^�b,�܉�j�{�����HW��RV*�4��?�r�K�I�P����o�L��;7'2�d�©�#��L��<U=Z놦6^������U�E��0^LO��rC�ߥA�Ab�}dW���j�-~]i
;�X𙉉�ޝ���Ƴ�ih�|�Y ��xv����_�f��}����"0���#��+:mӴ�����/������rk0gc�خC��ԟb�+�mR+������BٸR�O����R���r㚾��`k�E��wg�����7�f%�`������ѯ.C]��9U��}{�d�
_�F����f>�S���%��@
����J:�᧙j[���.��_�~�t$����*7�����)�,�l4͞����Ћw�'"]Y\t��7�~G��2""������'�G����c���Sz��*�t�o�j��C���Z]6PR�/�V��ƛ��7�q��Ia�(� ���t�|4*������00V.�������{�����ˠ��
w;��2�N�I��	W���j����#��E3x�ի���1C�L���m���[�Tf��k�mS��b��,�R@���~`��(j��&�H=�0:=Џ��"�bh�3��T�@?�Ti}�*�<�.NV�"Il��0�SfMɖ;.������_ȃ'�.�|�����}�1�=�e����k��n��uM_��fS�
2��a��u� ��H>c���!�W�G��C�H���͜���6�5��2A6T�Cn�r $X����e��ȽO�0��R�d���e�!�lO�&�����N���7�$,d2�Nc�l��3L!�t���Jއ�b��9yc �\�b�P;I=%�Ut"�_�D�")	3��`�s`�Vtܰy2�R���/\jO�{�߃r�rj�~������qQQS�� ��Ks�F!@
^�N8�Tj��V[���U��X�+%�C����OD��Ҵ@��|;��=����/SaIՙ�7kKG~=�yY9= rcЕ9t����Kv�N�a[@ՙ^�C$ɦkw�%�}���S=��s����BӃ�O)���g�݂m�$�ńm���~A%ږπH�"�!��U.x}ET�5��#G�vt�E��'Wi\�ZUJ����$��y�z���\���؀(3d��1���ՙ���e�I)�{h�A�$�V3O���� v��[�Q<&O~�i](��?�9��	ئ�#x�P��&q�߸�U���l�$Q���	���Y�5Y!R��]쑊��[��>R����@��jB���h�e������ߟ���A7^�3�Z;�P���a"��^�L/�Q%���*C ݨ(����Hm�\v�|G�yRsF)�T4�l�č�OO�:wܝ�T(n�kR�J��jmn*�w�z�l�y��xq ���+�.�΢���ul��^:�|���o�2���q�Kc�󫅺�Rz������dd4�萖���D���<N��>�c{��i�?���[�0���Uϣg��)�y2�Q��H����®���������ypz�y� U�����Q(h�M����D�m���΄�'�k���ӭ�=	�ɠ��8 d�p��S�tq��	�����Y'���dC��x��!W���F�T�.1��׶Խ'�����w�۹�_�&b�,pOg�6��V�E�c<U�dgLr&n<�MCPu,�k�ݨ���t�f��@R��f H~z&�w:����P�I@f�4\�ON�(�~�I� ��FMz�r�1#\����B��%���V��ֶ�i�֨���;{~��A���������V}��O{�k�r�H���nF�,����@�:��x��=�`�Lr�C
�8}܎��
b�e�pL�/�+�Z�=�E ]�����r'�Ux��M��S�_�����H��ͅ����싩	��C�3v�n!�>Wu�OB2��eA-|��z㫹2�0"`+b/T
���d�ͳF��ʖ\���{�J���5H�7�����<�,X
�]��-�(ٸ*+7h��j�^������XY��ܰw9	~�eO+�1\�E]`3�cc�O�W��,I�E_���a&�k}�r[EFz	���GH	\M}]z��L���zkr`�4>0�l�`��ELv��ee)]���i�&9�|�WC���ﭵdΪ3�����B���d���;^,�F�{=h\(����[�W��+�D{�h6r�Q����j����w;ʥL�)\}x	�(?iȧ���DՄE=��J�qS'�K�)�4�����i���Wk�D�͚Һ�It�&E��.���Ȉ����:��~�$K��
P�f~�`t���Z9&
�A-c���0����Sx�a�?@���r'�¤�a\Q#��A%�N�<M����(m��u�(}̦?��)ï��mY_��۬Ƙ&3IxB�����V���]��t � !Q�m��+�X�����,$s����f�%ϩ�B���	�ك�������7�P-�E�	�ȉ?�?b�஌u#ħżr�y�����D_�����q��apR��9*l'�'����$"���-l�� �ux]\:Q������I�v�K�#��W1�%
	�j>G` ��s�Rρ<��,�A&��6a��Yd��I�$t%Ԧn�Ƕ/K���-�w})y�$�af���ݢѴ��/�QL���>�%(+ɹ3��L���Sy0�Ӝt=��}^�����CI�+>C�K��03�CC�܊�NEs��a�u�O�+�`j����wj�_m^�.����q	J�ԏu|��A��'}��S��+A�i3����8X`V
ڑ�$���l0Y��s���)����2�e��o%)�\q���4��e>7���p��i%G��{G�SM��2��Z"D�`h
�︱�Zp��3tN,�g�Z��8\q��3��KSH5?��{U����r)��ٱ>�"mj���-"�! �'�䉢�n�$�q�rR�C�,����/���?����/ٵ�Wܿ��%���q�E`("�eL8U�����dp�:%�(��<j�?9��Pb��];z\�W���g�M�E��hUn6ډOG�vG��[��ܬ��_��T҂��_��h��E��4���l�Gk.`��pzЄ�'?u�W�R�i��ƹ!�}�!2����>6&�	����|/��B8ɠ�h�?�ǈ 6��Jc����=%~Ø^��m��Lj�Z�������@��W�G%pY��vX�J���nW��]�ɽ�>�FcЀK-B��/N0����O��M٧Й��b���a�Z/W�Ea��78���,�C@��K`(�]�d� -�>��n1�$冼�7r�f��a0ʚ�/}{��~$(������@��Ê�����)W��X�ГyG@޵�#��($�SУL�[>(�Y��Ρ���Nಇ�n%�,�p �������T�%�\�D��Ճ}�UCB/�ڢJ�h��ȷ�L��2�D{��(�C�l��8����س�[xۯ�� �_�֬©�}FyG^M����&�X{�����F��Y?����vg�R�3����(�k=�{���וՈ�uVIa'o��@��P�	�/E8$�Ҟͨ���'�*]z��fXv�R �,�
k`%oD�h�S�i�����o3����[س�[O�L΁
���/@������a���^��؄��G}YWՌ0��^�C4g���o$��9n�"����|T�*ۆ�(-�����\�Тb�k�-)B�vɏ?�?�L�� ء�[H�mZ�'Eo��fZao�T7���9pu����aRL���2*��t%�)P��o��~���@��{F��ސ��. 's۝�I��C���?Y�n$�~���<��t-��+�rl�Ϛ�9G5��pH�2Ċί��v�����~����hi�k�����@6C,"F��\q����*�^$Ԍ�W��0-��3=/�� ��>ag����q`ҙO5��GJ̶6�
���ĩ���3�L�&J�g����C�c�E��x�*y����[͝��#>��C.���U�G�Pk�d��o��]y�K��6���;�{�Lk�d�v��A�K���
R�}~�ڬt\~�4��vrf��5V���[y��������3<��Tx�0��IB�-�_��/u��Kf�L@ƾ�;�e�>|���2g���4�l�t�]��X���a6/���+AtL�+�I~�[����yt��PM�\�e�ut�`͓����
�^;o�
�27b��d�ױ��獷�xbb#Ut��yC;��v �����0wA�����oE%�ǝ<����	�%@��95��;0w��O��mM��מ�� �<6��m��1�d$6��a�n�\�ϣ5 � ��(�<z�|H�1�Җ�B���J�ˈy��٥�`-��\)�B�`�����S(Q~��s7	��)�b�����R7+����.T�b��2x\�Ɍ����@v�L��?�xr?�#:U=�vtW��q{�/�B�o#RnE*e��d��u�x�n��]+�������^hA*���)P�c�宎���m��Vq�ܶ��-�T��I��h8rG��E�!y�q3��t�F��҂#�<QV\���s,��+��Q�FT�fW�a�;���"
�?�2q���}�`睛W�s�>6�I/�@�L�� qS�TM�^�u��	��Y92��qGt0,�)|s����*��O��x�60�׋�*=�H���!�q9�;��0ql�V���Gvs�L�!>���*�QL��!�^`��t�q�Yy��:"M����VL�R�$@�?	�c�䴏�ط���	�q�-sĆ��2���,X4Y.bB�yFlW�vC��)�~iUm*���%��+�4���fH��Zd!n�l0�꼑���l �t2)'�Mbq�!��x�j������ܢ�$M��k0	�������o�$�o`X4�/� �V�3'�A��4��#-��'�rֿ�uZ\�(H��)"�Ç��hj��9�ӂ�c~
�����3��ҽ�f�ۉ'5Mnn��1�-V���?�m�6A\NO0�.1���Ʈ�9{����#՚�C����ytp4��N�r ���S����6�>�
v�����$�Ӊ��|QWr���>q��ĭ.TC�w%���&���N)
�N΀/��<9������Kfro6�Q;q^(l�M4�g�����|��x(D��P{hy��n~����5{��m9�1��9"<Q��B�u&��fF� W���6�^��ۚ9�z\
�y����'��&��i��E ��B�2ݧF_��i"��*�����X�ѵ�jsjS�����灿����h;�����"�{l:G�2T���dP�>��Rj7�O�{�,-}���AX�����LX� �vX��b[���vq��l��n+vN�s�(���4|�c  �~�D~��jχ�B��O�:���;��w㽢�2�H�`^X���MaO]ư�%D�,@�I*���D��i�좃'��F��|��T�ƪa,�g4�f��������e���9�b����S��6^��9lU΍
ɳ�*�@f��h�F�;���s��<��Y�ȷ!��`��'�v�Z�61�<��<Y��+��Vju�dV3�eVu"y5]�Y�ު�P\�LϾ݉�-��8Zi#��2^]S���D9p5E,��~���O�:��Yު9E�{Ve~W�B��}ܝ\�wg�����Tut���I��6@�ȀRCˢ-�: ���.ta�Bc����sO�?�U����L�����fȊۺ8RQ�J��r��to�mjӲ	�8	*-�CD�*�v?�]|)̇S��VL�R��x��'z3�zC��=7��6��3�H#gt3�������̪UQ@�E�?���0�YK1����pq��M�Q�ב�"�b���u��|<4�� )�O�N�Xƭkr��9�a6��Xa�>>U/A�Ė% �*��.n'H%#b`Nxu)F����l�W{� ��!�����RwѲg�L�!����,@��gݫ҆uSQ�He�.��3߇��-c�Y���gIϼ~*_=c?��Uo�	�nL�^h?�"W��vV���T�l��_��&/�'���X���G~� �)�#-�7��q�|��"�Q��7|��]�w}�c8=���NI�x������g�	p�uL��˛'���XK�Y
�H���������>��W��2��y=�#�m5~^%4�n襦&�^��Y��&�FT�~�3����d�(��޳�F����e�C�/���
 :���pb��[Z�mOq�Џ@C@�
-��'4�����®�m*ؙ������k�!�G���Bq��v\O�k��������јJcw��+�����DH��cz-ܝ��R��p�Pd�'�f"�S��z�ݲ��a>xd%/�Ү)��-��
���Y<����!*�yG��W�7<#tp�C���k�o���-y�\ ��	���W�^����(�W��>CL��q�ļP�� @U7Mi|A�/N�E�ؔ/��.3���*�� X���0U���g�5a���}��0��:6y���i]�}1Z�~>8��H��X�WR�6'ׄ{쵗^{���@�;,M������<�T�k�����$�3Sť�a��tf�ׄ��\��C�������_�X�� �3��0�J��Qh�u��bFJ����<5� �A��>������(XW�l�Y1;G^`���'7'�@��v7A/b� -�ׯ���:�P�ϡ�4�~!���Q�If�^���
�\jG��`�)BJ�QF���YB��z�f��Y��m�T�X�+��= LqfQ9;�����:Xav� ��ps?С�f�cķC��>��L���/֪�P�Fl���C�J�TkN�Դ��ܔ
��6��ɍqLﱁy�F�7W;3ј�ɟ�6���"ɓx/�*��-8]|���`r�nY��=�#+����9Uܘ�M+l���¹b����T(���B��)���%�F����<Ǹ8�FN�4o�\�,���J�/��޶N��5Y�+����*��`+n�i�p��Cg,&΍F9/׺���m��iZ�U����9*��?=�_��nU�U(�y�So��b��]
�6h�p�1%�ǒ�C�*YT�0���?��׫�ʏ�;�پ��2�B�Y*����in3�ӓ���N�ڀ�(b�YU�yXBa�f�p����O�������$C�o^�@Ce��P����Z~�&�_��w�C��+��_�c.ˡ�Pտ�v�H������?����Q퓠
�p��K���@K�>��0M�Z��ƪ%��S~7!��V'�����C9��M1��^����K�����]��I+h��q���OM����ܵ���S�L+}�!ٴzB#������ �''�Jװ8{��b�K!�Ek����-Pޏ�u�J�!�S�����V���֍"����UV��NӰM�ς&�[^\
������	�"��Wj��av���_PuWK-(h�[Q�C	c:|��*��J�������WB�'Ű)����qn_���r���]����x6C*�C�9W=�)vV��������`��\0����=Og��)�󌋠�52]@c������������+�hh�iU���)UT���x��������y�/~�O�H�R�����كVc$���\﭅"�F�#��h&�%{�6��y�a(;_D�lSͰ��}u�f@�QP�^���<���^~d���7J/hg	.O�⣵���e?d���'�_al��؂�u�+P*D�n+�S�6%E�ǖ�i�v���'ER��,V��X5�6|=2H�����g�4*Gf� �O��Yń�� Me�ӱ鍲���������:�b���_�e�K��X8F2�*��g[�����m���<�d˄3%�2�8�����ffD��T���BCx�Ts�d�P�܊N�)���3��F���_�T��*%�����'�l����Z��Ipx�fGMm���>jO8�9������1ة�T|����A.�\���Y�pҀ�^�A,���&MY����`]Ĝ��v{���7�Z���KDա����y?��q�[�XeL;FZ���w9��jv�8'�����l�}5�'^w�%�=[�j�Yb�(.�N��|$a�Շ�"�`�n@��A~֜<�8a�:�.����1�Ԕ�K�iYV����G�kœ&w�[��]��2�j�)�;B��S+q&5��mwKL<��SG��j�}fH��Sn��.������-}S��p2vA��Yh��/�U�����j݋i�E��1L�Z��~c]����v#�-���!xS������ƸN�=�>sQ���n��S�&��(B��������U�8��7��9�k���o�J���M_c�68���Rҧ�0CZ�Q�@��mW��|�~+�
sQ��睲?��Q.܇���˓�;A��U���dT��?z��'���U�קl}��gT�H�}c�OX(��g�s?��z������)8�c������Y��SP̼�c������t�i���+歂���7å�r�W�*�����
3V�������-dl�>k��
ْQfv�\��=W���ĕ:]	>��˭�Pd��Z�킡�]e�`� !�Q���I▬Cal�b�c�{���mF�h�/.��� 4+�u]��6K���jJc�Aw��3�5{it�gT�0Y�<�f� �aC,x��tD�tz����Aڠ+�A�ch�V���h:gu������{t��m,��YG7�!��ͱ5�����6v�G�u�B�ѯt�����b pz=�bk�ro<��1�䂂X�\kc ���q�č��J����)Of��Cg��(af�#nL��,��&Āc�|Q7�V,`�tV�#��z��P����b��
a�"$���l�7�l�c("�ZL���$9��ޅ�t�<��;�����,hv_͞�2T�~o�t�"Ę5������R�c񾜭��3�d�a����<��͡gP�}��h��G���C�}��q>1�}_�s��h��׈ɼ�BMd�.�-�2�������^��`+��D�ȼ�� V���#�]���ӑ;o�[�W-5d%>�D$AH�q�Ʒ{���õ�ǕdL7�Q`�$*c�_B���BI���l6 ��^�3�ֆ�WQ�:{Is��`����Ä��|�@�䀠\�ag˘wЀ��������,��c��

K��4�O�sq��R��҇�ȶ^�=���H���4K`�0 :%��╆�l���O��$��0}����И1�H�����u�����<1}X�p��eA�q�BG(��e)n?����ӑ�n������j�hA��0\kox�"� "�R��g�Y�Y=P]�`��u%���J��)B�s�E�"��F�0���&�mU��V�t2s2q�䤚ӝ�%�98�����N�H21�-��Iz��3�L޼����z�\�k]"(�M�7"ּxlj�陓=��殯�wf��\Q�L��Fӷ�~_cZ2z��[��`	j��[�{�L
'��A	�YO��0�w�^c
[S��ψ؅t��Ȝ�"��>�&����ޖ�����
$-`�6,d8����]��.,2�B� b��j(c�Tr�hJӵ����+7Ͼad�RJ�nn����G�n�����Cs���Sx��#RŢ�jY$@�0erk����t?b�S����{�\�Ī��4��P�5���2V��t!� 8�b���B'�C�.���ap�i*�1i}�f��ג�Wo�;D
ͨ��A�ۦ
I��
e6�*�0����f;�4:Z}��r�6�{�ܿtR/��=\[�(�F�| ��C���H#t��a\J��մ\
��R��Q/6b ��WK�ŧ҃��=0��.ʥ�F��7�1m�P�2�k�`ki6��`�9�}[^���,�$�?����h���}#T��@H#�[#0y���׀	r
�^��XZ6���X���Q�UZ�Jb~2$Lƭ��)�N{�(��~�*>�Z&�u�G�Moo�7O��:̪��Ϊ�4 6� ve�@�R��,ݰ��ň�A���inz�m~8� A�h�|(.;��֣���}LԦ���#���X��)�F`a�Gq'��cC��?������ji<H�4p2���9=��ldt�EǗk�����'Q��� I�OxG��䣖�<7T��;��S>�+��[ ?�@:�bz�{����Si��K����О#"�P�JG��侱�5!��`�T�����rN
�vA<�M�q��7�DD�DسEGj����<�E�m��Oz�Y�E���S��?Q�U��%(9�,0�6��C��X�H�]�KӀOT��;��!��B����I�)��j	��3eki��@��u� ��ɟ��ek��E���]Ȯb��Y����z�����j�Ct*�f_�4e�֗�Ѫ�脱��"�c�N��wJ��l�vH�m/U�"�����9&^�`f�;O��`�;��WQZ+Kp��`�KG�7����+�Z���k��*�;RVze�;�G�D;
�����3eo�˖����}t��lGҲ����R�5��x��3r;E�,��"ho�I�V���n��H���P�T���5PX�f��zЗ��O�X��[Q��%s��э>1Dofs�w��f:=h��u9䭽� �p������)����yG��혒�������4{�U��.���̏Ea�#���F�1�=��2|n#.����kZ��@M��6�͝E�'��KXq�_�q�26��J�w���3�F��@y�%TY��ٗ��(��,v�����%�]�9/݅����jfƆ@N�������"���0ky���m���0V�)��
/��	��ޟ���i�|�`j±�/'�hG���� ���P��4�&���_�D�|��C���1���϶Nq�D�ds�5:g݂����<��"ؿZ~?�c�j�88��ˉ� �ͭO~���U�GK���(p��I�q��Ë&�-�㒤"��j`C�2)�EK6}k�Tt���JGl�f��[H�e�����;i��ޝ���d��F��������1s���2����Зژd+?/�aw/�P ���Es#�]�S'6��6蠎7Q�B7��H�U�i!�/�6� ^Oz?hʒy'�i[}�\mgP��cC~��.�V8��X���M�w�YUd)������D�tL��X��%��@�@�����'�#Q��w����R����%�$�|�g�F�d 7<��9�SD�-�	J>���|[�&��׏����d�	R�\i�\����qu��u��?j=� �q3զ��o�o�1������s�W�B���rL7�R!ՔnўUL��*�����(QfpYF�3Emx�Go,�zTQ������Gb������%��s:e���M�J��#��AV;yurى����|�B������5���,�d���4�ZʄR!/֑��	xl�_��,��\]^v�<kuG�:E׉tu�};]��t��R=��c����,�3$�#�Ϋ@����#�㔶��;���A������QF�sjH�����߯Uۂ�%SP�C6�.:5�_un@�҆	�8��fĢ4����J�_�g�����ۮ��vźbvٝ��J�� T-�R�i�{�f��I<!��X�T���E����U��ǆ'����^g;��,���ơ��֏$?�������˲�mbχԀ4(��P�t��vt�8rVÆ�;�S-m�x����L&�;��.&0�8�m[��ui$'�{����jz�K�{'Ԅ�w�$QɄ��=X�^_PY]K�Y�����C��L������T7���>��b��j���j�����u�Bi( ��T��(8/���t��#�[��_'BP�ӥi_'<���CB��ܺ�!�%8�7�|p\�����
�K�z�,� c�o)</'�E�jP��e�,ɨ��`��56<�@٦��!!���Ir2���k��y�m~��RJ3k�.�6���h`��������vYqͿ��5��� ���W�H	�9�$8l�-rמ�b�I�w�+���xlO+�r3��f�p�㤦�e{c�ގ Z��U>N��-+��2��!�S���d�%d�����;��o�1}N>�0a4r��V�s/��@�>����o�D�t:����V^3�u��SZq'��Z�<1���r�u�c8����1i�<��)�������b���촒��������p��2hB4�3S.�W7�����Wɡ}��'7-����݉��1B���؃���uj�!�k@>%*�H )]W�����5n]u�s�L�B�P���GI>pז'�g"����gqu6��!�`YC�v����@�����*&c+��3#&��_�< 3�՜�A��?1�}Η�IF ��QU�o#-��<���7:\`�ҷlk2U+R��[%�˴�-�;��)(�A�H�����d#2��0Uo�pT�� x���癗��%I��R��E�N��T��2�����=N�0;�cȂ;%1ѕ�4�F`Q�h{�x��;�߻���m����MZ�a���`��rC���y�UU�N�c�����T����5'���Z�?������5����,���+ N3B�]�s��Ƽ/fc݂��֑ v`��%\#�{$�ÛL�69��e�w�$�Fr��� Ғ*	IX�_���;��*ڐrz���X"�@�*k+o��A'L����ٮHt��90��S�r�F�f�)\�Og����Y �n�9�LC��>դ�#�IлsSv�Նx��l�%�ߟ�B���{FP-�Dӳ�sL�Pp�F��7���n�6tz�<8�:�x;��*������a��&���Y�0X�7jO����⑁�I��,#33�S&��J��G�T�`-c�H��"h��vF�.����a[�ۢ]����>�ߔ�����s����( ^�S����K�K��t�l]�1úP�~]�e�
h(}J̦����RbUS,Fkw���`>
e'ˑl�k�_��x�c�
��`}'N�~��`��b;��I͌��5`�n�)�ǟ p\r�MO�oN�Lk�&a)����c�tH���@I��؏��ˋ������}��r��9� ��4�j����RŖ�!�]��u�[KM/y�uB����N�[ �R�7��[��n��� 2��6��vd{[Z���u7�y�U�f�O{Vz�bڂ��1}����)��v�=C&^v���9�1E�\���+���p�V�����z�Q8z��0���m�������5X�9d�/���!��d��=�A֙�����PE	U`w;�Ch�{K�n��)��֨�v_S���f�-.*����&8�^���L������v��0d��U��*
�(#.���Ʌ 	�������B����!�&?w�O]��a�`^B&s����2k��M6�k���wG(~��+��UV�%du�!ٟ5�JwЫ�6$�[�.�o0�N��������:W0�G�а���f�*�t��.�Q���>�U;/qZ�`���{����`�_s��U׺��Eܴ�k��sE(z2o�47_[c�G|L{z�5���^�����=4���:А*��|!a��M�1��o��_r����L������t��+�][m���(���>ҝD �w�w��}d-7��"�(�z۠
�ԛ��R����5��]�Q��B�"�g~��i������ذ��wg�dp�÷�-�LD�B2��/��@����)Vn1l�jÎ��=�����P�&�������:5���Uߺb����32D��w��1RK=���osD�_�L�߄�A_�4*l �_=k�ugq���$(!�W�'��,�dH�W6+5 ���C�K���_U��P=�i�x�[򇁘D5�1+�~�hG�
�Kԣ|9-�Ʒ�X���x�eڨ�w��,������Ә��Y�!y�a���o�77������)��K�a�~�E@���~<�������S�/�5Lx;E��>K��޶���v*l:Շ�xB�Gh������=l���Xt�w���P�H�I��uS�ԝ}���8G:�:)�|.�f�Ǝl���Q�����2ҫ�P�Eb����v�����9C�{}�ܲ���|�����6��Cs5�x��i�< c�#4�-�Q����0c�-� C�%���E>Mۀ3�����Ȑ>y��7Cm���04�ߍ��+/
3;'��w�s�Ht�Ņ��C^O�u?���بU�u9����1��UŐ�g\D�I�/|o���Qk�:����i�kp�9�ǗE��Yv�=/�X��+iJ�s�	-7��޴9
]�t�ɒ�k��~(��<Q��ˑT�D	�����-c�J�ݖvn�W�y�����p �].N.W y��#v�#^���Rs� �*e:�%�����~��8A��kT�B3�ga�,T��iO�.bi�<����'u��=l�m(�KI^�U%�jJ8�w���	�D�ISe�^����3'��I�ur��$
��t}��O�V�[�]�O�lw�yۭ�m��(�Iy^�ld�����J����_3E�*Ri��;�Je�O���
"�;�Θ����Pg)��e��._��%m�[���C���A ��4l�̰9�{�1Q�noI ��΋�"s���p]�V?����H3�^�_��n��V
zmȖ�k�[/<W����C%��c^wJ�f�1��R8�3��i�E����ܔ���J��ߏD�IE.i4�� �w �ɣ��{I���ߖ�B�_� �I@bC#��󩗤�O��\fw	�����^��Xjc�J��)��DsG ����_�U���Em�6;*�+~ӬnG?�q��q�+�v�=�(��.]�N (��=ȔN'ٮ#�Uc&��#c�}���oˊ�?=L�@bJno'ѯ/��T�s�Q4�[�&v6�_�L�;�"�WÊ3��}���m��d{;�'�]:�0������˄�詀C�C̔��O��'������>=(\18��.i��@Ԗ�`fǀ���<_��A���lZ~L�Nw��8
���AhB��n=$�P��;̸#��z�q��0�}�����f�L��d�{d��>9BH����>%u�`t<�׵�e!dk�Oor��Y��i�3�ج��.�>��nUO�Ρc����(̍u�
LSb��3]މ�ŲF�xv��4����:W�X�vHdxh+\�4���M���+�n�l���;�M�I����ڰ��G+�!��gy~>���9=H��6�|b��Dŗs��WFQRi+l⋡p��B����l!���*�8T�W*ah����m z�iB�A����>ɩ`(w����"���z���tJ��'�b��+f�5��Wv�%���m�eW���v#+��4Z'8kt��٪�־�q�x�\	�}���ht��&Kޤ�^���j8����*��h["�%{h�����S�gM�Ï��b�}��_�� ��;�(��AE?Q��S��8t$��v�YA0ㆅ��:�.���/4�����BA�j�e��(�-̎�:�\�Jf����ݎvb���V.��������B�(��Kb�����w/�xUJ�8�)��Kb&��d��X���)��57��|�'d���9"*���h�^7I�2��HY%7-��;������1�w��UO��+(���qA�Ց��Iv�����6q��ʉ�W���B�>�;�q�ʣa����Υ��`�K�d����F���
.��Y��MZ�ρ��1��9\/ jN5GV�$!X����6;����я�%
9��ao]�E$d�-�gc3�}�U��	eF]��O�q����j~EU��-h�x��
�9E�T9��ZD2�$�o�?��2ՙ�ŕc�ع�������oةN����X�ZS�LVF�O�$��S���F��w�|Ch������M�{�X�����Kn��8a�#ޢ.�$y��NX�{|*��ك��A�n'}G(���.��)h��2����U���Xrx2�&�V�X��A������z�pg����[-S��i =�A��
�s �ڸ!@)a=�	�Utɭ�P�}^\zZ�%������_-�ՅzǾ)(�{p�=�"�#��5����}5�H
QQ��Ϫ��I�Cm����>�S��7��F�Զ�|X�ũV�P����æ*X�w��YNZE/��F�E�*�Ƚ:P$ЊO��W��nb�,��_��>Gڮ��󎡈RӱNO�I0OC�ْ�d�.��vM�-./K��Y%����PJ?��rT�B@n����_g�OZ�eD&f�pP��[���öb�qP:��,x����1�hA��Y����N��>��܅	��Fю� �zT!�,�Ω������&讋;�ȀHS�׻�=�c��֨&�w�!$��)dQ����o�%d
߻�0k��f7O�ܝ�qƸ�I�7��)h�hw7=�o�4g��4/��cĎ��6)�jB6$21��ڊ�Q�Z$HB�USϤ$R=ݐ��̓
�����v�F�鏽\ļ���������H<C���~�+!�o����zͲ�Pwnm堏6n�G刴V.,��*ٽ���ABL���[	̪}*#�[�.Ugr��mwt��C��p$μ708�s� ��T*���)m&�����G�
F@V
p8*"��yz"<����yT�E�[�6�5���z9j8A�6&�E�雰�.�#;���V򝳊�T3�^^p���Y� h�s/u����a�$f|��KT��2 /��2��E�oDgF�g#9�jS���� ��yZ�pzn��NȄ�Q޾��*r<��`նi��	�v�㢥b�i:m�>�����u���h�7�A^�6���+��N77fo��մ���Q�7i�m� r�iD_��+w�GR��y��)g�_���0�G�a���O2>M�-�SP�5׌{(륾�H�qql�R���N�e����|�� h�%qb��mM z,�CM��(ǂJ��{��o�.����5?V����s�B������<�"�M��0�ݼ?��.�K?����5kK�K95ı�.`gN�6j�}��9"r3�%@:�������i�ۑ��y�i�Y����GvHI� ;+�LT��w8��ss����'����#I8���D��T��!�4�4�\mκ&������n� k���Ja��.[�m�k���~*T:~�S��[������3���5 �s0eJI����tp$|��o&6a
T"*~��!Ю�Y�[�z��Q�g�±�)�G���sqn-;ҽKl���)��X�����e��� ;�D����{�������çq���Y���1���`wqK�����S�}�j�Y�+�}� �u�d�?u6����l�
��?7�O ��%����G�:���B�X'D]�ȏ�_+�.W`���OG�_�hYӥ9ٴ�:Jc��q�H�l�c��q�v�k��R�]���h�'��8S_kt�VF�u�i���b|~B>��㐖6wƦ_�4�g���N����ޡ�!c�n5�0�v΁���t���T)ş/:ȶ)/�4:�T�a���S�'�"Ũ���zy�H:��)�� P�˵� �.��(>��|�P��	��}M�m�k^]}m;����"2*�X��o�d&Q���'�S�m���"9�TG��d:pr��q�L�Q�~�7u!���*��!(���i}��A��QE��]�>.�5|:#9�a��M�� K����lhScH��p��b\*��6E2=��zխ���l�F������W�Y�T�U��s}|G�a��Zv��Vdb_�Ib1%�-k�:dE�H���Q�I5�Q��`�C�Tr�U��w���\��f�����x�:�n-��Ї N@h��hק� �H��?�\|�V{�U?�sa��k?����Y��0[���j;�f�'
����ؤʲ�"5Ӝ����%(S1$�j�!�F0��TCF� ���1�E�ϡ�^_	�f�߆�f��ʽ���{�Vڥ�{z��n+�&�f��I�n�%hO��;lG�;��BF�"�q�6Ң���16vQ�h����9 /�ȓ+H��u���\c���,��k���'l�WQy�id~>
�:��W���&mGm��u�KSK�Ù;���˘�yZ�~�����ұ�!�eo�����z�>-�|� s'�NeΆv��U'�eX7���ƺsf̘��b*/�6}�̣��J�y�q㉝�vT_|2le�ؙv�bv���z_@j�f,�C_� �����m4����]K��������k����n��A�нm��"EV��r�`tE�*H0���!eȼx����v8}�K�^�. �ϳ��F���յ4�⻉�O�>q8�v�A^TDz
fcq�٣0䬑��(,P�X�F��������$���ƄIY�l�
�t�Ro6J�~�0���פT��y$ZS~s��g���ԧ��#�z�n�X'v7gy>$���~���_�(�]��bT�0�2�%�ksm>��<�	�]��%�|�%F�p��삏 �[��$��U	 %�R��6٨�QVجg"t�g�u��)�3��w�w�2�T+t3��>��U���@����q�c@���?I��?�蕻�����$�ѓ����rz��_9t�7KČ�AJ�;�� �vc#��i����ť�:knAz����%�=���yt��vM�qE��=�͟���dĲ��s8��}��	���S\o`�Y��r{��8��O�w��RT�O�ÙP4r/�
�Wi�D@#�Ak�jMå@��0MPKt��E۽#��!Gw ;�]��7���{	k�4��<\��sU;��B�?>�B���>E�y?�i��)��L*�kz�И-r	l��_�W5&�+Hj��ډ�8x���2$u�bC*�p��E<H`��n\�I�Z3���	���)V}Ct�SO�^�82*�����C؍Q�y隺7T6�_��bL(u"���WO%��؁bg(�(?�kg~����(��me�"�Mi%ߢ�s��q�m���^�������'��LM̿��q]�l����V0T+��f��)�]��n�q���:~-�$��p��=5DS󢄾k�wtVp�,����Gud��߮}7-4Y�26��� ~EqlOZ�߮�����}�r���ύ���t�W���\�*�a�����))�3({��ʮ�+j��7�o>�P��+p��xT�٭;#��ך�}���2���L�8�L��=��S���p�)�
���і�+� g��ޚ��g�Q�H`5رE"�"*��Ҙ��D�I���ɞ�m�5)��o���|�] ��^���i�;qL��Sq�y5�'za�
��=�v<�T����y�X!�(0<���,����ܣB�O�2=���g��7���b|�s�w��zSMYf����O3!&]@��Gz����^q���
��(c@����A�z���x�;E�%�07+*?,�hpL+�K�D��9�Kʯ��UNa,Ƅ<�6�z���r>-z���X@Bp���RG�-d��>?���7��(블$��y����fP���/��[|Bvb-�W�۽6�1�/Zp'�㵂��*����t�1���OX�oO��8f´�.՝���]�e�.Z���1э�\U7:�#��o�q�	Pu5��S1�h
n��ũ?s�~�	�i�J��%S��'��-�_�(Q.�'!U`�#譧�6c�0����[W)�f����N2�j��=>��u���"Ɖ.s�*�9�h>b�K�>���^vn�\"���_��,���m��hUJ�A�]�9 �>m��+���L���]��c��i�Z�����~s�Ij�3��D�_�^�Pb�[�W,t�r*���R�_UZ����'��Ko����	��~uό)�a�)�*"�b@!%�州��g���~Ǩ"��K��7[�0ȓD�%���>�Z�Q#AKȣ��?�TTL��������"oph�Y��`XOvu�q��g�.��5 ����@���м�eX����g�[��&%�.oY�u�	[O�4�Q��+N#.����Q��e�Q�i�G}	sX����[��>N,��y�������g-�����	���k.�|Az����"�r�`�ЌZc:!h!Fw �Wȣ!���Lӫ���J7���1,��o�����R�O�ɚ,A$T��v{�Ϋ�����]\��+���(���X�7;T)4E������P'M.�O�G�g�����o.j-�ՅN�(�K��Ě.���*C�to;l�9:Z�zߺ �*'A՚I�g�ˁ���Q�gg�lP[۵B�(���v�Y:��R�C�sCB���^�(F�4Prۢz.Z�6�_$L +&T������d�"x(i`��U�r���p������"ֱ<���ݝ�/�������Db��q$�S�U�V�y9�=��ga:t0����H��D�YfG�b��t/,\�NsOm��Ie�����x}!ݪ&DF���7ءT�{�zd#�$�٣?.^q�v��u�ݎ� Ԩ+����Q�C^�*����\tf���Z��C�X�Z��Ҁ���jZ�
F�Q-3t�@��L#��8/��0!�J�x* V\pe�H*�\m��d.�@･Z�%:�њg롔��ͪ�Ǝ���+�QM^���X�b0�{}�J�㠁�J�ז���Ϧ�_� gY4}�V�;Y�E�	�BXٲ�,d�e,^#Ч�J�_� ل���p�E �@Y��I)�$����JM���X+'�dY��Xm�TxO�a�[���"���5�Y����:Bk�s9+���q�B��@�S�Bÿ�h��nt/�����3�w�X���Z�:u��t�ڱ��˗��} ��>��V>	Y�c��d/mO�d&�C��^-�#})kL��B��S�3%�_��Q�u��! ͸�m?>��U��UxKc��J�H�h͔��2ƛO��ԝ$o �c'�(��"Hy.ne"�]ӭD��930�����`A���=vJ2���X+�䌋p���9r�=�BAO�v*d�J��V�(��� 8�)1�X��(T�[��{S�Fd���nۦ:��h�,���5��>C����=��>cB:��5ȹH'�=4i4ǽ�P=q����:K�:�A)#L���Tn:���=6i���@��ڞoO|m��΁.R{�a���
47{����V��K�V��>)�)�jE���1����k��5���*����Yܸ(�y	�D�Ӳ/��+�.}�_B���{hs�n�\Ș�gR�]��������9V*�@�����oW����D���}����w|d:J3p������M`TH��e�&�J�=��R��&�9))�ȏ��샶��I�7��z��'����7�Ă8���O0��Jƕ�F7_.����nK��{i��v����������hY%���#�Uy�t�U��o�X����϶^�B���L{Lh�����<^���&��Gym����%�ጡ��߰r��S�/�/�6�����}��o��G3Qhdţf�w�Sà�s&�#�5�m::݁o�)�k��^/��v�p'��]�L�����m6������ �� �$m�Ҏ��h=a�4�X�Ю��Y�sڹ	CV�5>e7���$%�*��4��6ߺWPTw�pC&�ӣ�__/d2KQ�L�ʅ����m�`V�������5fn��c�n�6�����~O�UX{Q��|�Γ��Ȍ�>	d�ZL%�x��A6s��,R��X [�����7��ah`o=��.�fx�����ޞqۿ}l-��<ِ�w 3>0t4$V�H���M���`Qu5%"�/t�I+�h�ʖ��=�9��I��SlJ�:l�U(��i]�����mH�RZ���_ˣ��Qɍհ�i��ӏ�VN=o|��}wԈn3O.�W~��m�dV-����P��0Dlp����G��]�L�)��禷e��I���C�Ӄ��$�{��e����o��p[�m|���_"���շ䛺�s�d-�AQ��P&�b�<O�ii��Flɫ&AN��e,ha�����e���� M������jj�_�b�a���l�osQ� ��\ǂ��xpi|6�iW6��7+��u	��F�����܋&^�HJ�|��^�����u�𱀈��=�}�>~�Ð�MA�b��FI�nʓ��� �^WkHНz�N�&-�{<d�)=P���\��}"�ː� $���1"�s��E�4�]!�r�6�ϻL��r�L��<Mg�F�e���0�qм�;Q���;���K�Y;_;%+��/�D-�Ejwp�2]�]s�w�(���3�ylh�5�rH�k���{���c;��6�8�!�x�=���ԟ C��³sn�$��\����]��M+#ϛ��nVbuQ��S#���"7��s|tL�H
���%0�+����a���#be �`��4���$�뫎6��T|U��s�f��5.zh��%�����/=w��e=��o�6Y�`��h��溄B6U>-����m}91� 	��90-�Ғ�:r��Oj���%�g��mh­��E�p��?���hy*��ɦ��BgO3]9�+��;�ܘ�ď�Of��PH��ϯs��|w�ڟw) ��|��������
!�Nv!���(1�$ ����T�z�8Ώ�lE��#N?ffp�\\Aݚ�X^�B�ִ���R~�mL��2�'��f�%�Xn/LW�FZ����2q&����
C���S����ß�6ԫ°goƉ��X�wS�Y&Ŭ�T|><�<Ttw#����^���F�q��A�J~��?m\8�$��~gG��A�ٸ�B�ܞ���o|	O���N	R:b>��E��٨������,0�D[�&*Gd�P����c���x%[3��9�u�c�$�Ę�a�����9�tRS��+�Vx���$�Zc�8k+v�Oxl%�BP#\A�30���S8�&2B�@`�B*�M.���u�d_(/L�?�����=3S7��M����j`|}�Z�D����;��\�Z��'���SN�@���j��f�(0憊)��7߼]�K/��`����Ai"�H�ЁB�K���i]���H�_kD����vqjP����&797���0,��Fvp�߮rđ��%Έ /���"Gm	0��b�����2߫ �:�N�~[%N��w+���ÛX���/�2$����J�k�Fy�����*{�~bCQ45������a�����b�D_���>�b%d��\�e���d7Z���moj��`��x(�H��C����?Nc�pY]q���6\)߹HAhQ@����f%5�J��{ǎ��Wg��M$�������l��I�R��~@�kUh2�e��OU��ѼZCr�]�����#�7.]ɬU��R͸���J���f��Ӏ�t�v��%�`�C�ԕԅ�%Cu;��U�(J��S:=^�^DD����e��~� �(�uk��
f1��Gav��hʺ��%x����o��93��:@3���!q4FE=>e�s�H��Jo���P���_jJ�E��b��;��8 ����;<�8�L'U��|�i�X�m0��*�gA+w�w4��i�G�bOs�"[��f�'�I����0�a��1�$�5".QD11ZO�o[o�u�!�p���K��ոu�I]�s�s
*7~3�䒰��!s}VcФG�#p6m	�ن'/!����$0=���C�ɞ�{�c��Շ�9���Xܥ����h�<j@�-���Z�$���,L#T��.@�)��{,F��@ij��F�o0�wɁ;I<�p�	�x--�0��z�r�(�>��6u�e�dD��7j�d�o���Q��o
z��}8<�����µG}�Z�k��P(���s�ƴo)��DKm���/��o'����`l{w��u��u�KJQ������-�d�l�������X̃��K} ��a����<���Oܬ���"�2���9ի�g �$'+?!��;��g�Qg|`��@P	�xV��p�{�-7a]��~q���+X�iY�^�Z�5�O�,=��� Me#g[��"]��-ڡ�PFh���nԩ<72_a�3dN6� S�g2��@Af���~�=D%����E��Vm��m��@܆.�3ְL�oj�D�Nr��O$gPsfQ�akZ���AX�琲��/;`���W1céD����(B�e�SGNR)Z�yY~�.�$$�����oI`W+���T��4��9���g�b=,���[.��B��e>ʩ����3�����$��dQN�_g���#k�κ��,,�n��;�S7�f�6�3D!���j̗%�{|o.���t�F��d�:;천��S!����_�&����>��]�zߐV*�$)/!,���+���H7�u� �M)�鬁�dy�F ����q�b��`�R�ICS�h��P�<�CW���@`�C�,}𖍇�Ƙ�//��������^�"P���s���6%ْ,�>�`�q�W-j�f=n��'�����q�B�PG�У_�O�ޕ�֌? ;i�Da�xe;g�K~����nD����8>�l.nÖN}�,���pt��Q�[��c7��pBV`2�:nb���#��HLt"�(0�spZ�b*@�`�}Y��Uw�[w�o<���/f�h��P����Tx.�;��+�%sX�<4oր����KaD	Y��ߡ��.��l](�"ue�j	5P��Jo�ݑ����(_.���Z��A��T�h����ł➩�i�� b��_h�'��~V���KJ�i8��5��~qv!����+TMrœY��z��8ՙ�?�:��}��!����;ۊnz�1�^(���L1l	�� ? �]��[�!m��`����bG��*[�{n.K�V�[I�ڏ+��iX�0h'��/,6�h�s�$��ۀFQ��R�l��Vs�/� �O��U~&B�}�`l�fW!I��C�j9q>�5ܴ��y��ÊX<#e>�� �� �4W��@�O���y5���w��*�Y�9��:�3;�+�[8C,._	V��1�����9�\��bSLsu�VB�0~�R0. ��9R n����,Ԛ���a��f�$����H�|h���V�a%�7����Z�$c�U|瑬�n�ʮr���?f����+2c�a5�V��8�1�妗L��y���1p��q��uә+1��ֿ�$8J1�?<�mV����@�B,�HL�M���)5O�Yc/���?�����&��^�m�D�F���0�I��W's�`Ρ:S����ϳq�S��X��{�y�bMF���l��+��7�2[�	`9�E�Y6n����g�-�K<�$Q���?q���n	���H��χ���=T=��0"�Uz�=t��^/�MRaD���5p�SήK�@�a2]�4~�[�首�7�r}�W���d���p�����O��
;\9_�Q���^���@�ͷN�1���-P�O���/��Il��Mޒ�E6T:ٱ^}ք�{�k���pҳi�,�S?���ס�vz��}�51(c��R5x���sm��������S�yQ��49g���R�(�~m�	)`&�����"}�fx�z�_d���_�$�s�Џ�+5G�cM�z����,��]+mx�)��e[e�]w_���f�U�<$��-�i(���}����[菰N�1���%�\B��%��2)�<��H�N�XC�7IR��w�&P:>1!̝-����m>wFY����ㆩ�Kۻ�!���/2��{wu��t�i�'c� �v�U����Ib��M�j��y���o!����c¤"����w:��O`ȺP��&��O�0�H�Y�Y�V�i\��c��"�LB�#�*�ag�
:���<H���s�u��:�qf�w��(RO�k�l+��L�l�� ���X��-�@�n~L�,
�M2T/T��2��z��R���D��
Mf��.b��Y�ٲgW�9�ەw���w��6�1/ou��I�KN�w��VN�û���0�{+���?V+�-�d������q����u�K��J�=b_�p�Z��|�q�.��̐�*1hq���/q�>�]�QZ�(։����C���K� ]Q�2+d ��R���ɦ�Xr�G��c͂a2���i��L��yN�������bX.p��\T�轓�޻��L����3?���b:�`䴆������S%�A����[�&85
�م�x���n(��h?b���yLƼ��B��/&;�~��6�eHa�j����Ƶ�
��>�O��}�K�D-���-3L�e^��!2��n�w�X~~�6��	&��V�-��%��$սg��+w�:���Ǥ_	 ���7��ح����q%�u}��%�ocp�M'�2���%�[*(�<��	�2�14|��X���� .�8��rC?&����Bu)ڧ�ʅD�~h�p��*�P�ܖ;(!��e���'��Ӗ�X�J/G��t���̭�ߢ���N�Z�mj�����7Td�>���&Y�Ui���&�iqwU����PA��/�P�<Ј�����A]V�Ԗ���gE<��:e�$ð�橩	DPF�?��WF]����w��ߵ����0.��xW�˪7P�V�3t�F.��=i�"q��H��8Y�B���!@y�rd�b��N�]�^9?t��9���.�FK��1�Z���i�>���caw�tL�Щ�s7��1$W�>h��ۧ�Q/rX����:�׫nA�Y�e˞�Ƀ\/�ĺ���0�L���z�d�;�U]�s׍����{/=l�T������n�p /�g
ų��i�e+��x�S��mo�<���E�[��M(�0q��
U��F�V�y�Ubڹx���aęHF��LI�ؤ�dӮ����K� ��\�Q�І ����4l�x�|�7�42��/�mڈ	p��tʈ`��c�/Qr�l����_��j˱+�.�����qb�F�5��A��)]x�f����/��ͼ�Z3�z eʺ��FKA�ACs�5���A�J�<��3�5v{f�N	2O(p���OC�z�:�Hzm�D#�SL�-��D\�8�;�����ILQ�xL������@�Y�lY��n�����/�x�e����T����ys�|�(5�oD�h�FdG����mj���4N���F����{	��g��z�wo�h| ��M���;�>�ca}y�$���p��D�Ft ���q+!ٺ��*�+�K�e�_8�����q�RG:Aw����}�3�@H2<[�և�5i��h;*H�O��_�y��Q��~�k��EF^��W��ջ f4��Uڮ������᫚;(;�4�a(jaPݔ�~�ģ	�ء� t:�h'͊������;�㘮����?�ǔ�]���/��RG��)Q����L�:+�I�,K�I�3L�Մ������= 	`��Dm>d.���d���5A3��E�����$t�h`�b�> \���:w��0m�㲄c:"��wD�X����o��ԗ@�o�#yʈ�1*鬣�ȴ�`�=۶ӻ��8�{�/7ޛm�9���st9��Tg�ٻ�����w������L�jR����+߱�B��'4D��S�K^9=��' Z��p[��Z-�F|jj�ą.���d��5��[�+֕�2���
�7����쁰�%N��S�T+}���F>�:��߈J#�MHH�rHq�!���v���N���C���̹I��l�`�Zx}��@��zay� ��M�Y�FbB���Ho��K��\\e���lN0a�Z�>gr��*&���-Uˎ��l�C7�4��m��Eqk�Z ���K��>\�b�rm�B�. �|�c�	�4�n��' �~�J��iZե��/���C�!J[N��j�4j�e�k��h�cn�.���{�z$/<�$��y#��hR�8��>���� h�<FY��4�u��7�Y{@��􅙰xL��G��;�=\+AoJ'��<�m����}3&�'³�=V.D`�)���B����~���Bzq	0��R� ���{���=�Uf�t/���~TT���eh�lU���Y ��y!鋾A~��u'�or��B��Ķ̳���)�h�k$y�$�WZOpU�+��2.X�S�N;��l@�6j��v��RDG���T�"�ٱ�c�ff���X���M����~���(/�L��6��3O�K���_;�>COL��>�AZ�q�|E�
��L1]�j�O^=��h�S�?�Ke��$;Snf��w�v~�+��Hw��ۍ��Fy����G�S+�;�G犯���(Q'"NXZW���%�$���sT�����VR,*���69'Ϧ;��ov���[�p[�+�n�\@�3�B��n��	O���bwZ�[�-{�_{��<�LƼ��P�����AA���;���j�>��i��<��vS�vZ����$5��p/W6��kչ��Z��]���ّ�-*B��/��A��ʔ�(���o�HkdЎ�|�PX�B�(�ߥ��{��юc*��.���O�o�n���`�:�����w{�9����{�����A�e��ͤ�@G�n��1Dd&�W�t6�شvp^��{�5��WG'&�T@�N$X+�%��Vg���5�	��Q���p|�����zd"�\TOS�3�Y���o�%Ӻ�@�`Ga�P�a᳐gwi� s������%��[ᔌ�a�6M�l7k�(G����֊�RQ��'���&��d��S���k��p!K���k���Үy�>�D�	=�ݵ?��F�k�/(���w���y���oVuZ��7T�(�"u뙝�`Sz�Y����_Egh��=sp���dި���R�����hv�|K���>�ü�3$��G��Z��ïBdjdխ��$\����帟Y�t:x	Vn6��_F�ߝ�7g>%��������C�U1xf�9�/����"�M��ئ��R�٩Y|�7��B|d��qi�C�����;r7�	�r'�$��O��~˶��T0�S�3is�r"�M�VO���MLj;��GU$���/<��^�m�4UL;�z4]���L�9*G&g��s�]��/��[AŽ�=��X����$wlm74~����3�:he�Y�9���NC��AYG�C[�"�:
��C�I���/��_rCSQ3��p��_Y������l�i��ʑ�cX�[�jؕ�bg��,��]����w� ��r��|��W.f�qow�+�r�3����IP�Z�Y�+�Ac	`��w��X���@'��:������	&��-�7��2�P�;�{>j/y5��������C�K*>a��u�f|]%�v��7<L�ڌ�� ֻ�#?y��<f�����b���+�h>�n�n��+(~W��DǏy�N��뀚�c�k��е��n~8���\�N3���Վ0���ҥ�$�nm��G����v��(n�&wy�l�+�M:�"�b[�a���E�����b4�W�y�J���������CVko���F������n��<;^�Ul�TW�^�����vÚ��Ki}�G7xK�O�/�S?5T̮��tez�/'�9n4��ޥ"Z��4�,juG����[��o_�6Qt���I���QBK��n�@��P)���;�-�����7�N��r�z�|E��ܼEr�� &s���&���[�I��xW�gj쪺�B��B�bc��d����srx݆04S������#i��2�+ڼv<!��6�.�� s�$��"�R�v~@rF(T)38����i��'S��koqY��(��B��{ֳ��~�����B�D��m>J�Oi��n<��=�[��8�VQ��ȗrᓧ�N...��l�Z��Pڣ��ߓ�b\k��aΎM���U6Sbl� ��C��<zJNu�t�Z���~�Lq���!��2������ ���	�{������z֮ĝ	x=� ��U�5NEW4��w�������s��`|=O<��h%g@�cQ�:QRkgiӡ�DWSbQz�BcΘ=�J,��#>����RM��ר���E��x���	��@p@sʃ�[���AYW�O��G:2&���e�ԩ^���=Y��n��K#���Y]M���J-�����&Bc+��rnK{v_��I)(3�?[m#K-l�(�1��A2D%������G��6�﬽��}m0ȥA�N���R+��"��Pp����z�`���a�!�#̡��2�^)یH	�7��&lC O7�T(�{B�3k'��"��6��p/_]���@.��Y�RXPO͍����[��	� @��CX]b:��[S�A��I�lK���[�I}90�mZ��I��s�7��CG�V)x���|v��u��(�� �sT�\�<c��-��[H���bP���'gg3.]�&ڮ�M3~�0�#4D�Z|8�vkh@��8x
MK���b�7�[��}�]jK�řGw)jңAp0��\�3F���&c=����#����-}[)��ckGş�T��sq�h���?(S�u�~�����Vx�U��t�,�,m�8�B)>�t2�g팬���yƅ�U�S=H�H�Q#���G�bㄞ�����42+��`rYRP�b��%2���ZM�� �Y���h��q�:�U,bܬ��q�d���v3¼��9oO��V�djC�`����P��V��h�Q3&!ѥV��,=�u�F��.����F�8�����H糟U�ރӾ��"b`ʣ'�<�������L���]�:v���aq��� ��/&��Q�����i{��!e���NHx�B�S�pg��x��D���!��]�K����vh�)@����3[^"�;A�~)s���h'wkm@�5�Ǧ�+�D��� 4����iv�x�/�/_C�͛�db�u���|�]�&�V�*φ0���<BLA�`[���{�6=��r>��}qRjS�'�E�m�����zZP)� ?8����v�C��e��5�EQ�'m\$k�/�0'Uv:qŕ�x2v�F�T�� 4�:�8<�Ҏ@�z��?$}��LCHq͒�-�?��Q�f,C�삖�6��u���/`PqRr��Lеp1ߧ��Az��@�ĕ�����%��������GW�Ru�g���Q��L�Ɣ��xyL�W������9f����c��\�ڬ� �cn�ֲ��oG�ΛΗ��?4S�s��Т������F���e�.�����$95����o���g3�Ux��;�<Đ
|r�^@C�1�N��w�:eh%#�S���*��Xt��@5�?b:��6}ʕGun�kh�-�("��-��O
��	z#)�J-!}g�#�n-`x@�mQ{����<< �O����AC(�d��Ck�Zj271�����)QK:C9�,|�*㝏�>��!����z�㧼p#��`�c�_���<T��~Wl?&��0ʗU��O�bo���O�ͭ��Kmx���~B?��Co%�k.ޔ��X�-�j�	�A�\ X�+��J�L�^�+�=��m�eFG�s����B3	����Gy�B<;��w�����d��B^c���mGs�7�>�T��5ODs8�fŝH]��s�S���-���;�a�������x��Ӧ̕c���WL.o͔�w"��ӏ���[��~�����s���v��n�\�����0YUVk�ߎy��SG��ĩ�t3|64��4�OD�ń�U�F��hq�l�mN�!��4?y�.Vߊn،H_	���dN�8��x�9���u��p�'4e�ERs b\0?ʱ�����[W�\��c/�HH�/Or�N���B�<�d��b$ϣ�6��$¶�������vQ=� W����KVQ���Wp�
��./�:}�Yy�J� ��27�B4��$�L�1��z��������mK��+�Ε�T�)��Qg������9����x��\|Qh�w�\�IF	X�2�� �"ȶ����;2;�ˋ�g5��i="֥	��Y�
S!����P�ҮP���ӫ,n1Z��aƝ	{�s������H^��V���|D�3�R�>��vS��w�Fy�\�.����φ��������JF�H_ʚ{-��p�DS��!�qQS�ή��\"{*�^�9F<e�=d�&����X\aU�H����m�>L%44�0�Լ����u�.$b�0���HD�>*C��f�]?~���F�k��y��8\�K�>?��t�T����k�gyM��P믥�#k�x�:y`�:�A�F��mxи��3�#�U�x}�H�z�� ��`��,��W��տ]bG�7)��w���ˣ�Qt�G�B�O�ۨ�4��W�#�_t�e��tB�����y#�.��܄P-�g�������ޡXf��8�EmBmcr�7�f7�cW�R�VP�Q��{���s�8�e�P{1#�㱅�8�&Fz�B���(�6�ȯT�="���B6
�	L�6�C�-���|�і��k{����N`evΕ�h���o��ܬ���adP��X�v�4J17���H��׬�ύ�-�����M��Hɺ�;�R��������!M0��G�Q�/�m�W�E;Fx0g�8����)��|�vo�_|y�7.9�>Xe�>��������1p�R�@s�������2� (�b@��XP���1*O3��=�_	g`��ثQ?��F+�Y��p����0�*�%-��S����F��/�1w�^�N�F ���䔶��`5YcY<�)HnO&%��Qs�q;��km���&(���2�m�23��N6��!v��1�nm����{UIT�a����M�����;�BP�4��˖ż��N� ��+����^t;r����p���r�9-a��m^C"�۶Gh�<����!�0M��㿣>����GG@���ʎ��֑�e�C��~�ϙqL5xL�?*�۾/����pYX�7 � q<6�R6�a"��֔I)+G��;mKw���oR�M'�aRZ�-��mc�QWw�@+����Nx��b�Jf�����������:P����l�q�|g�v},Ϛe�1]���e��g��������b. ��`�8���ۋ�(��R������
�Hj�/Κ:d�c�C���cc��tr��{�y��{��U��&Y�M��
���H����9�Ǎ%����n!N���#Y�/���] j�1�,m}+��:}[i��)�)�^�C0�g�><U����!hT���+�86]��6oE'm(i����J0��&$��X�EV��D��ޢ�5�HHDon��[����]mL�?���g�߫�{��"ٹL�H}2��ԝT(���Q�)����PNt�����T�KRC����#��VTll�0�B>�ﴘ�B|8NFE���/`=J��UE��}F��c]o������P6gW�O30��V��(�@N��č����HZ~�Z�{�Z"�Vt��`��al~t�
>붖�������g�1/�]��FQ�-�QD��=A��ꎹ6�*�:VRdEբ.�^�I��e!_������y�6�)�y����C6{E{��D��/�͏b��5^,�m-����܁�f}׀��
���(�䠄�6��#�?.����c��+e��Od����(��L�Ƈ�B ���9$��-!i����
��^g�+��kD���0<N(Dm�b�����X~��2�L鹹��Y�RY�$I[�|���UQqj&*�=�)�g��(r�u�UE�	�����x5�G��0�HЋ���w�X�֦}#�`��Y��>o|q�I0��F�?��4	��5�������xG�7��RJO�A����s��&�vG���"�}������`�p(�!��V�L�p���3�q��?~�{�'�+e��-"�hs���T'�(u��EH}��2<Y�M.�׫R�n�47�u<Vih��v2�zߕ1*i��7J� �(	R/n>gF+M�w�q���ڲd١�ļߩ��$a��r#�hk"[��TIx���&�[�L(�rd�s�Q�Xϙm�5��Ȧ�u���l4�r��h�Tt_�W��[C)eט�=��-�u���%~�at,��S)��1�i��om��Q��,p%�B�@2 �(ѢM#��}�Ŝj֖P�\�K�`��V\�R� �$��<8.z�ZJL�Z��2��x�_�p���_uz���H���h�!�����nty�J�T�q�����u�O���S���P�o���QFy�-l�W��I��5n�+���p�J�����ї��,}y�����j0�9���Ɛ��(��_�����{x)���-��ζ��ۏ�:Ю~`���D����T �1蛿��It�o�N����w>[h��ٜ�dpB�9l좀�{VN?Ê�k�_v.�|�i��X��9���V�:}L�/�8cSaM*��-�Vn�r�ɰ�ڬ��T!��ץ�݋�f��h����H
��u�B�"�����q"���'�ISmt��s2�����d
���mK�,����%E|�(���ӲQ7�u�R��}g�%���s���@,[hXq�E�(���$�æ��0�$�D�`�TZ!:�����V�=l�m3X�^�&��N{KO�o���ANU�*�f�,�bjv�=�ˬ�<��V��1@Y��Po��d �$'9����:�<Y�<�Թ��Ԥ3�e֗,Z���f�T��p�[(�v��rk��X�"@uPE�����W�#�IX0=�����FP����@iw`(j|�X&���ŌɌ0�'��������W,;�Q��a����ڋ�3A�7��K�^������uX( ^^����(�X��x}W-Gg���û[H�Z���DL:�P=}�t�u ���.�k,u<�h����O��wR�.	_20O�^�� �fj�K+oG�굉]R�!>P�CJ�?cΤ/�F����ԧ㸊��N�ڕ)^�P&--���0;�:ݲ������8�=x��
!�
	@�[�H�>� �z��=�?냍�=���q;�jԤ��Zż��m���n���{Qn�HQ=�� Q����<�j�!�IG:#@ӊ| ��*�I��Ѹݗk���s��"��qZ�/&�_�:*@h%Lͦ��{����xu����`���w�'*�l�Q��&����IKo ���#yYi����T��/4b�@>t��C����mLa����R�(� ���ϒN�?>����v���+n�dw��k)�w�d�Xf��"���T�����rU2؊"ec"� K$WZ�F)�k������7J@;Ro8a���rȀV���U�_���(�l�U�x�������'�>e�N�Bm��g����c.qԠm�S�����4�C�
�g�2��(6��|%��Y� <.�zL���-��b	�F}֤M���Z� ��T!3��Kj[�B}���D�,q��"_^��e2F�7	ɐn�A���"LƑ��9v����x���`UD��E�B5��?&�c
V3����Qc��<�4"��R����{E���	JQ�c��fozI4$8G�J�7V�]��cBK�-qf���mi�~ӓl�΋ ��,Ha��TЛ$��Ki�zT AM��z�����QP������C�h���4��{�j)�y�����m�����	7��^����ؼ�!/{,��A���]O���e���YB0��"�)[$�%�"�O��#�QF����a�Fʾ!����-�8�T~�_�w�#�n>#�NE��鉒�NƗLASU�wX�=e�(s!O��B�][+�Ѡk����C�m���͇Mʄ�~y�x�������L1�Z\�Rue��d��H�(Xi���rj*�@��e�Z���>�E��� u͆��yh4lC롗���T��]A��X���Dc/���c\�>��אsQ�.����oo?�u��SK�̿�e���R��k{�%�'ˌ�Ds�fI�ȊW�މ�6u���%<��H�n�h[�J\V��2v�,���rhP~�'Gf�@��J�@w���!���\)�+�H�d{f�%��iC�ۅw.�f�)�W��-:zo��'8��d����vLՉ+��Ϣ@�N<Cb� 0������1T<�Q��"�P/dpU�|���0�F8��(Q٘wN�vm%�Ky�H֥�Y���Kb0�}lޭ�f,&L�B�QC!'[7X���)\�?FK����A�3	y�����2�:A+1�d��z=	݆C���b"�u�P�#��IHC$���*6�'�Z�2�F�x�W�N���0L�{��.Gq�U-"� �W�����'e���b~��ƍ��R%{7b�^'�7�V�G�$��J"��5?�]�z�uԘ�s(B;`o9�o����`G�~b�����
T�V>O��cڶ�5�khP�j�oVID43��Z�a}��G�Cj�\����9�4��g����<C��Ġ��C���;ݺ
���߉��߽6��q�GL��Pۈ�3�oE���Dq��w�����2�](IY@�]⟣W]=� C���>��-*��~[���n���Ύ�Wۺ����,�D�nU D��Ɣ��V�N��P����M�?7�GvY;Y�����^�I��E���/Za�ӼG-#s��K}Z�CR�z�G��h��z�}Qxls�c���H�c�f�8�gZ�d�!SU�_���%���(�]�ooFt�$�
�O�qs�YE���cu���A���Uם�hKPo�V�N9U1=�8�y)���T�,�bM���tHC�* B��.�{��J�?))�p���fk*iͦ�m/���?�~����\���p"<n�������&�d�br�&���nt��'�������A��[�]�T3��0�[ޞ�Yk��n� �>�`\�}�����mk;YM�3��ͬ��?����[��zْx"�����tn��Mʀ��`?C��xy���x(W���8fs�}}��KB�]+50c��Q��Y���p�q�~6�ig����9'�����im��dF'�g���j�nٹ6A�һV��m;~��4{g�[F�zxH��Y�0j:�p�s��P�?�_
�i8�����m�/�Q��[\��>�Jh�Ѧ]o|R���{���!)'�[es�H��~�����ԇ�%��wB�F%j:f�0�	.��]pR��#�J&�̩��b�(��z�6}��������a<o�-P�,.8��7f��	��&�f�16\yM�,�F�%W�8<�_T��j�j��q)j�I(b�����@��G��tn7�|n!�C-��ӭI���T��*�tU������60�-��� �E5�.�?�x�.���Qї�5�.�$����m�@���7��j�!��w�^^�dw��FI�Gg�Ú�RH�<��ꓑ�AC��4��V�Nw<�egf<�o�A@��Z�RFx��T͟��F娐^�q�,���0 ������F	A)x���o��C�����d��;�x���w��0?����Ζy�7��
a����h2����ڊ+#��Y4�|��+т�Iy{{��xMw���_9��Zaf��C��ݫ�L�חj�����B?��(�T��\\�;!��Q'CIb�W�K%���t����
�?��^Wݲ�S���t��21���w�җ���9�����G�H4tN��VB��uCmח�kVW��i�s$�p�	�'�r�KkϮ�=p$ԈURx�?�;=~��V�t�� 
��x��_�N0ʢ��+	0X=��;A����Jʹ�-5~���z�s��ZO�U>9���m�Q�C�
A:�6�~�U�p|�|U�mk�D�/DW�!�61	�&�Z�"D�JnP����z�������9�hz�3SvDX�[�[)���oG�Q�Qc�b;��#����φ,��tȜ:5�Ïz��@�<)eop�K!�O^�Vjp˪8�һ��اn������<�:�����d��'�*1@O�}ϰ��Au��D���否��Y��w�������4d�oQn��FX+��ւiU�b�G���� |m�f֓%��頁���~�A���+�qsT�c9�Gk���i�6q&�_�m�`\A��j�=0xr�S�ِ��������v7���(������c���̦�>R��$%�I�d+s������'¥�)Ԛu�T>����c��l�ׂ<Z`���&�\�~��T��I��b���ګ�AT�]��;;�16��ԇ�f�μ����hk)���U�wd��Q�]�1բ�MO���w=�H|)()ފ+���(��V�-��Ԓ�;��������t?�3.m� �Z�20�_�at�n��A�?'%��#m�?�C�<qIwh��u��\e=��	��N*���v�O�`��f�{�-�u�}�N�\>L�����@��hV~�u�3T�C�^!QzM�4�F+��3Eށk b	%��lE�K1�z8f�ۖR�2K[ηz+O���!&��k[���]��&��
K�OX�&�hAK#g ��j��れ&��z;H8�Q�_�4*��k�'[Y����	T�򼚒�L\��j�퉘�N��?�RG0��4T������hǦƺLᇣf��S��M��`9R��$��s.��L�ኣw,g�f�EL��Y�H��<�s�Z� �+�n+ZD��G�V"LBx��{0t��hS�H$��\u���W9;/���>�ɒvķG3-���}���OmGCy-Q� S��u��Xw~���?lX*�w���!]�����zp�~T��<;�}	��۱��ܨ�����@�{S���qzD��'_}�q��`ڋɵ�?�ԩMʷ8��L�2$ �m��g�����!zr6uط`�-͹1�o��sl����t&�ed�cᮀY���JP��Dl��Z�ն���*)����r @f�9fȚx7��Y Y���2��CѪ�
�P^�*��op�B��jfPײY4�U�ۻ�r�$�"��C�|2�u�Y���z�D{j�����u�#��ݪ��U�0� p}���kp����aA;PoTs�Q��W_�ܻ*:|��y�LU��<g|���Ɇ)�Y�q�e4vx�!������:l�@^��[�egS��t�,T�{G�I�`0���i�	<M�e�m�oX�uo�1�@/ߣ��-) O�m�k<X���#G����U�$��BL��K�Wm3̻~`���r�6o9.�LŢi_W��_r���˲#�mTz�ܙ@���d����J��+RW�j�0�� ��险qCm۰�BԸ���]�i�v���=�[��I��f��k���H�F�*�4sȒ���&x���Z�b�f[�uV�r7}��©�XUo녀6��w�#&)T�3�����}>�H�w��N���t.A��D|�}�#96�H��&�~�4�$p�i��~���RE�\���s�Om�����'ըV���T�4㡺H#|y!�3���c���	E��iMIt6G%��F�H��e0`ŋ �5kD�?@g8�#,F�8�&YS\x%"g��sZe�N��v`��`�z�]R����`��0�5�(��麱�M��ALs�-������(P�����NO�1Έ�	�&#(.��<4��c�����͉C��	��C&r-�(
	A���le3vr݀�%����z|U�c���zq�<,}h��8	�i�ko��Is7���f,��qKv�}������؆���'�I�s����A�v[�E:We4�t�+��e^"W�zk�)�F�pM7�:�}��*x��l�̽�E� d��&��c.��"U��'����<I�_�C$rW��ck2�z/���қ#��Z����?�����+TM��+�Q c&�t��v��N0�D�GZ>S.�K��&�;�PdL�8u��ǖ>Sz��4���o�X ��*��̱ʼw�Zj�2��f"J�̩����P�æcu�})Ϥ�O����>����?���2j�3ʩ�ßa��n�/��*}�f-�g�`�>^��-��>������2��w��驓j����5)Լ��7 ��3E+�:��r益�}�I�դy�!ƈ#�%x���(���ل������B���T�,C�-���\�⏈ڼPG���������|
;ɂY6�m~ku��3 �/�A~I֖�/�U��uڿ5{�_��;��"���΁�h����"/�h��酥�� Y�_��&�����X��E��qSDM⳧�۳�X6�]h�|�[���f�5�bq=�P�>#���`�#��b�)P(	�hR��R�&��M��w���X������3{��R}�DR�Ax�.{��+�#�OH���cVXby�s�4�B��-$�4tiJ����+7	m ��F|3a�g�/�8�
���O*��R��	f��\��0��%��j#E$�|Y3Ne�|o�j;C��xT�\�e��md�[��� |����qc����z�Д^�^]Ԯ�EKY��فz��S/O�
_�ۛ��������V�`����T ��T�����>"M�&�Ų����*鍄5i��E�f�}Z�m2�8�+�r8K�:	B�,�,k/��eu99M���X0��ns�$[�G��G�6�X���z[�lȷ_-Yot䃊GI��6���i7����� ��|(X̹�RWE�4����z�[d×ȏ���1�t]����-OС���Ñ��0Go��M^e���5�c�L���D�I���n����*z��{3�8p��?��e	 ��T���]�hZ2K'�Xr�	i�Į����H�^�%Tr�/�|]˥0 ��z3]26P��$5pg�O(0��b}�8)���ߴ�:/\n\�����w���\�Ӡ�(��L�B�Io���珽ɉio�ɠJ����(v�{����i�M�yG��'"L� �4��z!ﮆ�$���o�Fg�";B�^\ߎ�j�K�n#ɇ���ސ\_���i �����w"d`�i$�+ju���^+5�Y&r�Q��Y9s�~�',��;�}kJ�x�\�qo����R�&w�o�B�;	+�E�CUA�0g`J��j��T��8�����K�(��X�!�S�osL��s�m-�.�����~���$�,i��궵2�2/�۾���[��}���[^㶀�6�E�l�;>_��́B�{U�炈�ON.���+XQ��&�K:O�!W��=�H[dz���<&��I��a��o�\�b��@{iQ���n[v�J����@�yܰ�^��Ĭj?���ɑl�k���	I��@�`$IDZ�9?r��չ�Ԡ��6�"[�(fH��ƆzA|w��|�� �R
�\����������LD��1'�f�� �-C�I�};@�a��O���0_��YB�i��Z
Tl����!�I��A�>������"�`�F~Ʃ��+�'WmC�Z�kq�mt�j�#%^�� *}�:ߤ�_t��V�3l��哓�����h.Du|�@����,D�RT��HZk¥[��oA��295<8�ǻu�9QC�,�DH��>^yRa�ig�DR&m���č���x&��"�^��(��O�QF�Hc'��;��:����Q�A5��OJs6
*�	��]m���Q�hk�a�\IJ*�X�P=@`����1�̈�Nʟ�iʦg��[���{��3P(��DԦ�&C]`I�nf��kH4��bs�&���B�İ�T�ɫ��l�����&s]��}�f�I,��"�/EA���.�5�� rذ4&�F��x� ���Y�-q�P%r����/�^S �iF0����0�V������`�]�N+uV� ͷއ:s�	F��M~�$_١Sk�mQ� {�*qx�=T������0�	��eS�eUd"�sŀ�M��?9���T�h���D��Gn�v���tJ0a����*���� ������]Yk>j��4�1�ukCǒꥵǖК�N�,�`�_����߯�|�$o��|}�ǜ]�Dj��r��n�i1�ý�,WqUM�xI��;s��(�	��m�?��d��PS�S���2���40~dq�Ҝ��E���(9�Y�/驣V%A9/�F�qu�J�&*�O.XV�ژ�'?�^>�U�T&Ɖ3��`�	"i)��kC���c�r�Kf����Uf�r�b��k��	��)��&&�!M�n%;y�1��N��U�T\#M0ç�u* ���Q|�LS�6o�h���8"��}x������D�(I?P��J�5���Ʒ�n����DBY��v��\2�j��2�����xuD'�m�o��`]S�+�/�L�}���Y|Q���cM"�Nh��"�Lo���H_Лs�]���Ys��`,pV�j���T�"���E�����\b�XF<��v4Ą�P�$~{�i ��)�P�����2=��\�t�ɩH|Dn��kau��䶅v��c�R�V�3�ؔ�}��b�����L�Za�<WgEg���V�%&�T��'��b��:�w�F���B���w�W־����u=�`�j� ��Y���Y�@�cǈ��9�	�:�Z)y�a������2�b�Ӗ����,��~E�ნ�|��.D�;�Mg��R�x*��=bm/YC-?*�c�d熵�b�w�eL�(9���K�f�[8�>v�����Q-4�-�ӟ����r=a�;��iUM��%���4���ٸ�0�@ҍ���#�m˃���1��G�H���R�M�Ok5_�ʻ��k���_�l[���!xw�K9Z��.|W�;��2^(&\�Xy�hfLV5̞B�
øVd�#��gı>�o�$�Mv�v������:���蜅��ق��+�-��G��`�8X�|C�-?6WY(sT������VA�h�[�$�)�w�u�x��?3�zVl� z���������S���v?L��ei�C���QL�Kf��r����z����"D���)@k��]��-L��
-l�Jr?��]�>����a㹮��z(�#a��"�/| ��M���z�Bz��i�1�V��N���+�A�{���ʬ����SS�p�J	�K��Vv�j�u���R����6�_�2$��X�P	m
��LT�U
���/�^�T��sU�}쿷�`E�߉q$~4���sK�U>-Υ���Oӻ�g8b���4@V6]�z8���䧕	�γ�s��_�lZn��#o\��� Im ������FT�aYw�_W�����,��K4�Y�b���=�u ^���9��,�1�^�7����X'����j]�����AR
4��r�[mA���������F�7���$�:�3���vO[0��#��b����J�r)M�����2'�5��L����vɤ��;��@.��g<f����>��
�����<�9��"��J�(nk�����b�:���9}\�Z�����(ݐZ�d��?�o$��Q&LH	�1i/�qR�j�����/�4�!��XO�d�񾸖�0�^���2c��x.�2�D	u��Q���x?�'bX�'�<�`g�����f�F��{�/h��)��L$|u�ql?[Wr��O��ԝY`��+ \�lmux�Ó� �h��P��<vIґؽd�揈�P�l������/�٤ ԱOF��Q����/٩��ľ ����F�|����+G	��
���a��ٚ?� ����duDj�:��RA��ڤ���z2s��pD.A�T�ơAr6+L	��7����bW.]=�Ձ8O�)�Q���6g4=Q��i��;��^a�ʒ��d|�:��4�pE�u�����3z��Z��>�8��gɺG�J��]i@T�'��E�2� a������e��d����}��U�֬�J��Oc�|���³l&�V�s�R��
���e��چ,�V�u_�o�����+_�B#��U��^�����pj�^E{�>���5������d��~1�u�a���^^��h���8��	���"�vt�wP��N�U��Y.:����b[^%��	F�Gqb.����G��f��/��c���~��vvH��<U�n��~�C�ܙu"�|>C��k�jx�`pЍ�_5��*~��  BӘ%=����'WGBF6�b3��[�Y�=Sg�`V{���`[�|.���ǳNne��!�<���g,��&�4W��x>٧i�O�<��.y��Ҵi,+.~&��3?{�F� ���m��f���M��<��x�^Y..�aJDo�M�0)rKQ�W7ڤPL���x �؟�_[Tv��٤Wf�p���X��]�2���ߣ����t�*(Di.�`�`��hZL2,n!�p/Rp�*Q�E�Q��4oQ��B�9���J[;zP}�(���تk��.�CuO��%�����V�k�J��S�J�Z����
��,��u���G��t���5a{Z�����L��5|ӷ&���K��VgK��z���q�A˺�2O�����Zc�m��z�Ӟ���İ��5o�2�-hO�$|&�v0�N�1R�����V�PP����j��o�=�٤�g���V�����ݭ�ue��� ���4ũ�Ҍ���a�)/�D��)ӓ�0'���H��й��o��#�l�~�h��ς�_�����@�==$�������_.r��C:�$��q�C���[�.�]%�'��Cy�d�#��x����^��`�\А�K��n;C�����޶֔�
Vf޽�� ��*S$6*U�����Lp�2��r&m	���m��z+�k]	�ģ�Y���6��m���X�[L�̲3��m�0[�|6�:�M�h��'g�m��=Ja;م:W0/������t����~^cl�_z*~���L�b�&ZiC�8c$������@�>�S~.��V�TV�R�u�I�Sbw�� w����!`Len�99'������`�,~/����@���G\xn�n"YK��%��/i�e?��1���>$��0_�g���e"]("�L�����\(���#X״
 z�x�����nv���n�Tx�t=��u0��s���f�0a�e��m<B}�7�_VU5��ji7l �Y�f����ЗZv,��������Q�C��Ub�!S��YO?:&�V\D���|��"��b_�P�=��|���&׹!�F��拄�A��1��B:5�v1І�A�es�}N�
Ȩ�N��*��-$��& �-�$ �����yZ+�`�N��PRى�5��N�ד�$�e�[�R~:���.��"����dk�"��ª)܂��0!b�bhW���B�o�r2�,��h�!e����僪�=F�	A6�J;�H�;�ڜ�6���0lX| ����8� x����$`�l^e}a1�/d^�ᖨ����S�m����ϻ��!Ժ{�|0ѯ��9&�,w��y�p�ˬ��<�V<w�+-�j��Yh�ĺ�m�τtӀ۸��$�f�A��+�z��U���(��/�:9�ѶźvX�����P��h��[ ���f8������ǐ��^�������x��s=ͺ��ӹ���կ`�D��Pцna�8���2�X�UZ|X�ro��Ɲ�=xF%�!_4!.���s9�3��H3�e� 쯟bnՐ����R27�J�k>>��p�@�䢼��m��ہ���S=��4��l�Q>7�RQ�v+��ªU�-2�� ;;X�F"'��^�*ek��̵������E���j�/#E{�"�$
X'�,�e�ܺ4�D*�D0�n� �4�/2����<b;�i��B��Y�Q�.4	�X8{����\526��<*��7��Ph�	[�n\���3NBq�h�y3��F�b
R��z���=�.�S#A-�$Qe�݆��;Cˈ��I�}����)K�v7B�>���V�sU��:��X|��2,p��W���ޚ��ؖZT�{�*�vw��թj
�Q���0Ú�����S���V����%�i�Q�������[�v^<�h�`O���.�%h�D�`��q#��G����~'�`�Iy혞��ۤA�@ ԁ�A��}�(U��T�1�*�Sy���r��l�YWe飭#O���鲯rQ�4�v��ؒ��~U�ըo�'�pzS���4�.ji�+���ղ����÷}?��^s�{��q�#���Bֳ��[��9����Fnk����{���B��E:�����A�w�G��ߢ�;�E�[�^��~E8���N �t̂����W���vzq���G�s���n�;�ŒT�>�m����	��C?�
C*f�"~�m�F ���ݼ}Yqúw*}��=�g��� �ю���ƬZe�o�s$��I�VL�y3���E���,^�i�:w���"�Z
_%���@X��ihvC�0{ܨ߾���y8c��S�y�Va�YIY3���ZEq��.�Z��R�F�ʎ�C�y����t�_��6�VW{y�����U_ݞəo�tu�}q��f��)�BD\mӱ��!^x�Nś���h���&�Se�z���<��dї(e�`�}�N[WVMً� ١=��Ѓ*�#&v��KT��BZ�o��ͩ᚝�^���)P����jTJ�M�vw�	�C�n(mg��Xrȋ�H�=c�A4�Xޒ�L��{�	a�˼wýӗ���J����&0+P�`���cUe�Ix��)��(��oX%�y�P)����&;��ShL�|�����s�8���.�OL]zX_�p�n��P}T�B嬚I�qT�!.�l�����O��3Œ����|�V�5d}-�<�՘VT���e�[�1r?c(D4Jqh/��JZ��HJH楖��,â},xXC���p�z�V���t�i�Jl������P�7wP\.���z2�?�DK`��l�nܴ��^K�,��-h��@��Y�~@	0������œ�Ć�L[��x1�4œ]�%��Y�\j~N2:��7Ȫjhw��}�kJ=u�Q��?SW�'�v�K�@�JPp>|��EY�/�	Y�U������A? �S���*�}4�@fs�q9�?D�"��I���Ž���)
/�1�~���ɞ^�9%6�a͖"ɷ�<:�.�k\\ �VŔêIgv��Q ���ݎ�+��^U��7�7�n�2�G-t�3��Z�8���SUr�;kJhW8�*иh��G�%dv\��G.g���ه�m�zgl!��Aq[�����4��f��8%����;���vu歭���[]�Fǅ�0�kL0��f?��FIE�yj�Ъn����¦+�Ɂ�{g@a��2��7�+{0���� ��Uoc�ђ��q��ȝ`b�s��M��>z�8��Y�g�S0�kvW�d�ӥL�X�����t�� " ��(�٨I�:
��`����Ѧ�<��y�����a5��TĘ��-H�W���H�>�>֛L-ڤ��l�ݗ��C�f����'�Z�ǌk�PY�o�N:I�zH���Vǘbw�t�AgH����n�Wv� ��t����ۄvj����5��"r��@���f����$9�h�:������p�6�g��imf�Й1r�0!�a,i�ī4S�"��/,~���*[��y��M����-�
� ��YaNEj�kJ�.o 4(��|&���@i�1���i�G<N�$����&�GˠV��0~hI�U�V��7��a&��#o/��>�Xh�N�I�b鮆?���)yL���c���#0 ��LP|ma-ˡ$�ߤe*Fu�u�E�N{���d|mR簘��O�����Ζ�m�'�H�N�7� �;,T��l)������ ũ�r��D�%7�m4^��<�f>��f3�f�no�~z�\�k�֬�쟔a��S���x��Z`/�L�X��:*��.�����em$� �d�-v�Y�a�)��6��G�4��n��
F�"��J�Խh~�أ�PtH>�����+�BJ�~�9� dE1��:�K�`3��>��S�g/Y+%5C� �Ȑ��
�Bb-�I�u��������*F��.^��2i�iVm�RJ�Z%$EIr���/@�2������D*����ܔ�MZ�z��=%=*"V�ˏ>��$�L���Г�s	[z���OU�.c&�Qe����[�{1�xt������9E��Mc�����"�c����Ϙ�H�G'�}�Ú��=��DƳzJ
�ԝ&��7�=��d�� ���(�Me�t�#�<�ԿÜ;��U�����W�\{,���ۛҁc�܅�ܛ�� �} ��RQ��+�(xn�%Qu�0�,��n��O���ƑW���RƮȰ�p6��v9j��f�B)�֫�"��ݨ��g�����,����NDx��.��7K֕Ǚ��1>��;|�>�*Q�ꁡ [�b�T���(�����fe���<�K�?�s�aM^mM��擯��Ã���<�O ;<5'Aݨ�kbh��s�+/ޥ#3�s�v;�J�'��g?�%��X���� X\DG�gk�Ί����F־˷�	P1팝��7��Xcjf|L�o���:�=�$���`f��K�Bq������%O�����"m�(GOc�i���1��Ko�9\�"��]����$:�&��!��94�����PrfV�b<��4�4R���FZ��n�ʰ�{��t�<Q�DҮF��麺K[:����{�0�C��qNR�-�)��2O;�w��>����g�����s�vYq���&�u���BW[ʼ�F����ˋ��&l��H_�l�F&�nq���/��HM�}
�����=K�"7�(��m����j�7O�09z��.�ҳ"�9!
����{�{2��
�����k�`�Z�����T��@�e���e�,�sj�#6H���h��!��%J)�O�LR�=��T�ϰS�ݼ��0�;�z@���H=(��oT��-�WD�`�����n����;�6xE���n1���J3�F#,z��;r�q�Z�!�J���J#q�dMϦ��l4�yΊK��ڵ�G�LO��1�p��3^;�N<�4w��%H=w�v����~�����f�R��]�.N[�����0TmM;�(F�_��f���bx���r!�j���6 )ȞM>Ec�O�H/k�(vZ�@y?n�+��tzC�]/k3�3�x_VA����z}w ^&�%&�{�T{/I��֝�����tR�a���MDz͑5�+	.*eq�6Ԇd�(�I�l��Z��i�q)+�Es'��x�ཚU��-kH��}��.����������_�h��\I������Kɠ�OH�"@�'o
��\������1��M�v�J�XQ�~��Ȯ6X�@�Q�,�Y�:�e<R9^��_��5�)Ӛe�4���c��0l;����GO-E��i���٭��ao��鰩Qqo���c�~�}$ #7Y�(�	�IuS/���e��`5bL����]��nNq��?����!����=�?h�OU-;¯��x�iw���Ua���U��d�s�q�
������(���s��f�Vt�^E5�G%b�/~>Dv�S� {�#�O�Qh��x4�M2��[��'G�����O*Fh���7L<1�m�4G�n��c�c��� �_T�r���󨜸���G�f����w����E��~���d�F�5���6=K�Ɵ1k7
l��NpX(��Y��������<�R�Q���I���Q�|@x�X%�_ +~Y�H�W�~)h֪R�N�3C�7=$v����j���=�vUݠ|A�s"��R�2ڤ�ˍYo���"K:rIC��I��Q�ʐ|�`���z۟c�m�*��]�O� XCu)0Ƙ�j�w+�`
~�hy��sY�;�7�L�����2��h���a�-����%�\!:�=5ȳ�2'Y��J����v�o��@��)��<#�>��PFd�6�@�w��y���(���]�\��b�	��X���	���Dw���v�?�NT���k9j ��հֺ]����h�8|��~c�<
��ky���z���e̔|���_��\�:��[:�n�F�g�L����z�=���p0A��E!�}D�oZ���j�kzc��c:ߨ�(�Zi5ur����&��&W�l�*�>T94��yΉ�9BvD;H��LN�W(;ZU�������.��9�1X4%�7�a��ծ#�[�f1b"����)�L��yD��K(�6�X�"u=���9��?���N�n���~�-%_R`b��2#�_R���02i���1�CF�`#Ct3���4*����/���t��Sd�}e���]�_�,���W�H�X��w�E�!v�y�<��;��l�5Z=�p�Yn
���m�]=4]n�	"��'��LV��U�M�О%�+�'"-nS��B:[�S4��R��X��X%��wD
�8���གྷ_�е��W�!�9�1������J�$����d��n�+�&e��K��B��>���=�O�מ���C���%��g���JV�J�2K7�*�f�Dt���a">�\�0�K��7���g�%�^�A�sG|�ۛʸ�_��ifBMij�}q{u�뼳'�W�]���<�V-6o������GB	s�r�je��J&^�Od
����3���E�p�%L�Ǆ#��4�_(�8R��5sGϸ�o �OQ�?@HL�`��� b�Аłmw>�����02�0�tZ�������i6�pT�/���5o|[���O��]@���j����fv��\�^�A-����<�D%H'�^F2���>UR�K�K×:Zi�U�ZO�V���т���\i�]<��!C:c/� �j�Дo�J;c�� B}gh=U���2T-��)dO(�:<������H��@,��I�*>����ut��>�>]�q�S(����))��iA� &�|�Ҏ��"̧`��
VM�c��ʉ_��t�k� �U�W�o�>�|�e�z�H="�(oS	DF:�K��/Z�M����`�	��_@I{lK�-�T�P޲��R��;�*�5R����o��_���
�7�.A�ٰ��Z_�qGŭ�=d{��l�G�=�l���&5-���JG�������)Џ7��9j�Aq�D=2�wVN��o�I\UF��)��������l�~O������v5��d��;�4h���,HI����|�WG�)*�v�5)��X����>�.��q�V�����2�3���ͦ(�$(����:��̎�
�<�$����}4�6 ²3+��um��y�q�`VN����a6p��X���d��R.]�l����I*���|��WL��e'/�E��i��GyMP���:��� }ş��9#m~�����&DC�p����8Z/`��Y�Կ�������|�E��b/��\�P[)G�< pefF�81*�}��88"2�b2� ���s��5 ���Vs�l�����I�~>Rz���&]b��E$��ﳞ���贳I���3��B��ѣ��v� ����(��
�����t�H/O+����f��S������_��po����a�!�(	�?��^K:"�c�g��j�d -	��%!`F"���d�g(͐�CM0#�Yb�<�<q00�Efm��ADLK�,0�$��LI�ҀE��%:�>;�l�/�?	1��_@P�&��IRWa׊k,��]9ys�+�S��y.�����ұƋ�Ƽ���J�Y�Q>�m	G�4	������˫�D�p�[�r�o�pg�|ͪoN5�����7�..۠�_�h�q�c�{�E��ڌ�Q���J6���>~�����)�NM��N��W'�|Qe�eg��ʼ��s�=�۬eES�@ߎ@�"���a���9�V������
E�krM�t���K��1��ԥ��/�Ryv[����s1!�N�G!g��Ae������~�$�	I�tx*vw=��IQ+�K b���%{T�|�����z��������뵒�f��Sr���5�d�����>2���5D��|�QbVj0�&K����ȁ��_	���ұ�9xF�i!f��X�H�f|cVoΒk�Xs+!�WXC잻C=-��]�a#h��q�7�T
-�[�I֯�ߢxD_x��S�b'5U�Nd��X�S���9}��[W �����^�*W{��"�v���9K�a��S�l�̢�9r���f{���=�ޭ,����g��h(��,����H�6������9x�78M!k��-�Z���>Yp,��fl�.7��~X�_}b�����W�s,�������Rzm-'|�5<��� 8
~j�*QS�=��W��gѬ���`W+�^�O�2�[���c���+&����,�O��Ď<�@����{��E{	ƿ C��ۯ0��NS�E��x�o�L&t+�Nݐ����	��l�읩�wWk$��!μo��QP�þ��i���﷊R��o��d��)���
+���� �?�l�_�t'�����:�''G�h�U��5�ۓT&�6�E��	�Zem�{���8�5	��&^���U�<�����pT��2��d#��������G��W:7��ȴY���K�n��z)�x��gal|0��T�+zH�X��U�D;�@am@3�8g�6� dt#�� �7HB߲�i���s`w�T��k�M��Wӆ�g�+t�ǟ���1~��:�_��88�So�O������'.HRZ�g^�P�����2|1c�\�c�&��}k#~1o�Ao�Ԭ�<M%�DJ2�^&���cQ.�GQ?7��>��m�r�/�{�f����k ��c�B~o����-c��d�0�:�rq�"8�Dd|L&��Sy��\��mC�I��Uj>|�շ��Q��ވe:6@$����������R�Ѣ-
��Vs���Y�_~p� �e����4G��!�_�gP���t2U���H3�Wmꪻ��)����r�;��ݺ=1�G��U]�s^&��L:To����#VT�ӳ��k�Ԛ��F,y��!G>q*���%�^j��ؚ�dr<����E��.��B|�p��5xs;=QXx� L|�
{"O�K��J��& ĵ�襞�Ȫ�)}E>&��ȣ��a�������+��euF�٠��?f���Q��#j�F�fؙ���iǨ�j�=�g�N�A���.@ ���f��ʀ�D~��1o����;_�ʾ�$����G���L���������R�J�4l��󬻎[��#���:d��_M0�����ܢ}ʊhG�KГX��7��x��АhwE�{���>�茅�(�2�6kaR'���o�zEq;��;Rd@:s�l�^�u�iaz_�2�����X�s��,'����N�En�۽ڐ���e�\Ҧ����?r��P��N��!L`|pb���w�,qo���z��{C��jу����h����\F"oa�F�tＥk�Q��(�5�]%fN����_D~s1�����YۅG#ڴ$	@\&z���̔�������?��RI�����������0�db��2Z�;�f�6Xm�x��w^	M���_W<n<cyA�qbl��@��[�0'Gp��b|�O��Οby�|�{;�u_@=s�jO���� �Ë�5◗!��D�1������=cOw�qI�^ �V�g_3��.c
�)M�O�%��[��Hj/88�{�L��f�vD�hY�ڃ���0
L���\�O���"8AC�TYunԟ�$oͺt�!�
b��&��!���2�B�f��m8�Q��^�F3-��Y�)�6Dw���:}���^$g>�I��+^�N���Sۦ������ ��p�@�<>I�G?ɕ�<��$�����ׯMAeK&]��t��H&5������B`��=����cB��6l���&ǜ��J`���P����p��J{���0�Q�2[I�7�˭ի�~b���0�w��{��I#s�I{� G�I�F�&Ȝ�jM�"���龃���u4�`i[�Y�x�}O��4Z����e�ψ��ն�J��|+�m��[pSA:K�_��ՐKX2�;�>��ZP�1:�a���= Wd�/�]��4x������i��p���~��s*7�6��3k�

4	��u㎨��Dy��\<4�U���v@�<Df��P"�}�k55�ҷ�~�}�\��jD�9gە�Ֆ��t�I㕈�1R�;g;u-�A�7����?f[]$�/��FV�RFW~�ѠL��[�ڲ��B&�=I]�<��U`�kF��t��؏I]<��!Q�~�>+�e�g�`�{�+Ͻ�mI��N�wʔ>���k`Ȥ�ݡ�8�{���d���H
�)�B��y���#�H/F�e}I�]rc$�/�����֝�� (̑[ �ʝ���n����gp�eZxC޲�m_�y���e�M���������<�Sc>{4A�J���"�ž bݘ�?X+�VG�+K@���4���Ŷ����ɚ5ÿ�t�5�i�6� ���em��DE�@+��V}�B>�A-.7��_㌇P/l���e�W
�ex��M��/�e��<s�ao �/ˌ�D/�
+c��Gu����NF!f���d�Q|;�X6�oF��V����[?���mr����߆����Ƨ��͐r�K�^(��sq!�"�ZcLm 2}B�e��h����H9fT�.u]�8f��k�sj������2a����YR��
���|=H�q���%���ӆj�K8�cw��8����K�/A��������WW� y���$-��Òy>�}E)9.�9-�k���=�����$�J��� V^�|Q�\�D�������&�l��~59�lo�����ֵ� ���;�F p>���y����υ���x^�Iw���k�2t<+�<gԕKp���M]:��Rlz����?�i�˯ׯy��U~�M_��G����E�{?�!�=պq�����ڊw�Pͼ���='�AЧ�2��r8=cr��a
ܵ� �&u�VI���Vj�>{ ���曪�kK�b�S�{\Rc���8���D�U��-��1�>d��ҍB�t����
*�y�n4�����njs���T��{Rp̯i��Wg�s���^$6/�u{Q���r�����=o��<���C+�
�M{(F������l�s/sE�/+���De��/����Au��®,�����A�s|A%�������/�����1f	E��Pu��p.�N�B ����I	��L�6�s
kY��?�W���3�����h5/�$u{��c�5Yn];n��8�ߘ��<�G����C|5b$|ّ$��������Kֲ�G�ӕM(Kq�]�x-*z��e4:k�������]�;�n4��ɭ�ik�T��x/^蠅��#����>�o~9Ξ��6[�-�8�7\���.ͪvғS�fX>�p�L4����w{��U���
6�fH���
ln�O���V0�AX�X���'���nU%X���M� �;Y��b�������b�����z�'J��O������&+�/�;���p���b_�Z�@���W�&����pI���%�����6�i$���|l��{�/�֪[�a��a����g�����G}�_���l�G�Ra�9Ts�ˣ�'RR�Q>�|?��Ge�o�2y�� �k>ST�r_SN�\�q�a���y�$j�$������2�R�N����������t���/�M�h{�g�'3��o�v'������ ���,��'�v�]����o2*C#�+��y�0<
���zd˥��}�|����Sk���t�d��	�ޗ���t?�e"y��@4X��M�G� �|�]`{�%�i��^z��|Ţ�ǂ5£��$X��9(%��d�������~�wԛb���3�L7Ig���E WKuM��r׋4	����]e�"Y�x=XH�?�AO:���c�kkPb��壡����V����}�Q�Z>�=���2�2�{�)|���a#N�spm%8Y�C��]NٮJ�rfI���J��P�F��e�U,A|��9$s1���!6��p�d�%Bl�TR�&�����X�sҒF8)�00��:ĄcT[�Vr���k�LWj���,gC�5�M�(mX���y��N~���-u����n��ba��W(G^8<�XfW���Բ7Pu�WGN�����2�#�S�8���,��m<��%�_H"���@-�2�O`=LJ�����~4Xp(��F���Hi�{6o�K�+�<���d׾V�0�;go��k�
���?[F9#��z,���H�[F9��Ir&{iÝ���Ț��/e�6��m��1bQ^~�����\�R�+N�t�9ڠ�+L��G�G��+l�p��e�:%Pޗ�5-wlċŋdo��.+5����>.������7HΜJ`M�#��z>�&���!tK�U¦�ȷT����lP�GE�Jy�	qZ���jC���I#���3�h�V��"Wb��lT ������m���\A���fʔ������]1��!+�ź%|���)����蘈;���e|eb�)=�W4����|>mO�P$��~iB�Pʛ�����J`��-�E�S+�t�'RaoV�����ԑ �	s_R��Y
ءu�V��B�jYg�I�kNPq_!�� �� >:����������L��U��K�9��d佐��U_Lw�$Hqn�y=H�ѭp��͌�<�!�7Z>U�,{ix�}A�����
��qp��m���`s�^�*Z��R3,dj*1�3��F��(y2�F�,�"c��}�{�/��/d�T���S�nG�`q���F�)(^�kz������^��#r"�A ۘ�_%ּՏ�%dE�WB�7E�ѝ�����<�7�G�}�:Drƻ�OAB�Y7T`dI81�0����ʛ�(jߩ<ǇbD��neV���r�`r+�����v���c�(�ء��������0|�R6�o0� -��ꆭy�:�~3�����tkp�U�w	H���l�l����95)]ۈ��%
���ïXp**.3��p�H?�N�!��k�8���sÏ�΋�"�t��z!8��6F��-@]L/����y�=6J�?��쌸fH���Z]��o�BU�ؾJ���H�����7�^�vk�Il<��A�IN��R�����9�MS�	��m:�I#e��}BT#]Vz���E�<:"�I�(@�!��a�C���<����F�5��9�6��.���*Wz+p4�YA§�&#��¡DX�<>�x��ݦ�C�5e�A0_��j�,V���/f�:n�+�P���ڹ�ȃ�Uf�.O�K�h�)<��S0�ǿuV�MmH �����P)K���x5�P�@` wu����/���H�p �^��!�զV�bw���3�h�Be*�ݨI�(_mi��� �J2+�#/��:�f��&j��-��^���P����܆���mus}(Z��:��}3V6IrL4��v��k����3��0ܮ������d)��r�&�-��ܬɁ������2. h�3����_d[�*Z�}���Q�d&��OF!�sxև����#((~��Z�}�!�"wfs�����g����iLU�PŔ0��B�?;|�z���F&�z�x:r[aYC�:�̸�O�؊˪	�kub�_O�0��,�M�b�O����M	��D����6wk�q������b��_
w�Iq�<��p��p����H�5�游v�oCk��'��	�qvOe�9ا�Yp�ջ��� �?��� ������X#aɂW*;+�R	�$ɬFW�^�q;<���xňo�G���aL��������-1A���/_q����cK�0��+h�WA�u�_�z9`�ut6�n�S�(��LOO�}-;93U��A��$��m��-+�m���6�p�B��8� �y�´�3$��Ï-�$�.>�S~}����_���އS�"Y����}"t8$���'�kW2r���)N?yy��YB72Aٰ`�|Ɖx>n,��|q�'n0R�a��ʁ~Ք�G��W�r7n8�"�{h�\BA{G
}���@Z��><4���_��׍|{��Y���KZ���^���.'��QNl��*��Q+���� Ʈ?d2XX=�Z��:h՗:����@(������2����)\#�XB%��#������Â��ꡣ�+��!��� ��^8|N������4��x�v;������q���������s_�!�GA��۵n�b��if���u�(�5�C�4:�y}�҄f-[\o'p��)fu��s��9���#5��-��W��+mEvF����N]�n8+�Ъ�R���z=�~�VO�7B6�i�S�g�%����%��:��Yvմ�.��$����ܕ+��R���(�s魄��oS���QG/ź�i��_���
����MX�E�!:�E��=���h����U�0d��gW���K@g�Ճ�{�\����W�b���9�*�H\ǹO�ڞ��:7Va�ɐR�#TRE�cA����s�p�K�N�����؜Ee �(:T�-0	.��]5h2��(v���h'���ڹ�Kxa6މ�b�<)��i
!a�(����U�G'm`(N���5������t��J��R�x��ړ��Δ����"�����au�u=�(��;hA�~l�N��9�x�NvQ��x��4�>nM�ܽ�橄(��+w�o�&��p�P6�k_�'�oX�"6���Dw�����6�����R{�Ų�\���a|�h*��V�/�	���01�[�m��,.3�/1�X���uS���W��`n�Y6��)�?|g�U�n�����.ƋI���d{��������0�E�7�~�.;'�h�/u��h]�ą4=�-�G:i4�!y_�V���V�O%#�N�r�W:z�q��س��; �D�d��5����O��օ�����q���C��qg���|%����K���-)��_�Ƞ�Įh�)��T}�z�~)z�2M��#��Z����.OE�[�<Ak�E���Ql+L�4���=ڬhoHO��w�OK���q�.8��S����3J��W@A���V`�����x��i�#�mSG�w.��M=�o6ٶ�O֨��?��C|�eZ��S�m,�I�UU��ʷד��l~Ty��{��S 3z'�]/	��*�ӂO���
Qd��?�GA�KRc/��P�������aP�&��\��\��Ɍ��3�z��>x52��z��m�&�^�4x�(��2pټ��gl�QYw;kx3{��{�09�܀�6E1j��4�G��f)wwSD��i�C#�)�qΡ���-i�L��)��Ip?���i�:�IW��9�d�$�}����B�@����`�(�*�?QI(��Z�}H6IQJ�[�>�e��K�;�_�����HH�~��ţ��b��%n�ʍ��Y	�I�cved@JIO,�!v�j��@K�����~5-X�� {�3Y���I��A���7�Q�ŅD�#A=�Ç<��Rd�y·�n=z�h��j���I*c'���>�_��
��#�H�u�L�}KA���TP�p�"�C������!�Ģ��B��[�Äg�Og����Z�O�	�)]#~h3���s9����}���{>���K �~�~����3	�D��x��� t�H�S�$��)HC�)*���Qy|����p��*��
J���W��#^J�9�RK6���*Q\I�dg&�9� �"$���v�F�N�2x<�8zdi#Nc�;�95�-A�~Ͱ��f.��I$[�Db�������\j���vDHY���V���ŭ OC�g�l��~Q� �����ϯ�=k	�0�m{���6t֝/X�yLu�>S�n�w�b~�3�4�?���k�1�d�,7䝓aV41��E�	W�v�p�W_��ď��@1��R��z�xܕ0O��4+�_�OP
��s8*Mj��V������w��eĵo]�:�����}	tQA��e� �O�V�����֮�m|�X��KD�oe�1�D��KP��`��y�#�� "��Ȩ9@YKE�GY!������(,��!߽B�H��(if�Z�^�ԟ3��CC	3�,�V��s�Y�y�)�$��^��ץ�d�l2�����͍�30��e����Y5�@Z�X&7]�~],]�
p��8�g���l���fl��c�Q��N|�z�fs�>���2j��_gǆ-���Nw���o9���K����m�;�a��*��6uRi��dp�7�4A�j�o�|ں(.�9C>�<s�m�b�Thc������maU��冇N����X��>.
�W��/��Kxϼ��W=Ix1����_*饆cWnh��|�^*�JC��%sP���R��g�ǅ�+"W������#b_O����9�q�l0�[5Ɉݷ��������GlҠ�/\��kE ଋh@�&�7w�:���e��ZCn魜�u�c��5!x΅Z��L�vhe{��<P!����g4��gU",C�� ת.!I�8�h����uט�
\6.q�z �b����6���.֘,�n"0Dj�+vg�,���j��K��|5l!E��953����ݱq����gs��1�̴��� �n�P�N0��J����iǩ�����W�x��v�;�Pf�8f�.����W��r��=�K�tO'+G�K�VUo�
��/+s�oaM�15���h�����]�Q����f�Ъ?�#��"K-a�Ҽ#:��|��*�)�8��J�E� ��������v�2W��S�@���j�ُz�1w�yY��N5~�Վ$�{����ߣ�,�����ŨC�_���ύy*��/M3p�.�w4U�w��:��E���Ɍ���^O6�M�C	�a�}�M&�d=BJ&`��D��������V�����̳1o��z��v�dM����_b�����I�(�#Jk�t4
��9.GZb����v�m	�d�h
"��I�m�Q4�.F�y^�F#��d	I��s(��U2�@�&�E�Z���-�T��<5}�,���8g)�L/'�]�R���d��Mƺ�9S�~���)(	�,%�,��Ƶ��B^�YR�ċ�<Ö�?��;#&�X�O/}n�wb���S�Jc�՜�����utkk�&zv�p�yLcҦ��č����1�/NK�E�=���ux	fx�25�䗖�(~�ZZr���2�*��R��	����Ō[q�t67�g&�QO��Ю�X��Z�BYI�[IF+��+��l��0���{Y_ˍ�n/�7`�ɰ�=`�&L���X#�u��WL��Á��R�Pt��~g����ݱ����p�,��f<�F]q���0 oe��m?AB�ֿW���l:}B&Q�G��_T�f�l[0AP��"�w����9��T�P�.x$��c)N޶��lV�����dqM'h�^��Q���f�O��@&c�\}MC �}�_�^fi݆�tl+9,��4ܹ2�cq�O�|�Ǉʮn]f�������2���DlXz�k��'i�'�P�R�/3��t�brf}�kf�����T.�}�a�m.$�Wr�:q�O���9��� �55Ӻ����k��M���|�yN}d�\X�Z��e���s��[���n� "���H��VUO�T�����m��PrUy,��֖�cX�{�g+��o��/U��P������|3�Ђ��S�i�H��=uo�Uu������7> &��c}s��ֈ#�N1�y�9��9c�0�{�8�a��4��dH���I��T����!���{����l������'�1�)H
@PI�h�M� ��1��>]�+�IH&[�dJ�7�R�:΢o�,WBTA�CN���S���1�kۢ\�F7����bV�!���'(R\�'j�HQ�p�(q���	n�yB�p�c/�ڮ�'l<��򡇮�����/υv��ܰ��-Ίh	�Gѥ	 gnV����H~��I��)*6Vѽ�
d'�~��9�}ʆT�gh��I$hv����`(ǒ-��	�#�#$Ɯ�<]�yR0�38�Ž�p!
><D	"�����[�<G�)Џ"9e�� -�)P��U�b���|U�T���7��˨��7�5�L3��6$�d��u����iv�A�[��Q^�UoW�&j��;N����İ�$�Е�HAܦ i��H�3���LݟEK
��o�������>��p���ל�/��m���#�i�-Gڛ6K���n�l-UK�Y��L�D9�Ο��+l۹h1�劁@yC/L�����F*�LQ�(ƋD�	�ni�Z����&w�3>82����,^%wM������UrXS�c��Q=�r����&"=Aj�aZ�d�oFf\w��X`ia��U�X�y���"����?=��/�G�&�E�9���_xW)j�љ��Ȼ+����3,kL���Bo��	��f4<�6�`�u������`�U���~��n���
��(�#z�������N=5w�w �5�H�ƀ(��!;d���B��)����m6�sǫl\�Ɵ�����$z�(�5�E2pp �׎�z����]/��6 �͸��b�Q���(t)k!�p���`���)����c�D6��A*�IG�J%)7%�@�[^��������O�6d��(S���JXW�Ĺ�rq�ʏ�2+�HX��8{�2v�;	��oH5�[0R��ʹ2?v	d�D�Ɇk�PնՊ��in	�n}��Q��X��c��c� /�P)�i;�Zο�n�I�����R��Ld3��D�WV>˸A&B��+�GH�%K�\,��sݤ2J����G�ѓ�ux�>��r�Pl_��X���8V�4|��>��k�+�Zv2/zG@ƝGh� �������S#���0�̀�!���t}82�S�.���\'�b�뷑;�w�d�A�?<�Q3�x�3�u��w���[/��rg�3���/�M�u�6s�	��7��/4g?�6��ǽ�oǚ��E'B1�̼>5��g:IU�LG%O0����W�O����*Ѡ����,�C�?^�̒��M�rE���zZK�У����}@�D;Tg0�U3κ�Y���i9h�	��|**`�}�(s�E�b��}��Lq��p�A=�|�nÙ�o@��X�G[�1lT`1��o���,N��v��r��ӵ�h��u+�;�]yLRI��O��8���]�����B�N���.ľ���Ͼx[F#a��^ǘK} O~�d�&����	�^?�G�Hv�j����.�U�$� (6�(�LRT��[� �r�!�YF�0�TKK�N4�'�ۘL0�_M�r�^��
����fY��ZC Y�3s#d�E���e��O'?fnџ�N"�_,"�pL��Ω�C�Y"у:rA��ѡ��e�����֝7�%8�U*����V�P�Lb������z 5��O'�|�~6�礟)�r)�̙$�}��X04}F��>�,.�o��	ۂ��|�\6�ꨡS'2V����S�ڟ)�3�ڊ�,
A7n�&�0S��4���hyk܀���g���4�p\��c��L#+��j��I�D߾�!5�<���E��$/@#D��+uF�r&�پ�;K�5M���^{���L7�g�$��mPk%�Qѫ�Y����ʮ\ڡ�zƛ4��`�y�/<%�|_/��6�s������G(�~��jK)��yf� ����9i!�K��J���z��.J�W���,o��]+�pv�+��B�!dD��PE��-�I��ThL�@%�8�5eP���kf|H�5x�0D�Gu�(��
�.eON���':*���,��b��O�~�_%>�%"�	b��T��1q��K�L���'8%�
�)��E½����ёO��eJA��j�0�v�^��:^�N냀�3!�5,9E4D �����*|K��NK���.hX�.�F�"��O���]���	ʓ��������)h�VE�'�Ak��;2� j��s�Z�j�թ���K�A�]�&%}ru�␝5̊�S	=��q4���V4��ڧ�'�;i)��=�8	J��N52�e�*�e�RR]�ٝ��4����̤1" �vC��~��/�Au�$O�����0݅Q��b����\tHS��c��e�g}bC�3����{�n`��d$<y���*��b
�x�weK
$9���Ƈ�tnx�B]QT*yQ�ڴVPA�Y�Sf6	_�l����9j]#�5� ��"�ß��7�
� v�=���98 �>%c�vܐ�Q9/�t7�n�m�fc�J����iEQ{�]�Z9�^U3$����͓�S�y�nP<�|��t��*��T���;���缩�.���H�=��zd�/VAo�$��������P�$�w<��G��<Q���e-^'Z?vK����'[y�M�s������n|����\G]�9lF%��'q�]�U7q#s���)	D���7*��<���m�&W��
R�q���e�b�:��1����򝉀֧ݎ�Q�x\1�L3�D�j�!�)��:�R�:�]���Y�߫r�d��G2��J\q�1>#�9��y6Qf�kY��>n�E�&)$�dB��f͹/�����B��q<F���5ќh�ɝC}��b����
�^'\�\H��vh�ރ���\�vpw�=V��*��Ra
d-�C�����&��՜L�=�$-��0k鰞������iAx��a�W{��E܄�{�R�ٲ9�b��~8{�[DCK���(f��f�mQ�?���W��zg\����!@t��z�@����j����^�������`K[��(v�,E�L��i����N��=��cv�D;���'�h׃_��`y���(�e�esi�@����X�`�γ�m�S���^�Ӄ�C�~h�^�0/2XP0ra�I�B�$���g���GFId�9���{��X���#\6ݦG�&��Up�"��0��6��G�i����VL��(�3�h��k.)���XL��z���`
�!!ݶgp�2�;�H(�I��>J�]�z����"��N��g�-s�R"w;�:K\��[k*��	����nf�.@��@ 2�,�'���L�m�j@�W~0d�T6:�����g�T������L�!G/��9����}�eH��h^�-�����a=)�$��ǌ�j��
l���>�j�����Ir�5X!�����Hf��������c�fj��P�i6��V�v��H$)��'����( IZa�����h>�����I³�tĭs<�.�w�9��i:~0����P-.�HD���P���M�3[X#���}{�1L��=;��`÷/>���54�T�(�Zp$��`�O�dq�'������I&�U�eBs�˟��/�1r���-��P���ڇF_D`^�r���P${�EAO��f@Q!V7���o@�4�͜�v"��Ԓ*2���#T��ψ��?´�`X��m�v^�\{�#��v)�a�lEE�(e�R�j�;����,a���y'�O�ˣ�z�'G"C�۹ * �8�B������������9A>ң|*'�`ya�6�]�{��D�e�­^J��Vg�Rs�噓��#��k i�Q.���c��:v�d��� LdT���*�'��Y|�8B*�B7�YFMM�R�	H�Z�"�:���ל���3O-t��A�c�)�+�}0�2��*FA#�t�@���lZ���C������xj���;��qX��f����.�P[�܍ �e�f��e߇��>nA��E�-�vgI�7��݋{_U�	btR�R��?�[M�`C���y��1������׆5gCCׯѨW����Bt����׸�G�ת�Q��x�&kb�C�wt�0&͸�b2c�$햰�6�����y�f�3kS���̀��&TjDvU�������B��5���>; �۵L��n�f���?��j���{})�j@1�eѬm���?�Q\69e�R�\&r}7i�ݹ��N����ZKő�x��D�,r��[O�BG��q��{�V�r
���8@_I{�����Hu�l��DG����om���^S-M��N��ِ\&��������A3�$  ����욢�Õ~��,�$��
�����"%ݏ�s�mq�y���We
�fв�S7�ֽ�F��6l��+f��U��H�����=ӈ ��sY}�6��KŝP�Y�������X������0�f�H�+�x{�σ#^[X@E2+�4���$2����a��R�փ���.3p��8�3w�?��:7�t����L9a����	x��T�u��|:m���%�7�ܚ��l>.�mN|n�k)eGu�O���BS���[8m�֣�Ѯ��F���J8���Y�ӂ Ȯ=o`�{�����*�AI�wLJA/ޕ(�)��"����$�`�ܡq����D��m==����T��{4a-5�p^��:3�'iI��3m��/�h�4�)m�h�Kd��z�gf�\m͍�I7{%�N�>Z���E:s��r׃����m�il�И�O�乺ϗ'��4��dEIqձeq�&\=��� Z��M��~n�/I_K܌"�'��ٙk�}M�c5�`�a��o6�:�f�h��)�jn��V�{a�8�7f3Ժ�z[�:7�¸�W/r(�[P�h�[�XC�^�a�=Fx��)"es��Ϲ�^�MYT��|��$;���Ĕ݀Ţ���'='q�GGؠ=QP�+3)�R���gb7[�)���֤E�U����̣lB�]�Y��o�d:�d���\��6r�<A�ܖ-^I9��!�s�\aK����,�'J��"�hq��W�?�R"�
��K�Y�)�'�gϼ*^��Y���^1�APF�q�W[��,�S�WLnj/YC�t��o�OA�ѓ^V�DT��!r3�ė�����pa����X��b��߭�E^�>�L�������,B�x#c|>H@,���
��0A�
�f�@@��%����xSV#.  � �;#)� ��7Ӎ���M�|�	W7
�#�O6�(צ���"B���V���jXN��5tJ��;@|���f�X�45�$�D(K��n��T�j�1Hͬce���I�.�&#g�㬛�[�U����`ZM�.!az"��d �R���\�?���JD��1h6�k�g.���b��*��Q&Q�Iv��
�s�ZW�8��q0Ȯ�`Шi�̅�w'�,�$pH@W- C��&�Rl�Q��=:�uW�
V�T>�(}�-��7��?�iKg�Q4Kni�Fݭ� �އVx�Q"1B�H41�Q6^S�4��g4RQZ���M_Ew�l��<iHF	����[���ύ}E!뵪ι5�4q/�׷!W��n:��	�3Z����A#����N������K��-���8rr(Z^�~\\�~e4¸��|�K��_%I��smŻ�yD5�]8Y��ڎK��b	��:��,�oB�%��]�I;�0��W��CT�`���� �'P�B���-�wV(9&I�:הѝ�LwҤ�����K���NqC�xjڤ�-Ɗn޽V��b5`Y�/���N��7��I>�1*�� �[�����IN�������
J�ij�m��d�gw�79-UOs��V���ku.�X|�/{�)Jdh�ɜ����PE\�gWVˍNM|L��x�j��x�h^٫���s�R=^Uj�v���|��$U����^	-ű,���?��b�|5�G�v�J�6zk����*��G���.M\�A��}��3��5(әxcU��\��8`P�ڲ�s ���z�2�c���.L(q��L�1��ѥ�H���Hl�Z���L��,����&���Q�m����R�z����o"�
?�C ���u��KN��4��[���I�?Gi�m�2�+��xVw�No����ӝZH��@��/��r/$����R���� e��8�k?Y�0�9��YL���ͣ���Td����
�T����j�[CG����+jd[��Lxq���v���$��4Zr�>���'Л���Ǌ3�n{��Um���q�@�1��@8ْ�4���jR;A�+�E��<��5]k�εQ��B!eC���Ὶ��o�)�[�^��q1�9�KTw�e�Rl A�g��J���V�O�\�ç�b�Z���+�|K=0/]�gW!r	Pe���0(�Xt�ڃ��Hm���Y�� k���J��S��.7]�-�U�Ż���	�1�!�f�n�p�,5,(Y��<��)�Ŵ�ċ5X�b��lur�-�MYq'��v��@91�#�>s恞�U�Gm����^ixΈ�fM~B�q��W`�~��w�._YE�Y��ٟձ��Kϡ���|R���'�r+!�R��nʛ��Ʉ0��2v�eƠ�����8��ӹe4o�?��PN�B��ϯn�ˍ�`���`֐�5 ��p�� ����3�"��}����u
�M.3�����b;B��0�8%���		P��2�e̱ˊ����k��%������X�����fOڰr��l�^n��;���֕֘-��#W�p�CCU`Όs����Pt��B��Z�^��oR��*[��?�p�!<LgG��6�h��.��*�|ۧ���c�l%���1�'?ey��E�n�30��^3��� ~��������\r�t�&:�����"� \�5��ڏϢ3R����I��iG�������_�wv*�Ɖ���u%�ơoKʉ�Y>v�A��"6���tx ���Xtq��@Ƒ�����27�k.�W/�ԂtZ���>F�!	���F�ݗw���c������=x�
�~#�l���z @-���K��H���<CA���x��0ޫ��S��G� 8�^��u#+EHn}b�r�6�ƕ�����`��k�#kii0��x�iN+� �h�(�%7�����(��	�d���`H����q����r��u:'r#�Av���,�MՆ�>'�g�kX~߰�\x�~	�t�)�H�k��R`�ƭf/Y9�+T�V�E]H��<5*��l��d�hq$v⸑Qܳ��������'�n�_��K�栟xɇh�9��I�=����[K�.:l�����j���/��	p3O�M*
^����9A����4'J?��J�ے���(N���WSws�� �V�n�R���l?�i��(LI\��׮�6�6�Jڳ�����vX^�Nv^T��ͿB�me�*��细#w�+}��E�
���Su}KG[V� �����N渱��W��'uyn�qd��n��� �!$5;3`A��Nf�,F�y���n`1�Pl���?���%r�9��2�m�鼿���@��k���!��KoK[��~��S��o��	���Q&.K*3�D:�����Z��z��gĺ�(����םe����)��
��s���������W<�>�,)�/��g;�w���12]T�ʟNlNK�;^lY�Q���F�m�
�/񯢊fS~����th�o���k-��1J��X��!�Mi��xڿ�yr�Q��q�����b�D��>�G�p�*�@��&D�s���*|Ў��J� �Bd:�qBB�`�720&l:n�Q�O=e���Ǘ�Mc�����Ļ�����7��;wՁ��K0X ���k����4�h�Sx�V�h�,���!,q��!�f�������8D츎+W�T��pd�v}�fBh�%4���n�4�o�2�g �(�KU�/�v����7��m�y�I�7n��m"SƏX���Um���(_�B6'�x`�l��w��X���NG�c�w���G��p��/���v�`k������9��<A���B���N	;�5���!K�S2� �|�He��7�A�i�]� �m�<ҷ]���1�F�TZ;�ɰ)�Ǐ dO8�MiyD��F2-w�������8@��9�[�\Q*/wrC@�W4�3}Fa�=.����ߪ�_��-c��A�F�ŀ��Z���gJ,ߵ�4,��͞� �\����®� �����O��YVo���k&��nS	���f0��h���z�}� R��J'�^�{m��[�q�*���O-�S�e i�:�ճ4kǛ�1=hNg�V�������7���I�	u��G"R���S8�N��
���=~�B�}Y��	皟�ͯ���8���G��/�sܙL^�q7#@��^��b�Y���h��DBuyg��J�(�����6��J��*�����5I�8����N�9��땽#�VK���.�]���AO��2r����E�Qe��ezɓ���풑��7Yy݅��O�����Z.��RN�!����3�&b��W�~�p���{jn�6�UIRD��VZ�#���ƙ�sһ���zC07r�8�p�?Ę������{��i�-���O��+%����t�*8)����~.���BU-_��y_����O���_��N.j�FЇ�)o���h��u��׫qZ̀�^��6=I]3v������C'��� ���UFl��U�uR0-�cH���'��,�I�?f)�x��T`�&�c���x?�o�O�1X���x#O7G�m��P��c�*�c�TS�@�����ʵ�	?���b��N����5S�o�A����V&Fz
�X扟%���>1��\J�~5L��ӿwչ�0��wl�K�� �(O��e4RDI��N_$ŉL�n��E�Ou�f�Y�ۏ���wU���o0 ��������v~L�o�y��$�){{�;��W�cP�sa�J�m����B��q�|�ِL6�dy���{r�${4X�7=O�1: -�o��2�vu�d#�V ]Ěy�7t�⨿��-��<d
��$��E;1R��o�+�L+������~���)iKuˋ�D9dy^۳:6BV��_
�Q�0�W~�z_x%!���	��5uhΨ1�O������U�F�HZ*��< �_��Ϟ�8?%�-^�d;*LfiF�>ыy���E"{��%���o�Rb#=�Ϛ[M���>#��mK���.��c��!;{;xH#u�1��Sp��Z�x��1�$�r����HF�k^�F���va
�D�7�p��j��>ϐD*N!G�P�A7B��/��\X�n��d�hc�p��ו &Yc�_ ��,�C[}*�SL�8�+������N;�wޛ�b����T�J�!\��@�@�K������{I;u�/Mӷר�I^`���SL`@b�u��D���gp��с�T�>��HO]�q2i��'��a �C^�l%�&T�q}��pklP��{�/T�IN���)Q��ؼ�r�S��ѱ�?�l��6B�T�q����|b�$��h\d���yQi�X��W.;l�-��pze����^f*��h��5MtHL����N8�C�t�2@�x��cGț��J$RTgS�wz�Lu�zd��S��R��J0I�#w��K�����꩖2@�@ 5h(⨽6y��ɂM�������1�ɼ�8z�?AL����{�{�>��L�6w��nV%r(�.lg̀��<�Zͷ6
δ	h�ZN�ޭ?ݍ�LDEY� i�}I�?ʔD�{���Uw��='~0̶����Dբ��/<j��4..��;�Z�īN9{�-�c��ǯDc��7w@�#cq~����uE�Y��L�ݟ��"�7�E�8~
�z�v	�#�/U~%�> Dً��w����2Y��q�Ha�!��(�A�f�]O�1y�x7�g�o�N�ȏ`��#
�F�
uJxW\Y�	�6�C|
�V�m^�{1a%��{3LϘ�z��x!��:18���
��Db�A�]��N��Cϼ��q���z�z����xkHt�F e��}�4Få��T�>+�F�T��j_r�+�R�6'MZ�:5�o�o�|�^��JJI͜����#�^�%�� ��cq�2E��O����n��8��Du��Z���R��&^�/��t��/8�������	0���0�`�m�"�?ݸ�8��$è%���:�R���i���a���Kö���*�H����F Aj�,.�r2gS�`��h�;g�,�Ք�o���|eL_��8�58d��`��%�P�w��w��ߴ���*��6T��]�l\�~�k6�xq����;p��:p�yr�S2�ߗ'׈�&Y�&�6�d�f�{c�+�Q��k�)Hv�$;HC^�ݎŊG_�1ύ��3[�̔F6���83ہGs�-�S��P~�Hj��G���#�9����-v�]�̖�I0�΢9~�nb���Gd%��i�8^�*O~�5L]R��&>b�IrP�G�m������7���Ȏ���BI���4�Ë�k����47x� �hwA��sj3+�{�ͮc�����u�v�y�����k
�mi��E��3e9�`�f�P7���Gʱ&��"ji��"��f�� ���5����VcSx_|�������s'�5`^�\����p��ӂ'U�|sz�x�+�ҵ:HD ?H:DRX�AF0Q8�M�zrej�,�#�WMN������9*�v��vC�q����F:��]�w��o>g-,��i|�ۑ�x���'�$�{��."���zh���}7<�z胾d�]Ԋ�߂�D��|(����+p�>k�S4�_K掣�>e�X�8~��N)I�e�R�f�^<Ԫ�І�}m=	ɴ@!���A_�@�Y>�o��^����Љz�5A��2,��du^G��M���v	�"��D�)��ڕP��: P��<m��7j�����)'}B�ZϪ�U�Q���`�)��K�]O�LS����z�� 3�l�Uѐ�:�ĢCR-U��B�@4$A�m3�\iVƓ�����H�Y��
�����E�=s`�O�r���޷�3#�PGȶ@Z�UV��?��ᬶ�Y:0Ax^�g�^��.��g5�����;����m�[T�+kv��9[�(��@_a攐e�4�4�WIH辒�{��r��bU_1U���$)� ����ܴ/zJpP������w�Q�V^�&���q��J1�/���A(̷�������I�d�ja�5���w����98ۘ��]ի����Yr5�]�O�@YK	T�SG-�B��+���r��ͯH[=�� ����qE��N�f�rA��5s��!Jܭ�/F��1�[�6R��A�Z��:������M�b�/q�f���g�9�s-�M����X���u�խʗ@wE�+g�l���%&��OMNLC�ܥ����0�N�A$`b��^�a���fHZM4�Q���w��W��pkGi娖���7S�oCE�.�l��K�����"�J���Ub���Їe��)L2�����\��Bf8��o�|4�C�y
���A^"�	D+�hK��s���^f������H&~3���_��G9NI���L�c,�w������G��t} �9-�T��~yV]d�"���sā�g%�A�'nST�>�_��l"����5��1���7�4��ôH�/�ۭ�S�:=�	�6�-�iu��Lʵb_�y�����WʃHl��aP�w�f���^�[5_L��=	�e騲0��"R�Wv������׎�ۂ��jk�6)�X(��OX���GN��7u�JW��/�INW+	[��l������c2W�������e�=މ.�$5��sQ$jJ3���%�-�X
x
/0��]BP��𼮳Ђ �Ӟ���f��ET�N����F�-�?�K��;����S��R7�y8���(����s����t�R*�m���R�,�� ̳
�	�v_.Ig7prr�7��<���J�U��j�X��'߃�2��IG��6�V��'5cu��$�sܢ�~V%�����zZv�2���7�ǹ��О�m�b{�}+��JX�Z�P�t��X��'�T�4f���H�0܎3b������c���mH0W��J�(�R?�]�d���rI�2i�`���aerC�6����Wv�E�=y�
\����������[��P�l�=!<���|Ȏ��U���9����<��e��
D������m�����N)�N���`��
e?r9�.�"s��I���6�z�8E6n���~Y$�����~�m36�T�٫����P�k�v�LD���M'�W*���>�Zo�����6�y�����	�Ќ]���h_�P���o�4��X���ŋW6I&�AAt��ڼh��Ђ�S�|����{G��y��1�\׉��M�÷��І����O�!�w-C��Ďf�?�T��*�`J!� %�9x�:k���b�	�����o6�as/.�/nP�W� .���M&D,�@��VL�x/M�֟�;:��<�=@rk^����Lf�[�Z��s�/�E�s����W���?i�O�6Z%��A�-���ߺ���j��O����9:s�閙���ڲ55�Q�3�R��� �r.6C�?�ya.Xy�ΐ�;^��������qe=}�*T_i6����Fd�Uy�NaX2�N�޷Չ��)M���9!���|�,��ha4�{Y�"�",߰?�|�� �^m��N��1��Ri��h�]�iLN�����olO-}N�9�$��F�v�w��ҍ�],�t���Zh�ý9G������FW��(LbpK���{M�:ĕcW��^1�@3U�VFC�����#`V������H��G_��?��.�,�b�nF�{��KJ��6x�N�iy3��RXL~"�|]ł��<��$�|
>�JʿU���][~ۣY?|��B��gVy_J[o>%�],���골+}�\}E����� {;{6~N%\��I��b���4E�]� �>ֿ��فt4��FC���LѺp>8�j\2X�)��zD�G-l� ���f0�f�j���J��Js��բ��	��/["^�m��}�m&��UлrES):�70u� � �w6KX�g*�>��$ɹ��_�Z6\}�;��	�|��V-�vͽY^����4Í�����\Pu�%����3x���heRx�zI�J.���M�@��$��UțE9#K�}�eF��W>1����
�Gx�)��d�L��jfYV�(2�H
�lhx�; ��Ņrbˋ����l���-^̷
Ҫ�zb(֥o�� U�{�B��5�f �|�˷��ٔ�G�!Rۙ�����Y��+���]I:�U�2K0������!��G,�^����"��! n>H���1[����ņF���f�8/�w��s%ݎ{R�<�R�i�Ci�,�&E%A�=����]�T3b�be�SG��f��Ֆ������PtL ~V�Ļ��h$��3�a4 ���1PV��ny`��{-��=V8����^f|���+�(�'����1]sW�n^i�[q^�=����M�6r���q�߉9J��(Bn�� J�+����v�j���Z��T Ə�@���������V��q�`�f�ct�D����a�x�6���x5��'���l6Q�s%P�"K��߬l�<��V��������fM�[Oe1w1UA��妭�0�Cq�A�M`�>��ħ�ЋQ�'{@+�[m9�>��D^�C�R�����Hy�u��=l�R.`��< oa����Ds��NS�lx�i�ݴ��$�ӥ��'�]�����G��7V�;�ܯ41Tu7Mc	�ہ��P��0�=UB��Lxk��>���'�c�v��O��T)�R����	b��b����};�2$���"N�4\�TuT����D;�̸�w��Y��yK
�$��s�̏�˻���dyT)�lq.W�x[��\�(�'q� ��z[M��aD+�l��������v� Y38��������/�Ý�E�������#%�`��l�U�z񇀵��%n�_DޖՏ'_<_���y��پX��J�g{R�Hh�S辘�.V��a��Zh6����:gG���__�ޡ��S=�憬ƊZ����|��4�8��)�8�Uk�ћ2	�`��$�Aܟ�K�-�����2,*_FEcY�`��w8^I��ɀ\v��ϦM"��d�v9K��F��!��8�9�����؀p�\���\��i����M���<|M}"�,��a�W������������Ҽ��A� �v�u�^�$.�9ݙ�E���8#H.`�{0:���Q�����&�?�~���OS����Bl3O{���� ��9O�7�N�8�u��5@�?)N���p����Y�XV�i%��R^TK�wpپ�=,lKb�Ǫ�@-|�A~kLq�
k`;3������m-|�5JEcw�@5�F����+�[3���&�aa���
�0�
F��u{+R���%f�t�M���_E��%�0z���"���Fts�ތ92�7�5-��j>��A�x֧��������~>�E8��9���n�%�@*�����][ɞ�X*���5�kbL���7����W���v�2"ߪ�gd}�8/��ٕ�fe�~��9�+m�)
�c���1z!0px�����]��	��v��!��.��O2)m�1��X�א�h�_��_�&�l|mf���� 
��4������y-�$����RCm�j�pX|wAM�j�[}ҩ�<Z�fz꼾վɝ�`�����-���g {��h�#���{��c����v�l*C]J��1�K<���=͕���i�~�I �JS���.�&'� ��n�)�������6OvC�x�Z����C�L�g�>��'��B�z�5�Q���R��=2�����2�ו�
�b���S�WX�S�';�E;��0�)��p���g��o:>� ;����b>�<�(�<�4INQf�M0�)���r��T�ka���G��	�>��b"��'8q��iPņ���Y9�L(V_ܓq��[N�%H��~t�a�^4Y=#6wnd&��B0"e�<�8�[�
Ԣ_�nj��눘i̫2�u��k��D�%3T��@{
�Bp���[�F�щL�du�/�F�+���Ѫ�?q�0�1nc#J��p��xWz(�u.�!��n`�{�{���;.L��L�;LYhG}�H��� 9�t�&5fp�ׇ�?[
- ���(��/֏��^Q�8����r�9.���\���o��/�h�֔`d��<a��Ñ����i��q!,3�o�3p"X�Փ *Y@�:;*�/3�.?��~Bx��q.�V��j��|�d�ٴŔ�0�1V �ƭ�9��Nkv��F��rM���ɪ�5d�J�A�g{�z	J�(��+�O����J���|��(F\(���B��`�(@X5�9�n��K���X���秬��Ń�m
���v��i�~�|Ȳ�m�)�2��C�IE��
Q�r�跺��d��iBrp�
8��0��7��O���>g����
:��-˾q��|�re��_m�{mnW�ߦ�h��1[�J[�C�x�`G/�6���O?�'h�p���v&�2�?�b�o�{��6�����~S��z�݀؜��2�`$m�G��
)A��+�� ���C��eP��5��1`����`~ �Q�ݩ�J�
�[Q9�-�H�<ӑWn��@S�Z�l�+T��*v$d��Fs&�_W�<84b����W�q��&_�iėy��B�]9g�	�9��i�s�6L�n	o�D|{>U��q�K�>���� ���u��˽5��`�����;\o����hӗ�Fv:����wIŋ�b<��	���u�W\����?sx�����qU��~.Q��NΡ�d����mov�o��Ms�L_S~�Q� ���=�%K�Qj�]K¢�/,�U}����x��43����o%�qXބק��]���@QNJ�ûN����&Ibc4i px1e����v��εp�H���@������+p1eYٿ���D��ʕ�^���?i�qu:��;5HRt��h�@����L��b&��DoRr?����l���E� '�L���W\="Ԯ>\Q���&��Uξ��LϷ5�IٸT��w����ɝ6~�b��fE�	\g���\��BDH�E.K��Z��w�H�9F
�<C؀����M���L�:7(q]�-����WV0���]��"�?G�F~i���c������&�6��&^�ʓQ�\��\����b�����������	@V�v����z�ʅ�Q�u���w{����k	�'����YB�Ё#$L����b�7��f讅IAxAӚסּ�ҧ�;�Y�"�8�DP��tF��5P��'h,���0ǒzDISt�&?�����3�{]<,|W�庋�r�X�+4q[�moTfqS�j������A�e���3�D��ڑ���f��`%?X�ŵ"SplO�.{I���}��<�G�Y>������� ����L�`���7�.�JF4�YF�G�ݗS,�T��Vk{���]�?T����웶���H|NF>i0�9Lז�7�@��?EӔτϒT΋F��q��(��[7���	:����k\��|��&|���(TK~A��m�Y:���1{L�,�r�.f��q�{`[y����	���xhS�ذ����g���:�%��u���mGVD�E�R	�턦A6��{$�i�O�B���|�T jӪg�΀Av���:9_��� ]���
yEvj4��x$�A6\7����n���v㎇���K�䟪,�BG@�®��c��U���eѝ۶vO�^�wh�+=נ�bb.����8X� �ظ%��D�j.��V\PeA8�3��	`�$�|.�N�E	V�ɸ�C�Bټq��Sղ�XG6:mG���f֝=��s���X!�k0c�vzD)N��9�sӊ��A��e"mN?,:���o�1pe��]��;�{۵y�D � v�t�g��S�4�)������zk9����Iҳ[�_��s�4�٥H3�/�A��a�$� �	�:��p�m���6�Y^�����T���_��z'��Ɨ�����'*D���a���&�m?��i�G�R:�/)%v���FǼ�n`����E����ݗyhKKm�󺌯���r¼J��c�o����0����1�(�[�\=�����Syf/�EZ`���#x+5�Tt����������f�D᪢c##�ӵ٦,�,c)���5i��upI�6H�zvSfB#[px-��'-�!0� �'w�$������<̍$���� ����x}eW �e~��44G;?*DgT�a'o�3�`.����}�"�K��m���>� �7 ���VK���b���(���UM�]k�2�=�v�e�T��b�v�o��¢i��%�9m���-�K�O�;r�r�?3x^<)�`͠jr\�%`�P:��"$5����jL�,�&_�Rv ���6�i5�Y �[���tm	J��ۑ܌���nϋ���:�6��yW����.��){�.��C_<�������6���:BO5�ĒY=R<���Ò�e'������,�%�&��2�����֕�^B:�f\�h'%@����M-�3`j�}6t@�r����*iݻ�Gg�!�p<L��c{(�r���32���!��垔HX�l��\�?�U�HTM�\፭�*�ˇ�ҍ�B�we2��ye%P��<��W�?���,��I�O�n�@xS��U�-&�tf=VRj�r0"<��q7�٧5`-^�i��$�)_s=��KG+�(��I�9�9K���t�^�+�g�;�۞n�o$m��6	��Hl��'�n�Uz��R�l+�ç���)�|W�g��ʽ�Ϥ�슴��hPfSJ�Q����P�W3Z]k�י̍v�[��3�iJ��o�48-�[_�E]�2�8n1�NZOQ���������QxxlյG�������|�����-9��)�q���~L�!T�F�&����WW���M�"j���_q�U�~�Y5�'3y��1�%�I9pMu�23����7�qs��7����Q����:a
֙�7۴��I������,����p�0�g����΄���q�	*Ǵ��Q�����< .m����S�E)�q��I��K-�;���>M���-��PX�"��X;2�Gn_hS�ѩy2����O�_հ�g�\�EqA�S�/ж԰[�+6�̻C\���ʯYn�n��u��~���w�r�}�HNX4��z��ْ*�k��g��^4r�\:��;~�8����_;%��ib�d�=�kS�J�\8�\�V@A��z�ooQaP��-���a���Y�=�I��C9�
	0�;d�"̲�ߓ�[.S���_��<���9Q,��]�]>�	�☀R��7g�Ҙ���U'Pl��Aj:�K굢��߽e��b�Rå͌4\h�x;1��)R��9<��ޟ�V�! >D�Y�f����ӱ�of���K�@�	��t)ڙєb)g��ꬅ��ހ�M��6�����܁�
�N���J��(o�x�C9��ecb��y����s���arOû�x�qUڄ15AO��u�X��q�j���'t�>���F��4�7�g�)�Xc�ŏ-	���M�?��P�;��c���~�ǷE�!ۣv63���^WRI��At���++��`IhU����R��a��k$͚޲8!M��C��˂���.'4��m/7��Jb*��V�R�t �9l L���P����+]��0�f�Y��@�*������o��р`bCtW�*���᝘N�4-;��\�.NxQR��{wGϹ군���&@[ţ��~DИ6�o��@��c�>%�b2���p��)���C�%X�e
�-+t��ڤ���Cyt֫ItmJu_���9����b�K��x8��Z��X�|�����d$1�GЫoԥ��V�؏t��OI���0���W2t�S��� fƛ��'��k��<�Z�^O�0�»]�ܖ6.���]@�55 �e*UրMڒϹ�A)�\�e��K(����|�P�زG���h��B)�9���Ĺ�RX��9�����+��$ǚoۭ�<c-��ʋZP����s[O;u��I*����cׁ�4��͡���{�B��k�X��9�W���Y6؞�w�MHsָS�8�o��H{��*E��E�h
Zzj�4���3Ew�|��j��<"��f���}�9)�a�9�j	sD|�|BG|�҆�p<�L� ��{�&�M}��p�$�I�	���N�vM��T�FK�u��M���5���⍐S�3�[	��cD����ўB��/�*��JS�	#GW�b��o�-:&���9Lއ�	3�b�a��d�k�� )�Pk�R��7��ʅ㠋޾KH';�.�w�@�<h�}O_B��^�j�aLM�X<���ac�-�}��$(& !V2�Ε�y2��F=<I�Eo<��X߇l ��I�k�z1������t�6�n�lv�=�W����yN<M����Y�L�����ʨp4�U���VQP���/]X|���k����]�ޟ�uE���)�Ą�Om�ߙ]6/��P݀�(3Y���6g�s
����� ^R=���AB�g��24񾃔�=
�l?����2X>���z�58�-��O	��`O��E��:(�J�S�N���aнʢ�JkL��tL����0@���ƺ>$zԖ��K�-��Y:�����?΍�!��p��z�E��d^�I$Of�������M"�9�j]�x �֭��V��գ�e��;����TΕn�q�JIT�dUZR��;o{ B�S�z:�Z�M���k������\}��)�\q�D���W1F����XX�I�����T
^�Hc�>vz�S>&I+<�5Y��M�87��Ժ�o=r�����H��g����Cr�.\�F��
\��[�T�El�3�(�n���$R'�Xߙ�NҶ���)G�S˺Y8�ޱ�1�,���]��2��ݷzx��	���UU�q�T��Y�	O�+��5�P��a�S��/�|�� x�g>t����N�i�O����RRe�>|���`9*��]y�H�����jX�(����&몿�g�*;�a�%Z�Cn��g⵽�$����N��\��2=� �-�v56KɩJmc���{6�A�	��)���~�O���ԫa7/SKip��386ju�U7ji5�>�mz�8o�s�qWt�.9�ɀᰳ3o���hF�^���zv��`:�{�o��Ƴ4�؝kd��7�}�#�߮ �RG�9��Ѝ�p�����L���݈ۜg
xI�,�0�G/��;C(<]�w�c�e�9ж��T��o��Ԝ��!����7eΓ\.�(���0v�[��@p���s�m���X��Q+E��ɐpt$�-�с*٘2���#�������3�����6�AX��t9�4�>���bL��ԇ��I��O�J}�.u��͟��+GWzjr�Ǒ������Qͅ&.ad� ��Gl%����6b]�VDNT�E�
�+�����ŔN����^*�S��4�ȟ`F��A�v�O}�w@���Ťn��ܿ}0���g��]�EI_5؃���p�rz�`�I��Ͱ��52�S��*w��z����YW5vE�*AӧIe�䩔�dL�a��٩e�c,��>��2��)+~z��fE��=��<s���>����[����o%$�,,ݘ��u.!����	�¥��h4"ѣf��L��\�0?�]��b��ʳ�܇+�j<��A��yWf��\cŪ!),e���G���!�r
^����h,��jL&�:�ʹ�TMyA�+�ur8�")7#bp���&7d�`,E�j����_pwJ�` T�ֆ�� �?
^��)���k�Cl;���
W�r �0v�<-����Sȴ>7��-�k�����C�)3�_;ml���Z�4pbe�����5`�sg��3f���,R��s�|IQ��'�o��]�N�g�M����t$� �N���x��4����O��Pa'ؠ�������c�l����$Z�
ɴzpYf��^cAS��_�"G��+��f��PW��jNO)N��� ΏtX@ �Sj�k�>��@�]�yU���ۑ�F�n��)�Y�@5�<�)<%�,��/�=+kخP��A��7TBv��i����&��K�ct�K�`Ɩc u�f����7���CG�TU���%�5�`��R�b7��=��Z�LV@���L]�@��7qi`�5`։[ QQn'�bh֮T;|�47�H!W�φ^���2'��i�C��'�x�����)\��J�_��GXO������Q��Yg�?~4&�u>���+  Z����v�32OM[��X�W
��AP�L�ݶ�L�Lg�^�)�Ӭr"���DT��4�����+z�d��P>Q��:3�:<��|z,�Н���vu#߁��m��Ԍ�`��[fQc,t4���Y��r�d�j�G�ܭΒ��&�<Z�cw��1�=�UHiH�*�s%ƴF��GˌL��k�m�AQ4�{Mԍ��
X�oq�0&m^,{:
���]�Wt� �ҾT.�+��`7v��*fI%���57��K�L�YQX'/��k�kh����n2' 2�h�rM04��9P^��8��"jB� ���g@~i����gQo��;(�D�K0M��J��L5�m�^5ǿ�VۤF)�{l�w���#�w(�V�>��u�S\Z-�3�1�xzűe��!?y����J�-�Ǟ���aS,d��"p�H������ �$)Hw��Y��ӱW�p{i܏(A���[��:!�&��q���7͌�μ-,����F�	���cZ}.�0A����~��K�0O���&n\Wە�9o���иu�����U�j�G��������OЫBcB}\
��6]�o�!!����7{��M���i�i����.)�Yw��m�])����_�M����wT�l(�$�RA��>D2-h�Nd&4�JP�f���@L����ƙ���4��xMX���A�B_d��	F�8���V����o�=[��&�4`1��A��y-�8T�B�Yϵ?H�/��Ge�3�����.E�Ay��h��.�]G�����{J�:� �����k���%(m��My�g���4W֏�-"���틱��s��qn�Uf�����<j�(uNT��cU����9�6�ֿ��W�����G�;�� �n���Wn@W#jP8X�h�\�~��]��y�̈k�eQuBd�������{�p���*8|�RR�bgL+øo�����MX�d<����qpȟݰ��l�;_<Ś�*�tt�L!�4��^�P��7�Z�+ �5|�R�;��I���9��	0,�[�6K ���J�W�5���VKM� �Oy�V��1@��;8=\u���^��sQͳH�dޓ_��qT�p���l������)Jr��["��-JseRL���k"c���$�Z~Qg�O�>��!�hJ�Ζ5<�{(�V�C��U��;]�)�c7��p������/��/�^�5��/a�Y��ʠ}(�A��ov�,������攍}P�u��ZRa��]�tP�e.�-ZN������מ�3�K���+w�B���x��s�f�<)���+�3�5Sj
8m�h��5��r��>�T-d���~���͵�r�9K�;��"�3�9�}�8���5Ɔ�x�Sv���V$G[?�>e܅oh��醫)|s��08ޚ5��%��x�gf��ꙜN�[V�R^�h"'+�C%t�r,W�^��k���Mq �%u���|RF�^Ǆ���į��Ao.�/�l�ѡ
�J40���!���~��+�<Lvv\���]���1A���:(G�RAb0������uv�y���t��Z1�M1.$ŉ��8��z�q��L�	�A�w��;N��٤s�� ���T�qWȳ�r� ��)ϥ}��<��~�|@Se	Q��!O�
7���Q@��
6 b�>���O�Q\����2Q����F�c74JR�Z��A>�q�����<q1�IdX|��&W�؁��}.(%��3���]����گ��eB� ¸bK�jb ��3�['A��h�ү6|����KFF4%^���{��F�2��B���ՏfX:J�b�a�"�2*.ȂByqH���d���J�lm	�����Ǯ[w���v�n�Y[ʂ����v�^CbV�^H��=/��X��I�������*��T���Z�`jt�� v:D�k��
��;���<=�xBE�̐�z`d�yѬ���'��}:Fx�[�n����D_���h�f�$n����5F˖�$.��[��+�6N�a� �u���'q��q����F�Se�fiWt���}�
��j��n6�ۢ�'RCUܣ�3,�:�l��'~rY�V/��c�Ǻ����w���:(�}k��n�m0c���p���?Ta:��j��^}kT[��>i�V7
Ue���2����@/����(n� )yq6���¢����a�,��$(�:��5��=�,QJ5��'Σ͕|Q�i_MR:��Ri�&Qnd�k�A�Z'0C��Q:!�0�@F�;'A