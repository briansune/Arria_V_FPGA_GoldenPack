��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t���g�l��8�8A��i���;������n1尲�@̄Ԑ�ys�J���VAld�=g�8w������B�4꧀kd�n4�n�z*swl��w��br��x�J�G7ؿ�M�!�3��];�"�fX�&*E��ՒÍ}��׷s��!��a:>~�.1�!��k����}����2���YU�����4�]#�/"�*d�Z�8ˮv�WL���=�8U��0~�D9e(���ypz�e��% t�\Ώ��CɃ,��eP���o\��Q��V�@�N�T5E�*�PL�93��Sn@I��(��l���6���4�{&i#Y]�<
�D����?,e=O=G��Q1�Q���M��zG[;�p����V�
�
�Q��}=I4��/c������k�W���/�)�B��8�E�'����9���K��qmR̻0�h6�F�o��?i� ���<M;F��_qδU��i:��bN��}�r�Nky�+�g��"Zν�b%#��(�5�����Yx�U����hO&� B�E�	xЬFN�޲������6��Ѽp�K�P^ ����AJ��6e�w�;����_>�=PV���R.��J�����X/̩�NX������U#���_g�}�/����FL��zD�pa�J�uJ��Ex@F��ͼ?���?��	h�eQ_�M}�Y'���"�A$q�����4�>�w�.E�۬�o��3f�^��U$�x�
�^��|�As�]��B��F����+��v�Dƍ��ʨۄ�����S����W&���TVH��A��ժG[_��Z�*��t�M���Ӹ*����4�k���c�h�4̭��ܼ*�n��(}���<��$���d��h�C�1��F��Ey42�%�Jo�*�G�A�R�,>+7G��4:��@M��Ҫ��L�p�y��B�{i�v���(� 1����	�-���m���nz��LeʪP+s�w����RE��a��� �+�B��X�%�V���� ����OV/i��z@�<�f�?��y�s�?���k=�u^y���ל;6�,�4'�¿����с\�.v�!���C,�V��c�|�4����1�'��.O�rN�8*-kW]o��t�ڞ��U����B/��cX�U��NM�)�R����
w8�ʘ������@6ILȘ���j���fN�Ӆ����Q�yg:�Aq��Ͽ[�e�R�
3M�lT� C�= ��Q�@�e\{Yi�o��qz !;"��z��ڔ/c�9Ư{MgMHa�oED���*���ޡH��՟7��-�����ҍ1�H]X+dH�uױA=0�g����v�C�T���Ңt<'�f��\x�̌Km���O���σ��陜.M���ۿ�FZ����!]l�݈��@�w���U��C�D�u���;N��:߃�����M��G�E{���͌Qԇ�b���ׯ�_@K¤���w�~�}���7�%YF��췝��Z��A�j���ҩ#%w����?����*������/o�zf�
���Ű�h)�S~���0���l�I:7���h��Vx|������(�~�� ��3���5�D�f�>���\�@	WH�d"_(C���l+�Y��Io���Qx��0[�6v�*�5��GL/÷N�&Cm�/�uEm��I�l�ڏ,��-�z��HK��p���j��� $�c1N����Q}��	�B�bWP^��=�,=�d���k����[�*�1�4�N��R*�)�=Wcg�B{�g�	G��jTE�.TZ���0F�ɭ�;=�+4`�q�.wG�1�Z������!/!��}���ii�C!�Eکcj�Z��+1UU���l4Ҥx0��h
�1�ζzc10{�H�=xբ��	��7kX<Йt#�yA����7�I\�߀xW=6/��4xo���j��7�;Q�rБ�U3o��e1�?5�� �"�앫��>l���m���}ȕ���tJqg����>O@SKe�u$7=��Q
����'��eި_�����OY�)���O�%Ɗ�P���,�r�؉Ȉ���8�]Đ�_��#wԪ_U`%Sr�A��^���3ֹ���w��`=�ۦ2��9V�� ��?{�~a5+��	lU5��M�ax s�,Sy��8�9���s�E���8�
�E`�mjͥh���
�WD�O�o�t�**����e2����?�'�A�&et��(3׵9p��p5���c�����p�Ė�dI�`BJ蚷�LdhZΩ���of:ƪԐnϕn��Ͷ *�:�t�.�"Z���%�a��:	��PR~�=~'Ѫ���ذ�d�P-�u�f�Y��(YkJ�\6�M?��qb��.��P�6/���X�87V��]�"R-���b�7n������܀����R:�z`�K�?臲�bF\ߋ|���LX�N�Xr,��]���7Fc�%�;�wnr���|=�t�,��K�����%b��Vꐑ�Y�y�ab�s��R	��lA���۷,"a�01/���%Y�6ϵ쪦.u�7�Gࡱ.ˌ����Z\�P�5��(H�����~�w��&۶��)d�f\�� �g��{�7��ͱ$.�i�s_�ɨLy��h5`ɤLH����X�S������ ��A|@��:p��y���J�u��ɒ������|V�����/^o�/�i�g�|Т�*��M�ԁc�<��<�.3�ݑ/��S#�U�����&�����8,If	h^�>�����[E!�>9�Yܴ��ȞMr�F��ύugMH����H�R(������u�1|{�����UMx�eR���k �l#�F^몃�>욼�:_?i����`�E���L���YJ��E�X���Da���5$K�Q�\�SG�a��6���WD��2�Yo��6KB�c��(E=Uub�{�,���d�B{T�&_k�=cR5-�r��)F��S�~r���)��lk3�m�N��81 A>��i�r�@в�YDb��`�1����mQ�2A�R%x���?��'c􌍶�z�j��j�t�tTQU��S˄�5f���b�*����PBLsr���Y�6|��yu�͚w0�-�6�7�͒�P��EK�|.X����Ґ��D��+�Y�pu���(�Y���m���9;"q��_��rW���Uޮ��+X/(�̡�� ��g�Z�5*=�a�l9����e7r�pk�P}����Pc�!����6���m����`C5��,k����2d�P�V󧁰�}�c�@��~㟊t���*��xW5=y�h���O��B'�ݴ�z�|am�a�2�.h�=d�7�V�w*�:K�l�O���� �N	@�$��j�I�ap�NQ�_f��������'ү���M�Y2S[�e�,nxv�k��M�N����T�<�m;0�d��	���
��1�+l���>|�����TR�]�R�|�ிrh �+���7X���#�]'�C��}%ݎ�(�A���:�kyM�Sȫ��Eǎ{�O	�8����:/-�J���W��q�+dS��^j瀿-��;OY7Zíp�>��$\��e��?rp��</��,��Ť7p��N��Q�ӵ�p��T`&jT*��=X\�S�S�����lD��6srE�!_N�T�~�+\Bc��i��q���3/��ǀ���A��aJc��]J�U��������;�,�g֍�9�T���F�w�S!c��H;�D��XAr��Z�?x'�������*��&��X���x0�=���8]_��\����Y�us�HPE�k޺�
n2B���Z9h8�ZzE �� ��L��?�Ǥ�%4����#đ�\";S������e��d�yy��!p�|3w�I�Վ���\~L]��;�)BEAN��PP�8�˪Y~�U,����a!fK�)�M���w�w �Y�P2d�T�*`�j� �y����}��'T�l���m���G�'Q� o��Kl�Y|�Up�5�E��
y�@75�&�ވ�� �,�#��/Ԛ�vWN?Qf֗q�{��+�ڞ3���'r@�����$OU8CE
'F�c.4���r��⺽AGV<dg/�γq̿~��$�a��R��2Ga%�'>Q������ؑ�兰հ�/�y�ɇ��Ú- ��-��z��2�3嘆IV�2�w�;��[8�{�Y�!�GM�0��~����(˵؇���Rd�����pΪ:���3 �;3��&�XU�����.��g,^�o:�2e������c��d�b���!.���2e��v��@Y�xr2O@��]W<��(3���W8�*�r/ �~����/b%��$��ܭ��P�2O9�5^w@7����cW�s�p�arٟȯ$�T Y����DC��7Y �����D�\��M�~L>��]ƺ3bfk=n�;�u�ľ�3+9Q���%y <̐\����?��b�\��љE�����,�F̯�	�-<�A�����{����-6q��z~4�w�;%L������y��/Ȣ5p�W:��>{������yz����E�c��^غ����K�/����ai��7#S���X7���sL>����g�ō%�1Q�������h�zc`��2��`�ʋ�1QPJh~17�^�&�F_Q�$ă��*I��Ë�ϐ��!�������\�P�@��{ڙ��/S��M��3�=F<T@N����֑��
��sB�����{���q�F�E�T�"�!�V����$��5|�� $Qm��"m;���|n�q�|E������6�������k,` �Z�f� Q�S&��;ր�3��Ö��p��z�м_���w7%\F�����(�l�;XL��e0/�<���;r(Ν��m�Qʀ�W���Q�Zi�"�54��׋S�H��ǵ�$h7��Y�DU����F���������!�Hq��'�I�̲>�<��TR�TY	�`T~��p�����U�ح�呣����;V~�.�����D0̯�;�>G�@�i4#f��m�]_-�0�_swb�{hX̕h���J��P����\��sΠ���P��W8��=<{�!'�����rhaQh�;���J�S�|W���)@�J��H��(�����a�nEs�l�S)�\���xd<�����2DH:�"�g\o�D�C��~Q479�7E4�0��N�?E�Ez�Ktj�zޖ\�-rq�|`�K���mb�}LH1�½�|� ���;SR|�Oe(�B�J�\����{�_d+M�>;0C���d}P	˞
��
�ݕ\DȮۥ�*Nv��a��=#�7P`/{�\����)$��DW����h�^ϯ�
Wh�Խk1�D�Icm���-XQ����+�u�эG�0�s*����#&����J�C
hɾ֗> %-A��r<4+�q.��+?��h1աl��UK{/��%lm�{�~�u�A��tiNe�l,�w�z�4t�#�Kǯb�m,�����H�ۛ{�~H�c	�
��)t,��~r�JőkG�����~uۼK����R̺녗��W��Wx:v-]�5^��ҼMy��<!m�KR��V�@Rx�@C�ĠMp��r�-��X^u��b��n��l��։�0��$�$�の&�0����qf��̑����c�Ͻ�ds�ʭ�����ll+�1�-\D�P��� &mt5)���cI�Է��@_��21XUV,p�U ��`�9�zR�8��F<�ym�	�)�F%������2#���C�D���?�b ��f�N���s��H\���<'�7\�)����
��2>/�$�7�&�L��7������ػ@v{�C1���³������U��'T��z���
/���o��B3�>�H�� ��1`����P��:��5�-٧'�K��_���j;i���l���f�m(���W��?�x
���k�2�p��0A��ъ@�]E���\͖�
7����=���,T�AX;�r����F�=����c���E�p��n@�>M�_r����p!3��Oc����xFq������0�>��_�V�#꯵��*���澰�|����e�y��2�=_V�~]+���j�9�1�"�ס��$��e����'yG����/5H���ce��M�Ll��藡k�N���c�ԻR�W	��- �}��J�[%xv����.D.d��u��B�c�����O$يr����g�G�/�q�O�s^�X�m����;ә]9I�Z���Wnq|�ǩ$�s	ج4ꋞ��j)s��ӻ��<��#(�V���Ţ��DC�s�>���~�-/D%˜�b��T|�ȳJqn�4����13=�%��]��$�*8�Y\�i��H�������ɪH���AQf:�\�Ν�;tw&K*^#�ğɝW\D����v�v4�CV��A'>p{|���r,�f��o\]7���X�m�2�����/zMx���4������:]�3����v_��V��p	�+z��p�CW)��R�hJ�PZC8�A��6B稦J�]�̰w�Q�[��s�I%��+0��O�JQ�{��q=��
�������*!,u:�J�>����F�V� ��WEAN�L��߁���﹕>a����3�9dF(�=��Į�`�r�ɕ௨++e�����}��̻	C��뀓q��g���d�:�wM���L�_�vj����{
r����"o�>/)�PI`�-�6s��*t�$�;m��B�O�H9�sM*c��ר��dex���,��|���3ZN��PD2(��[�UyAI������i4k� ���;��#�}A��8���g�`t䟔��[HH &��I��)I�_	m�r�g��4022�a �|Rl�Ozz���0r5<��D^X�����˧�.-�$���'?q�}t�ă��l��ԦF��]����^�Y�R��E�
�5#1��k���{S��Dו�蜐)�G՘[r�{�F ���l��v��F��F�J�� ���-�]ࡋ]�|su�O,Ѧk>�_(�8a^Dw�3�c9�x3�v���4S�*ٿo��� !�{Px��@��J���r�r�QS{_���Õ}�����%ܣ�):Tr��Q[�4ۏ��R�粿G�Yzؙ�=ےR1+c'����^��`�*Db���N��/> ǲ|;"��I�����V�BZ�]��X��2P���۳����+p���n/�D�0,7pb�6���i���G(���}��eA�O�Wx��� uF���@YK�0��2�Ȩ�5��� �'磫��]��\�o�a�c~zL���� ��E��6I+��%��	���50�h��E��<�����"�+�p�{