// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:27 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YcQCzgyKIxIcNkEbqUZLOJRgX4U4BDg/3fXQW7OvLRrLJIdx9y9JOjE2vi7D+/7r
1VS0wwe9iC9UJRfLzWg1nCf5iwcAEAYUQ2JEVyuGl5+Qd8aqLESorHd33m37svZw
F3aGyoub8JmsPe1YqbGbqvjNxDvV0sRXnB5uH404Pyk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
974zmo85cMx+8u5z6pvmuaheXp8iPQFzlbNrXf62v4hOR5TWJpE/NJYo8LFXspcb
CH+4pLmGmQLlHrkkW9aFGdIxJhV9anZoynczfnGZEgQTxD6hgm5aOBcOxDnKoYFg
PM5smIdFNE0XB9IRBGg/qKbtD4KvVMImtAm/o5RztjLjsAMDpjFnLENwdOIPGKWE
R9gCRSfRyu502yXvDKDDb1MmsTjYETsnwCGyvUPwiRepfNQXspWqpru3Gk4U36rZ
VSpT4nekFZhUddFkTbtLuwDjoVW+D9I1nva5mUlAQ/tmBftPK37XHKIN9ZK2Tzcb
ltfdOzK693vufJycwrUqKMlvrkZZbKqF/zlT1eI8XH7WON/jDK506DotVhENZOkH
DUGF8t8QZnIpxgfmFCt7rFeLesZhxdLxtE6Qfex1ChsyRoCKH0yW9xecFtClsH8G
tnChAYZb5kNT8e8RoAW3Q2bVs1ADrg6lTzi/nk5s2ROJBBslJBxeHvdDoLyWUh7b
T0B1JV4t1IKOwWovBytiEfmSC21UG0gIUu94/jZ3UANnCwGT3P58OGGa4Ps4FwDe
4Ui/WRgbcWiad0FqqCnU9Ip47FiXRSmNSCbXGazeDNBw3O/OcuXEgcFo8BeIdTmG
ANSGe2PTd+gAZEVjsnfo/saB2dURfZTbBF8Y8OcGkMaEhpeaASecDZxVK5PO3Y0y
0D6UQOo1P3V5AyXCLk88zHv99bAfMcOjxHMYOoqDjl+pwX9K4i5CajfvdZohzk8p
dtUWuYXKVbaLGlc1hi3Dl7QnmMMsPFj4Ulw/F32J+9ll6FsyZaruagSZ+cZJVZ3e
4swogUjK8eC1pBnfNlfYT/RNncTC/tF0qIrG4lpPlFK1F01D8xFn5jsLhJvXTgy9
5PRap4E/oOsixgG+iY02hY8KNK5M/UzPwM5/+uQFGdLuyBTa37y897tU/Thiz5NA
KAzw2Ug1Blm15oo1xf1r7cjbg3vL9yWgTU52U4A6o8D7NC1AaKH5p+ROYmnuoWzK
7E4cvIIEKSZaTsUW1Tv9GVeUbXt7sTvhgRN6flBlzuqIxegHdJl8d3cfDVANKZhq
WNwttJUynKHZ16UacfD5Q8TeoqJzYhTQHLUzR92kMb0u8lAkkg6sOwOAKv1aT5Ik
E+jDvLvjdBImp0M1jg/WVOjxI+zn/jKpxlPD6Ag25sB0qQx+mTIFKRzVJhO9PFUU
b85aDY6BCMiIeYC7alsIrr+SEEs3jfO+P/8GL4mSd7T8qtSmi2EvyYUZz/eGVW4a
medz72s8KwPhgwMLJrvpvOUkTmKBKw56F9v0YTa2cVIVHkQ97kAb5T2V/zfhkOcg
Wz3e3tFC+pvrtUTqjYXjLLBsiF6P1LBYTkvF/mr3asX02veVokGguXCwEF2ufqSd
40UdVZDqXmCKNj90jPyxVfD44MrhoNVDUTPelN2AnRlBrxPyqiuHBArK3JVBS+Ee
+fzepWdtgKGO7CFcptJWC3DgMK4xSywBgXMsMFzGyjk+t35tQiOOaECFTYWSPcjd
d7JjKUV6cWdAonJ8Zgd4SB17e3TxPYL3de8pn4vi0PmsYvBOeN2xX9Yf2b7HN9YP
GPijP1/yV7PZhCqD94zCwbFjZHJlppWfEhzp3w3Eksu56QUISI9C7LyUOeZ4ratA
BFdBded91g25IHoRKcqiMg2Ox+BNdhDBefeWUjAi1XstJVPF5WHW9RXK+kn3cEa3
8MQXkJ22/Ce8qbB8N6Ut042N+ji7m/jUr+Q/bvdJA2iIBhaXjCu9buoRuON+Uk0t
eKvbEDQMUpsy8UoTiKtyaZcriB7p+FGl5q0omyHCDGjVdI9QxdjSN0pYjPTeeQqd
cNOZQcn50Vy2cVXuOn2mV2ashS/WpjYSfz1LD/4Mpwe4gfSRaGIUYJZVFbhuN2c9
Nucl60YTclND61I8T2D5r3A5e95jJ0LGWnF6cBEyL6Zm9T8gj9cjgOv+hCVIIb33
7C8XeAFc9jij8PJ6gzIY5PQlsubWMbPlf+6glczOJ/lAXeeK9y+kbTQzU80fo7AF
U2AgnEALqgi6u0u/5UNSxn7AqwrBaoGyqb8e3x95iOwL+s3gA69OqszhfA9H3VlJ
vV0gOnEbH4xC2ninoiIrHR0Ffz/6+Bge5AVzBgC5ajCfCvrBIU2CYEPkmM6NaoHU
c6ENK3VPEhw3qDgeiI35OyUPHev1ziypcOM/LcUKtfGAAsJZzNsqDuHakxmh2xa7
dMNIU5vrt/xG2ITawmpyBtaBSW+U/F8GIbQfq+UJvjFLBieKHhU7KvrlIiqF5d44
zs9/QP0gumgd+XQJnxFCEXGwVzaRhWWSYpH40wBQDyf9ePFJTLQWXWk8rIYn54yU
xs0o+9GqzHw6RBQOptgjYfYK8AX3wIJXuZ9GBxo3ReBuMHZNqwxhs7Se2T/3UlBe
Pmf0baAMX1ryK+S5Frt/P/XsG1oWDlpZTupr6jw8ooEMJJmxCnm3M0P5ui63KXqu
3LSVCd4ORQk6hlNpMc/fjH7aJ/Q7TX+svgARRlHVihdkCsw4hM3gg3ZL5U9dejI2
GeUFnRfBIfDphlUFnKn0eTev10VJBBxRUV06bIquIm0VxNcmySYFybRBgVxKDmBe
w7V882/IgMcqtURTZhevZyDQAShPyyUBXkqzpHa2cAEXQ7EnzWn/ZDvbD7ykJ0gb
61jQhkY9wvCAcis6wuSfBppMFK55iDtns/IXagOqLGxd+NYd/IcfxH93BxzGefkX
4H9eEFwaLCk7C2tXTdlfGnbZBXo6irMw/8dmX68xbUlhPRTO3tG+dOMcoSHXfiKX
ylLxWa/Q1KZC2Yq/xph5WCPyTCWF/XWqmfoVduGjiFcKF0499EUY73b+C7AL18IB
F/9JvfBntkxYoISUT9ZmsNxiyqaPZKoViKJFZPyLowUd3RwdKLeiWygS5FHTDQ1B
n/l/HrTyy6nOfxtyxAvsRZuiy3dbhEVuMJp63Fq2QTW2S4uZsqG8mrqU7lcJDfjO
QqmHxdM03AAEsdlL4fg6K/i2jZp/LewsF9lFaPFuTvBJwvi6z9MUAhrdLEz1UVUA
5VbGRvwDSGERrW83y82i5j7cOdCpmlUv38CroQpQi+CgG1XoXep3Zn+q7dq4BRcc
Iep2xWwR4WcK/glSvOeAr7C01WgRLvX/AkDMJtnoxzr9ZEkMLDQJeRrLk6wnaKBk
byOIszVuMYwcTjKxZuc4gUu9/2OXKvrkknLg/ywGCpA0q7hwkDUCmciykJ1JVySc
V5Je8VYsLVTvwkgzi4bWQeKvnhsTU/00wos2SBENdl6w6XJiUoKW6gtM6CJMP49I
S65XB7vt2YvKXBoqi4mEyrED75FqhA/yF5w+gdZ4lmDayXW6d0Wzg/R4JUvbLYkn
ST4M5uMUxeKY204t49sK3X8qjIJctRFs/k51Jp+Xyw865vAxp5tYB8qlLbwItPlW
ty9VQajNaXS0rTm7w09BbfooczpGKefJ1cIl5k6HL/HPQdncA1tEAmk12MV3eNGI
sZM7ZmNPtZHmTagmnV6ZhlItoX6Tg/1baB3pSXamiG3KW+lE8Ju30zHvLIs+YHQh
17j8HGvvOywMbXqKRwvfMcMXWECHVf5+eLsNysUx8Bsy4aOHmTvrbHlmLO4tij+z
phtuihcEhfMpfZ9Bj8I94PfeD5rBghMjX7g+3bR7x4VVWDR9BW2smaN+eUeDp1bw
+zX1DCMCNsPbg3gZ5VAXXWcGnL7NVrc48KHgg927rYSd2pW6ojehX+RBsFSXEQye
pCkjOkRWJOb6X5jzXt7D1Z7IDmJiCYnjl4zcRf9t0ToStyQHybEEfvOkSVuIiGuF
n/m4T6dQIm1mKtlGF0ejFGqd61K2rhUiKYlutKKNuj3q67RWYjLbXG/zZby0+trw
qeUbHBkJBftlrasv9dr6dcgYug2fRaqpGCyTtNqyaLx/nti6zm4RuFUw5rUyGy/W
DBeN6c3VN4oHLlx67+Z5N4nbczPeNDtla6yxWO7TIlMuQ4NZMKgwf3K3/7ZEjRFi
t7SOjJuoefXxBN2O1g98m9D4dfHcgiO2hqcB3UT3w/fPJdZPboCCFkWuX631nBGQ
4GUrVyJ/pCk0uhQLnK636dfFKoKZ79f66uJBBxt6pdCWNkQOFxbBzzPCSOmrH5y4
/rORZr3lBE5lt+hcM4sqisqcynlAkf35cp7kMZiBolANaqNFkPZb/OvKpbQBD81v
x8wwvb9lJNKhzUbBRQQzXNDcTamz5cu92XtdQbFswuWTH7EyQqpWS7vwdDDlN3PI
W5u77IBTTl5gmirGqLD/MBcjHwb1/j+UKjetSxiXlamm9wtTuSFpoWY0B1AVUBsn
NoA54C5d4gOrecjRG/6B0V59DIFb1YPkY/Bp+0PORQkWONOcVZlIZjhhmtoqdC4t
97zK65IHyDGe+CsbMf1oNhpfN9ecR5GOWgglLVcyL1VzIAQyOJsV4uori2NJULYt
/JYhsQ5FELHw2D3/3gxk5JbOB+IzVwP0fa/vj/1dehLrctm8bWDOV+ohtHxo/wun
lV2LZMQd/gPSPFqLPvgx/MxuyLgIa+MRA6a+J2mnbEITRoTlOVBDitDg0+OmRgGK
gtW3r5+l37D3TjTbOkzVI+J1onXrE1Xw8ePpq9PEufKYQJJX9pNAH+u5MsYW2juW
zkPDeyGSJ9cTwH4vraUjBsFTTKR4I7Cg9yomlVYOgRem7srBBW5S6hTZ/LYx8kBn
50M2CjRJBHED1Z/xWBGd6L50g7uloDVVfISO6kNYkkmosKMHzUEGgkLX2uy0gZTC
HdeWj0H6d9XOf9i0jsQogpyMax9s7wegFK/d5/G/ArrwYjdVYMg8tNvF3TsYWaLF
rZnezGFqhdoLXkKyYYOqsGHq+0yyyP/0wPuK8yBtco+xXY2mVcP3HlXRqTp0cAsp
yKx4Ds752mNcNn127JPZyJucS/S3nw7+SZ9tBVC9QK78lBqNWgD9PYkpBeOLrYL2
AFQMQdn7jOnyUvo6kF5TKpLc16PDO9+5eoGEsA+THDR7a3YWeiwmoI2UYEBGleTg
wXo1Mkavpc6ZCn6B/cPPyFnmqQNYAj9NMlzKZMUETFD9yuWYEesG98tYiM3OPEUn
BmT/aWmhhj46pN/5E78vNPU2RAe38X2qYk3oVnZgB8N1iYmBvLg+MC2du3PhVI7D
GGpIkVaCBIhXVKNQwrwdVOGJXcXAvv7jUwakVWctN3BsyeUNuG/UI3G9D8hrHZF+
KfJkDnniTvuDgupraRMyvBSNkdkouqPWsuoate1sYuh0CR8GlrCzfjbgEqXm63m/
GY7JTOoN9nM6D36+nCJU17kYmaK/6eAFzhK2+muf2wUxXGesxKcj88O4nCpZKIZH
vfdJJKIPj/XJmt6vN63FwALZHsVpEULX/6OoVmygvKj5LtM1DMSQRnlWGDb/jd9q
sLjkXzVXAQnQU+6zhMMyEVR0GtjvaMKuKxhEubKL89N662UhqVqCG8o3Ui7wxpIJ
I2mKSTB/Pe06AhLIxOBG+jWVLHQcXY2E79bTSP7lSlWAWW66LvyxIQjce1IgsMzw
3Li5itdx/+pCpzh0LuS0bywkJqh9//8FL3gIJ+fYsPNiHB/JUUyYi1T2HJQJH8LB
o03if9rQ/leeaJNFhS8rljP5Ceax3k8zLp3IR2JAypar5EQ/1jgujPt91F8onlVg
h/Ul2MTJZ3ljaR5Llqm3MUqZYYfD5/6ekaL2enHn53RvWl0c2msRRliow/Nhvmks
HTgZYnaU7aR+jj5Kd4i/1pu+oSNt0HChvrn/6PfCkGgZ4qC+NiOvWHVJVDbK1uot
5XFYFvnIzx1cF5njrnD5Cj4XVJVlQ6vwBvmt7S3L3SzqfCY3Hu66ScadeqGG6AL+
V8PQJvjo1ZKPCOwJcdrU9VtU/IBjfDLVGoUMm4BJ1iL4jNOQnfHbpb7j8eLoKt+z
cQLu8C8AAEhVj2FJwoCgJYI7U+NzVljM4jOEzqNcq3fimWOW0XPa7LUYyvI8jcTA
FfvAzBotxuTcvqbOVagPscr7su+NnGGbQBvoB+g0rUwpyeUYxiOgpjXjJ1sWShfx
jVUZ8Rqr5xRxEFpxLvKDZFhnGLI3TDISBpNfW7XRBhYQNXB0+zEQgBh1tGBgZX55
V4I31eJfJDpUU2lLVcbgCOT5u6tNHuILR3w4StRnEkkyE99NFwbWiC7++kvv/vUJ
z9Gn1mZjTO+c7NxVOrXjhI5OQXNb36Z6QNsQnrzKBOPl+KD0BIi+IJI6hS8NT7Sy
o3trjB5ueSGbapCihoCVrSL5aZIHAfsRy/w5Gye4RfXb4Kzq4i++N6jzGDI/MJZ8
jCPiMNQqUJPtj9jIUzMPXRsyhXt4ibj2Xw84tJcKZMzFbvduAz3gFsvEiS0gNkwL
evNu1RZK0410Xuq1U424KAW0wDSURvSYoHuEUqbs6HuzwY6Pkg1Is3ZkMmSHWhC2
6ereG1wovfF0sOYCEnax5bjv75Ob1cP1P+JDlBhuWGrglWl+Mi7JfKJJYqShpXLQ
c3tr6QumzJz3UUMWlxpH5jWsSWri8d+EVlbxwVZetYnQ96Wq53wDI4flvIn7Z94L
Gy7OiHBXibo0KX8D8G/VTbUgY1UPiINlcNyIoAEd3avN+eKolk+q2fc119FXoog+
MJQ52kH6xMDKadeTg6CKGjWb4W3ZX4oXjEI+WMv4pWxCptvlRtOsxxfwb37WEp/W
zfC6eUXK7FxJI9aJj1KDszvf+gRldDfXK7PyIaRSMFf+iZKBg/MU5MMvLbFkflU5
Pgn1nLqnVOGAzmiTFPUe2ByeoVZVGtHkz9qApUwL+fsK3AKgah078EwTP2Ke+rMJ
da6/mkGC2xoNOY7hcEanM4Lu353bhIdu6+21o/nRbLEMuOgGMNc5MVv3DObALm/u
ZTQyTatTggvCBHfPtdj/7qf/g0ksppG9q3phuGSrZLiKdubAGR9iElNpVBaGacnv
8kr3LjBzgFeT/rFZl/yP0rv90ZWK07yT1H0wU8O52WscuFkA29dyuYEXFiZdN5VV
BzXquHMLnIsxr9/Voq9hGskEtsuMGiA9Qd53hPgoimWedyVoJI5FZRZlAWuYp56U
LSMEub7D1rA0B+QQbeLfi/97Ed6dJO+fPFY7z+idpKs9+1gSh3jLVN4a++AJj2NR
6ZNnnh/pDVSZ5+g0Mpaf+O7KhFJJrx4FsLV3LnAPqa+9NCpktyDGYNczoHnPwfRQ
fmQTsqIEWEICuU/59AbMywRlfDHxRSKQUBr46QKBZc712nMHKUj4t3g1zUpl8O3o
NKDrteNL60t6Q7vhWnZESk+NvjkFE5hO5EkTW1+pV0CWArvFf+vBtmUdeYDmOwik
lPmEXc0Csaw2JGsjtJu1j6zcjKGHnr+E3OAC5K/BqTUQwZlAXXBPv9XiVvVjPFvO
lhlro2mBxTtHFF38RhxjY3uj+IWnaO9qy3DCy9C2jw2nZSwFiFt7Tfa7CXvdx0aP
WnepCv00v9N5rNJupdO4Hj59Z4BpsgHmPdW5D8K2j7FvbkeirYb2pj3ZrvsQR7ke
kU+HKyN2/YBK/Wn/cikNSI8IgFA1Js4tQxFEiVo7WflhOfZljo7SdI+0TPrbI1mT
`pragma protect end_protected
