// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:21 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GyJXkwExQ/0kMkCTA7OS+3LhPPuO3MIAtP/eXh4aeNah9dzDc1+v0DkDbzN5s27M
T7lbVgziSWo0t9PeXk404vmHFEULW/hGXv/fHQk5QitHmYEYhYhzYbnQeCN4W+W8
8Ft2KWi6m6z2Lzb/A6BLQgWT/wRVZneQ6pNM3UNpukA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
aMzzfNKYW0dLC980Pr9EGDztdbWjR+fWq20AcoDl1Apa9AprRzbCQ+Jea8OTQhYw
TXeYX8wgv5QhDpl308vte5yJCBtg3XIxp2hA0LAinWPks1+SUb3PlhBXvXLL+NIV
4MBR7zgk1MZCSE8toRAFMKNJkflvxSNjfEVr5eq0W3IBsHwAY5MjexWrE7I8zfUV
HrjjVxVl+LZlEYONiwRlOXu/TIjptnj6eVLrnE83V4fgCyxViySkiXyPpnBF/9IW
gkvr9BpO+/QE+vz/3AOMqRAnno83/+CCRNBWcCLn7wkzp/mrPMyNIndESN6CZzd1
77FA6xl506ggfOI+wUSr0SFM5NjkDFLYLcYXiZlJvrcG7AHs0Ydu9pfVstQFmo/M
ynxIql0kTn0WOsN384uID3+EtEMNIbP02xlBYRIYkqgzbggEdXNcl+mKzR6TEpyX
Txo24/wAmBFQiDsGXdGj5xEDh1M9/V8Dllkc3MX4sLcRGyzxRlMGiNuG1vyTxNBO
G78qWPNn6EwPdi1WKyh2Xqh5M8Ngc3dAZ1LGhEVQbk0y1acWjXSPUyNG4sWYjK9L
T7Akmr6eHU3SETAOgee9tZQ2bWXHMEvkWuC17ASrnFqcZvK4xRKzD9LMeXLz84et
GKFBYs7+QSFtYBpxluzy5J1h6E487ukSzF2MJbiLYyPP7oqgGAJZ1TqaTkHwZ/8A
GS1R1/U6jztqU0L6poku+x+YfPxR00q1fDJn5EISbyDqpxl2jNkpvvmLLwhPQBDC
25Pe/Cspd0JvwALZOHGUY1SlPL64MVmE4DHReMYFRRvCvhgBtsDrySMZFJCxnp11
sO6JKzkRVsK5QsI9OzfOy7XccfyFFY9vJpRmVNMWPhixozxHSCEWzVz6Lf3Bip4q
VuqoeYLvMG/Q/PwNajqLkmG8R49/wGmhnxYodrH+U5LJBCN5WgZR56lubNF50f1/
NjLvXUHV2lY1PJHJ+rhx8wf+BM0vACiR3112LJKFYuJafc49Ef8ze7Dk9vuxFq/4
1/EfFXYjlc2Wg8ijEAsBLINe4/+sVeFxMnTpq6hhGTqrcn5Pjxu1Mw3lSJd/AX6x
ZVXBoSecfRfIrJQLNTOSp4X5HyHbdH5hRnHxrDkbszu1fT6g8BkxEon1QqChyZgL
sz+rRw0xoY7CFKhyBx0B3IOHbGD4elBa2niHWqRC/hIZ8f6DqUiD0pZ8ExBqrfOZ
Ft5ikwHaL3H22D3nMyZPXsdhQZ1ilWmN2KZsIeUPJkpxSMi+OPXbQNUEgEAkpqnE
N/UbtipDqXT5uBDT8etpAsd0bIzLGA/T/kyFDAevO/0gZUDANSIpdUS2TA5WEdmr
Q3z+52qoZV69Pki9Fq07JPzwMaaJJq/28i876FEkf5Qom/5touspXwhbSOqikBnK
KO9jtNJbBTCCL8o+Qu+lXZX5QTQALbTWe77PUBXptwEq4pEF4fu51EnUxRzFHtgx
MDfUwc+UheMoMK6dJhjgiQX9xJRq2MGLNqkCYPkQPs1BZ+2JqUjYH/t015QLJrAT
C7ukPuL4mc5M3LtrlmmwZDqbwxEqF4/MK7w3ODDiCWgTZconDcnwVkKjs1eLuOy/
3TbZ4I1cqlfQIxjSozvewvNAEAwsjBj0Kg9dmIDLi+snHTFQz2YJokmQl9cPnPEr
E/qZtYRB5qKqOgOpHdGRGBcyIt2EpthrUnIwnxnf3I7XmrTUYgGh/2KHJUoBgzrq
SB1f6RiqlcwwbTi81/U0b2CvfrqhGbjW0O2udniRYxUJyvyHepuzQggbMKZy5+wX
SfyH79k/oAmO3EMXGDP8DkcTMVeYhZOsYEyung8W2n2rKwLhdnq1/Hz1SxhtGRA9
+HJFRqv59K0wutzfp7G3UlPjXBZl74WqVcDTe+hkK7UI1Fxs4i28jNYJb91hPOGg
Ty+RcgwZSnnxSsVC4o8CmQTFlqxvGBDGPWJBRMOPgdy+Rb63Jbnqs8jwMD2T2aVf
u3zE5HmEQeksuOvdzVTMTT9HywXCLe6i4xHVMUseJxJ75tO89Dm2PhWqFdeSRf5d
5dorY9d7kqAN2D8BGLg4giSUvIaEy5QpsAr/RfWlUCah4nX+FB2pvRY7mI5f1SkB
+C6gYr40jBUuGoer4HDm87vPGdAVcNWfOtGLatkUyy5uVzOjMRFuppt1/cjBGC8l
grikAIb4oJdr/Ijes546KAUdu9orwbN9denRjSQ5wfOYER7K0X/Dsahl+muT+E9C
AHo3DZ6AHAkmyKp7Ss3BN9mXrLAMffvD0C0fxocRxyMzjBhojcUXcd2DX9Zdk/dl
sSIOR3yjpuePhfB7a36qOhKtXRjb9GiTNKVCV9Qc0ZRET8YIz94m2qVzQ2p1aLSx
636FhMDU6fJ5qQkKJu1VSnvkB7wBZVBiWkvOo01NYj1/t2PNtcwrzYdgNqtDAIoP
mtGw+fKEmOzbOnpmu6TUkHgrTPlRFdkQBB1LoaNqfRXr5go+4xe/SmRpxfjpp4B/
RjIU4hYluA8oSAA0G+Asj8XnkUC6TjJ36rO6uybCrCtfimq8byOl24kE+EXN7TeI
xPyz/OnKmZ7qEqMkFRjsXnmQNCuYgfdDLn8LMCMsijG01ed29deUCXz6Z5OOHLQD
3XhcF9GclIGCUmv60Gsb3AuoQyo6+sqmqRgmZVkSkOZmfsartVWX47G3WYpTobLW
hnvNdIaC/i0lmObjvV7XxWGSKw83lnoimlumwUgoJn5lorKY08bqdO2RLKfL2VRa
rNnFu1ntje5Q/CFSIvh02TdBo/OXTHFvnORs4g4MN4dNRl6JosWx2SvFvG12eNda
VxlCIIhRSl8S7B/h5yUuKe3qDiaYdmr1pbRkX+nC7v5Api7lI+APGubN/IY0tt9b
oR+L8WkLyDtB0aCDUKJQ432iFJW6qHeNILCESrsvSsEH2UOywNQsBID59f7Qxz1l
KXFZQ5d90Vpx/om+SAR0fIBk0i8cHrlQAdcGXuBRKyExa8LMSzsRZuC4Q+XBWiya
KkowQOMfxXOv0iyYLa/SPJceVJ32h7saDaV+54XHKEWlW1vVl9Z6u/sB8BhT06Th
vLlVCozflXYYFkAU13F7ETkviVtETvK1IEDJ/Kknfzd5IsfPAOSaWWPPpYMDkhR6
ZqJWsCZCiQzpGGzay+f8lqBVVbtkF7GqSlvcpW/uQmg45vyTu01EDFsiIWkznmrS
eQnbhH2ZKdeYSRMZkMINn+Sawe6bANyVBdGESS0ZCu17s4sVaTsCJq+Qb/auKt5Z
4e+JEDUYBO9JE8UNPZZL5qP0OCuWfM/fuzGN5DFn+SEtHsGqSg6i1wUQc8Gu3xLI
lRPsgVydC3zUJU0SiQA87jQaMXYl0ZE2j5vPHZZCYzBvGqTFrQ4kLZX/52uOgV3K
QekJQq9tXlC3mLxWDdThXSSFzHAvqDAzAB886NxGcLECRqBfMbdqrAAodhrPahVs
JwVmRYbfpifpygR4ta2h3PZHBmIgs8Pyl3yH2cooEuX0X2UvnntBWPWH8Jleoium
Y3O7aHhralrmpOkgm3Hvz29mfxo7y5CEein3KkyIMmCTE09LmUsoQ4yhw9J4jbYV
+3tGFdhtveXmDLBneHG5Bc63wqeBR7CV+0cK2/UXJMy52MNjlI4q44WvgkqNR94E
oP0RC3Fjezo100eNWNkYAmk6wDlZdCyv180V51rqZZibtAfAhNjt4YzARGfpvQiR
/u1O6YOJJ6tN8E2lWMkfx5SZA05JeLMVA+6Gsai1SX2psfmip/LizA7oIQkIoysA
2wHLCV9AxOL+C8G/O3Hb188JVAwSx8iIMps3c9wyNbDPClAs5rNArJUXdOu758Eh
/AdwwtOZlS5S/Pzwg85v1mqbsFVnxqn2BNRYgEnLMbrrVJxvu+CAzj3Ns2suAtva
vz5HJfkmsQPIKqMsJ4nZZp5LV4nJj2TlXcfyOiFSNziXnbzXT++q9PELQLjw8pmO
57y6ET5ltj4R/HeZiliZoeVQi2ptSHbHS4rm2gSo3WQPNdqnKMvLuhTPrNHNCWJ1
ZI2aky+Ol1lK/UwWCzJd1gbcwUxny2DYVYH9ZmvzKWG12XYynA1b5MWU9g2OELZa
2vuBwnQL7OzYFzGA6p6qAls4pJ6B5vfX6iqe/pioxTN23/40C3AB0XVDiDBmOMmx
pdrimOdDOgF6HSxqBP1X+zLvRqtsdujKrjZQopwjVdKcaTN/yLA+DMzym7PThzp1
tfVftlpeT6rBWTdtiWlkmnhAJpuUN+fYzoSOT9603ag7+xCY4W9cfIs4jZ8TYLj4
KheAx6alL0OOtBv57CmOr08mRUlPzAcRT71yD5LcpLhQZZLD+7s9IdtzWGzoq4Oe
UNcbMaHMZxuLgFANA2UvJ3VnOcQ8BrgTubM+fHYEuSJl004kqS9acaGwmkuvn61X
oKf5DnnGoIGEmqc5O1H7t2IGt3iFRosBum4pdt/MdWeslsCbrzLsefTCOa32ntlI
D3ITkMzKg36nRgdeM1vTI1dQwXWtk/3XXHyf1WIpLfZBTQymfIS95E5/P9izibgP
fUrKULMwnAp0JaZK9G+FSO8iglrzt0ulaYNnV77ootblpRBQ/h/eDNDaaoR2lEnW
GTAuhYP9TBdr7d59C0xBhPXdtuL+Pyn06m/JD9wgzl5aXR/KHMrAIjSI+O7kEH6H
hmWmVsTqyUkPdEFTYnDqUs2brmFuBZRD7tLklrS5v4lehDDgqgFv2iJNRELmLSp6
a3+3MUY4Yp/H+ToCzhGzD2svR90aEojT/uFgxZpZ5e1HSLXu2XKH245zszl0hT47
A29icvp0ocOJqHWxKeYIzpud7TnW/1psdOYyVXyvgXwU/UiXMfmqKV/FmohqWe4x
+Lafd9QO7+eVde7CjTi29t3z27Z4kUUY1k8KuwwXYc42Gh3AbYSHjXpVk3CdRD0Q
CFxiWx4qwlUVC/42DRQJqJ5HWJxon7HLcU5kGSCkD95ouz9JKA2qgUjKkC9eDJiZ
oYKBLfVxqrAMVD5jgQtNIF4YpmyblrTjzExSQURgQaEgu/xxcNMULoxNRImBJSLC
OR/TqthxcwspIrBsfTmeBTkRbG0+ROM89se8d+4y86IsCip2PvqgbxeIQrS3KVgu
tzphIi6IT5UdkZl1GzN5EY9I7kC5JxQNYOik2gOd2HOvDKcTc9b3zEcwlgG263uj
8PevEFwwYJ0A2FXnEkA+YQpphTpktJQYuikcxOqX7FQ+Vz8K/1TBp5eoTAKn2OJl
tPi8mm+ivrGoHKN4EIsldR1rvCDX/0geiBRRqSNWvXHC1LNesyALwNRG5IyJXEF7
k0tCuhnTduVUi4ovjPPbsbedyocmCfAxX5Jz8xf9yFOToqOuWAbHWjLikwJY0PUB
jOcTMZEhYKvDKJ5hJi999RWPD3VmQ8O54zaVi+J98F+UXMM8jUwkgFj3vzOYQ4gy
q1q/AbA+iOLdm22i/3sz5vMAgrtOYR6T8YtjVKNbWaRWkWpVBNGIzrZLI3QrZ3k1
/f6BFgw6c8w25zcJivt21pO+h+5Yy5pZidyUXZp0NNPUXs5epHjT/YPyDaTs67zM
yEODjNO2zW1IMkwzRiruPpXOLtVdVG+WDcwCSsuOoU1zJLXxXgv1OHJy4ynOYhes
2DqHNWL3GmI1wPZRNhgN6eeZD0xiR7AOPbAWxDaEiCjl9pMidIb7bcOZt5m1gCXt
ukbobTQ6H2t8dnyeLU36NjblR5o2zDoPClg5/EJNwlpXmm1si6aEQpA6RvvkPIQw
talJL+457R6c81bhtzGd+F+OsTO/1TK7bG2PBYnjTaDnYu+Ayg1vAs8L+QLtny/Q
ibiNPmFxL5m0/hqj6rym6ZknvEL79fBnhcucFDEFgvvsWRVVYxywtTnJ/uE7jh2D
NfAWAkHUKr9wcEqnzxSpfudox36symHBueYEjR5OCQz0NLr1r9VLRLtY8yomwKmU
dcNPjf7gsRVyW7VrDnoUBdoBWrD6Mr5AaCmMq8hxKixXXLcUTWb5OuVgdmEC+C8t
/nKPpPx17NJcdKZdHRlSJQmd+KwD3JyTEGh3wy7Pf5os+rl+1JOPDpZufchtlq2h
PdSkYFAiJ60SRfDHUlSMdl7l25z3yNWWk2LnjzoPeCGm3jtZ6Kd5Lcrd7K1cpAwE
TDNiZ585tiOvYfLPPMlgDIHB/b5nztqdiYsrswfnfBuVIoUI1Z7ctUGfyRPqr2tc
uvUGNaU5hkmun6524z1Ew/mE5WcaA8yTXKtIjODFN4Kt1IRtspLgkpwp1VqOYpRo
eA+qM/lGLacA6kJuD0dLEplzO9BOjhn/C7iBtzBD+BiTxjnrpSXiA6QLtI3vQf+D
C1xrTG3wfLUasvrMfK8RZv9QCYTVjlc6FkVa6Fi6DmbTJ168bkuLkHqSQx/2XwBI
FdTb97nZCSKLPAKnD5pHQCwlH06W3b0dhel9PcVBDg3gLL6NS/TpIccbqLHLfzyd
Tq5UqWe+KWXdWODyaWey4ZyxG1KfeMo7OB1ZKm8MAYACijbMbT1fosObBpB9Y++m
3WgmL5Ht5n8NEUkH2DCJqw6zKijwzB1YwBoT7F13i93W6hKwT6s+DRPbmP7FQFVc
FUhCvFj2eTThl9MsQ1wHl73QF0RCdXtpoNxdWABmSA6qe6006jj86f8dDDfgT2AR
Tq4pwlAnmQ0WqvIB1DW5xwDYrpfr8/+uyGcpOHvepciJwwYwAdrke6MSlUNz3IR3
wvPIQ1S8O2kH5C5m/iiiC3gOhdTu/ObNd0cCazyyPH+9mFNmTaV9HhZRVhGSe7b7
6Pl9r7dMZ6jvImqrfP7XB6PM5Dl1fqFAxvk42Hwc35qQoRqY/kYwYiPBJuua96yq
XPG66PzexQXNLvHL9IwF+gO53E02cDqVZ3POnAd/5rwNuMZXo87ChAaFfe7MRajB
Y7Q1h/7e9gIOzs3bmrH4D/psA6Kdj1oUnXLVsDP3l3B92M/9WOHvk6DIu1zfTkrg
ky6UKtEiDO4CHaxESHYYDhATbB3hHtwRw01WXsyphfnj9lZ/vvNmvFhE5TzylDk5
PjVrIdDiPTUXS7L5OCFlO48HHonfz0fYzZSb9NIHN0SsrVxL8Of2DwD0k8bWc6wy
88DoxioT/p9qDe1QOF0Tt6kBkBfaJ9fUMejmnW66WRmCEgEE2UKTYo8fLHI4PziU
QGkozpeskJ8AytUSFD1BaVO07ekWEQLN+PjZUsjl2aKQNfOCH9hLJO46H72lZpmY
JBAi7djY02ueWxeFQv1s7xBk3afjwS4wIrWuWzccr/qXfxtDjGNsR1+yXylCBIvC
ktxlIovzKFsHbDOL+XoDiFmEqyQkglnQyvQpMYFhxpeRnHsjpHXKo5Vx/msjwwGr
Nknl0qdPM658dPe75xv5MCTIDgIqpabHpPWGDDd1S1IvC5/ceBY8qv1j8tys5GZ7
GYmV5SvrKIdhtCk+jpScJd3Ve/DcHsfLcVla9cQVhXk0Q2kNXjSH9qpBe6t55+lO
TVGEcWANIdfTZbHPguCOUGDbjuMOpkysu71bu38dPNJOFMjOrVZzS5fs02S9so+4
qYQhzxZ0lT33tx/m10ZAfNp2zotRx0+nSq8lMw9FJ6GuMJURAiJxmX5IypUxoCvG
QA/KuaenL3DuPNQ662oGTrKCoGmYsxfRFmCtoaO24qR9E2vzUj1iPwxej5PZCout
4c7Qyp8fEpfFM3sVRFgszAksf2hGR8VbO3HF2Bm1gD2eOfTj668BTcRHK6hsAKwm
i647k90CRTLNVYltsysHkseiHzQ/HInlcFgydFnfilkkEzDecSVWjSPlqLS3T4yM
v3aqNDLn7OFVysHb7qVfxDfxqydaPHtHw69gS73kf3Ja9tWHPXsrBlWmKkr7GfFh
Vhs3OMl0gThBH/6uQW2tWQQTkbnfbBpqiVTl9qAImxHhbeJEHLUtZLwyWJrQJzN8
ldAPlwuMQ0NdHmq8jQ2+fbXW8lOF2xOlL+gxb6wMkv92pzVz7UdbkEb1TuPfaZ/9
AS/fEctXvZ7jsPY9+fQfV/z3jTlXJ1pPCPWWHZr29qWso/H5LSukM1rUJA9pW/h+
1VObeyXaGinFNcWp/HVHWPgixWzm6U8P8bLk8Sw+adTffABpLwD7yEm+uUX4bDsY
jgiP4+iPqcRtBero7at75VWLJniKOulFYO18JKcwf9eYPoKvOSUupWOVXiN/FCCO
0BT/t7lXPE378T9twxR6BMB5YGc53OmgR0jD4ayTCAk2LL7W4gr34z5OL90bM9ak
Z6sxoKC1ZgyQljcWNLEo/Psf/Cd/kamnK9HFRHflKzp0GpaR5hmRHidItA1WQvNF
xfoPZdD/5tOtq2uBrwmFe1RHZ0mmC4EAtgXRxbyVYwZrR3kUnScQSn47M+0flpME
IITVZW4ZuogoMSL/kZcpKY8KmYN3gWBz3Rr/5q9HZMCOxHklq7zgjbdHPdyyFvYa
J57vCb5HUiKXkMtE4dvwUmYh28F8R2twGPXW5SfJ7ACPG9hBHWR/oTqDGBXKOOA7
5QknU2LVOeDBAHV97RMfr5UnyQAlojx65s8sRsnlNfAPEA0316iCpkwJt+EaxhLD
u38iewyfvjcshsJw/iqIKTWrUtIwGbtp/PA/IO3UpFZoZPSGzJSUDksTLGmgAmLR
EH3x84ry6A1u6RpjvjBJQOY3LFubKZS5BsZ012jqKnZrpX/P1oJLm7hNW0/bVe4k
leL0CryiYqWTcHbWa8U5GG0heeYXOYI0YbghVtWUtX1uPnRCSiPJef/wY4FlNWTw
lAJJzyIZ1Eyeb5pGQ8BssuKNpAlmIdk78MNU0SL7+MzGmuyFzhfGBhdi4cxRNU2B
7qQ5xrCsVjij9GA3TeWZFYX2rrNpb5rfqjP7XZUbEWRYaP68K33X3W2IUANa6HPz
p3V4AzSI6aaG2sWhPV24r/7XLQQuZK27jqTb+L0TeDPLiCpub2RlYhe77VEtcTsc
kO1i3dn8sat1jaU/WEDe3hLCzvbsGSJs0zZvI7R7Ck3A4qVIzWN6EkKq+7zzaDQt
t/eyAVq8UR7MeL+86n/OkXD2THQfIwpHVZavVCBUhJlaDXqFdA1Eb9Hbp6laeHRu
cyzzkgWDzPJsHekz87h4eCWbF00LX9UIcdqaBEK3ThrJCtzP+AhsE7HssNCfIybs
TvYknEF3+Syn8dbs/7zzqnzjoPO6buabcEMFqkDPpVTOkD0r5BOzDsURm3zciYfg
C8t4/HVsV2/OBdBTd5GCe3k7Ndq+jdEDMD9xgFLJZJ6LwsEoNpkBadr6JpBvfpiH
7xRxggzcl1DeepMm1MxjWuvzsvwIk3vyAHn/NNPEMbweZ4LdUa5Ho8Jm4BOFIwbI
URoXFwQygHiZfXQZryryeodnYRoyITagFjIAf63K3uM0AlpCevyvbg9qwF2KoW4d
Gzo+HDLM5s52wp8t4Ist0OCdSbPAuqpRO+PrOh6Ib384tqeGlD7fTcMbAw+dcJBp
EJilw+dpG411wMrC72Yl+O0r4B+lst+FLarP5GONM33m3EysQW747OWBZFc6owEL
dzys4UmAU3ib8Z+HlyHMlt+l/weCaxqrki94kRoEOLUUmbOTI0KuDfngAdfg/xIN
OhgpvWBviTgd52e/SR63Z9Vg7YGUxWf2ldqXlxQjAdws49LpzEtnRcmew+39H0pp
WWQ9RGYTW7D3ayMUnfVZ15qDEA1tWv8/+gA2sLMblrwSrQhc4Drz4XSveLEnLQg5
RfOrI6FuTg4N7jYO7FZLrJ5iiSDjEPrjYVtx/Jbj0WYWEegk2YmGZ/+hxDsoOeRC
4H/U1zUz9DL5krY/4CRldDi584OA+l8mmH/57igj0jd7ZDCxQ3AxSIxL0JfWKBTR
mgCj1c7Kwp3Zwsw6yWQ34aLaLRRPZy+9qV48mYWCHUwIP0fIbg3yUDNHYD1yvHXv
CBy68l33d6MCGxgB5Ey8xrzQ3LUEvoLfQrUD1+fAPMTIEvBI1fYOE0c2PVTRJV5N
de1ToxOv0YBCB+ZsKVhFOVw31AYunRsbNYfHTxIa/c+u5STzLnmPMMHnH6RouxGi
n5qPzLGQF+xW2F8oZqFagGRulZlCql8YSQog1pT+/3SdPhC2sx+Xj34dGptMBGRJ
zocqFRMgieLtd8nCJii4LDIhhzfpn2xpy3ywU5XPIv7Nyw1QfK3uMEnMUCj8C5EF
KiQ+DY0iEFClB+Bu3o+D6sDHr0588XBA/61cdlU2jKwS/XW5akywDcM5STIitZs/
tWR1qFKc/BcFMScPeXT+Cx78TOQ8s4neNSLo1jpsvg6w/4TXFHCuFCTbfGPgGMXF
YfAwRqC/3zJyyeviKckwzFFnMhaaSSxgVS2v35vitxwrb8mVu3kxTE9Cnet6Spda
qF/OVz/FvwZMAQOdEJucv399sy71moWxP7b6hQVhnjdFnURAy0TL33WggHai/su0
PsXLSjgKYcqWtvtUFHJEW8+l3ChyhbqrAeWiJKdGIKD43+7DZCOdd2he/8ZA46zz
WzHSxXvEA67o0GdZTBHNweiXS+vz0gYdoYVWQEIi/BrEbCSxQfd7D733EUOdFTO6
fvFaD95f36Y//0MZ70sykoLH9m4Z3IgW2Gh2D5lceaqWyBvoQYij/Ba9vezF80h1
+z7BOEyQeXCdrPY+27wEhq8uXSz1ycUrxeBeIkgxPQ8a7AyVMvnf0FEy1EjFkaK2
7VLZxXTBB1V1CUHoZ1oUw7xiOH9m5E7bhV07eY0aY0fyhghAArMro3g+RDF0/PTy
yWtSzLcZWrZftqZXOngrP3ySmGqbm1FWadxivhFNHAQgC4zyXxlqZLOSNb/cNAGZ
uafDNbaOWfqisDBDkIhlDmru7Ls4hi0iGToaapKORbUQ0qKIbzKmDn1hEKk5IVGV
PBKTFJl9Au18y9YxhaRudETUKAvqKWHXpJvVnJz/GoUy4n5MTP5kDUdgzKoYvTJF
/7NXOBFABlSxv7RYISYwPP6dW3ejRZuo/8oexHkJnb9sNPqWkcQCC54Sg5ZaxZXN
zrIj9PnVinVxmiXthEeXk5z7mLAYOgmBZAPf03Te8S7ETowsfZDMGyfFx6QzDJS7
fPDuJDnTcZwbOfwgTq77kdN3tJRH6isfNcH5tG1L/dnZ52yfYDsg+dETWP8qViqP
S+UuTMHEeeVuDqxb39KwOFWkD6rjlz6Eh6vz9Y4+0YCTtQgQ2JqZp2y1zNkp9q+A
`pragma protect end_protected
