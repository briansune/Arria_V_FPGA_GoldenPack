// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
orGx6E4QPgQXgrwoY/IYitEH8O8XZlsCZ8sea8kaxVzlw83fbLY25PjJTzTwkuel
JybjaIP1Jjc+WSUHqNTMNn0d9jF6V9gN48wrXluRqUDMj95QyEajvFw3gOkTxn5h
TRSwsECPvqtqubI4s/wCgub24EP5ZCPRZBJ/Gs/lEo8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32784)
xziobqLEeJwWcImRkX61FsWfg2r1KggN4K7sp846y6xoHbZQzvNUsewoM33yKrfI
PGwP2iHKcus6ThyI5qiIBSl1gE6QemPdBLlImLvpyh2eIHq1wqCkWOrolRdVFRAO
2Kc7fp6EcBam1akL4rfx6+Fhvg0CZ0pFvbstqeydXzWm2Tep69Krj2aRYegOfBzU
PhODWi70KR5x3gkVCyVl8eWc4N2P1TTRW8MSn+0RX6YCQnMwslMDYwR5i9qfw/WS
BRwIN4+qJ1PwBb5XgkXKg9A6RTM9ehkFS28Gqban0v7YFAFelGGqsVafQKXf1tv3
ncEqclwW48vjTDc1VS5ZxoQP4xLjzPwruBmMQIKXwqpBwryQ0OA7Bc4lr4aoWkaH
Sa65Zl3LuFXXzNbYuGohmpssO+F5Va/5iqWBvRjZ7QL5wFe/PtIt/NoD+Kl0sdjR
qoZi5hBlMczQeLx/JlH0wgn1r8CbxkjANMmjBhJPyP+liUIa9M9A7cyqX3ZeZkGf
slShioePxYd2STygYTAG7QSuhrLGK43aV2CUHWggfvw8ciFaQf/WD/gmFxvt3uF/
95ooPSazWQvZINK0gGM8y54F3pf/m2a6LYACUiIVJGb1hXbUZdT2eRHh1GnUzWoG
6xgrM1TxjvXZaoxyhEB3vycLAU+0M5fOoAUb6b70Vc1pzhN0WCbpg7iV3RKNE/j+
T/kgbGYFT0W+EJW87o9cYPDo4znifqlkr+rR2+5lqTtDnNBBLM+nFJonW4aaMHfC
vXbJFeF/Wq9UrBLjOcT/GOciqw+rgNn6oXEmuQjtsjBlH5DNJ7dZuZq0I7nicKDZ
N0ny3sftu1WX/+8URdB2QtJsP874kRIU0bmwLBBsEWICZ4Lzwt7/EDCduWi+8O8R
nV/zy0Nzl/WLke0Sp2gLt+zOEkSJC6bwg41kc7oc/+ifeAWCs0Wgc0QaG5JQo1aT
B8KUJrSlwYrsV6skiiIELhU8jRZQHF9rW1gymxN8HpfP823ytTW1W4qwtBuK62Uc
1NE2zdppVPM1upCKX3/ibekkOjEfBrzah0aB/A3Xo+DbB/mAkTrnFfs416JSa7yN
MaibXuNL4SxtnWB6PhUWOMz/FwRJMZUucm+7C5nrlWDDveHP4m6pW0Jpvm/XdkCt
OrB841e/MtJu7T5J+b/8sVdgrUNvd0r5yrq5FsDp7Ce/woKgLO07l3vY9PkrAIfe
KGjwu8mhqqLiwrz48P4q8+C53UuzciEz5WoBO8E7Ye4nT6pzDwOqty23zOj4c4Bg
N0n0cLQr8fJRJqkl4K+k3tI9IuQ/RayGtCFG5tTlHbxut0I16Gp2Fp4jQQoIOEKK
O2uslmitSCgX3xdJYozs2CJnbdcBgJ/2BxZR5F5VyOva9BNvA2zQmA39Hc2l9bqS
mCbQh0Lc1oH/Z9nBP+qObE8A5LncWE1oMjms1/DIZEx4W/KDBCkGlabmqk/32n5k
A3+4GVmTMhZnkMhuYTHgUxncp6WFMOxNZqvTDdNF/y5x041TLANglSLiMLHpt6DT
21VurJg5T9+tL1ea5xqBHwa+SuCARbua2ezbo6PBSjyEMYlOK0Ha170hUhmRjCDv
dAagIVcuJBhCjUvvlTZYu8yOtbc4hXge3lNr3aJWAdQfynkNtilQiWbyDjmioVjC
2qWMLN81wkENW8wP6t0D1oXfan+LF1DjErQjn+vhfh4pO6Bl9m3IjSeK9Tnm1E0x
JDMXi75ef0Aez9q+/rmEjggErEOqI0CKamfJmtyNJVGuQFZPU1Pv1INjgJmwOHSR
zWd1IWGDzaqum8V5RFvOSC/k+ol6+0yoK/KusBqxBsraFCW3LeP2QUclKQG9habt
0HMQbJcEJxf09Rqo2+wASMK04jCjtLAtMu2VeOdz1pSzC8ColrDHxOLgQKzXKAPj
n1Z78C0e6li3rBkhQAJjkrVG5hJhVPCbUzgMBHnczWg75pG8Y0I7/9IytHlhFdqx
0OGQj34DdWzP4kizbUMZItPIJw1sPw+AbNctAStY9fUZjKfyUBAPDdzqrWAndf3g
rPdkdNRisUgWoLFJXu+Zcz2mI72Jh3xkN4XOdL6Cp7AM1cT3nQdfpmCuRZvttzgk
eqIBiwWyq2ESDz4THGwul5ZleSJvu5X1gWJ6fnoE2IO9YrOsAeszK6IxffLJzVKS
Md86wSXZKTD22JkNAjB+8rocD9FVXa/+OQdU7cruq2ygbbjL5YqttRwF7r4gUis3
kTYbcNZonlN/xDS5UFI/e52+9Xd/XItCQQu+C49g8pCSOdm+fuCS1hm2dyIWiAzl
Zg4WMQymclUTYf0xJkhBV0iaHQ2a+RFpBgsjUh8tQgVjnhPntgu+n0ayHGgsehiY
R/pTFQM2kSCzY3F+XVpqE/02bxK8pYXTmQDGjXEHslCZCyyH8LB8hX76XPrtGgw9
JYAzEpqDPtMHMRkWZzFKRH1L9qRq59MY3j5rPQDyc4uBnjOJS09fY/V/DTvkihmI
QMpsFo51hR62MFYz50pNs1iZKtknMry1yft+w5PPY/ln6LYoVC6GmKpZGB6M9HhZ
YJozMXdLtUCBNlNkGuiamy5K/seUKdBdHDYRjhJVhDL1e8sWFx/ly6VxyGFOJFgU
w5VkLI94OZvg3KtcERYYUvnqE6J/SEAHOxnjAZ1i4LoWVWooITO7PVNcvQ+NMsnw
V0PyC0A25ttZ2gK/TaCMK9Prcdik7a1fMK64rMWCN3/peKiZQt1HMLLAxFT3Eg3E
9BAFcr5K4mOghZwMdweN/YHnNOe5GXYoyFbgSDnaFXQYidruDuXxs5xXwiex33sB
r6fjLtXDs9NQ4PKBgkeSU0j5/4qyCtXrrEBtJaoQWoTFmf4wymw2lu4B7ImAPorY
5nrSoOcc2WumTNABD6h0017fus8/19xKcuUCdr4KZF8QRif4kss/L+ESrFJI0wPr
V1Ly3WnRbjG55APl5eOb8c++GlDZInLLkUSyFBhwsZYx08DQIrqI6N/vlMa3cl9C
I0JYGSN54IH6ZBGOZsfFXOio3zno6ArEulhqK8NuEBXSl5JE+/ef33+f/m2pbsmE
qsMl6eMC9xRWlo5s9p2iydlGFQ3/6ESWVTnNvoamuSmoSlLUBqJuozDNay93u/J1
FcZja+AgGKSlGTkQDmvg/RT0zll1v/wc2WdwvP45ud6zHCmTbwNh9DrRpVmHwxsQ
NmOumaH7S1Ma5Pj7ZdG7U2X0l9uFDnPvxxqu89nKf8IiUhsEPqChKFfvtl+luSZ1
T7HWK8Y+CxQxfccaHsnDaThJGEBt9QkZNFrS9YzjnhgkJWhL3hmsnzitG8PZPvZr
22dXTX/nkHGs6BakfY92WX+cXjTxLUVKP6VxJQ1ZJBtetXxxiQc6JUSW/90wwZ3z
KOp0HV9vfGSG+sQ3qphgx23khYOQg09ji+P/CrZ0Rg5Vu4YbML6raKZczdhdhBeZ
kBAkceb7MmY5jMLqM9uJ+wyHtC+U2awVyaGi53l7zU0FuNS2E+HwX+++lEfEH7g3
I/dbowUvqcd4eFaqqo8okKEFKY9f1xxNmslFKA6zTSgkRtmHcilXVmPCa5SDR9W2
aCOZuPDxTHaG5TIgTCpVLfBN4IG4SVli0LMkw5IvgMSFt9PlENu/JedZ8u27E7tP
y4SD79BeBYT28bUY8ddbTxrXdxpPfnusJQ4X4XGjBaIM6z8U7seVn6j6BfMEtj34
2Gg24whnpFX6rQivtTSBbmO2oLibHAfms1j0qTrJ6/pUaEkkTITkVOtZApQpnR+q
fq8I3CmZSQRHiYG1GK7s4zSWHiwOg57WNlgmPy+aSDKON0pLInu4riE/z80C3PsB
qhZQZQnntL3QdwiCGHlAQCmndHj+u4HnD9pebSHtWcjpVwpWmhrRIVs9IwCbB5rZ
P1mT596PCIIkSnEEh94cOOhlZSTbYJCazKmqqznrDZ55A5USc4HzpFPj8DAA9RyO
LzJBMK6XYy8lflEFqfgAlUfqtZ0BQ/RYz+0/4LTH1IngPYlWEHSKtcSbFuNK7V8T
tGo12cjd1PjlGpEaD/finrvRcsIrQko1TNYhOEGP7ZqsQNiGIIVxXHFzfTMIYHVq
0Id+c+MiEW23VmZuDpg3CUjKJ2QaKtlaXefBSZYOZi40a2JYtbqkJ3uAFb4Qejna
h7lU77+LcFCQctXDzAJIWn6VYLs4tfOR2DMlo2Za+AzxbrV8fVgCiTl+GP+PE0n2
fXQR457U2mQ0COzKrNkDH82rqzpCAb9vYjniezs+af2LZ7JOHIBlY9XLvfuFtdWi
aKtlZbHcvLl+KxVXjUVrcPUslfuTr3nWMY2x9IURG4Y4izqve1e+QijQIzaWyq0l
ZCY1gmLcXf9TRdVI0Ymuslj4qjjwWfQfYndPn6JZqYI1deFvGUoDkexRF+c1SPOA
H85qDrHaXsJBVpNWMZu5vaCp+Eq6yJg/oLk5uXStJCQrl6g3J4P2RyXAWG8FqqJj
4ab0G9guG22FlrnyA8ZYJn4vqWw2fxgwyN3yioPoixMdq1/AiZDXsl+0/Fc78XiX
IzYcmFd5UulEKfxPWf5GS6/rxOyueKqZ19Km4mxjkPqkPSCoXXpdUaYHbukV7mYm
aMnoMzQA4W7mMkxYILEkOoAN1KqYSAVsDDX8GkYG+EUKwCYGE8dhvWgxmPhYlyMy
VfeW1e4fJENws9dTbGsUKsaLnyvke02v29puM+t1g1BZsSx0ejY+D/uCpJ6l9Tgt
oL0jlSrEaQUErnVFtaN8ynrM3YYGITE+lsvnzJM7OHez6T+INSY16Y3VjP5nGUx4
aHfhdqB7fQ7f95JUfGLWGYeIilaqpWWhdX9DpqDgFK8uHzw4/r8yO5PunmwoUA6F
8BjOk3agkhl0dBGuD4LO3I1oVfB+rVqB2Xa5jCuECo7EAQw867LcfpYGOX7zyEwF
ER2WIewBi7LuV1K/4cR/afjX0X0mouPB27qsYMiXTe0HaabMplEWpQh2Ej0eRF0+
xmLOM/Lp2RcXUjcsdrOvHpaSokw49YX290lAurl2kQItY6x//fFrCUO4AZ0nXtDE
6CCNogIMhz1ojA3B6CZupkuPM9lKD+sGQcyvCzyim7iNi72A+4hYlm6ufd0cK+fr
BqcvqEaELQ4MIx1x/WyeKUGyRo+O5oYHM3jW/E5GG1D00zUgpoAHA3PHOJ+XmNqG
aqST1PzkK552d9ZUF+K0HcC25uaCdHyzGpvxzjwYt0EHlgktIb8mzLi5WlhpAGDs
bdVQFdPP0q51GRaWTxLz/J0XT4xQ0hCoyzuYoIG99UJ7BuGaplLfALAPbSsrZ1j2
MuaolwWrkII0rSsSShibhmyr1YGAbyRsMlyKwi8CfbouGyS8vs2QG/XzvfE0hH+2
qJ+j0LhwCCHMZGHWUX0d78MtEuLzr2h4qYA7fAYujhaCU73GhV6yiJuT2qrSedXe
os5w817yFE4c8gT+/D6ULvpddqXV+jrdG8I5pghGNsGTcD970QWq/U2mT8bZ05wb
22+Q+gdW9PcrBhAYnZCTyZxINjNn0etdQ1Gj9uO+pJnLGHe3jMYi6a+Pj+S8sx0n
x0Wv302mxJHHb5qwGSiGsRNiwWqR/kGAPUYxzkhp5iNk/9zaDTJwkF2TJsovhor0
8pNYfMX10jrthAdeno1wGoQh2HSGiUnHy1uA4K8XlqX7n2TqTlCU2Rhaavl6OMdJ
fpR+CtqAiJXlBtzDipEZZ4IbUxcD6vNW8MdkPXqTgkjoGH/CxhWEmVCQLYtn71L6
qqTLH/pAny5oGjr0RX6cLkHpdbPfKNdZGw7zu0Uq5sduGwbqFsFxCNWnl3lrbNkf
LO+oifXzjvdPQQKRfdj5LsXAmalxcluYGoZ+cF0DdOcuSk6QtLqj4Jf21aoDOm+e
z6UYAPg6SY29/eiwtA37uZz8WmzYcZeWJ757i3tHowFrn8qf4yaZAdXKJ+ny0cd1
3uTuT9GHtprmPxEGgEa0nTT1Q3ukyIGapzDzGa6IfrW12BjUU7dk/GlhvaFSsCbT
7XEeDMIOIJyeEh2MGOkU41/UJ2TyHuJb8aQ1fv3O/e5VGnDG+X5YB1+Ir2B9MmUF
PV8uVD0j/tWvqQ/R29PIetfbJRove6NM1b01DS7gfMUnudu+/+RptYhF2Cjl4Atj
yx+cnYLaaF7vdvfBah3IxCM4eq87uHIV5leYrieW3jPIRIUObLsT1yLh+zMdWyc5
M8DyToOI6oXqTPWomqYwc5IPKgup7JwIzeODVJWgDDqV3STSTJorIZGUHU0P20zn
eHCSuU+XyrjvPLRMtko+jUq5oEqusMs8IgD2L48Q529EOFniEGByG9xq9CEmK6Y9
ZPoAFeV//M9nT3wJG9FNZApA0Dm35kIfxGPnrMpuWQ09mJw3fvoEO3A03Yy0CnO4
DCeem50J1van9X4jEZ7r8DPVca9LX9BLABrSwRtkzGk/nqp6mXxXP1Qpi0p1kEdo
vcb6uB2MOmkPu7mM0ffo2OiLzqJ/K/69Z9Yg4Kagqwz+LvYjPbqXoWkEpabPnLSw
9QjSkrr9I/Hyx0b67DCIEAJOyExjAUYv6/DMVxF1oDzQy6nQc41T8CLdyGVakndM
2PZDcNL3tqk+EwYfXN8z9kgVUh0cj8m5Dm/qGK30+gYFCfXEI1uBjNQFRtWh//PZ
K6NLKrWRAVJI6t5Cao00bK0iT01wQs/IfptJLddxQuRqsyWdYniHel3k6xF5qw9T
W2ILWHlWJluam07tsnxVTkRWOE8ft0QUNkDRoEXAU3umhxS2x3Gf8vZGh6XIktO4
4I5wsB/J4RsFO9jN9BV3NNcao10A1m9XHB8cKbWqFdufFFyGosM1QcHG4/SzEgni
qQn0vuN2Mx+N4Nwy6KvbiDznOxbrSKegYvxnt1zht4dI8bjnDIlJFGtgA7/fqvLS
1c0zmubG0Gn2s3774TXajpzCuS8njvxGmBlcBAoHeldpsiXVl5vu+aRQf2HZmbRN
DTthZ/6nEQo7D6oxC9S0TQ2lCvXPX1VUzrQPSaaVQnagNWmO3dR/QmXTp9Vh+64e
/PX0UT6Aawi5deKqQP/YFftoiOvh1/yuhuKmbdhLrJ4B1TnSPqQjkOZU/9uJOPWP
cPGNxSxfTHdxyUTW8ZTdnq9eJiIwqoerXErugZVUCRfi0KjZxS+1PbHzs7jvW7bw
lV2pDa5Tlnvb5xk6hHMMC6C8v/ANqWmW4beD/kIhY841SsSi4p2ZS3eNoZuvNQl+
WsVnfdRovxvm6jruDSvVvFodskKLlXqaGfieN6yhSphbMvc6ejIfqyDjYbCpvOFA
uxa63Kpmlgc3LScZu6SQtWZBXX6d690bPSkwA+cgVGl5hk/wO+5hPpa8rV+8LSPb
bGzXdYzCLYIw2d+fyshP5lEbmlXauZepTeRM/8ku2l99LOrWIz+ZIo7rRKCt11uH
kmF4zVVRygfnL7/0VHWicQ00UQKI8o84S+80xEkeUsRWJNWW90XKtFleJbER9f43
gln34a1xdJaalwPIBPN1t+T7SedjR+N+LkD/SGbCBY2Gsv5FreN+jjS31f8vREMM
MFsxoDQqScaD2hJaTfb+me2xul3KmkZpkvizDfyQR7xnTpZiVQZAwskXPkB78Ms1
Ihfinp8teWJZHHGaETvW9usGbuT2KLIcoFw7NoJypeq4uqrOrFkhinwaEM9XG0PJ
CYYXACXF3FVXMOAzJ68LBTaXdHRKmwhPMqsPTo0ROl2/9+cXoCbEtnlxD/zGfxzV
oyc9VWHXjxEGq9BWZugZNmgpqpIJHc6q/ZUIm04J+m3a3H5H9ceJU1diyxs2Bd9P
bm+uXoPXHJ1B6RS7jzQJIIrQW6zA2sM1oBhoKRwL7eXGnhJTSUClBEOfvoYARLft
Dz4RKpjPBxRc8VeYp7bDKsU7KQn1m4zvkO7GGYpUFZ4x7DXuEPRSUoKmeEyHqVd3
6yv+v3nJ9Ub5k7PtCAnL+kcnXSX7NrciypEoeR+s0JCfGOdpLU+vQ98iMLb6xtVz
0IRHI0b+nGd77RcnU4+ksqDo7SLO1IJxPJ+3r2yXU3wNpGkvGIfC7MiZN12lvERk
f1d84ZSRsuRh+Ufsn+Dyojq424ZDfnkb+SvGgvlt3hl0K67ErEdPuInj9DAebWek
/ddaRqwgN+aE/Jozr2NsgK+lf0NBzq3WB99VIahfYv65XmLFNo+p/G87DenE6DGz
+W2z4Ovr8t904BrITahP4OyDQ+8U8Ty1OyBwYzWd7354hUB1m9qbfub4td7V2Dsv
k9tIbHRUy2C75epvGitaKbchZpwAow48fgHAYQ0OkRJfBuuUnoxp8mYDzbcvLpEz
UoMl879QgBS1gDZLebB06w9fVj5wP0tASFxGtCTp9GPFp09knEmCVl1IDhtCooNi
aUXpkNNwXB2eeHFZlss04020haOCniDNTdNmF7LFSRWlj8wurQTjlqdi10XJQPtU
uxyBZAOrQD/blQwwUY37AdGCBMzMLVune8A1DhfFKqe34qK8TIdfPWqCZRkHKcUw
PNLU36GhzlJeezH8WMo61k3WhhhKhnl43yc/li0nJCzuULwvEyPdcAoYYd0YHhrO
SLI0XDAqFXmHgPKhmL2fUsntdvsgOaqzLkz5bBbekkE23YFM2nbYbiOno1cgR8gE
SJPl8OsSSeXjvOvPUNw4uf+3CPHJ2olmZMLobLSq3H1Rv0P4BalD523hVLpQDobX
6H6IwfgqP/by86D86es9bPkmua07vsMbjEn+A+sMwVf2Ob52OySHNTdb8QYsl9Xy
nBbKmaPc73rTpN+kiJxVjmJrBSnqhb8BUJe1qbslDZ/QBDhHMHb1w9U1TyGyuMm8
3Q5LRJpjlw22oDQItgtYfKvkLQJ6aw9TQwRtB49KWyR4FxDpEZCxxIEWKt42FRUJ
uvPNS1DQJAYD0urAXCEv1MTzlV7H9N2A+AQPDJgRomYekdphiyhJMw4F9lZtWc4p
GgTpFs1+cUU/dH7/DgA/97xJ8YK1B22SgrD2QGGZZy2yGeOqTn4dtB4pz+ZUxI4+
FWdg/2uN2/0z43kOzv+k5A/8Tv+3yjTZpt01rvJKV8g3AQUoXWAngrr1EsCR2iss
ZoT1fLFBL2GzjnLMqZoty+cRLqJzALK+4SvpK+aB2uioOaoh5Sb9N193MJMg+brP
DWYl3cvyl12C0kYDEpHJGVi9ZCnLdWVsDTvU8RjyXPhiy0iVSAdtZtyI6wXJSxKx
fMd75orbvd2rpWSprjRK4ZXTImWccDzKmpZLXgIynEDhfQt/n/7e9Uj7kWHF9uUm
mhjdH1EKATvSOJkPl1dMSc0/9uF+MoRsYSn3r1hi+YQnlsBgPVNI+y3ZuO3B9OXv
QjbceQxdE16DWckQaN0cSTRxHWlf+Ta5hI6+n4QXbaHq0XTq2ku4zIpZDrBpkttj
tcVbseo4cWVtbW5BIngkv1tgk4YxKjogeJqKqm+jWPF/pyHlffYXCGeCZKXNAuUV
hi4CcRbZvUmRX/SKxJT1UYOJD9zbi+WiHLj4IuNpcZWSM/5dvvtiYdRPsOp/Cbdr
eNtmwMdAfOltEHcktT6awXfZKYYZBHQ/iJcjqrWakUBVtnG9b5NQlMexjF357wnw
y9f5/NdxlTPEpgtcMOAgm1fYTKkL7epJtNAMOR6q2QgUH5asbbaCFnpu2lHDKz79
SDfcsXzfqTWUgpi8j2AybvPxQm9eHVB0dZKOj3a8V4hdpW8GkFPblXDesnF2Kjhy
l3A3Y1rquzwHT/0QqDp7eIUbwMSxdECGzkzFEMnct2z0bSmlkcFEQHQMe3w9Nk8f
eai3yOv6RXoRjxil+ky0It8bPT80N7c8cnp5sYPnpNZj+sm6sSEJ+rfMaEphqrLO
/vp65XJFS5Ty7wKJsVRYSCuFNCQQZBNcXMYBxCuaeDTtNlWdGTY678A+QOkccP2k
dyF18B0+hnc88OmHXKXszFTHWWuQTnQGjDnJ9UWU287KOmJTszQpK3DrNYA8BVlv
q1JnvPoXne9M8QjNFEbCLqytHqgvBR5UA/jdUrX9+qWv75zTzQBY61zM2RadYoEy
bBbHVqVbk3jI0qe/RGKpj8vq2FdmxbyV9Xf68vUuPjyXulb29Iglcvi4isYUk5sG
XvlOLbcZF5KjcBJDT1DIDxO0F3XDIO0bS7GUpgZ0xX3uxvArvy9GYhgMW8d2Zvrj
OHhR6jQudCUQ178FOMowrAHpW3FMVT11DehsOYIjVH+So4X4Z97dRMinkTQWgxzL
JBaUeuSYB0V8TCfRkbd9CEU67ytuE6+7UcWloXIkPSMHjTTUysK5nSkEONqO8cTh
xEB28TM2qKMud5UL/hyXQf/Buycf3shjptCrHDSRiTP3efvshqBMWCq3uA3wQZAY
68JkAZUwnua7G3uX/MG/Gou6QJD8ngdnjtAw3gXJSIyFY9r54q4/7lrBQ10OzV3W
2IoR/eW9ErDg4Tu0X8WI/HfNdEkq9uMARp9i9vtV35iMYmxksvn5CwXEL1abO/bD
p3nZ/sLTn7UDfiO0c8GoiWeXgMGKLxjTt5FbSurhkVmt0AiVlM4poIeX+26BAnC/
2U9PQFO5B7qY9nO7HH/Zp98Vnt5poY1EAKHPjotI+pgjRos3tU8aBSmeUOa9EqpU
gNoWQFmllCudD+KQyJUG3aMfxr+0Cq7znOeAUyFLpjkCwoZShAXGM2uDoSJzmVl8
5+HzRRkXgVp0PdkQPrQMITS0DM8whzMuHjSnzvNBijoA9tHGKub1lgq3hMUvhQ7z
4+FF/DSqxVPcwGXJdaBZi/7Ur8tEiC9G3JF5SjWXf5C072QfXA8gPL0SceeBSElS
1dgWs/mv85qXuCgGeof1V2Lyxb+QhKO6cmTJYL+Tye6Uex2iK0UFCG/w29Fpt/ic
gzOHAjQCQKVM64kTKCsFVYKj3G8EfKyAMhqnxL/IJWJ2xE+obH3UzUT85YA4UyDo
SAgfCOvGLMdxGh9vkygY7IS8ZSoo1PXfj0FEX59QWg9Rk/NCdVlb1mywr68tNGAd
BZU4HTev8+AfyQ56bV/O3aSbyX868NGK6RxZ5N8I/rjRjsIbYLAbzRT4ZES4e3J4
nXkud2cMi5IrXzKMTmN1FsOeRouC4EvkEaq2mp7C08ymmMVeICM/6kp8QYw1jbgf
yf26IUI27K5OMKIK0ytFMv1XVY6Elb5FfRwT9o36K2thQy769ji+PWuAGJN4eS8f
v+JwrdVGyFNn/hYR1sZXfLTRe8ZpW0ZwyY8jTaPZfkeMuKb8VzG/92KNFHRfJYUL
ku90mNmVWAKUDjsKinv1GVFLjxIbN+DCXzjdR48iec9YpVHD3eCVwCdk4Wtc5IV4
UOg+kKd1JN5VluiDvIAWcNO4IGAqzGZI6Xdz7ZpZYGcKIEZMp1Txs5Z0aBINwkd5
1BSL4IjTNUmVNC+0szPK1JkAH/2clnEveqJtf5vE3sfxSWvPuKordYynBxs1gjYK
hWrf6TR0vBnlTi00UIWd68p9YVxavyJxSlHHxU13ZxgN0liSFTxMFXFFju7CYaMW
JIK+pf7tMacaK51PdlqHs493jtIOkUzM3PWQXyFzvWuv4juxJEc7cGnQ+EeY0pwQ
wdbJUv2ocgQpNHijviU86SAnU+iqRziW3/+rJAdo5Chvq7dWgftGs38xF6s612XH
F/KsvyKMHtv19yoI/Wxfal31P5nTberREOZg/BccHdugl6ijF53KKxIyjHxpbtNo
685QfoVM/vQj9zak+2aKPgo8bbW01W/2vRzUW/Dl0qp7CMSlLzz2v4fWsmvud+w1
3XdNraz96EA3iE9mOGFTmw0ZfN7TPxgTgnWikqi/WFuZj0++2wIE9L78gAJwzXno
j/qJTxWjh+N/tKP9D936Lw2PBbnzKhcUzTxyiIDqrkjsxf6/9we5fdbM9F+zu0kg
tKKjQfquhtGnwlkuzY+e2/Vp/9gZrzJgAckKkX89uKfvTVkH63HzeZBI/J4b0n4H
PCZqU2Oomf1PbjXbLlXbbetbAHCVHfjydDsUlAtCisUbtS/vb4g9f7MPJpT4O50v
0ZoKlSsCrv+I8TY9TQT6bAwL/RckZTNAg8/UxH1BwVI/Z4CzjouY8xPgy1f0qE18
LnbDTbdpLZqFOi/lVYl9kyUuGjmnR4uiYBcdgEHsVKRPL7wN0eEj/XVmW6Tm4ohv
rJrXLyw3321G0rtx4eaeqUBKnvOOZyO+cK+5eZVMRIY/RmkFBBScNyTQ8PNwKMFt
7ydgzp4SWR5WXZ14cVWwXmqWQXYzvUyn0nNo3cgAf+JQ+hnB+Cdx4EHpv3b6FE1t
/CTOFQX2RjDLGy2S8H4ENUD+MWGVaz9VcHBxswEfQrVVI9sR4bc1IyS23AdsrdCr
bafKxxuiGpmZnNTUk32dVuQCD3l91rrUfNqG4970ZuxzitGIqvE5l4Z/3JQJsHZP
WCg/zpUjUf5RFnmhYFHMo7SwO+MAtXwlEQ5OVMyUS1akpoKCB0uk05MomiBUC8oB
7QBq8s+A7rStiXSZP1Tp6H3N1Q4SM+uxXbvIgD9vVIk/ByyughYIMwTgswR3E/AT
PYysdNR3jntmr3Sb+kaJhSs+DxnGVgt7MdUGsQYJRrTHO2q6hXtQCSvYX3Jx8Zcr
FQL1oh1EuTuh3/NEO81Ukb8yg9NBzWLgT1xtKcBhzWwoJqcrZOLlmHtjSPn8xGuF
PTJ25gHQAicKHJ1+gBHoeV4Wt+GWcOqabBNoUrUISdf7ic6h96RmnFvqqj3cpYNe
iiKZj+0Ec/4Hlgn9xxmovqOrazY/Ka4zlKqENKORhKjGRTcSkcqRNXnmnAfssDP7
7/bWZJndPU51HO7p/WmZkSPvxJGwoA8FXAsGNKvdx/OuFVxR2TkJaBWU+vsSo6jc
VpDV7OGmcVfXANgDoP/mGnmLNbUm75gHFyy43h53EAEu55GheOPW7RPRplzFQgfW
f/s9fZyIcPTmvTRIvXfkmrNz5tIZsU3Ao0lZ8S5tZrY6e/agQAe2PFiUB742a8PW
/O2oPt8Ngf/LDIKHEZ2U6wrpMyPc4TOZ8Qx0/yTkpdJGRaB71O+cI4J/qnntoy6H
iOCxQf01xQ6ZvAehQjFGHBX2aiI4wS22t2Ed6RIl/f+PE49H83ZL4gtNcOHGtHik
KVt23Xf8QjI4vy68bfkrhuBnT0f9H8HWbLI3FXJLFH80EFulKmUyfl3ReANp6b/B
db3BbLYBmpRFjbb20TwI+UO79ObR7Sdvli7wohCCX0p+vAf1GTYDuFKHQMiLekV4
h/RT99jHGOqfnOg1CKk7RakPRt5HTrvOh7aqRY+LywBKlPQsaazgl1MDfkIpKKwi
Wmln9x0V0bz3WNW/oQeJMh2WESG/ClN8fXHGVpvYCAiB11RdUXro7VNwTVkPeakX
hg9iOVljw270X8zEp36I0zePLsRRS0SmeF29q5aOprgjFYIsinBLOm/QGddxk+7a
LCERVKyT5JyNX8chePrmwVf8t1/6MpzbU7hvwB3bpivssDO9Dsr/vKQUTFdCotW0
kGgj5GGsS+3qp2S76AIPwb0H+k8PPll9G9GLG086Hv0/EPB4IUwNQkrHOdecdeLS
5gdN769ehOkQAk7WVNsPw+6j361jO1TwBekWD4Poz2a2oSJNfTKBlZ6agKJSrhNP
DnRMIXdkZNJph/crNyedIsa8oQUtKYJgrdbR2Vx9le9iRQBIgbcOks2H0iCUHweA
nMqTTj3lfH8w+dQ2y6lmsivSEXCraBSF629h2t8U0aO+Ej9YmW5BCqXnY5zzndNL
zQysGiykLp0bLnp1UTv93HySQrhLqlDFdp2CwvdRZUBXlBM95bmdIar7zrm/kE5z
UQc1sAfZ5XX7HMJcmHty+9u+O/vEdKb5L7ugH/x9AGHulnPs/T1OTsGQGQQIlEDu
WtAmmVSsrRU2UILjSDtpeCVQfQm12AP42SMahAoDF6/y1HO2VvgP/PDy6iv1bimS
S+rLOpVmfTaIepVjgQ2UTV4HlhjiJMAnMgj6tiW3bMJ2OW2Sfp3uIxiAe5zmNPYD
tDimUQKmg8Vw6K5eTfWr20gS2vcDqOMJB1C7au6m+vRGDWROum6najXYbcEsBJlQ
3HZC/PRF48ObrRnRh+QtDWqHyxJcDny0Vlk5wcQ62OmcZUVxPxhCGC0w1db6q1BW
6QC25Q4V1TUlH2rLXnzg/CtI5ZHnBzCPr92JnulMPPSEEgOTIDdI6w7oUmDfcBuC
EHuy1qQ+KLcysnHegIk7AHFrd3LoHuZcfY32MTLR4An0KLFKyzcI/1Oeja+DvfTN
8HmZRCBMEXdcpytAYjPGQKcaicj/MOTOEMiv5FhhocKRiXLb/oDchh/dYitLP9pv
z+35svlQZfgOECP/JW5CvhLUljeRlWwBT2IxwKDvQE1t5ko548mv0nvqU3zLAcW4
oaYw2wqdNq4IEPcwI8wlK5YTVrBroK3bf6SKqdMudkFf9bPIiS8j5gvyMZ1xCAsE
MiRjUymOdU43ycc6NAo7wPocNKpHjxru7VBoKG7YsgliYAJcrh+p16Qp8nckLTGt
lH18lKGlsuwhSHtQ8xQLpc4LtSuo3TY+GiSoRWi030i+RKzTsWYJVcIQM0l16iBb
dfu07mA8SS2LBcJHNjGhYNk85HxDceyQUPgKOWPoqBpHZz2NbxU2BM01jyB6mJen
Gpy9BmGv5oBY10W7PUf0K6lk0i9+yHHICqW1eZywsneYCpi/9wj6CPbEcKSL0lL9
y+vyikdRZ39qLPOS5M9jf/gf7z3PR6rQUg1/AskSEqIkrsKueYwyI4HES6T5Jq2X
eMshPR+exnZf6H08ZybbxOq7dvq5PRvbND/5L6SlcL+GDxoM8pUQtrNUxrErlpR7
4ZHPm5zCdQeo3flOTB9TrRSXH70w6RnKePEH5Se6N233LVxBLg710TmZllxVYQ85
9G/0vIs1tVsyMz2D81ob5E5FK0rWGIq5nda/3IKIpwhjC2XyH6zq1NxIeIsrrItr
hoYPPrh+trTycVDq99Cs1de3X2ezkYkcY0HTKGccm+n6fC12HQ5BptPErGukEJug
/88FErAvE8JRk63HlPkxyZ3hKB+Y25s4bW9QFKN//B8U3gLsCik+FjDxzEkaKT4H
ar1V64bRBjGcCLfqT6cq1UcfyMSVDmasVUyq/rWnT/ws3WD6TLuaG59EOyreVhGG
V1SUeCICO6xRq+zbiouu5afE6nt+o/4y1unzmszH3YFnqIOTXkr47Fm+CEs2yHYu
c6T0DaPr3di1/yGCXm0L1ySbdwOyX0UXMe3QLhx59azWtoL8ZA3xU/dpXtlk80vB
YHEW7Be0JrCQXGkRK1RBI9nL89bGO/BbPtZxko3b1nFFJFDtXBlHs4XnvhVlJ6jc
pLlIns4tgH+w0LCwDaThrsllVhwgeu18rfAr8F0LoZEd+JvgvKuF2kXMA1HmIhli
hntliIxomlu9ZHjFUPGTt/mvAzSmPgkIlKpuCy9HTe7kdoDzZchBV+hvsEcljJBR
YG3EkXbiXRfYqwoXpmIrunwq6c4ohrhCW36N5z4I4V3rIRcqGeLKIODtBbG4RaBG
mRSzajG1h6cwSjl25X2ocptRqDZUCUrZGchsVyyBmtSg4lZphiCqsRlyzXHjPHSB
HCaD12gdjFBT+YrZfhmzbWAsdZjQNMRsHazIkiNNBlaVyTidz4Nn8u9x/fYdexAH
kN09Fzrv7XBddijPoDQ2r+ccF7UzDAqItFIcFahtUB0THBqxiN1e5myZZ1vYc86Q
yJoW/9SRZi1b4BFPOIOV9wqwBwqvhM4OfweX7j++MP4LX2CAxlVzbQqWECCCNMjb
v2X+MN4w76kGPfv8rkuF0GDt/SoGkL6D/X4nex5/nHCQcpA3IS28if3p6eDUiS4O
M60aTJWK+V+Cw4fxhBNH1x60MOYuS2/JPk6FCIDLnJbnyXy7F05jGClCafbrg2fz
igIdPmKv8HNFgY2+OT/tB8XxWXxF/VNzRPokTwye4+5ccdLfchNxEdXB+aJ5tXZe
crPm4NYZq9Rc4OLzpNNEUA5yc/y3ImB0e0xXftYZnsv2B8Rtvs2a66mB36yAXqHz
Zf80eFQJOrKZetMRm/Qr7pFWxcDoLzan7DwhzNxknYe+iMk8KxvWV5802q0h/C49
JGTYJ6HWXCtOIbcRMQ1afx3n0tviW3IrqSKapv8+943PvIyLMsdDWoA6TgAmDpv2
iRjwujxT99NnX3YH2CqK4PBt+XAA3awjEkmh54dfblUUnxW6JbzXjTT1zWpT568R
9+xk4NA4QkU4m/FRVizL3ca26FA8e0cTvITMc5HFiy2s8clv/AQ9W06rrE7+00rT
eU92x5KdCr2OUez7KWNXlqVAqZUe52MYBZCw2t+KrfsaMjxtw8mArOLx0QTbm0eF
kL9ARjVBn+HDXSR7SemFbdBgrJX3TZZdbszB+Egok1Zd4GS5X1kmOJoI7L3ExkXp
hl2cJelLzOhM5TWUaQqMiY8zOzGSSOom0OOeR4OcWaZMEvCzVJ9GsPuXO3D9E4Le
VBMmMNzKp6UgBYZ3CGleKhvc+pAWjURrpkF4xUS6TDyn+pXT4a2/v/bjobZllVvg
ECdjnkkjMpIrA/kx7CYnXWUqr0BHqa0QOBjJlx7G3/0HdvgEQBHs1xuwRWbjyoQN
knzw3vDw6OjSbWy4eEiSd4Z1idi+8+pTv1nfXqwr54iz77a4UrTEJy4TCJQ47tQH
/0mejf7l2OU39FiX+aHwJpcaql2Uw3jiIuYOe3qy7wVsTSaTqMH+bJiw2WGM7zYJ
/3X2nrPWoK92hB4fKi7RKk9CA/vEUoRl+wHr47y2BbyTs8ZfIa3MhQyPNyhPHPwu
Ddd/XoblObmuTkx+DM7t9z7zEQBHzms/HcwQYecfb+bnXdTmZgEZ0CNlzUsMG9Tk
aB0OkrShx4jNJVBfseju2loUQRcpuPk/DoG46355nESgOC62INQyurmtN3EwsR04
6AOnoCNNW8PkwAAYdea9KkJZqds/wQEDepEh0gThlEilzwS7PSXTtYfjA7n6BTJL
heCfYESDOwCih26ducpocny6wDNYyXwB1ewf+L3DWt0zUI7wWiQ0fKVQYcnQjVcV
DbLg+6cHZJrxg87VuMzPHhkFvt0UJVRixdDk2nq8n7tpXDUHduG+dntu2beGAj59
gYOfzGlGH07r4mbdMJH7OOK3O2NyhB0sb2RmKVHzCXX8fmzxCfx6t0sFlEs66TG/
Y9grTAol29sEyjLxTAqtFdY/mW6JgMjk4kcGk2PMsrNaPk23CPgZL/OOyIT3uxn+
DhkpPISflK5Nf8zwxHs1YfD44JMG3uK/iGD/ks7jrrGt6P/trli0HhyGVaFUsv6F
TVJdPtUnWy7431jx8aomXbPwdq46PNR8efuKYAqiLAwTTOVaZDga4LCKWb3tJb+/
WSfJCalErkKvi6CCmiqGXP+j4RZ1v4STYSyNbA2uDCnGnYU54cAe5WpTi0smB/MA
vZwyjv3NZ8XGOgb8p8G+qynI5eNT8ZtPi9QCuofDNNUNlTjESxkxriQYiMwIgQ9B
7OmmE0f+Gl/T+LRNHDQd7pDwAohXLzAOMqdeJREVu8XhKCIlkSmeKeusBRbOUaRc
cu5SHjj7Ic7JrJXkE2ITdFWNBL7f9j6m43IyBGcDtyoH6wSEtyJtw4Z0CvgUGgHc
neLwTdQeSkfHGctrO8hAKmaSjkgOxePHuHBe+cH3WLnxOlsbHRIy9Jyz5ycyUAi4
Gq552m+nZed4MZR9ezbNnDxBbYBFb8tt6cqo3d97a56lPW++23CmPfROLyXZ0yCJ
cmXr8+fq5G3VmXyYoqBhvHQ5pwWjlRqTrINrCx7tCy2loXSgA+N2ryanhlvAwIev
LBLyYsREl8++49dq3RV7ZxVkLk/KJcUI6wahZXidlpjTyr7bo2ezqVGdGpkhpE6O
f4EvjIBUN2FEXzTKmBueF9B4lzjn0/kChJkt2xr1GgO7weV3xu9QgR7iurClsrJn
QfD6lr3jaseF/8MRzxVkTv06y10hIU5GHMWDsIOh7159ox6VIHAg9shVqT1r8rtN
XYGvdVl4VhpdQ/dquH6MTk3KPzKKfxxjLhOhu1b/EHxllTyhi2PvB5vd6mbl8HKN
4UNysgaexrr95Q6E9jeoQrcMtkG09XOkEVb7qK3c9pttTaZ8eY/XF32DU1HpwH49
DmqPkc4GFh63HpWhFPd+PKX0RZlDH+WwSOxyCCJb/Db4HNu3sIDRqWrPUBVWXVGr
51yYV0x9+E6Zb+VesvkxCYoIGLaty16lSqqzhsNjfCdOi9mrMa9Nh/uoXPesQC4F
+Q5HXLWOjJ1XmhGOli/6i0m2pYIZYyspdInHzs0JSXfenFgyCq4CCdGwDqKZn+Zz
sNMZ8jB89vrcFglz5e5qagayEPiz5xJGYZfkkmszA+sk1UpWgmsVJgcFs7lucSzz
k4VUld3xxyFLUEqJD4OqVjtjmwJ5430WNETckHhKWrLEr0kHDYmFHjkhoTJ5/8YX
aOw9joZVcOfSSbqb3lf5gBZu1kBl2qepb4fe8k8o15YhgK6dkNMrKG/bS2xjRdhE
/rY3twoAlX22yoEE3GNpQ2NWuBQ9YG+02Sk9K0x3iLbRCRvoes6x/3zJKrkvLW+i
JO4nYtT8FycBBPxUEEUCX5FPlrsyUQ7z1T4Y2B6/oWD1w2j0KV/cJbkqHYwCuQU4
gHoe7J9+JP3pY8fV6f8MLiioRMXP8LHZ+nf2qHaeZygFC4ZMtLHRIKoATL9XQUFN
LXgUCx6kEOmWvbr3LHziF7TTq78lX0MJ9tVLXAUxOE9v+F13ZzudxUvyJ3eNezpL
OhStedbWd3PwFS5LHUzp9jO1auiYWfHARPC9pV3oxDUjKimgaHbhgGyuGrh8xQv3
XptQ608lbtSnxRhw/d3MXj3rAHHSYCJ9rZBJkv19m3bwuAhFaxOkuGL6715jj1zu
2rZ3dGwO09PyQRdzTXuGPWyspqm4A4YexyCFgjp763hTS30brP8IvolLOCKi/3XZ
NsuqJ48+LYHTLPiVdSqqoySa3/WNSlT370RTAZyHYA1617maE5R+sVQyGlSftnzQ
0yDj9eHl3zOovFYzAMCF8/YR3sQ/Xb+LOOUpMPIstybPHU1a7wJRCxEt2hp6ytlJ
maqwDbD+sj9cjVKZekx2gNlgNr7d/xLAoz42nWmABTsj1XG/Yozr3HNExZ1Tvh+M
495e0ts5X2EXvfzXD9W7zkI31OdIb/R1qy74L+qqU1tXnrI0g85mgkXCZnE3LInG
gdIHVDyw5m7pFg0twfZS1Nf5QDmioofIDmXg9hDSK2XnCmX0kyeYzUbWtrkpC9cu
z7NBy3ikICyXMx93ul10tyBxgZSkV3akcnTkp0C7aiHZPTK60ft3UnJBU/MLAqnu
gtE2IUnpS1rArJklTB0FCpUDMW7DxDZj+ZDQ2QbGtv5Rw3o3Tc6OpcFX0yiKtyNL
+UKbExUgrem0RfWf2Yc/JhHkk8Tt20o624MvOCpW93YyGtKuAiyC+GB2gtm+lLUW
Bq9BfZKIAYyXn4Ih0kFR1ur/Jkrw2pHlaCen/qbLkdtiLOAET1uMZIJ9U8Cz7wSZ
uCZIHDRy2n/5sKfvFAIRf575yaxvgpIThRhDUg4FrooDL3RaJmeeA77TUs42vqQ/
4Kdzh/LU7OY0Lev3KGB3dz9KXfojlO9E/SEBgjGIhgJ8P9MV+ndum6wFrT0B1ODa
QdjXFqA76JqhJ1anI4asm3Uag8JDuxwJfoyvsX4mU3UfLIIv7SwTL9JaVRQsFo0p
PdIWmKEF0kRL2jkuoumQitpCnhmk/oxD1mbZGHM/um0UdFMu9VfrygWIRs2vcoRg
zH/ycYd5cFOglgdOsW+qWt960tybVdiKZuMyh8Mu8epV8UU6wUMpU4ITF6tFrrkb
xwFczSjYMgnxajXICX+IZcmvT5raSi92YsiRwtxRDueGWLAV1oW/PoYl8FFW/xcw
mwRHZBTdOYrfZPTzlov+ZOciUNmMo8XECXiiHl+R23CGWaIKXQnOjpWaa4/lseg+
ctvs1E8hDd2lSKkheAxdPk2Woec26LKbm7nlbxfguZ7qDaxefHuQSuMZ93hGiErr
Xo6cYYCuBVxMP17habS1izkZrTEVJIHRMhSk3Fbz5KqztrSrthZLP+Vy2GeIhG2P
TdY/J7Gw6ZZuZVAx38CMjbQn39kxNEQAk8YhG3kwTPs2D2pb4JrrgZhgUtQa9asZ
/nIxDX9CUuRVYGC6ZOKnVYIDxWReHIwD2XWuThZ0nfAtylud2VpUsIV9n7z1V4od
wsXkBrb5BUYD7S5wRkpEZt0rADFEPPUKOtI3AT9iy0LN+xXciRuL5a9Ayu8Y8vTB
6uZ15LEQcKWD9OBTSy7Y2HMBzob3s8pnSPKlyZgW75hdZqVKRq+1JJt9YepGKwz4
Ig+6j5cEZNqAid65L90YjeoYPLFTwCjPU1P2cJZCPp2gnWOTuX5KkfgUjawx7kPm
fg+91AlF02iKwmeo5EsawprHym6pU9ieh+L1SXHqIyS/ZZniDg89hU041HBTxv0h
/mYw4sgAQhwvCeST99CWn+FKwGWJVJ+zuZh4d1CFMraFgre8xXK6A5jrTwTwcli3
N6FiSlOZBFXL6gaZuKtMDYlzML3jdz8MJEqT6zS/x5eXnSCgkfAh6IThvT53WC4z
09balUh1OJcWVoFDbDPem8ERiHdn0YU3Kiwjvsw1HNtXoyvext/r/33JOlMg5VZ9
ldpEbfIxAMk5AKOcxb39m6C965daec+o1IxbdTIFffss8NNXIpM17omARNQM59YH
5oSaymxjGDBl8XF4Zx2UajeD/WL8aonQnLBOzgndC4JW4tB07rEFsfXyDl3gq3dq
13k4UpFvwivknI9rGg+TuhIXNPM0qYS+wM896ff79D5T1qlgbx3gNBn+WpihGTLU
f/2cMnH0rqrHLRo+t27IXvQJ0RsjLtF8zmyf0iz70yd1jv9PFrBQmcUvV7iQl9q5
M1aeO0IGxwJgBzUYpvOfPzhIWmyd6vWSX4U/6TDpsYEK2swExuYc4VV/Pm5CFZeN
bf3OzzzbNyauF53A+Elm6T5EaFDNC1wKWOEr+WrZ32lPpL+Z3Vf9ecwgfhBXlMOP
Zo0GcwfV7jqriesuLWvQYdrYL73eEXRPGUxK5nbXR7C4ormMktxuFQicP5+QS4dF
B4+UbJ1LpJDp8bqraNWuhyoP+HRC+bU8cs/UuxAnKZD2Jfb8/enX1P19WfYoWdIm
W7Tx/ZNW8aC9RCuKLNS3Y9KxM1U0BvV9HKv11dL1ZMPCjvYyrk9nHUn0GMPC+ILE
HHcdpG5lUHbE7c3ZstGsW0pWmwE0vUISU0IrGcgHaBzC5bwYdOQ0JWg7nJghm+9d
AAQWtQlHHxsl2Kpkv/pzZUXSDsqFQC2CJXoKwcj6T3VR3JqzFLFK0HtsIhtjz2VC
GDn2Qp49YXRMpLgfEinyLCZVkmEVKLFT9K6r1PUSPomIdOaganJoEU2/ntr9LWKd
osJPVDK0qF5lDW8nahahDO71oOwQ6LGcHjWk+2L01096U9T4ipOWGmln0HTiglFf
1WLmLsZv27CmVa3Geuo0puTF2QTfhYHtbxFCek0EKBNP8N2rC/ID/+yR9Kl/aIN3
258qtXE/oKSEpoHVjeRMzD5DnkMR7pL9foCHN1IkNSeaQkiM4fyD08rSCYOH9mjQ
Qs6SRCQnx8y89D5Od4NGbbnBeZ5LiD9qO3IIWkpXn+He+7dDWHA2jimnHhZRBZHk
Elqn9DzmtzyewM8tlTKHoTWJFYTxZXJ2hyzKkDG2LPk1bZZDwPZnosN5RWOTxerv
70eaHvvJl1WwX4WVfw9QhSEud4whTYjY6l0nuops59yKRIpPLRxkgZP/SL6Ags3+
IdMnips78J0PeAyqYOtKwPfj+07TCUSwrYFji5G65fD/iFtCvJ7QvM9/p4uNryR1
V5hZFls7tF4pHG7p9atIq9HR3BgLZzxrqoWlu9CLEAqB8ZojEs1dU27MXEb4WVS/
mfCcU8I0LqWarAQ+QZjw20p1l612kUFu5qls0Z1kvup4HsNoDJecL89sVaLbo0Jk
E5mi9AOqDOxGQB8KkifySpwlQcI0GlA2YIYjMNlCnKompPW8OpKr8MIhKTRgmOjv
EPXTfZmJ4NBIwwLlSA3guAxZqNO5Tmr3tigGfSKb1gW6DOrb5hTR254Uw7jp+G1h
W6GA358+qEGsGowDz+V58iQCM/UJyqZdYiYidsTCsZa4QGj3qv2j8LEWYM79Is7x
BVzH4pRCX6G9sA5rrR46z4xGw+fEI/jJvDz77pGhymtzRq8JrneKpVNmEoG7wYLZ
ALbSFf1od6/vwDWIjeNTncxbBJt/dTOQ70jTHRvXV9DTJGl5spPWnFfwAVzDzWwW
u+0+qzaPFnJJYR/UQE4DXMXlblM/umCVfcZ3E0l34t7Ov5AvQbfiGsvdWxGp/ei9
gLBplQ/oZsJkQRccWfO2xC8bBCRQiNbrgwXG6NUWQKjHRWw2fQ9WT3dokfNdHN5n
t+XvQuc8xIjIcIQkCCshvBgm4UXUNfAIkdzJFtf2YcAWEDQetlHkGYNhD7M1D4pO
bGPUSKcTtkL6O3HkkOQx2tC8+QyM495zABIQ/0vr4OMi2SuIuMcgWpvllWlKBPED
QdY1iEe+U1Vd7Xync9pWhXsQE4+1ILJ4n4ZDnyE7XFajj+2K18FSxklwC2+yOsLd
F6H1Q4hq/rx1MROMsR2MrJ04IrR5dseP2jnKhL2EErw2ZA9HxsMcA5DdkqqFsEMS
njptPfW8xFJOSQTwZq5nfJ+5VPUXS5+Xye4HkATdedvsFs65kCvWeE6xe6C2gm8o
X7q6FX7E3+GaaVG0YWpRhSLUTB4d8FtlNMs8RBFA+irTyCsi0Km/6idsul8fzE4l
SDHcDIyqMShkOpPIhEvN76NAENslpEx/k7hmfH/xXde00sER5dAwX77DjG68/BSi
BJbdGaNnvCTzq5Svn0/zLnLMWUdgwThUJqYzsgZpzjI1eHV57OnwHE0GlLeDXP/7
45UFOULAk3mTWUtg0qtFggwjCt2z4J0hKWKk8qvIoXRgDp+VviC6A/bd0ZpYWtB+
Ob00ZY/BgE+ld65cMQMaw3aUY1q8AXz3t/mK6wHdkQCN4IPrOq9xfqEcmknbzQ84
hN0lc7RTtuZfRhRiCxqcp8dI+SfnKcvE+8T2zzPUUF/rjMKZzDEy6AXC+fb7mqOC
xDvjg738BQfMAvtsfDS9myLOfmHpbqF+5HwfBeGnottTIxO/JPCXAwpv45GJXyHo
oCXaGrfTXloqhjYzcqJar0DEzFYPCCeyC+9ND/oKGlyAtNe/YxVpceZhYV3XMUDU
rR7MJZRuoQAdpUpY/A0DtrsDnZz6NnH7KQEKy4fUx0b2OsA0Ntg6xFYZrKqNSaw2
zCzDZ0POI5KedHFCKvx8kBcgF1CWSkPN5fOugft2ZnCnb+1ISGKhpUbCR4BSKBRC
5Em0OUkAQuDNJ1NsRFnkPnT7VtALdZg/NJNbMUH1EZZJk6zk4hCH5OEHzd7vXmz8
JXGNlqztLkMjPAwY1hrr+fgq7wClxTeZAxRZWQK6GImtly03ebxCQ5zWRbpN/M5s
60UG7ytxV7aL4ECZZFg4QiHm+4OY87CiYFWRuu0EWWqnoZHxqcUaHQebcRazux82
KFnUsbuF2WZnWQRTMiCTrVG6X0zEIy52Y140ekpdE8pDdbmFSmdfz+nW6k5+/mly
4xf61KMPToiYYN1hMshcCzToxYE+HPWFRKsjJBGIubqSA5mRRkxdN4qYxvLEy74l
lxLVLIrR8YxgUdceYB9HxBlFkhmZPwtKSIfHkdsCYZ3X0oXR3vBFJp0dpmTNPTbl
7uwHRxt04JQJhpHTAgv+zqucBxr7Xu9SSVgB/bNt/9/yKQloTqRa7id05cdqEAz5
A6J4pKLbSXfJmn8BPNbl+dMm1DmsWt0wAfUIZFNbx1AlOGDOIHnDHQ4Xsfg9jBUQ
et/vmfAvqod7GMZg4XRfe13IrKl5flm8ValKEE1hwX1SOUk+C5JkAs/QvJaVVDr6
U6CTrgipUjAYZQnOF4t8ZgQCUWjn4GH879bZUngdY7eRIm/aMDkCHSsg292xVZHL
bzZg1b/tqWUT5jw5w2BzOuwyFMVY2ca/c2BqjsfEtbbzTNsAKAGjQe8OfnQ+vuon
Wfy8xWcVxDUjEuqXWNq4c0uM8LP1Phv0WuHP0oVp6R6uIK9fYeUkC15g7R2VTH9C
9k+REdq02MHvS8WuRvMqtmRhzo5CbfVPTfEYcKjcEwJPK9fJNpGdPqIUsxi6MnHx
a6r8O6fAjftumZfScxe5O/BwSiQRbhA7jVt3aURPSK+m+mvPZZcmhlCQPAq4/KbF
L5rCE8tMEUo4Yi9NymID9kQHqWyMwCuVcdXGc1mLOw8MVn9yS75mqkKqJshSghMX
hpCs4/ldXCDiC/LQprKAPIQ0r/T7oHoCfeprOb4bEQaVllcJ6i/VC4e0PKkGMMz+
dgddwSAZb7/UYb7l86P61QKuw4xAEBXKFn2T6K0wiTF9TEJXej17KM2fjCasTs6W
rR6y5C5o/MG3wODpyl2EvfCOi+xE6ZpY6qcHBBRFF6oDrBFYUHzOw/tCcf1X3KmT
vw6WwgMFFXEJZP8jObRjjYXNCSp3Rn2GLQmLmLDuBzF1DAdzLycv00SjiayIbUY9
OnZnERJufE+b9YVz2lDCV623SAcOkP2NnfkQOsN592rPklivBCRIOjC9OBpj1x+O
YM9lxryQv6BgVMY/veaqmnPirhwKCIV3SLXo/x4U3D24VMUgQBSO4gZlY3NjQyqY
2orwCNzDyi5ypXwGFAIe3BtjFe9eOig8SSVNuk+DKzr3mCkJbUQ80O9CgL4W97bd
WYQLcOlFw8c4wXPuB92vqpxQOZquGN2D+Wlwxlic3Bmq3u3lDo6Vnsm2uQfyyo0f
3UHNF3Cel6WYytm3U6bfVQ4I1Qn6yyhh9/mrZeMtxmJFKT5bTV/ABykfOeb2jlg7
PeaQIv1va1uuFoxsovXYJgDbyKwflR5UTO1iWZZ95j0kfI7/ZmX0YR6sBpy2N/dw
mMQ32QQq8NlDTAw8s2I8kgsSIdc5mR/zceUWv+Yp65+sqnSMSOsYDU7yOZ2jYww6
ix9a5ptxLXTDTmt7FlnwbdGIm5Ulhawg6iEJJ3wJxFAeQfWUPg7QhceR4sLtq8bH
GWv326NAj63yUwMWNlabM2JFeO3Y/aU7bBoAI+mXx64wJ2o8reGY1Q9RouR2NAKF
JkhVOHO5wzsN6jRVmQiFYmQQ0rmlPeUASvZRYkfDMJx14Dix/dyfu8KweCDBeBe3
o7/58KJCDK42vbE7Kv2ocmflEYmflMClSNeNWipha3Ud889pnOrVjBBpVsJ1rw06
3uGrmiyPOs7k0lfBVk+pEqmKCL3LLdMvcDjxJNciYzaUFQtkt6PjifvtyyBpYUPB
iLtbaE1Jraplz9K28j948PdJB+TZI+6pFJc/1um4HsOfCb52SICHP8DDaQBkk19L
Xwi2GB7VMutznT5EuWOD1NucvY+wMbLf0gDdOK5j84jYBidOAfTCwx2vRpiq88OM
RggQm0Mu37+Na7j2fCt4jGzpSIeESJLzHN2VeYUq+mnjhOisVR5Ugi/MaReN4be3
WrAnrMooYQZWt6v4XDGNzmlzqKKXI1OLzooi+1FndRlhqxZ5kX1tAEFiwNHkeCPo
6LdVYXBvsjG9SwB9RNGKSpJ4ktgQFeH5vkKfYF19h79XbIgjdS469Dsd8oQFZLaH
qnCYHXbkVzM0NeSgsG3jwj3YlSJ3f2Emy3clg5JoPHuZ9tUjaGW4muLHNPZdLP4t
KT8GutYOL/uEMrekwPQPuvDhVeI4lX6XkOxrfM3h9eZldhpjMRHBkrVX7w00fBSg
PVtlNYijMl+8qVhB5IPLl4y20u4OIjA2WR83PaWm/+X9c9+DEU2exPHztFUevbDU
sbGEv2jYuq2YmM/te6oSxarOnCoMGnxucKy1h9n7lkddHq0opM9NJ2925fg8Ufwn
padSEjAdJU/HDDiuYPlcfvj68EMWlX7r/hn9QOna9AOf5q3JBk+i+0ypYHjiYd5a
AjwhcA7OluFsS1QpAeWBGD8DSuvhaqk9zIn4RA9RF7XlfTNSyX4c2QO1/Ps+bofk
uf74YcrxRQNckTgEUVC4YOO+xwFffMPgKkwSytAQYZFJKVvybbtx0Ww1fwfqDou6
kmggM75DEBNorjmEnevOqhr31lcXIBJoRE4e/9DiwXvazscbgZq1H2XM7UX4OCD9
MZ7vkslQgqIYMr9ypbD5W4kE+cBmG89Aw0z2WIc0wBY+nobM7Uj6dCEasMZebHCA
M1j/Rcjv8G7vxEGfphV1BDadYSlbzlO1+q/SC3tM+UmAObmsTiWCUxrgriJ1CQVS
Upy3n2svuBF/EyQsaKvzcL5FBSFUzyVBm7mC/U6r7QDaXVP7gvUGUgTuH2agKfHb
PNfVk2pzfLzvsFj9Mn0pcsreihFF1GKO2OaV2yEjLthXQ3VnACX2s1yr+yoZbq2j
QgOVOnUHYTut/WfSPsZsMbr55wWRGbZgwrNJY2LddMqthEl+viJ+kK4lLNbw8S7+
zhGCK+f/ZPLdUInxeRdF5AROIqBQp8M+EkSHJwFNLiTrB8DGDfgYjbWawAsX8NkE
9MA0LMGVavkI3LDpaOjAH/kqTsk5+rskKFN3QwXkG78dreDCH94oaXIfquhbbhdX
p1I1MDQgqhr5rdliHRZ2K0g45eSuBn652KNr3h1La3q5xDk3+jz6AR4UpItsC9ZD
75CdCPKGjg1IlRbofnhxU+EZCEgXjob8uXLhow0e6dh13SqMu9+6NzxenT3dC8r3
rv42RrCr+iRnsw50jC50L4L6hs9KRCxGSl6kX3i5y8p8XEaHSV6g3Oac5WQzZ6Ip
9s1eSvOezfa6EfLIpsBF2PVC9MBl8fAP+WMLTiUEEvum5dVHOK9E9GVL5feLF1KO
oaksjCCuKAdyovOir91Jec6D73s3UcWymCWZ3L+jDwcHdWe8SjiVCnNmx93QZ7ea
dhIoHHlspCe17lutp+yR5NMBIabScVw22xmQfYhsOf63HLNTdlmdSwAZ45eaegik
3Wf1sGUtU2oYpzFx8ic6xty/6NeWmX+U9ILfiQsJBQ8NsG5rcZc+HOXY43KSd8nW
iduDisAQVB9v1eYOjdOmzkkUUj/2y1LqxlR6lMEuGi+szTcyK8vUcNEeVzQ08Pxh
h7stjZu0Zpk3a90SPIHpjIoWOHTphA/LPa1Rk+YiekYibVaSx9lRD1qm4RYobule
ww7Ce3O3qvYo7mhD4aRDa2nOzmUyfreSmDJU+tDHNNN+8oeYDav3FRJDwqfGdGOh
pd1uvhXo/emYetT0xTWIQxJP6v2iziSmREx4RuefrIJI05rtVZFQqzgHhNiAJiuq
44o57vJ0mx2d3OAvRd19tsPhbmhNJhybNWtLyHW/EpwniMeChA+gGyY7vr4vY2Yq
GEVEIlAaPsaZMmIqeLSldYVCSK878KGJDj1XhB3heExf4eVxkB4HD267LO6Ex3XO
KoBmagchXPktcJJpseh6otAaOTd2+BvwAfSd12VObH/yIxwDye9AMtKP35OWsqr4
mn2yfOvaAOeynnIAl//W94ShnQ19M6OGVvME2r76WsA0AwQJCZbn307mX4zFOryW
/iOmWq67adGz4BRxFp6qQn7W/5yUNV+jPjJFhBZ12X9P7pdhSATSNEhvX7KtkuKk
/npGnxMAwTshYmcS6+N/kibdpyia9V3qF42ZPrFbhE+629rFLtbI2DFu8HSkKvuK
Q5NQIhFvmJO0RBZTzDSRszqeCHpSGDSIOUmi+JkEV9/M5NQtB7RIE7gJnqXaxG5n
DscnKHEF3wvR0tYv4jHYIuH9nKwWoPEgwYhCaHWt/ERZreb/Hm0VtdGM1LdGp8IS
SGRo3BXJgjY5lbeP2M8j381E3EjE3AgQPDhOyK/KJSQQo/s/hCRWSHKydpjothB/
xWNp2qwCddKwlXw7I9LOvb0+DSZZzDY3U4GWKSQNH0Y9w7nwd3MgjlEi4sJtUEXN
tvJxP2tUEEdQSUnhvGLpKHqONzZZPS1bakpgB8y/sNmI5DcB9UJE2xzPy47BygPx
+46bcOkTHDzKL8OsOVS/KlMqhzzGOUMDhDSWdI8czWowVespWFup6RALLK3ivrNZ
a2Cr0TWVsc9zwM0MN1HTiqNiNAMthmRuvMFI+RxaA/Z+9tAplTMQ5oHLUTucUlpV
4Ic6ExD6Q7ptrm8ZDDuTcS+1Vfqq40TITLJXVgzqdDcG1mO72Cj8dgDSXR1tCs77
p2Y7VNqSVsHMwovrEa09luDHmBdW0MBqHugEs/CECz9XFtMJ6ATopsc53qPyVl0A
lVGivhVViQYbZ2AtjAUCyU5AAlfK9TINUeZLn+Dpt8pJj4yofYdWcOWwrxkBjkEQ
vAgUi7m7Nv0iFb8eyDO3nL1nZlDLkWe2g/Y51+bdaTtakGVp7Sss8KLqdne4dmyY
oIBRiAI+Ay2wSqTw/UwCLNGgl1OcxC5+lTe/Ta0TSubLtnJDExJ6x5SJfFSqrufE
uQ0cui/I+C8qZJFJCd3ljfvQ/OdrXuZ+MyGJIzJe6fED7I2m+2jYSViHRMvAvdlB
NYCdjZGF2F2rrR0biL/dpp691KJY3TF+HHWytLCFMekNScCigF2g7Wei8vFF9I21
znVOJ6RZxDaGoLoTZ4I8yVZFF3qAV2m6dlssoAVrmLcgVnctU0TcfDvEDga+LMbB
FC+IA6L5UUbBy7ZuFW7ifiGRKulwdciuc6EQqnJ4nI7h9tDK8mfXLMiU/SM0a87l
upTnwY/mvg/VWzF5bOredj9YE6erUZjVKDHnIiB0mATXoTPTPvdVGMYadifpERVI
G41GHQxpgzH/i3bHWf/0HPSxR4zQTAwDumj9qCj6vVfgZnjGtvB6oyOVk0/vyu38
uRRPEualh6ucRR/B7PAUSsLc+E/HLmYDlX8sDVfUXdZUrFz6Nvep8y8tN/3lQX5J
IB1b6mNCDgGP4Tx7KWzNc3kUDo9+tEVLjEK0nq2PjtWiQhj8qI8COy8fhH+qPrDj
6dvcl2byyLn0KEitPj8PEJdx4PzuUKbKMTUQlEkzVJZXJjDIwwhIxzyPgNJ2BjiM
4uyqtdzLVYNhkXPI27GvDPtThv+UzQFwZbucu24mX6TrsnYLfZCDnmuAKgFIWKIV
WME4Qv+eJuG9TIsfaQvrQArkU857n3Y+mNGk1mVuYkxOYInYgtZ1NS5WJtRDEq7r
ch3nRwzC5QtdkW06pEVkxI78F+PFoODGEOU2RpM6kM0Ab8K+Vw+tf2FNQ9AVWL8z
pS+wzjufqgqZmGtKY7XQQrPthp8OZRHRDpxh6j86Tx50D4ST7o1nR2bGadamgsvC
fYKcEiV40b8DX5V8iBRipTrymMhiA8rND0Qw/6se8pyg9SI2hGWsFkTZjeDU6MjN
2pZ9JYkp1paYRnT431qgWw4uU3yHVe/8wt4uT+fkRyYt9NJsGRAXj1+SUo4NOzk0
B765clZlaGj3WfUXq9D1JNiWcjY5FokUlYe7R5amBblHzsV0ko7t7MXaV8FE5b6Y
5C+s1jSjDG6kOKrmR3zDbD46QvLgZtT72RzdzF25WOSJa7LFsbZotYMW7RY1pK5s
G0D1u0RGUI3xweiBGsohsaIA40y2ATvzJCLJaU/NZnFsb0qdcFBdwhcjJ6Qb1JB2
dqfoANPeCM182ZNJUPRfuZn1tqv8PVtvz/IF5E3ikH2BNJqwA1HzXgQAflMSzz+L
NCxD0Yd5bYRUhYQRNYEvJMw1Jky/tV5Oa6NmggtZzwfnZJYBZeDEbQNPXt/VTYzK
EglwMihVl4AAsDikmyNl5r5d8t/UzAP5lU4JxWxEa8WY+2s8/nDY8LPF7lSnou+2
frh6phiaAEKGdr/vqktE8vgIa968x1oBu60N7Lg5gbo31U6ex5rYjE8ggnngnJQF
fnP4tweDQADq+8tOGHyQAazFGQQL5UPAV8h1Fd4e9EFtvhFM5M084iQs3sIk+QXQ
Y+9lXk+nKqp3Gxc1DGoCU20FkyaFKTF2o6l6gUFSuL+RApC+XTtW35/4ifmVDikG
ZcGztObYNbZb9IHdJp4134hZhouaUNrxBSKLd8AOi8YpDk5TV3PniqX/QMz3aVt/
fGSHNUzlGz4Cdc9CR2gcHR4L+4ixTqGD0B9zEjkcXz9fwwumY3iIyy/zBGDYbTJb
wfl8InaZYtkdVpxhouYa19YT2X2mxszT08wSltSN+ypsBjeA14TJRjX8ZWWnPpjd
VtXgcbTdkSeIlYvRpv7hTrPESQdbJXXoDcT3LLne2fEcmkzkMdoafWBbP1M71N0d
jgOBwoNmJobvlI9lyJxBfxFqxiz/IvsPFvHkhKKlA/BIWqKydfXlYl6ZEOJSpL4H
Xj93GJpWT0GqBPw5ViWLjtdPP0cXCm2b3wSEXNwY/iUNGxwy9pD5pZrrxqZd/7Qi
z9/3qGuMZNoDvhYiPCqJXPr9czOdPUH5dSYzxv+2Mrg5b+DpLtv/5TRnk2dQjs1y
WVATK1eSOajpxUe84ex1o1UQXWsdu3Sohyfu/+wg11HXiMZQN6iCiRw4ARfZUBvX
pmrYuWon8J0rRMGvIaNPGqw+/ORmWKPO/+Pwy3QT90B9vUnMUA0ye5DG4ar2hHTJ
6T+09yR8L+6IjfDakuS7e8tLi7dORNPA/0VKJYa2r7AkwSysdo07LH7urZ4ZZ+Av
5sPzZWGjG6hXAI7YNPGe07jSafChSkWrIvzMsmGBAXDrvrAMjMjo5/ZZDmipRZFK
osmGIkqQNAGKCWK0FjfK+1RIUi+9h3SuVU/Htm64zXZrNoe/5A4nAWb47iVBYvIs
fzEFHHUEHKgCM5PbOsTCZvGcDJw33OquXEboI4MQqy2r9rezy/Ef6S3nv9y6UsoA
ZyFUjHfW5sNig6X/D+qsgcUHnToX8wMKyq/zVKuFnfM4R5Gurn5g8EIHiu17iAvt
dmyG7H1r7ObNhrtwiC4GKyLOen9YxyhygO0eVZOuLPSgvh0EN8OFfOUMVJLt/amk
CrgMLFRAZTaYvrX8+xHy7KfpN1S75dv6AEQ5hjrhzUFojFxZdRd3FRBCxYJbrNon
KM9ij9znPJ2IYMe+2EKFqQQfYTnd9U8aFuDkE0iQvYeB7o7cd7djdfaqBwJ2+Fwf
mnxtexBBbXEoiQpt1nKHn9APnj0j2iRwYsCo6sEkbaNHfW3qjFVTJR/pwrspKQ2v
bVDVwgqkJl0D7kguWSA72obIfjgItGMEEa5v536tvOsPi6U5+SA+wQSfrfeRnpf6
yneBjTwuU1v2QgYpYFLDpFA3YBHte+QC6BYwn8b3FP96bYsBHzWtQ07iuqdKaj/x
LLnPfYD73ceWMgl32iT5ceTWdl+aVpL+LzZkRYIVSW5CLpkTqm0xDxfjbpX3sj7S
ix2rW8PiDYKIS/vYhF0if2YURSbIsyAtoqlVJ1QcD37r4MY/BdARZcc/lFoclt6A
sb7IG9/NC7NAAYMfDQdWOXjcfpBKscaP9tNdsS0JYgTXTfHJ2TRKdL8GovBXcEh7
01amOqt7FbILZIT3AUVn+4lGJWEc6jxAruMyNbIPAhUIO3Sgv/bvhBHcV9PK9hUN
0t24kU7BV/aMux+FmOPQrL7LqoA1N0f3GHM2PQpd7BGbOqzIKeRcPraJPkUz0LGP
1hPtmTEqiB1i0c5VP/mA0H6CHbgm1UjlfX9D0Pw4ZOEmKcKUz9akv5I6GY2LRzaN
QWqFb/evEVFXwHSO3nbWBqozlrFmtOtjrFx96ygrw6wf3a9b9A4SocPIHhmGgKcQ
STgEJr5LQ5XEWqwngUPzs+JHscISP2i9voDD6Dj0pBi4Nc/hQ97Zu7a1K9Um7x5m
EdWo8ILicBksI6zwt+c4SvpaXu++sYqi8hzhvLP5XyJT4wiQHiyuZn/0cqOWXSL9
f5XEcIJyLrkwPTFrUZxlHRvujWDAaWRt79OLct418zKv+OIQRZzr/7Lt5PF3EnPo
WCcG5SskTuf0aXnyY+UeMXq25IBhbPe1ZqYKQPjWTlnPf+WxXkUE6RUredwBC6rx
fD7pb34VkSBSlNXQuQKPNqWklsnxZttJKIREUQLNy2fDIo5X9OjzTba7Zg+Pu3Y+
5CqIkpkUdKzwSyyaKRUpfVnmZuz6vfgNVm74lOA/QvG+IRZ4FTRbTJ2sKo6Rya5V
9Y7CuNRWnxTzH+lu+Awlhv+GezXMqsjO+WakfplLTlKrm2oKmwtgrCBAP0iOG2Wu
eHYtj0uoOXzFtn/F0jWB1FdWSGE+NjR6KDi3HAmpF34u+rBlpbxJJRpJwoBtldBr
zUuP1rMrAUzP2MbDzJ0ggDTU2/me1YTPMVnQWhHU7cd4WDFhoNFQzK0Yij2yFx3e
V+kBOOiW6zCEW6dAwQ/fPwmzApVPxyqd8txMZXfXF7wg1wUKB6/2Y2g9HextazKF
hQc5EMMoEt/SP5BJZKXLBYSleGe8zGIGtS5TKRE81xDASCkPKt4Cq1EtHzb07NTG
82O2g3i7H+VBxxcCEVUhJzMrTwVyLYa0Gz2wh+mU3sfkdUO5FBE+hjWwEGhzHAOo
aOuT9XuRokSyW17U2NKShAgFYZfTl7W/fShWxQUlAUTtEUbNwvOKsM/GUj/PnGhP
hI4gZYIhIGqZjDy/gO+K+yWHylKbEBXc+ULf8SENApCsrsIKoXFQhhauxs3b/PGr
50pbe56J+7wkBqVBxPp5mIcvsHFCBK7hoWhTaxNog82C5hnOsauyWh6amsVkL7dq
5o/rtSFQdE6YbwxpgQmwq+RQcmWHKMZam7zXTFFH5kgpVZEXAZkAuGMv7hSSKKuX
lfP8XqMdwBO51YacDSQScfT1rNy7rA1XBIwkerje9Mr1U6PkPH1QncHkgatSiOIp
Ax4SZJOnl3LChXjHt9M7vf0/LoLPrL20/PQkYrgNad51Ol+5GuLUQsZ6Jn3Sjl4L
X+ZHBV6CGqJ23SwEOfcLo7qKQKiJMW5cWnBFXGk3Z9PSQbbFvn7WsCtX+2b9cq1I
/w8IYzOSwqcHdSK2sQwlLH4pHXLZj21nUKJYLSSEZM3YkGJar62AMgjwvXxVP1f9
JMddQaqoTrAeehcoxzlgRFKVpc82S9jfyK6CpPkc4hNttB9Dj9J/X/x+XXjqfZn1
jeAu0y3fo/rrB7e62ZbUtU1QaCkh/byWGCazrPlI3LmaSupmPhiovTaPvE1qAumk
RPbUB9SByoGBbcqh58/8F3P0ih+FSYU+pVxI7lPJXNmk5UnFQG7WYh+YUMWL1T7r
wAB6h7gMQ53ijtrmMOt/lP0LS8REixLUEzxCEjl1IZxPGZI2YnEJ/oP4QJTS6das
fXpR8ll0KpTMk3cLcPofTTwMQUEj6BhgqdPAHHdK0yjJI7wwmR3tg5nGdJq5Wt6s
htupClGFd0haKtBdehI7CVR9jEC71XaP/mZq7DkN2mt2kq2/MshrQvgRYYpGobw/
emj8y8zk1vfw16ccvpZPs+q5fLSMGGXrmKVarBlvdiYFdq9jFx+DPu7N59eWu1N3
+W3ECQpmEh+WB9WuhZSR+j1MsfT6YrfifWsIPExZ1hVV5mYMl/kbPsqRpLYzD6q2
nnJI3+u+cMkCfkUpThZSA3fBlVY8F27/5JqJir3BtuOdHwrXTLw7XIsjcu3OclK8
vTZvRnDeaxmEAdFoNYGsb8YCYW2nlEkkdHhlPaFGEPOccWp+4j0ZnAwzzg/ORJzc
R9dbqzQxKlNIV4CuwXLvwOagoGewx+JHaXoxY9/VE/7x8kinzl+MqRc4vPYigYUa
gcOyTYRCkIw9OxRjvuEvzDLCIKuMy6pbRzvIiW2s7kkpqgdny9Zy3OJSABe09XMI
AOm0borMRY/yLqYU/FhLX3TKWdE11xHp0kc/dAMXSxuBvd8RHD9RRLsMNGc9rZlz
uYXKp+vEYT/HmoO7a235Dz0ZRbfEeTINsGxhvKdcVS/er1ggEogR4jhduInE9Hut
5jNq9QAGx/Hjk+7W7O4lfy25SrX2RV+DazDYfrOY3CWGYklPOwr51S1SD1JRxiHy
fh8jey+9g2l0Xwh+SyEHBE8+NQPh30UwY9Jx69dOXQVFpIpMKFgc1JsyW1iSogBF
mPxz4hPiCey4zxNvWCpPI6S2APKzgf0dpG3rrqluadb1lfAcgUGsIXy6/bWsdxrz
0BqNLJjUSSpiRivaW7/iNNosF5AQ6/8zSyeRCoOmnsZp9/Im6FL/rB3w2BcYU7ld
C8kCnp83nqwVVCsBTzp0u97m0dmZP0jhlZyHbXnqGWcSxp9LTFrcmNQa/5d8DQgt
H2cVfgi3l7VtYOUp7sKq6K0xzvmsc9XvgNahn0MaTeA62E2AOdorwez5DUxKQd4G
mcX9IcRVja0AFqndA1vFMdLoHZqDs5UTOG/nRdjGiZWaicPCm7opg6GS3+/yCMCK
xlKFBjlpVDfPX5YUy1Z/lhCKLw5gmp/6w9oUHhqVofRaRxiEhy1EEFSmtIf7IfYR
9oXc9lMb2N6ZFoUmrHPbaYenmJohYhxlSfMZuSD9e9BDDLR1bGcHH4uztj5Mz5GX
ICU/qCmtU6M6TyZopZ8mDmFVVYrSuOKUMf8DeeXdDFrPlLnreDyRSGZEK1uYWesH
tDEzNVj0B9ezgK/3mcNQBcwgucEYw1IfQ4H3/tLqo3FiAIVHkeCmNY1AjCtUTQcd
qrx7qPpXPRLy18DMLQ7vptpae9CiOGVSIsF9CHs2xF24hZCcKrC+AgmpkLKu1sZ0
+rHyE9QxKIrOQB6Iy7D7Qvu8uzXxNX6Vt1AwkCl87+qYIRpassAM7OHWTFCLhRx6
cVuL1iDBMdCdwbZoSbYUqcXvRftEpuEjpmbfWuDNV4uiMUMQGUlO8kv+oRbCjRei
01IGkabjnZKaD4jgg1HyKx8ngEjCg074G4KHcuGy+bSj9QFws03d9sD0voMzNLBr
pUYiPIS+SJ3S83VIykURLumENL0wGATOLhGhEcG+4ppueGpeAMSJj1jWNFNkF6fP
qqb+TWLqUCjvvTUkx9W68g8F5tkBE4/WWgooKJbqK7EpNo+L48Ld6v6XNdY3pwaO
2swSTpmBiQeaCFNXYU/YTEaGiL9QJXGWVV5GV4aOD++SR0Y7JWclBElo2LVGWZQb
Nq4v1m7Mb7Z10upACpVrx5cxlGEVwj0qLsVAhNHtFlCRPcC0v3EupbsllybFxi1e
33V3IqcnR73OQStG3rbUThcfiwofylj3NZ3oJdEV59rBhN2ZtLYEYCCt9kHaPsOm
B+u7BsKXdqwUOFRsf7vrnkLq4pkBHWAlWHSW3OK6MKt/yAbBQPUEhy7EYUh+PEKk
Uh9LqNgqzK7fRHer74VBAAx9KlM8TvMH+24L5BZAF1b+LEg09rmwuioJgM1mUD78
Ox/mChzaTajsCAt02PLlcLhaUBzYyap13GIsVdui75Ed98CNVwBIpkwXvpDnzc8h
byH/CKOrf7ASNWmrQIsLRpcmBQ4/OUSXzA6uordpH+42U8LJDfSAp9uzkR5x+LdX
QLIEqMLJd9ihssF4bPapMXBSYs0JsSsE0K8S7i4QmpYPHAztHKbclDiIHsq2MTQJ
m6wtqmjG1oVtsrMZcNHPByCG5Ph9N+2u3aMEWp7sn7VizIPlwoU5gP1gVGaH+vhz
hkGookHrKNC68Omlk1cUzPgYTpI8y4kvaqAiNe7C+3LQiGrTI5sSWKU76N/7n91f
jy3IHKB6+LsfI66VZXs4nqHMY+/EsrhLuAMbCDEdoFkMGeVqS0kioHlEKuZCDTGg
G+jCkDNzntXsdXLP8KoklbGWJPWQSmPDkElrNox20Gq5eQe+WxFQX3tpig1bm1ZO
vf3UdFuGwI4JohW2+7m2iYXmdWKY7Ivvz5jZQli9yPCAlnTjilOwAcW9q+kbBQ3A
wvsxtwYesNLhKC6f9t+glTyyQiZ9bGPhc3hXapavXXSemr6ZNYs1k8npm04RFvZz
+wRyQGJRPM235yw9YNGnQHDlpiCi+DMSJtk5hvI2Xs+gb5y+f2w4PzOobg+HSgXF
M4xIHrXk4ZZpFaR8luf9ZAqMGT0V6gwsxGMdaBpGjeXim3Y554rzC6YABhwSqUaF
0OdkQdpA3omVLRxD15I7ywJuiDWknY0HLxeAvnwEK3uYNa63pzIST1NZIztisCWK
3Xq7MbHpVZmO2rmke5GYQvd2cFnTqeZrNoYyoBffoRNN4+nmotEerZXONXVsMYHA
gEIGJlTSERycDfPiMvxa0S5G6y7gF30HmsV95PIBZY6hAck1CLt8YS4fotUifOLm
Q8K6aqtErlG47BVM/omV4xt6Plt4rIqJwXoq/NJLEDsnLuAhq4J3p/SIq7cIi2v8
5Ih0wemxtlOJe7GI1mUkXcFvLlq3YP4fxtl8dP05W1zM2ZYminflV/Qtfeua8O+c
C+1ccIHLDd7rJ7afG3v6zuWh4wsfe+A/fOjarpZJU3mLK3UAj8j8s1X3fmGpvjKA
rjJjDyk6gf4WX5n/wJCVH2DDED5cRQdR6V0qFZhdZvyoeAky2dmV7NudE5YDsw9+
cTG1zUieltuK0TT/I9TGrA0FyelD6HYrLshPsJn4KD08xkxds0a9hg2WjroacJL2
hu0X/tZFUE69mH5oQwedgvcmcnKDPdxTg2lNLwU531yHT+gnQsVAGkr/9ecah8yI
Oe23EKmZL97KyO6P5PhyNCZX0ii7T7I7TJ1+NDWCJUAP3n7uBWSni1CLemem6p2V
LtrO7x30Ghi8eZXPTNfsM1OfAEBImFkqx5SVxVInviv3AiNOuwImYz8vm+RnKmxn
BtEz8HMhVDUkMQZRetBc/c04r2emvoOAI2QmQemAZ53K1IY/Wu4Of+Ep1FJ4Nd61
kVAg+irWHNmp0UKuK0h+UmEhFP17j4aomDFqARredmXJ7lMROlVbuJmrhc5OZ5I5
iwqZF7gu5Pt12yqhek60sOig4S8pobVt8F8czjuqWxB8ekupmPxuJa5DIXjp6pj1
TeHIj1ede02iFXZ7HJ5ABz/ll2RMFXe6nWJNsQyzzEqzxB/rCbn8mb1SeIywkMYv
Wr+JWUubjCqf9UVMs5XrKinZ40REBHITH7P/Qohfa6tjOn0+YxmupWFM9S5pgNym
NUWvTOvG4SoS/cFljb6G51uTfd1eSaV6UGBCz/fQFSJBYs+By7ArWwHSnRGvNUpI
3+wkg5+w+CydIsVdw02VM9IoT6tLJbQ/TsSTlK8cZiHGKOczYyhb2n+9UG8nxbfS
AwAOh6DZOkyucjhcPavbrbPs/AiZ7QvwIexWVBWPV/2t2r4hlbCNN0+buRd3Z8lN
vYZs370/teyfbW/gwTjTBcKjCwK+SA2xW0jFyBq7670e5B9GHmjIVX5Xylt71R2R
0b7xplpuZGB2pIMe0boSPpQN60uotTZx72Ef0M7IgxOSbXwbGNoyda5qSd1DE8NH
9s0BeO+qAiPsIExVFck3sYfN27i1mK2PNRXg5Ca3V+WXlGceyGhEkd+ULkXj/mep
vigbNcjilfET4lGo1cY6sH0aEs09klOaGbbCIPxTDU6bqywoyCnPZjHynQnlRYM9
aKzGMcbXpv0sYa0fXPtCrEtC+A3tf9RqLW290WoEjijYkmyFkucwoDnqX3gIQSy0
r6fIqnJG8XwC7VFdcQJg+8GFc6Q/6Lk6edDs2VtQhEw3eoirO44l0eTrCZ4ri20K
bAKycBQeJ1Ogw+WYOSHdfe3hzxNie6Fuvvs5nO/mLugCcJ4Sct6L4KMo5Wr/Lzb9
IX41uqP8ti4so2rj/WwrNfDFp7r/oFypd4n2eUn9SAVg0kVCdOjPqSTvr8Zplq94
NF+aMvaq9HF/l2Idq416fHHOU15zwn4zSN/YVq3cZ4dFt+RHpwcUwJawXLSjPdHb
eJqjbUxVSQbtJRi5+GKK3xNoDIvaUtfYhwM/pZ6+Y3K3eD3hppVNAJzZxB1ARXBy
V2OOe2VasDnoZEBNx9wlhV/bHvjJopFcNsbfs3u06ioFbg5VSTMflFreBAy22Wl4
0XC9RRYJCm9GNY2ziA3Pnwz9/AO9Srl4ld91487aoqstZXORltK92o1PmfWhTQuU
acJ7nRqgY4j3CL7jYvAdYXnhnU/STuiExwlZSir2cBFnzFODfQ5JtwXNgVdv8GAF
pF14iYXT6pHkNuRCyCIicVx62stOAtLqwg96zclRbP7+tcMXqHSvOU+kAK3g74oZ
Y5/XUyZ0hPOSUR2cEilkZKZBCoyZKoOpahbxotzgqKv5fh8Kx/OWeUv97qNeiVJJ
3tLxyY3PvGuBu4NuTVoZiSvw7Swq+dK4IB61bMjyV6aMAy1Py4BmeUWqdXCQR+YG
djUaHIwL+3MRyrpTZMeJC2qafxBvuhHAhux4jLkNpI4uFDRoY3uSGtcVBdKVm/j6
CChmUph8p5WdvtE6RZGAfv1Z3A/7zSi8s84lgKnkzg5RnCERoXWiDAQVGrtEPaHz
BkSv1RWatUI0z+6veDiYjRGXBJJTCkheUUFneSg4sbTieWmrxE5vngSwQTR3mCOg
I8Ins25g4vlOrCjW0WcTZQNJjvdcTRVwBzalNn+YgXOZ6bs4e175x+zxMbG3pKem
shqV23t2Hmw7ScvSTKcgW1gJp1Wj9SlxfMmllUPPjN1FITYKNCsva1tyaVzf4I8Q
eUQYllQee+AlVUviofLfEpPkALIJGwVkAy0d7TZWAQPUAifKmzzohgyzOipIZ3e8
yYKZTwllaOj9vNQL/+1hfUARKsOSUKla8JhQd9/VuKUsjPE4Pcdr7i563UarIC7x
bXWkJN9ZIUgK/UYX2xl1i3KreGfDzRML6QFA1mYU+bc7Czd8aYJA5nUv/k+BA7My
Un4IR2up8TtjiAFfVgvjPoOtXQ0byHD78LHCo/xuqvORppCVNRhWLdAtP2AS5/9g
971PDme9iRJDtqbuKom78SzgcLteuPzpOyeXRDLJ+WrKNFX4GahEfiL5hGB0PfZq
sPkl0dGWXaqN4K1h9wGklCouEDGjjy0CL54xD4j27OtNUJtafOl15W43dDdsSi7C
aEXem+9FSk5Zvzr5Q3eGeltDVhRoYUoZcZQrxpNWjcrRqlNmNRVtml32qNqPeBmb
IT8pigwl+DQVPLhU0P3djwo3Dre3rpW4VfbIYoeOU6+QOuxg884rf3JZLz5M82gl
z3b2H9pt231JZWHbNCe0LNeanR0L4XTqXxQPhqLbd9/aHFhYteFgFXAENYN6FY5A
2247VU9YpbodIJqmMkAwN8sGpAeOWg9zzW0JXX/gSYTBAYk4F6yq7eNBkVElsRod
uXYhBsId4uRcKwx3tgDbJZQ9VBzxBun/5JBZ5vMKlZuIaQqB/+LjdgG+1GiZBMDN
7kqeont7jF4uYJ4oZ7U7KzL57qN8ro0hCKPugSVh13cRdD9M8gd4XrLYLpGHCWzo
8DTo0hyt7NIR4WkuLq3rR7VfE99sYlpEF/KTDUIUg56gzaf6aQh1yWpSWhR2f668
YUR+ExGLx1WHKf/vInYlwDg2zOOEi4dPnJF0iprNb2tRp35bWuYUFFbsQWmETd8V
8jNYJ/OfrewjOWvbSm0sQLWzVI4nkuByNoXctBOofzj2mDf/oe30LYIfAU16N10D
HpSiDI2jOvgQiwLt0PZOY3R+BidVs92U8t/Q9pwo+VEh8ZJshtFR0Y7GMJ/u1IBo
Iknv+nO+aWidEByOoPH6toiklSp/cE8SgO+nfCY6udZgd++mSawxtk4BrEy4+/pM
epA+lyqTthDXNz2tT0jWE8c+l1RqJugsAzpROpnLpG1g3+jupScLw8otkGf6VdPf
S7ODgqzyHZLonZW1CXs3E16SrGo3ucf5q8G9e/yBH07uwPKVqF3zr5NTVsVV3YGZ
NK0WQliX5hsZWsvBEm2SBYJdRUokodSzWEze3sOqYPJ3DUlZOIaX98GzwGhVDU6Z
Owrnxvpucedv7gSYPhl5IWoRsPSqIco1lqE9uVtevgqxUE8CvFEQhd0lKfIJaH/2
hqZ8cz0JnprsbkvW9+k+etVI2te29VQksQjeY5oLPWaFPW7wsjvSz33O49lFB1Lm
WXdlUdejO6y20YeOhS3ZIb9Pn7rBbMp/i0biU8LVfhhRzxI0tqUuMxj8E2jdPFyj
f3axHMKgI0NIOunltSYd1p7vj6FsL21f+mdI5fyO/QdJHiJ5W2me7dcvELn7RhbE
4SkQXniLsedjRHjZS6DJ0rjk5MhpfgcLs4plAQ6oDzhyBSB/I/7OOJY5fxe5wk56
Coh43JhJQxEfVoYiaLb8v9TOq9Urjs5UZGDpwEDykO7rkcfbF2XNH8udYkdabdRC
NlYiRZrP+cG6Mgr8hLFjKn0tuKCavhK8kae9WQGChtIdRyRK63s7TbDrY9t7jR85
wTUiWc3LOi65jt3l7KwnmaQYoQx7bVIjL21AYhWH4q65+ErIBwTJ7eaV5xTHlYok
te5liGK2BvoiS/WxmcU8wRw6jNftQ2ebxIjGg7+3jNYF1NWFB5muySqBvnyyxOPD
EN/Hf5CzX9mGs8YfRhOnFLsBLLp7hnndLE6wDiw4adBaGM0tpKZcnQGcbBVeN0/8
9AtKwCBzfnm8OHT/hzV0az2MBANOZc4ZFwB6EGrE2IKJ+UfOahb7NJ7H4bSFQ/Mc
+90lRfEXpxdZ4cbjbwhLpAwQKIk/9MlhGu8hAAlPAUNuFT/RZr76hePBMycxfNGt
prId4eMTRzXQGwXYF6nD/nN88TrXsOoDKRNSpbBV0auoCk1LgUZi+SRVE+Lf3dlh
QbykPbolm82iJV4VF5LE09buPjgRfFGaoTDqVgLbvIed/KuOOEvoXihx/IkPrm2M
ei3PgcB39pLQYTAPiRpM10UsaIwRR57Hy2Meb9SvDT8iEO2w5OfYDwst+Dij0bU5
P0OyMqSlzpSt5B+QCenahydkA4Egk3gm5hh2vL7RaT/GNGJe3r1HV/4DbEr25+EE
M7uRwrFGNANOqwMXIdUo92dZBMLH4e/SILjlrbmtm1M+Q4aMJMBm1DnecHM4S0Pk
Yew1OId/ja3aOmjscqHJl99JfRbRhMzNikPEDJr4TTeU7Rs+T1lU+pj9sfwDm5mP
HEZv8UcJ7LXH5OIE2k4Qt2OL5z9W9cnzeiMcFgK0AtTOiiOWEAFBvMOXgPKdMWj7
mOptudBKm2ZATH9bUTNblUAbenORTQYx7veW7nwVISmZ+1+kTSoxj4jw9cLF0+t9
pfTyia9Rp/ehQvBgqXNcgOindIdxZb8yjapzAgxqbDo4LjPYqjM62tayeSyzfuMQ
Y7nLmB2YtSi4bbAeFK5xTo+0kYA8Og/YhnZDRaOtLUa+qoA+p8f6gEaJJ4DPIrbG
OQzENp0MEncro0VjwJDjxNaOh6mpx92De5C0SE9Mc5YUuigXq6qXI9sRsw5IKI5Y
nxJf35d11wCTNDXaC1a9SrWpUq+FOq6yBcdlmqmCVM5VwkjKMezM7xw15xoUuuw4
zIu8nyuzwpMam+cpEn0Yn1lU7WopekS76fehsnXfjqvD+9VrOy3/5qmM6LYXs79u
kpbEE4WSFkb0a6It4FZKurqQSdWbqyEh1ZEQcEROW+hDvA1Z6+1TxaLQA0hhPNoH
fNmz2+JEj9Jd++v8DaF6FcP0plAF2HSytp+EnzrtidR8iakzfgtOnEeGIYkXFH72
zPrySAS6Bd1aHkwWkRDsbgPDhXexck3xXRZuQ64l2df2b4QhZYv9CM0cH5xBsTWK
vVuZApMPEY8Wu44GF3x35nk+driQREm5wZJ4LBaxSFx8Vj4NF0+Hy+j8gdWwqTQd
tKiZRQxkcQpbgGoaoBY2e4jBFnws7dGLLotnvyrNCStvJkChoNE4Uzh03RjT0XL4
boj9WZbbDtgohz9L6s+TxeJhuY3zRvDArzdHPxdrUI7pKeXT2rRkcjLJAjy74MiX
9EYLhHRqfISON3gJmsGXYwa5b12mIQ9ZFB77nilu8g0LllAyr4bSRV7jBCVYGdlE
K8I4mP1avKQ9rhr/8Ugq/BjYODA+LMdQOkNrFcrDvVIV6B48NEgsDLi8rYGiAAaV
lHDedirExuzBs5GRjZhhXWIwyaUcyQ5Cfsk0MgTO1XTjE7AtNykQhYbWXTzyk0H9
mv/Uor0qrMh0uBu0Jghf9qguznR7CuJBNDhT6G3eszQHOZyddHgKgsNW0MdcUPzY
2UfHpIVdvaMEy47QVWGLu8hRHxsSNKWMrYA65mxu1gv3hyDqqyh4Aqx0H3GPqtap
iUQ7cik5HupRfrsPliPEU+xZXt4/07QMtnYfktaGHy3q/cRhyM8JD5DVWlD2QDtK
+87rld81FBGJcg9/p5cK04HUprRtcirsnvIcGNpC574cwucBZXicU+fM8+xlZsmq
M8+elB82nQkrohHu2qg8p+qX3Mr59IS3R7k9g3vl2LjbUVCBl9c/9AbBClpnVks1
OHtPy3+HrHzgcUU8IS1sTGdJI8ueRujM9rplJ9jos4MueDaG5ngi8q8BrpefzhdM
5paV5UkeouttvNCdrQmYshkQV/qLzvnXmNPYa4Wiz0/cS0Ga464zb39CSDCk2eS/
g+0Qvwcb5edfMqwME43Pp/kPAreKV7/GgfolHrvDyLDKywgcQtCwmAPnfZ9UDKVZ
yGUdb4vk57JWxiPr/yMN6SFj+Twat3W9HZ+YQGiV6aM0LNfEjr56UnVIlnHW4LYY
FCnk+n1CuRe2uoIsbwZLoBy9ZD0EF6iXWtO3WNcmNkSD1zUAz65UvMG5Vo6wlvyc
br3DPH1x53u+rx8+HBFIkX6yO6nwbSKSfzAWOoQ0Z6BXWRUuSwny7XmzwCo/Q0fq
f+Tbar9EnAei9jAcO6bqQEdLFRRiopmRwaIeytYbZf7nKV+J4fG7ZBdiG1owbr3M
R4WfnuEcAPR9PwPgb+r+ltIse76l/C8bccMAbOTA7Dlhcs95b/ARMk7ASjQhxf3S
z1hnsDqKjTRqlXYz4xLw/+ZQU66hY3V4VbkAMl5NQ4Yim+8zeRSY6io/Tq8LEH3C
1Rhb4qmavSvZMq6QqvjY0wDDkVsIlnUPtgLWs+AoOKPcrRoSPbSX0UoSL3M3essS
qG8Bae7c/uPFug1x/n45InwN0LumlBtEFMhILlT1yhIlhlJe8Y8S4QXRwIK1ssqm
60ZBQycAJORaIEdDzjpRp3gI/vSF7FBWEWZu37uWjZA8/VcokuAHDkmIaf8YpTSw
mc0VLVTkauGsTASUjYGQl0Sff81TFdI7yD0JvYPqgg8YYyHPDp6rEQljIi4ywpNW
edRc/OUFgBukTBoeipooyRvnTaqDtuVRKxXv7J1LDYh118fH3IvJ4dTmF7CPJ7CR
sOukKnRe+RikhSpRrqdDcNQKqBEGp6NTbJMt0F4QQoKDm0mDmd0CGzcq0T9oYNka
Ot26bqW5T+7LZpvYNBG4T+/++NHhKSCuPavRZ95uSkZKy8k8E4wVW8mk31r3g9Qi
DFWhr+ClOK+Rjx8fVgFTso383mQruh03tO92yaDPExcwbhaJSp1LOdKYj6ic0fFE
Dgw0J275Mo+1RRwY42VatJAnB74lCJE5HtOH1ggeSHBzWu2vF3t0RefFEQElJ141
zVjt0DHJb+K1Z1zGZSs/wbgVwwomcoXYfY884dDV7I1QX7h+o3AjPYWiQ4FpZvvE
`pragma protect end_protected
