// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:28 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
drshYzqOKkycIrQRULzSiZMrW/rRbXgjgviPVg+GWs99sN7Drbunhm2s3l2wHu9S
TktSPQQohg18/CDVsj30Fkx1EjrykLwHXbpvu3ZSMhnLHOM/hsYIDmax1TwiVa8u
AqGf0HWE40AyNuMmpVmVky5aiOhVvv/YeNmzI24u4tY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
RfP/YHyX0ZQcgMcnNe/iiH88iUqxGBDX4B8cEe75T0ghybyP4ZxhrGFtp6kHUTr+
xBCENf/RBEeFnDUx8jIgnJgcu9UJVjXMJcpLlOmrteJDJ2pFxehEYFnFEer4PKgx
C50QlFK3oJTHsIdWmobA4Cth1nhmlwPflF4Pezt5Q+u1y6f50Q4vSQ50yQEHr4l5
r0cgBPstq0SRIl60CcF97//PJXLk+aLItxP/iPN+Aq74Q5/+8ove7Vl6lB3TAteb
2cIOfAKX/QDbk4kQBW45aoqoE3+yVRyOIFiNJ2n7Lkz4Okv6OxhHAZ6HDX7m7pDt
2g7mSMzimz1c7vRgA3DmWDL8dNsb4lTEKmHQHtPfPEYufCxY2UI8id+825DbvR37
gSuYElGpR7ddWe7xofR71qRIktN9027R33rSaW6iU/8Uuiw2Ho+4kis0MZqMYMX7
tWCqGx0RRVQkELGrjBNl+9pIJeuGuIzBg2uzCOjCe6nE0CEMthw1FCW+7uoUzfOy
e0cwMIL76UmgNuFsAKROMwIzCvvbtnvK8CUYw5HTGR49a82IPg7wfBfk1KiO7Ypx
bkPmi7SlSMNW42nN9tIkiEqPCEVqh30EDw6WqIOqXaRpGAkgtH0+IoNiAhLWsGxP
iO2JZmLNVS94zb6SoAzxvzxxYXsCt22QE39+cA77PvxXriwDQcz1WnUVt1zExX4b
p4h0TMLaUo6doV5WTr+urRx+xGnAsv1kihN8odo7aC1QAyewv4OzbUSAj5kwAwDl
jHjYOt8wb9CHwkgfGVz6Zs1Iscad4yNaqpqC1D+JrbVAxB0beNKTZ+KuNGhWV/lQ
Ov4j5OjMdEbSaJ/MvYwUE0Eew2DpXTx4R1vNQn4NSIjnuiyoLJLzDYmbX86d0y7u
m9kwnL1nzIQAbp5a3u5fdU3m0q1oV3UMlW+JYRIT/VPIytupR8vABLt5pJdZgWe/
vADcXEDO9cRHgXlsVm71garGqBz+i0wgPakuDN/gZi1zb04UC8VzuJXH2ckS2sh4
BWUFl8/y5L29iOYfUK0U2a07zk6wOCtQgsJHYeJZ4GdoVoy0g4bqXqmlw5DJ+D9w
SqvQXG42hUNHk+0olWiYbRTcJLAEIhXKrAiPWrP1cUC7vwJUCLLOdAoweAfY+GN8
PN2Jw+lmJzBfMafnPN+CzE87pQurcWcbhIaOKnJpNPM10bptx7M6cBf77eQOWPZc
bRfaDRx8SEPxBGUgRMJOOKPaUFDCdyedF9NN8mioKHhjFb72wqealaRQ4UMoHYYV
FQjPTowF7w8gaKz8ohgAiu7y1KDNoI2axpi9fFQIAjxBQ9DKE0lBO8xxGCKsBX1K
NfMHRyBYDsVpqo4IG0wNFQeKJO7kvjEk8l03H6xeifX0TyFiOz30MqarqAuvPMGc
yJCzqSe+Ysvbld0ub0jAwGiJlyoudjBMHwzd2NLD7qSrqqI44YIsAMaKZe1hjj15
616+m0BPW7jpWR8f9bvnz+5Jc3yLTwMyhQFMSchsVk0oSfkxb6hHGz6MzakErSip
rdIzXffhdnL55ieVPOv/iq/SiiPw1UbHH/P/O1LVcsSI3p1Sj/H/ALDYdSf/qTuk
97rBgK6ozkCFo7n96r1kgR9WgSe4+rkw565Pw2SlFljrGRWtlZVq8O8DVfvoXGey
o9+rSy39Q2KgTZB7GsQ7F0WC3DX2hKuiFz8FFnj+2TJFmbubnMh9Q2oWvmyViwpV
DPDx0UilH6Aqz3EClQ4Ra3GRQzisBk/WIKqvdv8LztSWTi8hL9PJGp/IpYo2oaeg
kAkHAkuq8YJY0xPFcq+idjjtrIw6HQdrecf6PdpkSrwoqz5gMhIbc5POTIyvrI3+
gVcL6qxb9i2VsaBwLLKIqj3yF0zCnM0lbAETwFaM2b1/gT07IHsS7B1zJamNPS1Y
AfwZ0+l6qTR7pOjroKhm/2FZUypiJGYqGf0h/XB/nyzSXm7A5kKVmM9hwx1QXFYe
5QsooxXFGfWF7aYlBXUzJQipFZ9huQvao8mkv0mfIiJ7zX7PoniY4mVw5oFpnnX/
u+Ux694ltUfqQri8sIFlFWf+xvnczSyibHuo+pVbuiqzqOOf+ZaOsIt9qtiyCo6U
1N4lEUGQbgFie71QVbpeshX0mRpmYsn3yRKFUn8fkCKWegrROCXW/VRgJ20PyrCE
SHC5nAHdPMug3HebaD98Im1JzKWNk2JRQyAtGYTApm5uOViqReHZtiQbzkpd7rol
MkRly8vEHUS9Xe0E0Z+HztwkgXxYeOlxp/6kcldDNMFu8CGcJZ7EJpMBgA7uIrJe
ZOUpqJE8sksuLbbvUJqHkI10/nNIBeK4EC9nHIsQFbf8TzNeOhW+BvecYr54BL+L
Pad2RkzXAFiZtorMeiOf7+2Y3MEPeWIqXUKLV0o7Wk4/AOQyQh+iB61Kr0w5GwZu
csUImVk41uJD/SULH6Zt2wLEAEPlfNml85/ilSq+zi0x14jAgXH5TcU9oXq2uD/t
WhmGNJqNVm+0N/5H18ya4xzPewdL/2n6q0tTB7/lqGs1cFiy3NgNgfJZSQc1hbz1
5IgnEeTXecwKGNlqIvv2/Zb3FXtLxw+5nHZp+wgq0u5/oxMggBCtYc3dzWZJhr2E
AXXUjyMW6Q3meCb3TODzO5Y3lvvnb4FPJDNzNdrDmU+vFSuc6pYh/0f3G2dvFNQj
O5+Nz1WX/MlDlUvDG8YIuIslPmMlFuJ77KDRx/i1Z4o/3DKlMnQC9wvq1ZQRwxK7
5VEEUUqU0GkhY4rckOiea+RbOQnlxJyZAZaZ07EWQ8TjMbj10DadL+uWM9nMDqeW
mVeHsEjZCvRmIYa+x7PElSuo3Ry6J3i9Ap6bAseADzb9pMSr8MkRGCA2L4R3Nt+e
XENvO6tv/NXHTDdHo/QGeyzIiAuUbUJ5bl824uTF932NYhSFrFBThfwIMhHKd+s6
iNjaJHj5OcQUKYrtoqX9XSXJ1wNCq95zB7YXiOsx3fY9eS2qr1m34kHunxSp9X9n
oa0KumUlJrwmKig5bZJol9Fqe7E3kv051VCp2xlEEbI7n9pQWXU3POvh4WzQZrbf
tfUoeVrKi+JkitZyE5amrAMgccOdYnSIwkOaXYhzkKfQ6q1BGR5HCZJJPPdEBgtO
lcv+e0s4TyqwgKyxhniQa16C3Sloh56svFja+6rLGwIG6tw1WFRk7qugixcsTdsR
RxSrqdj0Pk63CNMK3laABq1zPQZYt8KjVyjjyu1CSxzu62xFhHNaQwFBtkZZbu3B
ButGCfLm7jK7mvKEGmGbSEk/K6o4ohpnMbjXT2WHYIGVYiKeH+bQ0ht4574q7LcE
6K5ESSb0zcFJXQ36VBDJXevTjya1aY8Sl0XtkOmgv+UpMFlOc8pX1tvwnZc+uOGL
pRXZcnHpd8CBN1/KPT0VM/W9MyKQaT527uKkb+iOUSFvZP6rVPLILxgAH5d3lTOF
GF3FR6u841gIgSffWT5k0E7DsiWmXXvmzPmjys5hPlimRd/LETIxoMb0UI8t0VMc
Wz0JhQtcXt5CQeYXhpXJsHt1fZcfuv9WMs7V9R1JtHE27Q+6MA3sQu16D8EVAbps
zmXht01vR+11Pf4irbnR4ICl3X2HRSNuCYx2G2Gamh2Ijrlt1y7Dy+Q/EFQpRzZ5
jUI7HEPSPHnjg82COxebokLcJI93ZYZes7gsMqtvw2eMq2nnC//lNTzqX4KY4yHW
7fNY5WqcNCVE3+C0tSiWWeTT9H1kIe4GiWdZsgEHy3q6ED3HNW6VsxVYu3B3O4nM
7LNyyGa0jdKV1bKGptcWxpBIXmh5wan85PSsEkbLuaQL8Qkue/uu4vFCjd1wQgeh
fKmo4SaFdqXqKfOELGyoIFUxFWH6hgq5d4rOKmRKQvoCh+aHJawQBtL6T7uIj8fH
90xoeJ2xvN0StSV4RIh20ifS2byqopdfgxXo6MAoU62tJakCFYSfWfYdto56D8Kj
goVKNCmh+iSkx04wZqulIXRfkUD7rfbs+RAko7OlJfjVcXpobT7ohvRJrQuUIV+u
jm/X9Ybktfve0x5AkVQ6LwmqcgFWRtVTc8Y0WTDMpSFY+zFRS57NYnPpR+Iy7gEn
bvLadGxz2gud6xRkWZZZ+i9BumpUHvZpsRH0CTJxtmYtqVkY6jkMcNb5RCWkamoB
6rjTGNMLrQYMkOkWoG0cwOt+H7yDOAY8EU+Bv31a5lE5IALc/aqz28ho1WzGurZS
yK1ylow5kUo91noAYvwVr1GXSCmx2+bcc0x9+f58hCDA+17NttZiAAgFjOycbHF7
utnrDSdOfZNbZFt3FXcc7fk4cFN+KCkWNoaDdVB5qt1qasUUJuHOq9i7+9aPSxSg
Thcf52unWLKH0acAPaDWO0bNeg7Q5cZ9GYc+R1CjRUUdncfqVvWu1596nHwyWq75
zBGzLK3boNU2C2Xit9SV+XO2fvFJIWoYGe1l/OrzSVx8GbvHuQNOjKX1y6ejbvX9
KvUX/7FK8+BaT7Ai8jRDIvYlir+zZL4/F0kXhuk8+SKLAS8khD1nEZBL2gOwcP/Y
ZHD3BnBcb75nUUrfG2SsFlnOP4TdMe0n2+Fe7SUIdf4SUdPdPjGP2/Mw7UDrBbyW
4eOIyisYE7lcrc59Q3P+U/nZdRkEgXttYtS56432udf/9fj2BYtxlWr4jGFeyEAd
CPu2DltGmk4WBxm9b9ol/ZnizpcINxn6/70IU8WtAo96eqew4MYk7WU3KWqYuv0w
1axX1MzKTEeF54bkN5QH3hMRxJ4RPXbtHAlFVWdGs0UkIAFDLhXs6gBNcDGfuy1U
qox9EIsn4lIXcdJerJsxtURtJv1kJGJn1WN0CNZPLSJPrzv9JpBoN4vZY5A++UPe
9fjo+EYqJA5s6rGUKao3ywf02L7eiKgyfsnjwkTInVrum8R9jVvbRLb9uIaJOI1e
CGZFsbYnwy1/S4i210lHjlifTTOuITkA7IqDq00E27sLFuGmA7Zn7Vi8eQSqCgtC
mpL6hE45Dh3xkN+By6vySYo45Jl9iW77hWi5QqtEPbJE20mCix86/qmiUy743Vm/
IL6n8qL/r0KldklsNwntw8nruIq6Mo+pKmI/U+UUswXovRLl83GWU7+hxXlY18u+
/8eH5PUMIOex81fkYj9AKoOx08eYcIgZ4lU9ELIoPsZ06iWYTERWd9lRqO6pZnvb
HMytSqfG8hREZIn7NaBKX3jT9SrJ/Bmj5/BRm9pFz8FNVrU9HCFJ1XZDiZU0g7de
0uzkCE63sUVoQ/Fy9nfWyQY+jYqEqydT+VdIzYCWEie9xLEU0N0o08iScIMBERPJ
35S4ULKVMSn8wz1oUqlpGbXWUQMHAji9YIgtF9ONc2GH65amG34twxhwx4HvDrFa
v54vgV8+xjZRXw1/3x407xjKQsnQAZIY/NJpvkMpranHwI8ntF3/MJQfaVXfhU0d
acix+jpT/d3hLsUACZBGf4XihaBfI5GJ6rVmoWinvNGf9lEalshgtM3XyikuVpxW
7JlxfC5U7mC6fXK+gQUQTz4UEobnBuc0dw9to28zelaQiTNp1VxKqtBMFQgumQ5n
Y0P2SHowVNgRZUTTiNSte2RTUq8BtUmKvV5ynOdWbZpiM986LSzr8W2I8EMM555i
vMg0AbFSg528IJTdSSaPv38IcSsGZnVNsneMQslko86F599Q7sOkPJkovDlcx6VO
ekEkFrh0KgXkjJVzIAffRanJ6bhV9DbmJsMwQBqUeD07YHplalgg4JggFUAvFWQq
9Z5QbTih0n5ORlKbmTRY7VlqWnIK4Mx4y0++UtouxvEURlCnQ1X7vwBuXGWv3UOn
vN3IZxqB3vMsCy/o0q7pQYEXZbHZGp+nN3+ezrwlAXd2xxB65TjN79XKsqZjAQN7
FYA9VA0cgZI3l5KTARgL1p7eZuZEUc8Sx471SWAhNHIFJjwrbyKz4MCZD1+n255c
fOfys3NKqCWsGgCRHztB727cY8THzFLbNCLnLr4DySmyKldsIFRGIV/mizyYCQnx
tUiIdm2TJPrLisGQNZE+pyG95WbbuwlbhzCB82VDcdFwU1e+uYXXlktywO9bM/KJ
TG88+4OlfSysL4nWUX+h10KZBQms/ob24xpZxVOnFCvB2oILO7dxrUKlCdtfX9UO
MhMa5cdG2kR0jLgt2cKmkUAD47T3hjO8AlOxz01lvwPHU50kaxDenEylv8jeeQrF
433i7VfMiL0gkrOLeAeHOr84c8ie2FGV7rh0uaqe+2uUaLBUdMOKJAXex24Ai8WI
bwRp0NYq5mnNX1GPel9epoY3KF5+5knL3QG+RuzwakFmaNPrJPFtJS9Wj2u1I6eg
vpAtnrFFQqzH7RCR6yR7e3e9o1wIjwYqO+/TlGLmJvnJrWklX3u0ywSeauhrOf0+
SUnivqeX3riYO+QV+wbEWhQrFbsVImtOy5U2APLBwMoQCVp4YKu9kiTQaRZLi4yL
iuKnGUM3/nvDC4cWgL3SNJdFpR3UlKBxGhut0cRW6h0AvQMUVVcfFGISKOf5BnAM
/WxcX/DX5A9oF/P78JnTl3TWXYUMC77ZLbrzk+WxG/Bv4NmCGEGWUCC6I6907s1K
PrL6wzxvPZwlclrr82EFGOcGUIIVRIDFplbUqdH82Agao3K+Ezws+zgj46dJUWmh
mfVr5ghYwIIMWs6mwzJGfc/qvDOe17REyXYG2kxZFLsD3fzHTR97dWCJYseyWNGY
UezPg9BdqB1QjSYzG/G3LFHRn1/PKq7hz7fUdxvpCGpR9fWR5+iBe/el2x54AmNn
t22RHXWgUhTT262b9TAJLsQCXZTar9X93nASuud8U5jbCHIZ72M+vujxxanM+IE4
lxWIlE3myyCVhlbQ4tEFYo6UULkPkaPTTIZY2QD6rP74It08nQ6bZZ8M+67upQFh
o5mc0qw+Vy1Qx+H1fSbDiW+1bU5nWNWsRU3lN/GpW1j9gmJp6vofbMs9FNoz080r
ZMFXONV0ZOV4EGYAlQZ1RQsqNSgBeyipGvWBnRUHdciAPEPAOzC9O4XKTywpVXXK
H00xxKNxGbZZsqRFMB+yKJRAnxd+85r2vicLx44EgGm8RdlMSRhNVfml7HtlU5n0
R0bjxRdcZ3mJsVPhiqMfIJoEgqwv4nEmbSxqjPmkthkFs7ISAV3pjdSBMqQCbHJ7
NwIkZa2xOQUyhY0pRZS7ZL8cAh9lLL2xCr3PX7POtvnW+cgBP4tiX3Me8tWnC34O
qbnONObjeEFZM70INWM73ranY8P/GcZPTr7npTPJ2YjQyNuAevQ/PCCfFkKkmhGp
cdQI1MnTxQjLh4b2zWE1i69aCs+drC1oaUb3z2eU3GOLLL22GcF49a75y9ZQgJqi
QxJZRlK1kA8jd4sqpc1vBAwn3nK9P9OAtJ1RCNZakU+MJejSDLW0AuIOQnZX5g8A
ayAg+6LHrGHM7ktV2dAcnRgawt7Dp5lh/A+PBwesvT4wwm0Tleg/s9ZZO7hKY2GZ
r9yIPvyYG6gOzoRUsN/racalIdeR8G3OUE5lNmEMNVtsWQ5K6h/XTPIdzsM7MFeB
LnWgS2tA3h7MTeq5xDxUigYjSrJ01fY4oeF9kXIisE9fHiU7igYNGHjDNUFRmJJw
mwbozCDbJ1C7ZVLqIEKTzpouy29hYAqDV62wE8tp/LQwJNCDNRToOYy4SE8GDwxL
2BCyeknCq7N68KxPWOe+LmcNum2T38NFmvzUD3/9qCZ8vAYLZ02RNowV75NzNPMk
/5kOaxR/IDhvDw3i/kI5jclNONZKQjGudedudMFL+TLwu2BW2SYEzuewqZSE/M+d
OZFtNlk17pAzj47WNJMoD2RiUwv5usqWMS5ZDiS0edamFncZWZk1QqQIiTSxSPop
J62MUJIiXxN9hCcVFUEFAig+5MhKlo3NSMocWXLPT9xxUKd101L/ziGUekWVGxwF
HbKUMFZqjtAPCZAU9Fv9GUcFS9OrAEDIq26UPzmvqrBNorrgUfCrowMY1gFW802S
ZY2U5ZaGH68QGXI7k5PVkZkFKtlgkFnxnmXtFw2gnJJnU2fy7sXAUpNrgFqezlo5
NZo5dZSFlVVDn4Ua93Paxpc3weF0LSD27UGrSmpK1VS8ztjKOrGZPf2m0528akrR
IOT7bcY5a7+E9d/VeyFEw+7g264U86pWzDC7ylaTMAopEqjoiSmrEj+gihpkj0ds
6eLRhtaJv78YPIAsDHTq4jB13IqiaKm2w4Au0BGVX6rLEd6PGs1v8G5vAzX3tq3R
97HEg3XubPR+ZuiYCbcRTqu/3R+JTep/y38BzIwmN73LwxTeXUFbMo7R461EHKHC
A6Quh/ibWe6SC+ggCstQlaDCwGOS8YwA62AYKoXYSRtzi/DRzW0hNDRSpKfZzE7G
3QkE8kRV/8FAFFS693oepR7IVuBEthRPhvz2p+G5IzCAVmRZji+jALJvROFRA37p
CHwQ5zpfjQ4c+LOIZB719L9Q1HIxGo0f9Heuqe1dcXscQ3l3Sn5ABU84f69Uti8k
zF6Jchmj6zsnxbEku8wTxg8SkzT5DFmhfvNAIpieYA3AFRrjt/d7lEExddHGH7D0
hBXe7Th9Y2tEMUkv4z8yjPh4DrY30yoOP6507AYrNMDaRrdSze6aLrVFXzjLNoI2
huuibt8IsMIGGrAaWBd1YHIzj0Gw4FnMNO8NU75UM4XZHEmyFqRlHC1c7zRE7yX2
NyaFu8Zml9wg0JGmICnTnAVqkm9s7imGJeK4Z8KOUMYdsrBIyVmuPYAK75/8FAsy
wrpvlkZDHRAlcIL2C2ePaKQKC1FVme2WfYui5khxpJPuDhvjncZCe1Hn5N2LJHDK
vNIohyJLfAeDZ7TUBQiIqraskV3xQbhin6aX26ftG0k5uHcfpGm/5jA1m74uNtLc
JgGD71xYOVuHM2SaafoFX9xHpHM+qbhO5L95ROCroRSgiLZARuDiHep0m56GAHd5
c2aFaBU1biiyMmyK8gW+vd+m9PcDusWelPmy1VQpR/jXuyfT3bqZBtwnEkFrsCQF
YiSU34O+ZWAsJDT5JjlQJ6WpuwN3QVAxrfUrmOmiKwNVRwrn0l1MeNLuwElXzqLG
NSTvACWsjikvI/4aofGRNmpcRGVKGh/fIBe++fHQIFMdlnYeEXKValKG1VGbLULt
aRRnhx9c8DZCReY0DXp7cdKiUcvhexKGr/knCmJy6CHpbnWu7aycSTOtx1bcJdDt
7fsvHjl1pg/9WyAFug7+uafjZRjtcaGaq62+POIF9bPWmhFsQc63Qio4rL904GrV
QtSEUzkfvTXD6oRRy0Zdq99h2VtbXpEXbHQDIRCMmByDo4/R5X+DsWqB22afUtEN
y0DtealLHUaDxPJxna+JE+MmvPLBpwShzLHcoK7d2sROl1pJRakcFHIydusblOwe
PHp4U3QMT3RIA1+hbz5CwHwEuQ8uUjlzlyhzrvILI/Y2U52hPAsTWN82DSkjhnbD
pHFJlWHYAvJZE2VWzD3RKVEPk2+FQDfckG37VMHQ2er57j3mDybKieof0WpqKT/K
Am3SzsZ6kKsyU5PgEM5OEcz1EVNxu3xUmc3Au8v4dHJN8kaamORfsYUg5awyxt9W
xd8u75Hn1RNSzRzDm3th5MWg5xNovRjxBln9JoR+SgTB41Qk0T9iItorvdKHIprk
uCwMF2B4190TsQ8ybFoZ+L/gddU8IBoyKcgPJKIBs+QuPChESaZQOIla81q3it4/
xbSoKNhsN7vdTvxy4qpc0g6Jtd8nFGufcqn6mdtYZ3z6gx0cau9qFUv28tMvAz7f
Sfj8BHdHYl05cKQOmbKjkjgahFzb6GHoODI8zc3rah5rIpB0EdHSf1HgiMnefvyu
nZQPVtYFfVOS/FXIuoXjWWLi3t5AtziejTZOSeO9E5u+X9WgAtiNHMYfRT6ZYOvL
fKTCji6kwcGn9WYuLPjlGBdRp4kf5ka2mYksPAnvNabilNSBHqC5fmypXrT+zg74
6AtYOOnHq6rsdH5rTVt4pah/TuBw07kIUR75Lqs69rkRtBiKYs8WRcLQNd5T8Jzq
75uGXx/3i5DcnyD5Q0Y3dlcglw8N4aSIP/jz98M/IYhq97EOtGjaGUXNwuQLGt/D
4c2wUfpcz3yHXxK62a0/1J+nKn76UsncWunQ6HEXrgEAxQaQHv0m4GV8IShZpr+E
Wu8Dp6HEfsIKC8Gp+l6nxWoYoi2AG8+JVwK35//Xpa5kvdJ6o5QwT31tkN1zB8T+
TRgy57G4pyEMLaMSHQu58cmaqGttyHTKCmfO2bdvHnohfHr963xhpYbOJg4pEJm9
daHn2dLVWrH4W2LfgqRLQI7pi/fRm088sXX2WNymNRW1zmY5XD3xzmGj2VvxH13g
Ut234lZQ7mMevgK51CwXxj5Om4sgVJu/ii10JBsF/A0CwVc3m3rHtH3aX+jyao3i
906RgHMaePm88zmRa6LSFSR4AkwwhrPHctgPR2JuJBLBZ4Zj+S+aFTEYQnMXyNeT
qrKdqaytqS90bm9hHo6ZHwXafxpNHWaK766+qKZDT/txZjyAPz54ZB3MUquYeJKR
xdXETRvl6k3FvOX2artNYbk/kknsr18A+cBli6F08Rpeju50TdsnENZmJ1WmWOym
xYeVS5fgSyqQd/cXPYnz+UmGQKHq9UkU7qhadrJ/U6s1Go7zxwzRYh30atI/CFI9
WhIzHOvgB1VUEEpb5A8knvbHv0M1ZSqgEobGFT6F/4sSmEYl7ZMxoLGayYQnCE0y
G5pRQEaNrl4flM7NjfeUpnZzmmaYy/U9xpSrl/g+mkGCFYY/kxHzPB2h6vHRVSnr
GVz/PFfimRLPxfOvaNN3yi3z8raIPj0Yll8l012TJL6x6eGegc6YDb2XW1u9tE2G
HjfJ2N0oV1ERQO/3R/4toMBSS7STy9uBevCSzRHHufDAdnBtmxecUhkhSyyE7Mj2
I6I6A5N5rqTdDCYZiVnE/MoNc/HbeQS1j4aGYugxHguNaTfwvBKFxmqxMsTF3f23
S/7rpOyPFHw5KP5HtAPTFL/qSm/lFn90Wi0KE+mvn6gqPqHYIrLT6PQNju40tePq
fhk/TLxp0//t2UemEtAKZzY9CQwMlptBuv1A3AF7KYymc8mRyq0KFUtw0vtgG2h1
KoLe9x3vPsHEx2PuqsnStGlJfzqiJH+Z7/jecldkuuR8tNzo0hs7Mf98ciTJgmtu
aAaroNE/u69fBwAgwN5bFLH6D++6tmcGdXiARq0lCxySy5WXoATguoC+KuOc3tLX
p7a9STMUQwkUFIjqPEPyh8rbw6x5bxmoTUtR4JJMHQmMjlfYVAlrQuUchh5B3ch1
1JD5oIadsDcYJuzBx/nKluKquejKNM/ymyI6mV38bY65GJ5IMjsDLljLv42LGYSC
EBURprfxBP0rN8/VkJNQKspsE2RQ7Ysct90e+UAJ4vgtJO+6j8NnU8McAKt4TvJ5
DYjFVYtJF6/KOmqH/E1UOonV3KsgwjytVUilrxsr7kyWg7PWXkzKGs58gax+kicp
fKXyeu3KK4fKv6ZKza4neHilQttc4FvmneRBsOL8CtrbNM6HrgTbv7Bwu+Y0tPyW
5FsCh4FV8khL2NKiwpGLcX/RlDtFB+J4qV+Tn+yg5ja3ZIir/RqBBp+1tWs7+zMA
5GgPKwSTzgsgLc7mYuttg6UVeI6NUO27LfKoa1MOivPCXcnGqRhbbeG78tdKNmOo
kk8zfqQVj5WWQvgMm29O3slildhPy+e3b/gWXkwKLVJkVNZrYES30wUV5W0iJp5d
vlkFJ54JORMik+by5yP+xXHsdxwtcjBdcDhGkDopTxZertN4saoUazUzFbhNu1Xn
OejRKYad0AjudusBx/YB+ktlrPVlQNd4LcHduDGNfXoRSrhE7too6eISAYlhzP8z
P3ORJU4Aao32siSUj/mgKny5axnBYlzea+O8JBqZL2qdZ6C++W7GY5sJytB+izKE
Mnib+PpWO4OfJgZVrAvd/3Nezwir27qmT+8VqMK6HjarwAEHRB9q8LDZD3fjEaPE
lNUZyg3nWdu19h/sR5hg+2CTCzr4iTbnNK0MXuu6Vt28XHn4IfLnNCQbBHhk5DmS
7u5hVdYo6dZDISrT5aZSt1YcaaemGcBS22cSgVuc9BI9O4speTXn2+r1vKpQCFkB
owcpPELTnafImtU3PD7Xku6Rsow7BpW3rrM9WJDVmzyNwoXb+p6RUXx/L30NrVEk
QQ4TQBv+/87QjeJoSvkHw5WsuPhdYlaxBeNiAHAJyUVuQSTUJASh3WwtLw4u2/J8
GsHGXYqUpO2F9gzqgGOx6klz/3oaHuyTYeyvzY7BrZ3XF7YhUdy1FiR93nVFRpAO
3ymuzpPMfyYb20hdoad1iyu1S5C+IDoQYV8hun4h0X1hRuVYr0jzjgH7s5DMqmhP
C7duS0zYR23caX5OXUz9EzoAQXhyT6THVWxbOCokbLGS7IU0/pYsf3NqCMSCOeSZ
uP52wX2wBHCv9xz3RHM2m9QmwKdy0mwrKOJprYvdB8zwFjwmuIR2jQYBWwXBXDYQ
4bNGdrAGD9LFhWcJcxoqQgQDHKR+6TKuajXAgz4fTsndWnXRE73zmLKBdLSSuGyy
0/iqmXWXfN9otq0G/u179p40A67YMJcNDO8KZnXaZCL+VCIwpcfhwoHTUZ7pzH7S
wFyJ/1/G1c7jJYXmhYRWwGAc9rijN8NkX1UZe4E2Z/N8ucU3Sy6NYXj8NJPqs4Y0
Z60UPiD+Ii3BPmlM9VN9NNHYD4jdWj3uu36zD55O56D9nIOG7xVBW7SvfmefekLc
PgX/EojUH2EJ/3Mj34WaDRadB6Qh5BK8lHV9G05fGeKOa5O/ipgnZEe2yIE4qID8
NessuJHCg4u+UgX7Br7NnpDYDDyj6OxYKzZix4iCBmFMdk6s7l4wRnzyIKRxlZQ0
WXEJrBi7t8vPWaZb1U0nELwCrraENL1KIXRPsCnKxznL+aeYGBpiP3SXQM4pDgbN
yIJCa5rJl+jKEhmj2LaS25s3As6Be45EdWkzNmLEoDpYHItHwCDivCUDjZ+dOCuJ
SXsRTm7CjiRejLyUOKJEws0BuKc5H8QfIe3BJweM6tWYEueOw09ysGui8xqWhj+G
3T4beZNnkIYQIx3cDzJBaumIQulDMtNqf1IyBT7v5WO3lJzF4EA9wsuTzU3UHzU2
ppjfF0HaqQ7QFbv4lxhTk6UIQqJlsFsvj2W97lded3vFqdDaNh3cIMkMhWOSX/EO
adNKuOVqPozOvududfsZlBnOOJgx9yBwiBKX26h8kS1fWt/D6L021ItzQ7yWKh3c
H6i16dX4i1eN6zPi2PPctYE0CQ5WzmqDcvraZ5zBK+XiKzOBYfh7I6A60B3VgJoC
5osHf0xj0a88P+joYzp9gP2kBF2Xc8p1t+jZyPePbpoDE75tFsSfVB972BwcoFEw
Bq0DzEXAK0r+4Yn91jczxfJMQjT78tO+xtOA/QP+Q6hJvjWzWL+VcC7+VrbX9VT6
vAcggW9924xEjh9VBF9bavylfh+a+YVZEklG3NLpnazN5Ttkb9wfyY7E5IQjBqlL
hQ0dExaAo93V5pECo5+gZIfrx/XHE79QegldD70/lHUY/18murgZdQcEOtF/9I/R
SJBmPh8r0gsEdLd7NH0J9fBMAls8zosTjmFfhKotBq5kUgQzUUAKgJDnVgzJvMZW
Olz+HkBu0UXqUjeRLepveL6wx05CZHH9Fb3cXFAVy4C2pN2oQAVOoy7o4hYHxn88
DsiatNKSgLSJitRwrhnCcPQEM0qIImOGugMJ7Sl4UKxNX+BeBH/S45Maw4cUli+p
8QXf21Yv1S6EdrO+Tm7VlGnVQfr529OwkqUl6zg6IeTLmgWyCaJshkjokDaUwxwd
2F/KY2v/z2z2WC3Hz3Mj6W98ZNgmZIaBZRSjaI1pm3WGXjWwSX27UdvvuS0t4ggu
I2tv9m/AA84IdLenDGaQ/HWSwzp1Ot+RCgQexYsEnyGFCiXOfH+CTYnYkhUgasMP
5V1BlPP7n/zlPei/Umm/08+yWb0fELdPlO9mvfMJg1W7rTYS11xCdgFPxq/UtWXW
lFEjk8h8u05SwUzYl4CsJ69sAvrJh6W80UwEHaVEQ6/oeFQKCznJbfqVbiDe6tyB
iBaFO6n2RrjQVdONnG0KySbNo71ywubaRSlJt92GrZAWOxIYs/M9m75swrg5apT2
13kh8MU8G5ik78hcrP9CgIU3qGY1Y+ZFWMElkurSiIM6Mcux7pJSPvXEmg2HOfnF
Ti+sIjRKhnd32ToNa7MVnkO66e3RP+YkvGMmPq2wrlf7RYHx5ZFkzKB1ANd1GTPa
EAisqnqeCkPRwvujg6httqzLDH6mX6+6pFbkeiJueLJFzQu2BMHz+GbwoxlFEQri
ghd/Ww4QukIzrvFd+j0Y3jN0HKsDuTXRYJkiqorY7TYXyfDU/qnf51+dIeyL2iYY
rSMfDLCgxSHViEYh8+tJaNtg3SufXs9qOuTpRo/hZ26BzY2E3qZQsxdr7x1ZctXp
U5xieyPsZJoGdUnF6Mk2h8wqyv+lMk5+5ESqFLDH84xrSeGm7FNrXr7jadPQrUK7
IcNqD/TKXknGTsLKAXSfxm8oLTBs0niw/7coyqtLYUaBy/s69Y5yFwDzmbYV5cN1
6j5KGxMeYDkTL39aBUpuEGbBQf7Ezu7C40S3x0kBFXfZNm9ZLTpTlhuBn/7TfWWS
0hIWsU2NhnYJKYw4ZeSNpYP4AFYW674PPiP3Hi6OHpmIqPXTFiF0da0depCuRzpD
/FU7/jrMgiI+9dNWBiQEynCs3E5RrVRD0P5Hr7qevZ27ujMpWi2s7acHVCkt2gxK
A0ktZ7xyoPY2yhX8z7SEmDlR/B8mgEL/O6BNMbx+5I4T9pt8wt7J6jyzrPrjSAvg
Uh1pg0AxG9dMJr1TqgxyklnvzSCuOyD7E7ePb1HtMAPh6IyZxV4qUdVp2N5Bp8Im
XkvJPIUC7xWG3sy1KI6fbifsr90niIURWZ1gcopZgmW1dFURID3j0pWaXtnu2z6S
S2VFrWsZB92xeujWNc8GIjQOZds7R5TGBsgOm3l9lqF4oSM1M0JFycWaHvqFohBX
KJTl616N9c0CKoRLtEiysXZ1wKQnXkYbfZIquC34ZHTcIauGLhBaa+jqGd5vzdH9
Fh8KCmv5kPsd2z/gZmkNsFMibHmDCL5MMseb5q6qlSkQL1/bmW6nAETD9R7Qo7Jo
ArvzRFZcX1pyiK0PxbcZKTFIrH/qMNwCUEsHIqpHFoXt5xIYwxFdM/SryfWV1pFB
0PzpMceo0+fmtrq9VO356uYNNYah3vICYf4VoInD0UELEiylz1qnfw5KRmPNBtu9
mJeCcTYyPKt0vumDa9JGQombd+Lf14uJmtPs9iRpOJT5+9CJ7oYCSZr0CDtyD0YO
5fC1tCiYjzYZhazOG9mQUWTChftlcczcHAiRl0ODcOg8W5rXairQ8kMtYaQ+huMe
stJNnPvJ3R9J0IjWSDKBM5UY3CxZn5tv0qVTOF7xPVdRhctRycSVwA4qD0SZ/eo3
HtEjrv4BdIPahBh+LLNvO9NYH9InXTiDgtr8f/j/NBu0glEab3I67h+S28xLmPGu
lLAcMcyRcQa3fLd763TYFoE5DnbBgeWwSbSq+j58WIeGh1lR10Zy9elF2kbPheCT
e99GWsj6kRoAfG+sB/EEezlX0m935fX9ZagEEbNro8+ZvLQwJyIDZWVUfN4W1rV1
PkZ1RVkfhbnKiaUuNKK6Bno0Bpwg4EseHE43htt32+BDMB5SF+LwM5BjVDyt/lRQ
NqlMpNZO24F9Y3cXhvWpiH/BKAceAkgWLFxKcsDCIFmNEQJUaKcWbnLVJ6uIRQ3s
JliZT4e8V6IARyqQFKehkBtavKvj/1Ri4K5IHuehwiegIPaFnJzLAndJFGlkPqH3
DPWA2K6xh4x+sJdBQmM84tzr1dUBvDqUvGtO+qfQRqwIvF7i06Mt2Rg3czS5kSX6
a6m0HYktt47mAT7h2K7ERskZari+LUEa4YWK78DwtdiJpZXyjlJEdmTCNCpd23Xf
hg9q5XGUPYmlUZsjsC+V6J0cqilj6uQ2FCEyi3ZH4cjNa9jVD1j9k6FH795vG90D
rkeMlmrTeToL0UmjD5ySnUuImcROe3X+jpqC80SLmC7u0fMiFyD7w2rRwlkipv7P
Xujcj2+nLj+HAoKDty6JUbBmpHOWuTAUvzldLEZkAt38mdTrwzIQEWOnvowiFAEq
6eG+l7IBjepFRNSkodrhttbtI6AqtoowMPIjBMwSl6eQIK6kk3Dfjj/ASqpDHXZw
W8oUV1VwOuC8AjYmAVwEL2s1taRcg8IP9DVd2jgYIKr8n+OrT2BL71YbGo7/di34
OsG7f35xfBuaVBECNM9+fezRfRFaSekqGLvSNxrCn8kICU1Cux6MSdImf/7HiOim
QqxO+dE0DUZD+H8rqJR6BqPcjgHLDAjBvMLXXRLYy1ZOSJtJI2w4wEBUDiCt0ST3
euAWRKswLjFGQzmVix6dqwEb4DXsPsDnwfhF4fX9q67PhtTnx+Pb99LMuVcfZptW
JpE8DO+jVrvPwqc1vUvHrljgaCg61jBjFRAy3UagDfZiQSySgnlf7UBbYgqNsRSX
MnbzYhsnOc99iNZ5bMkmZMajq61BT1QGGw6fDb7m5fjRvG8jc4JXpPzW1XyO0e7S
/M1Y76quBwVI97/NZsw0a91WlTV7m0pLTbJ7eUmoy0enWndSM5zfEyvJVPsEpVkk
sPem9N3VwgdRuZi4wb6BIX5PJ4Ho4zYwxv6fpwvsTmofGkpiXSGaGB0LH/CoJBGo
G5Poxwpsen8AJyaKsCT3A6bcs2x3Pz8FYBJAmRQmNNCHBNankQkFRIltN3iZtRwC
lShsx1gGN9HZE/HopQgyhygKiT5WAd0oj+Lzrng7y/PUkj5PWQFrM0R1TnTdGtU2
GLmLMDsFnqv+11YdZ4iXRDJxDb7eKnwDf5id9j4kpM5aE0T03MEIblTIAQRKURB3
tJ6aikIwRHit4zZKf97nmonL0fZUJQHLuvqOjhHTGQ4wYIVbw6NY0ZuaWFCXpIAF
4HYBi1jWoLues7AbayrU0mMwQRFcDEBKuncS61FC/gbCG0aU7PzOD/KBgETuaP+S
JCbOAb25N6i8sN5eYvFtVQ0hpPn/uc+7U6uIZMsO5Z2x9uomZzhoidEI2XnCIf4F
Np/sVR8ozMsWn/mpxh9fN6cI3q8KOC2gk8Bjar+O3kPcDYf0AdT/pZXdf7OvIim5
Ia3cYPrHAztJuOsJPeikVft0TpVXIvJajX55RTqyAlxJvfyyFUKyCNfQlCjv2SDg
uN55TIvRMGK5Fx8Fdxl0EoJHzUW8b6h3plZlqe1ki+P/1lMeyQEQoqxmX+BMqh5n
xZhCJ1oSagRcFwq7SIPBmxp+2MNWf7aN/Ti0g9y6WtsaIurgvWupYfbHgTzKKdFD
9nwf2T4PUxPDZjzmPblsuxKi1JtJAfbfhfPr9mYdhQ75oTd7TQeHu9vvP90FVGHJ
4E4V3W9prpfVaVAwGr54PnrCa2Kovx+2BityoVnLe5p3Nj5oS6hVPDkSPBZFmYOV
Wh1Xqk1VFux9Vv0i9jb5P8MVM1ZjK5qPWA4V8IRpRi59mQuHZ3286jk90R/nvi7I
oaFx7MYLQneQTg3OqmKfj6SEftE8+Jvu/8OlPSfIrMbMNXLYoBCkSFFD6IuoGayl
Oo9TO2DqVBpi6Ag2Okjbrj19xgODB5hmmgFfXQKdG/U0/XglBpV2DN4A7O0dFC4i
`pragma protect end_protected
