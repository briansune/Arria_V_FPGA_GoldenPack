// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:20 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qrio2+/qvEd0BNHVKn0oyuYEgbgpGDKJeTARfWlAYvuCRefG/rgF+MSfHMEC8ahR
5ggUX49CqK49BQjGOjlfrCe6YNBeXbRGgdiS90HqT4qXHcmYc2Frxif8rueZ0kW/
2hnS3CqQkwBUBYAGw1vXLkijR9L7LdtX/WuAaOWFVYQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
6MWOpRe80zTOUwfp/KTsBWTjNu5TzWX935Vab/afM3DQkpYlneFMHnzt3Ieg0Y8G
someTlkHZPI0ew7+WKWMywtiKV36XVZ/1OZ2ER3/P0prNzmIvqDL48BG7Q1pC7MP
Mrjg2693EbWidg/37GAdlpqPfPJWqahX2wilL7MnexlVlvrQUZs76XAD84OEGaqY
kjOGaVZ38N3M+dvyWmTvBlVtwbNjqHmJNMzLe60cWZyn6t1cGsHtlwYQrUkTncq4
ws8KL4y7KNEss/8C22idvWbUQv/NO/wFc4ZkZx0hZtgejoMFW/ylQ8svx2smtuzy
cdKOGUD9ALJdvewWJnAKeV+d6rBHbaaddKsFEr4LN6tkp6nljOLp0sC+i9L4099x
EVjhzEERYWswqh1OXrffD640//mm7BZmokkfVnm+GOWkkA14mSNPgJwaCEflkADY
Ve6GiWWjs6D7vE2WkSK84UQbW0ukyG4D1+c647D76KK94PQVOVjGjJo1TgDU/Nca
TL9RxCpErh1bbEOERK/1Vob2bAHgJqnCQUrMJ79zpa1cFU+UOoLHEcfN+He0zkd/
UR1rH5W+fzFnwbwBYbXJHkVgOAeI9EnLXhJbPkFwQAwG/CPYdBEUCUx0TnYyy00D
TBNqf+g4QKuBcwQ3vmVRl6+a/DKjKKGcV/HbNlJWZaKliTzUponwh0Jql3+DK4UD
x+f4ByTaPPepLpooZW5PfB8iMMc3KLRH/gjwE8j8mOK3XJ4ubwGOLBZ60ekDO9Br
dz1dBrcYCTtMLuazrEKLqlKat9r5gC+IDW6lZ+saCQHxlNe6CANSESKXe6G3WiS7
ZuegGJkHzF8dTLFaQdgFK2BPeMAAKRKHjM++uQkk28gLGrvKICEKb+GsxHakK+nh
nuNSvfM2cyJCm1qQmf3zhVwsiYbPN6fIWZvMgWdWetwWqiS9kC73GJvQTPVDR6sI
vU9gzccxAKFx7xQKfRXqGUxdovvcl0neekMpCsq4UNqnqXJHNiCZqwelk1PX/Iv1
p98KFmarO5wyj7Ksrurzn3U2R1rh09mWRh02w6rtZf6WYcMSlBurEvRqeyxs1T8k
uwhgpQnk1rbJCsKI1dGnTg/i1o0HBac53dHku9lz3MJDVZTgweM14O818LmqztYF
6GxeGpPe6xfUVJFq/pqqukN+qASJ4i+R85J1XJRKioDx7Pw0raOO0e2sqvflK7Gc
mKqWEU6HiY+r2hZT0bTklUSbMntJIKcrfSG5teHawI03YUbbV/hZ3WAVSeVkcB01
rNs9Gl1NqNxsLFDkn0WNgW2mwQNSZR/nW1z4Ff7Tq9bp8KzHpkugCZ30ivj0tgRs
pZgB3tXU+5npUR8s0lT1l/3S4H1TSisf3wVjgE6x9Bks4mTVwB9pLPNCqK/VUGw6
8yjLWIpgUrkARH9Pd/dWGSdisK6uMkW+RvyTQM1YB45Tid6PhCws9V5PMtZi/kbM
2bYG2n+dxHjbGdMZLEPYsMn48nU4FhIqIJDkjQ3TfMXgVB0StDOGjRCfIAzTFyhW
63gtwYOH6e6DLi1YJFSp1OaY9uBxusR/i5NQN+AUJPdz9FTN5SA0edvmGoPt8Wdi
lW2hidBX6Q5/2SzOKeKRHoqu1I0pgojSCfld+MmEw/2uM2Lz+ZHnTvffxACLxYS4
YBaBYyIKcJxShaiDHVosrsxRMiMiGhTHvoR0u+mX29Onz3gMj2lagyvBS8uPRAQ3
f44LHFHC+zpHZIod3LTV4QUf8CtyCVPxDA/AtQyjgBTGWiIUvk+S3oIGp2Vr91WU
yCLu/Q+rpfoP5gXkKTUViYuKQszZEw0iD3Kfbz1IFPTUu7TJuiN8JQ5/bymZWn/B
PHVd0djQ/cJwSQPkyU00oZv4ocj/1OfRT0tNVg15CqTMilhnl8OZHnmOOGqnPUNf
UZna//sspIEbcv8VwdT26d2Q8GyzoqPBk6kZ0W2S2igdCeFlWe7YSM8imbTcr8A2
CjH8n/1DNLB6AKBWZ6PLEF3i5fwMvxwt3kGOSJZYWF+qoQ38WUMYKTnomEMHNgoL
6SxkIQvHtLH8CmvGHPF5c9B6CkYeZ2S0QLx9yNmyXZ/xJGQT/J1w9tV1WJMfBRch
OXm/XrEgxdeyZJMJ0SShUG5HxMEjhqpO7cxq5IjJkfVsFI54sdr7l+KvDRcBGime
LnlXZ7rwqkh0McSVxh3SqWPAV2RoqGUwUWYn+IMd/thOc6JkzQ+blNFmsTAN+QL5
Yaq0YYLZVEEjPAZLwmSNCS1TIbjrsrLweW+lUMlgtF8x2+ceg973fkGuGtQoZ24o
Rz/+qN5CwjrXTiP+DV/bsoj5nTAPU0n588EO95YYMouEmKZFX7eamCyFe15YMMHT
YHYg7vSEsA4g3ZtQX6+eGT/LSEtL84APvcEwhqT+pYx3giQ+3ra/ecEPV2NRcRTv
+AtczMmhwcSGcAsgmWI+JumRhWqT8ZGo7O3V2j34UbfIHUU1Nm26rB9TdsFxglAA
IRVwq9J9PJGKCaSd+8J63Q9zeI0gJAMtksZe4Wvu1dA13AnNiYkhnuVlTqU+in8C
qRnqXKBaiiYIjd3Io0ulR/4m2Ias/hx0pPcMFu5WenViEb1rC5vEpEKlWNRNclRB
opjRYZyXI4+Ut7OfYuLsdfMmVpg+qGP69x0kZviqE2OqGGm/8xQduF/Up1VkI259
5J6vvVOO+V0t2sHIDZgGuGmbxT4fpGfw4iM4UEW+ODmsNywWfr/grvBIMlxWX+jV
mqABtwkjnsfRqoRZRXA4BiBeLzq1Nr57wbL5gFtgeYD4SaGQbzwlDNd8MdoyRtHF
0CbDpq2Uo0HKSBPStkY/ItH8ua+BoQ38detD7PQixP4i24uX8YlvWR/7XXW1g8Bp
zusji4p5bvgVLJzHb57uDbAeP5XlWau7Zhmv//n8eoGMgaJI9Di/5xtxXwvBcdYP
bNrbWgTVRR9+4C2vsmv6dRekab48my62ju1PDPPxhzszxbQ+zo55k0GPUnOYt8Z3
BivzP2vIbejgFb40InuzYpZiexofj60gvMcPbszZqwvkl022PoN8qCpUiyJviKkR
3Ghm5lDgWEyHAeQHNQDSMoZlJTI4+PSqojXbNjYjhbm39vbR1AryxEoJH4FE0E0J
A+Au22hOcHe3fy21FWBwfkpDQMgGqpzlhHRrwriX2+YTHA7qvySs1QwzR+lL7OMD
iMBnQUzhEkd0VBzNNACNeD6WZ2JYsLNgHSfEOIaFUtC4QaGhOyuxpFiT6rMWmfa/
TqwjmsIli6PPd0c+Y95ftAmF5TQyqc3m5JhqNIOcqwIQUEh5JXPfb2faye//cuvI
G3x45r6Pn4Af+jaO4x8KthUodRCUl2cU6ANeETCiXknuKu/2jLcKOw+P6WA1MUKC
X9UtmDxjncSY05jtY1wawqFEyq2f/FmOF02a4WbiINp8vi4Z9NPz2DUBB7ihN/yB
dr1xeoxDQ9aZQmM/yGuT6AOWjWNPvAdzOsrq6YqpNQd4ImD68nVS2WWkRNHoe/mT
77/eQvUnkJWeFLIKJmkfUPN4/dvmDLgqRQ761lfSH2ydlrE6FS3oSFEcCcB+fKZu
F0IAyi+MYrvJAQSCuBDBe/DoIbM4sCSH//G8SNiwslCqaYzz/TO2be1nPCxUOwd0
5YU9VVk8WpNyyB6T46GMeE6HN+xxNBpGiia6Le/YPCT+pDZdz8VrMaPcIsV6cT40
FbF++KISUOoE7oZfQRSi0zCaiQw6xOXTWnIu3t/QL0L7BYa7x6qUARszd7ZQTEhA
LmqoxZ+LsNSSuMZN3m1OnfcePH46okVfMgJGHAAviaQoD3Zww+jdyMOW91ax2umn
6M50Ogl71Q6l9AyCpqiR8T5HIAb4a1HCvJQEpTkn7j69cw9LyW2RxAEAE4U+2lYG
C7nx3I7FlMdOVLCNHRJOdh+6R+MUxal5h1c5jPLBzot+jkHcGl4WKKqNTkui2Vtp
oUyq0WgG5CQHr4JSIrjYWQ3feDaodFqSmqiISEbCBomt4duu6QtyZ4Cv1G9+BSDF
WukgYaFZpZfLs6LRihxOE5sN9oJVrB2Z+m5l0MZ5u3LkVHADnYCEZomI0bIbM/wg
uUm7pk/ljQaBgvL1Zcb/sjzO288OMZO8agZA8WbIbsMHxefsK46CQtHw7/e47lYk
2gzAHKiL9j7et4NfkX4oQF/QwN+DUtxsZFDFTMLAJCefiY1sKlsH7eUP4SIXwc6W
Yk4tjLGQzPUheLB5RbzhwaTF+q6gfiaLHfaU1miWK4lzCAR5L6H9wvC5KA3/wr8Y
014neU2OyASzvtkZ5b9Rrp4u3ZuzGcKxk1sgxKWGLAh2ELz2tgksmvxEl0eSGVXB
xHRWAbooWIsHsvlJIYNNLNohX62rcefwonvSEJYdeD1MVlYCVAoWulhXrN0fYj0E
W+N7wXxa3MnWNHkP6dvPOB0X+hXEq5ZWyGe9RCmBDpODPWz94duTwcDXqAB3FqGh
oOxjYL8JCs+i0krSxpS5BuqLuokkgNonCbbiv1QDgOlDTsO5EktmDFNyP8FSzIVZ
KwVYEiXzJu8JxMwM6XBE3Q0vGaK4Y9rWA6s9BLu4K+Skh1TTwtjMVIi1XtJhbVLc
qIkaCoC/TDqeyK2iDslE+jV6ZHS3JZGRR22wAk5pLcHtl3UURpLDLZcOIiNn9yfu
o2Mqik7tzkFWb959p6NQBP/x9VPYbvKN/66WiUwAGRnKEq3S4dwi8hYakqmEYqtN
zsMmqJ4JPGVOgoZLmbP64jAZYhFgZea0LjHruu+sDooIHBnEyZHsyn3j6otsvJJ3
PKHIgcecT+GwqfAJzaznjkmgxeSep8pffOAeXsgSH8QNqE6c8Hw7SjEBDVSrdNf3
+adGC5WFYk7YXsKeOFmSALq5W8HTlQg/O6W8Bnz+k66vY/1mJdvsKvdkzALqmVHn
4OCpKNtAJD412txmmEE7IDJGjueXQetQApYdTc8fJJzt5bxun5kyzups1LV2r87N
Len+wylkmaYN1RoFyF/3cNUxl0WvmXtNmS9GaI7uvLHnTtvYzVulbSV9eK2xDJQk
ymjobDoTvWhTUNzmlohALZlXD0uuuZAbQTuydbdtHjtbwT5LGLuaL0EkicCHeSGU
qzX7cpimBALeGFP6AkoP69pB4LiLQVpGQ4P3KOzOnuyFDyCRzLSzNB3NTk0lx8Ns
dO/gj4mLMUVEentjkD5bv4peQQe+DQrvGVSQI0msPK1J5yIa6fAAJB9SlDg76De9
Hk18B9oB17ONtpcZrEKa6NsECuzWJMOfejPCtaw3FPWCqLXj/bemYrYFw80fFAVj
G2GcjbSgPEaPL+WUKO7Q6tZwtQR6qLg8i4iz7+K4t1HBJx5RH/4xCnHSBDF295IG
FmBcxi986MLfQCzxmo9EbNWE/vGMdhB3IY66MRL5Za7GDKLccpvWPD7Hu3LhcvKq
CW4pQg/qHI5mOhRi+M5UjWhkuoFGWzO5FeO2/xmPtur1kLgICe/JlfRtAqKp+kvN
AY4x+kapyNUrhmzjvCOQvRm4yc9BV/KGqFICA6w4W95NT8idFT5EcgssrqcKAa8r
aYNOarc5Xe9g02HjaUdqIUeyVpXUrxlcHS1mlMDm40Z5MXjSbQ9fr2zxxfBFL80t
Zc53r6Cs0jB7yYFmIn6VMcwU2/Y8NmOSwE4njClIdbtocGPzWhKVXCCyErANCcaM
Qy+MDrdPrgk4ErQCkT4Ude32XRDs0kP/mq9I6xB3xjUnLLQs5yQW2hNPvWadUBju
s2T5WaJz/jXqsDOK1Q65bc4TKZk0xXfKiOULChIYICjDAbtQgWJMSasJAG9Y+5Ea
Nooav0Qr2/XFZMbztPkzC2BOX2cgAOei14BeMzY6jz+3VOaSX8Ce/u8JUXO/Owt4
yYlt8j0E5OcZtb+zacmmf7EVOaRABezFodtLSJWb3N/xrwindf5MqQ7pBY4yxLVH
ox9uWDS0NxUvArlvcnBcCjcrofPJKOl2XLj6Ns9HIbbBHK7ned0z/8EalVxEXJ9W
CHBW/MS/+sVJFgzzk9M1AScmZpgWmTsE4DT9exvQPCHwDrDZAmHo3A4ad8tXzvqF
AZHRpuYkri/VRA5KTHyJWARwigdgnGHdwOoByhlMZ8PMRtJ09WD6+OCesxDtLvu9
xaeDGnoXt5tMG9oH0VVRwYiiDv73kZXvTxKlU2+16vNBde4W6lVq1AGDXLACT8ip
3qsJ4BM3y3slj0z1gqcBS5ZiWfqY30ERR2fb0vfGdCjWkn+qV8Ao6HzJQwUygX3Q
+LwvFfmPrMlkU8fDd9KexbJ1SB3C46Rg0cU9kA5IldqDRZ7RUuG1o9YTCysV1Gp0
rlvvBOLvp8Sm1mnV/nCCzI4IiOTp+SPYaxsAfSsl1Kip+CRasSC7G4+MFOg6BJka
SI2xehsAvIcziIRNZ+FHgLkwPvN39z7CIVT3HPd8/zfW89gmGjWlbcdLkqLaMsxq
eYlkKxy9xGDVgPaQLWrWqHTL9y5SIUodAjDcTYgjKoBPqRRLSIa0+4I9tY+UTjFm
G5t+TH+DX2CSfCAVN6dIX7izTxtHeexzdW24Ze5ty23NKq+euhmqxlrKXeRw4ER1
+Gq4hSLQzIvva5EpDZgYZ8h9khrMa6FHTPlrWOai74yz5H9dvJL91hFWsB488YUL
AuZV1bw0GHT35Va4K9s6L/oJn6iFJj3yiOhjEp6Kh4qiV8oxoYUEAnmDcUyVuQzz
E2qCcS7QK2M1XE3OnlgIuQzzS5IlZHkaj3WwYB+tzNfhEUyKKF17nMcuifcn2x4l
BZgd0ffOboR2b7Q8QZhCpglcIhQu9JniSu7oZ9pkt0SFbAnTlLuqFNAYW8HC8cJ/
Mp54lDaUbGJQO/3SVbqD0fJthcQ83z3u3QWyzhtNmcgSolnilV56Ddpf3BwdQNJH
IseEJqSSSOQMS7s9zfR9KzHjGY1aBbSNoCpIys/BUDIkDku3MVe//oAeDlaJ3zQT
BZnaijVSi6N/1sD9wLN2qgA6BhPnYv82sLC4Ked8pUnUxoT7lHfL7pNzOgscSylj
WmLWa+4f1ecW6KCfiUTugHNkf7b33uDlKwauYzo+BxSD/p6+UQZuWPmp9MmY8kFS
scG0Jwl7UnM4nt1wrHjS81uCtznLRgwN2arNnmxQ18m4wBonBHvRdOaIiEnYajh7
fqQsMUxfYr2wQyhO1n5m5ZAhwUx5Bg/rxuHxWmFFCFGIg/GiP3fIMbwxNUuQ1olA
rBPdNIMluQxsVEONu19YbKn9rJU3GduTFJ4j1l0XmZjH69lUCQk3rVcWIyOa5v1x
PqiHbJd2OGaU8BBaPVHwvEfDl5u44L0nc01qpMxSu262qVZyh1l+iodbsM7T40IJ
I7/PRNWEu8ARwW0dleP1pnAYv+2sJga8FnsL3XahxQZPrHPKRaIkbqZlR5EkMeHo
92eL5Oh0fBpukhk7tSzHnEZqne1ctCRR0yUjdvIy9F5d81lCaRtr/5I8FBQ1v0mb
fXjGWcVEBeqPXfClNg9iFR5Zdef5quMFGRFXF2ySbVhs4qgKeHEbvxxMiVFpis6t
ZhMSn7lRchVB2qkOeKPDvXT1rwz6zYcPTxP8SCeh8QWYNY33sL9+BohinrKyLPg/
1NRc1BcQ0eiuXfjkEWBeNS7PbWhzrvmdJo1JfdRhLldbUy5I2LuREE8YNCgNLwhw
/D6yg/6KWUpfakF6eHaxFsrVX1wH9vZh0ykFAM2clwC0uCIOEEBvrk612mTr9zYl
mZzWdbFC/MuLRWTFEjL5NaH3PPJv51TP9he6/4ppPtNIC73gFx1RdIA+0s5RmfhI
LN5q5onHGGrc+JWYlOdT6mocOuZVint9yTPLG2lQ9VeahZ56xSNkaXGU3ytnYhim
znJ1Lxft9IC8eemqGC1bNQ/Uq7Hr22dXeSN8SxzwyNa2lKcHiWR/TLN7LFCShdWF
hjjWxVSEK6uEXx4xH7zJc+dKNQ7XqC97dL9msjIw7w7Ppgvx/WbLFZbsnvJSHm8/
tnbx045mr8B4x1lMG/tF/dc4JqiqOugB6opeGJwG/Iw++8fikGwXn0DqOpTJP/aK
m5htrvNR9oUbn5GJpWLlxM+BwQrOrcg818jHT5jipXcipHukD8tAWPmz2OqoadDK
QVPDcWWJga5D4zo8YLUHA4SWyykOdAkndOlSO0BGOq3zr5udrBamnicPrAEwz7fw
khsZFC/34BWpW1JUnZEgCAYICcHL3naz9w005V/d8Hj3ItG+UdzB1kPo7yCRWGbj
bYPiSyLAyyCInzlbYeRjJxsSHnEqpr+0+gvy993/ODJTdemH+ehRE9my0noHYneH
KzM1AKJHmWNrqBF8DCvr2xjDhX2mJq7663KQaJA+IvDWbacy7jvfSZc1hdASTzlV
urd4ONNxRiP45Q70aU5eLrjjlm5TcvzR5HKcKFclCWsAYYQkQbQ70eCEVpTVflb4
FYAhbn8oO77/lE2prr3GMtxYrjWFYQw78mi4iNTUv4mS/Pp6GD+FeGQIpX1VK/tt
JYQ+pPG8NGxxaPwZXIqkvzx7m+9COPwj6HyS6Yk3pzmuOzCjRM2GeNM1N86T3H/c
BsGtrLETfo+YFB7LgoKHvxsTeE15O40ToSQbWyqZrXSlG49lr6apfB1M64u69pS3
vXmakoRVu/Ul7YFbGDSPdL1KotOMQOp6Favnf+qLQBWUutdG5dnLJWlizBvnL/cy
hE46CqCOF9CBC6MEUobzCV7flf0djwBNFcZUql/BMF1CGgEuQBstOPRO7AmCyenn
mMWsfvX2V2XoGGopoBC8mJv0C4G63HCL3pyHXrvgDEDp41TDWX7BTUe61r9mewdF
hKHjFcN9Ftir+sPepMGRR9BbbJk1gpHfwQvbZoFc/C/NVjwEHkHfklzol97WYq2b
zNHZxKJRSDOejTAlMtNEvdokpJ+zquA8gf8bUHxyO0MGfLvYZ2YRWGu9plnBK7ss
F5RwPcaI0l5KdThqUCcVRvbZ2gZLYiHUhvopBRbeT+XJ4zsGHGAdu4kYS723eq5/
R1+TO71iBab5CTUTBmLuecaV2RQHI/6TUxrTnBEJeYrRFkgY0gtUzQl745vGrQ1c
gv8eNNqS9iqFhtm2Aw3zxg+9buJKftGqVxOVSpgBPfU5uuGeQCbu6s54BtytGG2Q
96S/7afMgqZ3KBwl7FkABYaaj8J6+A05oNufBNr19aP5NVByMCv08XtYjb0TtVmR
0/1HCw+XL2vtI11e+gAq8YxZVKrsojA+lnwB6n0tsrezkqz20ebAD2WBF2CUjXot
e+nGmBpwhjlOVD3trnghc9+Uq2jo7d53y6hLNL3c4WPdqfdsouOfqUSJ1IacjyWV
GHNOoO3IcErPdv1/KxB42pT+5fVcmgMv7W8EGbhplJNSG1riInuKiuoAHxdj+aes
GdKfIfl7GiErN61K6NYaQiBCdld8iloCUSKIJ/l3w0+krkLlgDuxwi4ginpKF44Z
U06IuxcHF4tH2Sxqjv8izF77WJHWyrWFmDcc+WBeR75M5EvSoHnVzs1zkbROJMoa
emNCiCrtjdtBNGZEF1g/+R1P+loNKi/TkzuvBnhYASqQLiYMBslfT1qTLVmdh2y2
ZjnMPFiD40Am74NsvVh4Ac74Mw14B7HKOYt2jRn+j8gXlV5wK0sJMhgDpt9eEHgj
g9U3HyudsFhf6XDZjv61sj81QpjjmKpsTjP/6aw5keQkgOPngPZowSpDHbvYfyLj
fjJF/3Qm3q8zKQbWWEokN2gM+aqb5Apv0vsRYkHLPn/ZyeESTy3aSQ9bYN4RJmtV
zwZP3fLN9W9kV2Xnbxuy8ogUnCN3f6uPQ63XtM4oeEeJaZ2w0g45bv72KzKJCAAM
LPu/oizDDPifP12tEGSHfBcbGyPB422XwNmfcRVLGikBQxwSy82gdApkdZPCU3ae
SiXTWm+S90T2+2CJCZLctz4XtwpCzhv3zDlLpug2V8iH/MA8CPrhOaARiosreK7l
RqP2KCKbuMLWfF2SgekKsGsz2kYUEmgEc/015ggjWoWzQZYvhQbYJuscmUZsmE6p
2SfzqttcmXK4pS9o77cDMiP+jQ6HSQK4Q0QtVn3nfdMP5RVYaLLiY33kXcdmTaig
dKkbsgEZ6SYaibtHMCD25ZnU5YfcXegjQoEWSSb6y6wepBtiZ0wR7MhXxnTiUXI3
CYHQY1NL3n5CAX+QlA3oQZRFrsmHP4N8nILdervq+ataxBHGdN5WpanlbbHw1iGR
yZOXrhOswlhE+PfUXz/uOoJk/0SYQ44kTJTFjtyDtJsK8w5qwJy1rsYyvffwq/P4
TOnLyD6VyhHUMpzEs7QMpw77hJsjrCxAr3gcH+B6ks8eg/OsjJI0mIofj2mk90/C
EeQj7NO7AVnrf/ppXQkAKge/7shYVc8HtkpBX3lQtlPNXHgbM3nN/GFxbkZ/aB6m
08aIbM1e0BVPMD5iuyRtJgxzkB3/MIcSuiEibuIdYBGFMC1fcQH60yOR1UtUjDil
8vo+MxmuIxl0CI7Vl08zXdcr7HOudzN8UpQUaL4qKyxkPyB1qchP8iN4Wi+q1638
YUUbROpVtDrIPHHuvIh3ES74P2BcPIa7CEw7JDkgpnUG2HqccfaqPnREGHG7VrXX
kyzQdulFZj8um1Y0bcR0TD4cl++sCgelcAQdnGY5YTuYfPNvCD/ugKjpqy8Cx214
zfMBw18rCEZgk6+bQZMxi+WgYwEmt2C0267CZR/98LTKDYq2us+6U7u2A/8Hsjpb
AeQNmcR/sCsCFWFVpZA0kDCFLom0r/tbt21WZwHFKZan91AiRvQxn5yE9PzkCbZf
erV/TtuuKYTagf4Dfv3gTLQCU26qBF14clt3tbWG9/MQlwByBx4RCcG2ZByNuOkE
yfarwttc+bH/ce/l89dwoiw6fV+QqNtXpX9iK8juukm5YKLVva431ndx8w04uNBl
yTdcnlV/qh3aVc8zJM98H9OXEgoyuBLr6LjhUCvvfX+f1wi7LnQLgJ/4YQk81fnj
DC3bS4jIRvEzzjURCQbJseFZj4VqBqnmwUO6QRg/TQaLiikz4gq2K2dB/aSjeJsg
KDxTiMEvg5TaaReW/yexXvyWydVsQDZySfgwQvg8apeYhbsq1cIVI+0ztMt8sEg1
Vf2JMHBUc+tTXHXpFrVno0Oo+9TC/7STZ1awRXJgP4rTmzpj7txLjSPpOrdom2z0
RJqB3hGwxnJlrdJVWNWe/kwiwVW2LCkej6qDSlnQn6JmSKNdpu/IFLNglflWj4E1
sQjvxmaOFzgdIrbLbslfHblUGTn67pIZ4KTnZ2Kso137TmgkPfyUjpjPZRt3Rf8R
3g3EzfiDl8Qxivj47wSgLt3plXx/enLJ+8Wf93DhoQJu26xsBxcJl0y9fbDOCfYA
ObP0aafYQUHDdBwdSry3rznEphEpfjJZ8wTGqw0bkx5RHaxcf025uNuKfPIFgl5M
8cOwxXv3+QkEOIEnRX6smHE0zdCVcaGa1nG+FKVH2I8dFKBZaJz+G7YbxUUYRBYM
Q2vdteoQR3MCAPgOGavqF8DKmp3jw7Qo4/k6RF19OlkVlmdufYI07Ea+luZYFRm4
AStgGJynIvuSZLd+hpdXij22xzAxpF5leCeB4Oc8s4OG3aJ5QovbVNJMuzfaVS85
LW0p5mWOjFiQDVfJvDJ1Pio9Iw9z+iQ3ofZ0WKrqd1V0DzQVOLSD7bqtb8jlluNN
ou3M+tZYgVSTStCN/TL5GT7G0+r6OHqL4eIdSa1ixbEcU+Mp9S1tXoaojBTPS8RJ
BTTwRs2j0yzarEk10RECg+ZmMM+ckvsjIfYbsuSLU8x7hfjcvxE5ckF1YCz2xEHE
nDMOSITlge7IRPFp9CCWsCqd7xBt2iE2zA645tSx2XsXtFbrlJPzpyzxmL0gi3Vz
PreTzVPgbmIqFm2OTFIT22rYUvKAXAO4rLJV9rQ7vbtUzezcyoo8aFdiRvfBiX4F
xCkxFh/qagJbIjsCVPwoOJIpPzK9itvnpgGiz5UHI/zXfI3+GsXhWvadCusi/Ubi
vGFO8UwpSFIPAbovXvDYkMzirZkne10eYh8nLPnoHsedLOVNCltVgsWBYGQY18xt
ZjDCyvW1ERqtwUEeHCVbke51Fdm1dSs+gtxULXYySE8o6uaMfymwSj5RMjOyN23r
zubnwcCRtg1BaazNRloxYfxPNVw2RmMLvg9wZiUo6AoqY5RfPpsd/tFb044UayBD
G0lgH4BReHo/ZQkq1TChnHF6Fdwbm6/5HWEjMNdxi49TKSESLwRfp3AXVvxdfNjv
Awm+V7BZSvewe4X/LaL3z5VNgBqTa+6IRLEGrGveJpkkSBU1ajItnBcvQ/xMF8LE
ia4I3uqCayiY+zjsotTMydt1U1IPZU8mbd97TsfIUoZGHwN3/z5LQMkXBWDMmu7P
kiYO9rrTaCLWYYuWe3DSVsP3v95Y44/hei5O8bl8dSGJXmmY3UZ4tJhoQzHOECq+
r8WJ73aQLnigVnWMx4CArlj6vXCXturgonDgXyetVL5qhIOgApaGKHrv6zM+0nM2
wKQqM1MnCUJyN3h7V6oUFJ7oYN8HzsOrSh3sFuUEMceLAonHS6sSJRzI6Q2zLpkI
MyaSNFi9RHzNvcQyIWzABhnmn5ClTWR9fDnlmvXIliqWDf+pzv6rrdS3YsSYfSNQ
qQ+ee4HvHhxL9uLMyYOWOA0QMPJIpwvcJDlzBbUL8tJiWnW9+U10NXUYUoPsvcvb
54sD5ZH3uyO5VPxwG9qg7vwxB1j7KDv7hPuQpnwskPAjP15gDYHxuR/ElH61XXMk
wOAJ2jTB8ychdwOgzwqLUhzwe7GVcXh2X/mL6934gCbT+NMW1DqdLq1XG8yxsIsS
xjskzIuFuxtMu3fcxWoYCtAqqZJUIhNDoIdVDl9rnCxYk4SS31pEVQ6GXYSgi5Ca
8sB6HRCxOJINxKoJhyosBtWtFZFtgkZqAdLgsMvGltR/t7aYBMbe5jdvGsJOwDZy
KuNDF5z15S2jPG9dL+Nu4c1GapxqGBXLbTtCTgd9TLWsngzJYOwQxhN1n5ykYQO3
D1OzivvLb6OelR7q5YZnK4Rl88Ag9il2wIvhC/Ota2VEywKTBnEz5uz/iotkd4dz
lQ89u2e79F9MVS2sEfB+Cvezdk27eq3IXFoCNFDlf0KgM1xhZ7NyL4T6UVCY8xXm
loSKXu2yjyF13MjoWnlVnhsEzoTshiDITARQ+8OdF8rH6mFGZ6SLzI358IIKx/Z1
sX/henxOC6nRCy+xci2mtjlp91VwxX+YSADMd0+yvDJdv9BWzmKJZ0YJgWf+m/+A
yDQzDCKCNPNk4DCRnaIJbYJ5dpp6QCXOJTffxX3oFA0MwTOthLscJHKLpU78nfKM
f5lJXoCrEmjGqj/KsBqn9F1C9I6/7/a4nSYac3ppEqYg17JyjpmDxM2KhL6UwxnX
SYBytyOpw0kp/DjNyMMlzYkPHgfw1kBhW5DIlTuqz/sxbwR1QRN5IIWaYNCUDsqD
R4ILQdrlcytR4NfDSUnKXzFRgHTSp56mRIf6sfRmkEemo5DY51i8b92E3uvWF6Kr
yjMF1tshYk2C/bc7+RIiJmUmj7TcwrekSAdXK71bodSudT3noQVARTrHczb3kQDm
2F7OZFFaxYZrIlaepfXGmVgz7nkrPVPXXlEVULX6+fUI+CwXNFfRMX3PlAtDf2gX
635I3da5AmTHIhAlPT+UeLQcsGGGlLU0oP58smYEFNFI29sqVD5yPHOQpJz+l2q9
q/Hrp0elCscpuRG9TJWTTTslnJaidz3T/lNPpa32jgv7ntUE8SZ66yN8dSgRWyb5
ycXMoHIjRuTTiWvRpRwD9Nv+0WMCC1Zq9JG/5+UFFylXehhMCdxrSv4qKCravLS7
7xjzjvYLLWhKdrLugrEmr6W6raGMsmoN/Yco3ZQPv63j1QtG+TmN4HaTP4lkkAJv
IgmVyAJewJs8ozdfEy/47rCXghhccm+RofMIlUZE9PEwQ1Y6hjiqC5deMM7wG10W
KUPtbjsPkg9RhI3TM6Gnph4LJ8kkp4+FMIPa1JsGofLDN/QGkly2xb7HJfkdk/p5
onMOHpixHj7ZwS3JbHYQyEOMiaAMIWjvPXRlAqfIiP1WHSYhnNkaz/BvIhGNgbAj
niWMSRYqISvXsqpkuezsKQuSzdyiKkjy+K3nAxqOT4X+d0gjmvIv70B+16Vh9VgM
vEDn6UFLNhwO9va6VwH/hXKWnXoHc0nUBuH2j9Mb6OJQe4bcFKmRtpMnZxHZ5fI5
Atu2nL8yj3ZsAYqVg3DXvRJNL2O3JS1VuF4Qro4XetyUepg4JWDWt9VpAXW1OAzQ
0ZmtTKRn9MlbFpjc/qlePtSEQqPbeId1WQw9y35yvZD5D4PfjggM8sCs/6zZ2RIA
USlp36FHUA5QulIBaChDP4aVFr+IenhPQqCIeYpeiWvhPSIUX55GGBM3xxX0gFZw
r5c8zdyZyMSEDlbqHCPsaXAhYZZSx1cwayAGb+IDWpLxig0hQphnbqAop5K5LSv1
c3CK0EfjTEPQjlvXWHWpe6jDiDmzz3uVff2qA38Mm4Xit8IYylmuewWsWBJgbcjP
fjsbmOn7+uQgIWXEsJTOY/D+DGbC95Cxi+CuOdNVAKRuhbr/L262i/oiV8PDqrQa
aie//OUhrVRaF2tHhFnH62Sh8/rjDg24sI3NOynUnXYpFTjqAPdmK2BlM9tWJOJX
R0joHxX6pB3ie7skAh+GwK5qWhTQ7a+fM5HLXcJ/Knn2sgdF5/Q9vJtpD5Fj4CAv
Roz4GGGnTsebdU2ORIeflJ5yozIlpIIPcDz+M5NJ4T+9HUpCKi0Khhz87oQtxhhP
k5+Xna5mounUfj/s3ATxgIsrc0I7MywkWqicPWZte1gPNrrydNyx5MJ9Go9wAAZZ
noTeZXtnjTr3KN16fJEiEggTYNkrOPw/25QEMU4lDxa8ehUGWnX74LsTU8+izHZN
qCTHjuQes/hz/39VKYUmcs33rG8si6QrGI22SW5ISKd4OxHXzKZtivuW1Hj1Zi5r
/BNR1ElEC0mUjyNHrWnba7LERy17nwi3UDGMielPIuZs/TnBBMA9ZrEKTMkUxByK
m4XtP5J3rBLIGmpPfv6csish3ApoJGQHvLVchL+tnhU9GubFo/XY2BfeP9yx6W1Q
KcZ2K6f+RjCfW6GDhrYcawBzNl3aYAkhd80u2VfeIiAOt/EA+S7xg2rur6JkESbx
HAlDIrEKpJp3bFJhsTJFzrMML/ye16Z4NvarRWcSB/GSYKXlzevfGB6j7HmO7TvP
Z565tqJB3FCC3W9aRnopviZ8tEtVTkbZpltAjbh6pTouCvVJdXpy3jKRh47UYrYP
OAPQwqEGRgjTqSH86cQrWg92SQW3s4kflteRv29UlqPW7GGH4y6Z9qUOeDdiJ36k
rQ0Qeb0ym+pfappngWmtY2MoCVd/V+1BxG+Aqzac+3eAZ6yhz4Q16NY2as5DxDPR
UA+G3K9lANzOB7wBRQNfjDtFt9FFDTaY8i0akCppGyaviPw98MFH6nfSJfFY7jrG
WLuSauqrFVPOywzrasn8qZCxLBRvMKlUaXZq+JR+dYheQlRYmKKUd5vDA9vieg0S
Y41iZURUsQ/ZEEI5Q7q14Wy60r04Pijs39Pkdwu6L7rDBYb/DVNdqteBt2WCLhQr
iN8O4TASO4ADcTXbEDx5yXC1+bSsVdSo92lXYBmDziWXJTaRlwzeeVaHqlUZ20dd
LNqBo0HeLMWCoqqd7Ka/SwXIw3+mo5tlJe5SIIZUqTFrja+me2vrLVKmc/Hqz9aV
jsb6v6wd7YIkZmVmJDc+4p6hy3me+BB4sIatfnXc1U2TPdksl+DiZRuDaCK4emP8
JVBxmDhORPzlRYlXryHbSA49SUOFrq4lXIVrSXRPfe3ASDexZXFKqNJIoMpMhlJL
EE+yWbNt3MgT5zr4qofUXYmqTbvUKqJxFjZqWEtvmmydnS3B92NiSoEVUt+s1zFC
fNmzykt7UAyvs15HGJCCb3DpsPB7KCvRvtxzcmw9fCtFPgaxZPj8DZnXp+Nt4UlS
ExTRTu3vCTveFcH3H7IOvsWjZGzaIuY2upFW3tE5nGSYWxxQj3pffBDHWUkiQV13
UWWU3zQO8JB8WWbdiHOUIwRjVlYWwSKW4nmysl5DLYnjKkGD4Rh6glYCGtUGxbkW
Jjru+cbkvZkwUxP02R7d65rEityoY2qJnwIQr1o5kaxFeRZLVWvr9tzEyB3ExWE5
qppXoaLF3oahduvfiKGLcPhlnmPfKoi2tYZGlRizmVPEHDWSCYrOP1IFwU4Tgk45
xmFFgcaBiKfzFQ7Q1wA/KqI1Eubd1AZWRUadJtT6xp7tbTMQEIDtKiBamMla44kJ
13hiisBDlndnPTj7ACy5qw+TAstfmb7yagfKIyckOCmaE7OVb2gROwM0rRlmFsrh
JGyHeChArpkRET5ykxejlvXy0E3QhNx9oSLVPBB1HLhe/zfbtqMVoPD83glv+7Gc
eTkft4+TImhAUzJUhEF+UaiAUjnXq2sO5lVgvOXsF7uMIhhPM/3gYNRaGZCK2KCe
3rHepmHT0gSomCwzpSVvTEYGMs5XGy91rEWccskSQpjZuCbYi/OoIHN3vtbf9A/x
HsiugNW2jQ11L7q9RD6iXDTcIfmW6fluHqYU4fwJ3hCt6Z5GoybCwcht1lVXVFgU
Cg5C5W92RyuPIfA8n7g/9cIIEqALH9t2QQuZz2Bn1XB6TuL7KW7U7tXCMANWbMuc
hWAQzUjq8QPx+8P26PCC/ZRDr5t524fJwxaLiQCbjIj8AJZFLvBZYv9vNIJmFW6G
Rvlk5UhuP8AJHiVZB2QfzyKz/E4dKtDuu0UsoTNn6kxRjRyoPS2ZJDNZ9GTYIu46
C9f28Q70LQ6VH9BNdn8O7zm2YkuBUHe9joUlUQBTwmI5VZTeKM9ItzJ/J55Zvq7O
kzanOHSoy25DZnem/GWn3XcyL2th73e+MHGpGdSj/5vp/gqvJH9FxTqKym0ckwWC
WjHOUL9XOQmLLTpwDRG6Kutp07qPkPHLX74s0VYhbd0b0e2eK4KgYMdzs/vpl6tK
z7B0fmDN3IHRVQRCuBP36TUCQjgtNyb3qTb8rNgmX1bxOzR4YjhqKv556st2FtIs
Q5G9UK5Dy67f37cFseV0+v+UaNFNv6F2uOqZneYhjW5HEyfGGfULzZXIIhp4Ndzz
DsyZLeAuwRM7GUQGrSV5+SICIFQtty1tx0i775/kvC9281UtSDrUgXmEdOZjztqG
uKCE5Pc2eGuhRKSt1Ffk32BF/+ZxFwfgQJSJ1pwvRjMlGoiFxDYN5T3yC+eatfuy
m7EC13lPWzxx+sUMebm09b0laAzjueYduhMvvOpqjBBxdvPy283OLkkmb4HlhzGK
eMRVcQyG9PMgtAjPcnLsJoWxYJWMkRB5oB0tkkNrFZ11NN/vRkvuS2fXAryU0T40
nXWCPAsHkUiYY9Mve0/IArImistMk2Mw4cQ1g2LB1a/A7WuOJZT6iJXFAgx1B455
hE7Iehm+TnMlYh5wOhrkfnkzcCFuCWlFKOWpJesYgSTExYweqQgSzA+118OQ92K6
/oRjI2O3cN+Rj3WNTlKNHeyV9aHtR9h/86A2cTHms7QqOqLpor1iGt/r32aZ3oft
MElZ/gbOA9K0NcWA5J+m+dkpljiTaARaY4rRofsYorK8Ks4FBkvVvP1fobj3j1Vm
FrdC9pzeVGrbMRLWHwTDPQRT5K6cguGbb+FM3RJ5S4ZZbgaroksrqz9ufun4BNqS
aY3DEInavLHJLHU0CiXXYZ56lzrfVOxaipRJ/j4tigC0lfHu0TgZxfcnienODBem
laqNa+KnbQjJT3kKFo0+iWRoGKsCs5TuTWnV4/uIexpfix86HmbRFzzIPLUvn2xa
p557TQGR1UdsRcFVcjqML1UM3fUKPXzhA5uWJJd5fOQBQQ5MrcKNwL691hQUa67+
REOSA9bOAdwfFjgdsFz7PGi7ZYUiWDbLUZqfKL8tXxmt6OLXUC+MxccUIhniG8Ny
uCsBGXSMGi+2MRCSEGNZlDHBSzv5m/hxw1nEgOLIaBORkZ9BQQb2ywJM17ga7t2t
sg6U3QCbfCW+WD/wp5NucedwJJRuspj2a33irKnzT1qMIhLV25FHXjRth3LHEug/
ZxCuX7NintruKvHw2vZW2XeemYdjTYYelhx6b+Ge8rFiyUhCDUMz410VnciqKtiH
JfDbOcIKC8daJ+F9Gzib88Jc0NTifuUpfmMdU8ttaKxMPwWKOc46fHTptlHijyKg
dNVHol0pvZI71jzJWLeNw0m8lJm7b32Q00aF4e6JcVIO+qqAUj6zaVV7Su6eVKRd
qxKyfjbrl7d5WtmB+pwKbHPV38HRG79CD2RdDlt4K9h/SRevGGkl7pkIiHfzrHGO
wTzv1iv/F1dyoxlt3od9+oODjJKQpA2YBRKT3eEIYwp5K1vBGrG89uLSnqRyQGoM
g7cfbOJstXvkWxAX5D3nidEifPEvKd4zXsmBrWPXhMuMS4XC2p0u6v2c9NQlF230
wgB9N7brO4w58x2teauKsf/eDZg5jIyMzdDZggSaITVX7x23pVlFbfTzVu8ayj3E
judlQWt1fDOmrbU1Oawv2wmBa5LC4W3CG69zSEp65hL7AjRtL9k7QmrGGv9yTdPa
fMnUFQRzmgZrMd7sMwDYFS57s8FsPPDUD7C70EOUZa8slO6gkRBQX9yPoHGOl4Au
+oZ7OI8fz7g6fpjPtpDLfdmZkff6WRw4dciZqS6OH+Mdo6QzJIsmQwFnc3QCGqMq
FjNpE1W6XqkDERQvXOFMXHC22kSt6hRgDsiemw3alyFKxBwUAWacqZffiRfkeBTO
FTxkj1NeQmtcB1fuBX3JaRnnTIm1pArb9Pbs/KXlGGYkRokjXofN8Tk8XxGU+0Pn
L8TPQyCpH5OR0+SGlNjlfqN1hHKA2QR0jCoUbQUO8bXEmBrhF4wfTt9zJxcH+3al
jW1vup4epCMebpMD9fGECh6EjR/ImnbwgeRYRvQ7QzQ9/4t8xiRxm/vFA8YtFOEM
FFQA8B+TDjxZuL71womklCrfsAHtyG520nzSHB3+OCMjUdPWhvBjnQFXGLxtFoxJ
XO/4vQW48giQgkRjMJJiyKFxAb9eVunnxtnCH0XXMNouUc6yOEq1glVDdCUvKyZf
xTGZqO6UuEVJZ9ATGmuIM036uVnR40eTMt3K85LJPXFei0UfPfTJykj483RzbDp+
WGKzQY0oxEH8bZ5G6ab/ALmsu51gwL7ctshfPhPsl+d+zKNccLMYS+Hyh9dXatXw
BXys6OuvXhlRYUNbtuI8D/9tLOKx5v1/H8EKcqaTmENTaVg1lWPzxCNqdI+wR3Wg
zKZQsoTD+U0JS2h67HADvkAIsaaK1yoc3APicdS8/gczXAnWNALndHwU083wN4Mw
Yw/YizxP8xPb40BHXU4Jm7LPow8zqI04k/3SNopooeRkHiF1nJb/HPSQCmPLsFEe
T4szj1i6f6mHgVQrwlf7vdpke+qcGdbGzJqDQ5x83xiQfgJh46/+2crhRMDt9Gqd
kCe89QgRB84K+5Ns3Hxr9FWlrKb99ssWeFkid8daTqKN2NTW5XFuf4exPzYowtVM
0m2Cqt746I282jDn28RrRIRyTobsXLF2xWJW+y8wTQokrlNfNzzoz7XAhqs01kMk
ZFVKsERQkruYMFytZaHd+riiru0Jy3j7q52rVy/Nd+QWOjU4E3Leb+9vwTln7oRz
Idk8195mkfC1V0FElZ9KhTAEa9PwCIjWsLNk1RB5qLnB47RI1awBKHQ33twKBYSG
jbxukFkLr0xPCVGpYTTv8qQ1elqvUsUJbRDJE07Og4SZgOe8RIp58rcqd/BUakMJ
MQqmRmP7BufuVxPudRJPbcBacYgBPTt5/bv30tICFhU66WGO3c8/lftywknLMIfN
bTsTI3Eh1u0c1qc27DihaaXbuSVNE6eo4+rUE0bKrYZCnUmIAyQyUXaa3AYAvjAr
6O+iBSgqOaQMKQ7SOnHCzxYn5TUcjlDeABqkKKjfnSir6m0u0UtBieczaGTImGia
QDVlmo+LvKzKCszfGsNihQETC+UfErn9kn7GHwppF6EXUkoXDeRSB14PhIaJmdaz
qZLsYps6+OglX+4wYIh5HRgYQI9dLMK0XLwnshR2MxWPHU3mWeUhM6p/1LxP0G5E
eze4RzGfXUVqzBqQBa4OpZi6t6rNElQcU9cjHz0Zc79sMUP+HG+cqbRTBG40Ybaa
Frr9xikDnoQMXx/KrOVdd+gIABkTGRMPhy+dygb9PqH4f1S5ifW9PHyTjjCnLv7u
cEtZhu20rcuug2F2v2NSOC2nkAZQDtI4Qz9byHjd2Y+p++CdNSnG6yURkaZxuO0q
48WTFootRPPdlGZ7YqLgCdl85TawDO/vi+vDxXwMP35HKRfmKpxiSipbMgokyf6j
PO4YVBuY93OtX7ojS/VTl3ImYLCXOr9MdvQiqZVr6yK4nsk1kOFObBRbrIoe09Pe
PXBhSfbwtI6jaNzVbvmao2bwZ41sDLgKRlQnCWhNLR72cmcUrCJu7aQiABvLwVhy
MuJd4LYeo4Lf8Kld7JOZ0NgUhWR28JRVxOPt4tRc3th2IRW7nHK+zZ4YpPAhWcUk
+oUHANXkhadc6Oy5aWbB59D6f9eW6y78lpTvNVxUEWAC17JpV28dyh4y28hqM7hC
W6p7XaZatcnVjaIKRAOe4bOW6/3aFNWeZBV1AQyaKL+J+Xf7wyOIMNtxYSNKUu+Z
BAmELwUJFdOWQlTNPWL8WWy1CcntIn5Jrt4hYMkWRxX6joK/Vx39d/P9eV4CenxT
tzWQMVUvQ7kFr/cC+jbK10bZP19QCcKxWkH4OyTCTZSTzOJbIg0yhx1Ee8WcPBZ7
/yyEqXVK9ni55JGzMEif37TF6Dbdk4RLGaWkIeKCkccEJa7dDMY15ng3QAIdb0aC
++oNM5wO74iZWCzJ4va3TJebO5NfuZM/icYUlzDsOsapknkRqNGuytymRmeizNtT
qctU8FzxjjZ6cjrEy2Tzf9esc2/lZeTndnUtqxj1j7AJkOcW2hdiuliofu0WFiIq
tof/LstGjV8fxYVhBrNxT3spLHhiFyvl6d8ysJ7zgaqE2RPTgcBDhfFf8j4fT3mZ
ewdUgMuPCMdLc6qY11dTz9S+FKaLkmZIbTrGnCchcH9ZqUW4o8lz+Z/YHjOqwhQw
GN+AYIy4sgu/wL+1UUlXzMd5Blv/VHMLNHz6N2uK75qz6us4HhX71JGmmdLf+SZO
Q8htjFWYO6smoczBo+DOjQIpvtbeqX6wFCpY3JgvJm9TGRYwExc9GZyHmZTUgBV8
C6G6Xqu9naT0TpGLSgdk1mGUMtNxB8geO2OBDu18UzBwO4eqK6tQfV6Uhc3zERlq
ZlVjMScL0XolMHlgwohBIntgghoCTUJemkiy+RI4niJoW6muMA1vFXwp1jHVFaSn
hRrVkAakBCbbFDwc6nhb43eeu8cIZ9fGtGmsbTdSFC9qeWxRALfaiuYbV6X9ILKt
2mhJxdmLV/cyzXtt7l6bzdvZE/VYfiYKAkqssaH4ZeEc6dKdoxFurOTYdgapbu2p
0E2cO+cFZKvHh9/3N/AKJ17l1wTo4y8CudwShgLl6Stae12jb53SeYVIPPBT2J68
+oE2i4+H9ko/TZ7BIr+++kQTcaQ0KrvFIHhoL8Lj2EmhPb6pCWEDlQsVFl94o6k8
+b+vPV6xQ3rXRM6BqTNZr4Df+ws4VDDwFOm/YBu10ipUFIMyCoqtTa6Dzriwu36B
jPWd/5TSflL69GuF/9dzNzrch1j7X2QMdZb8P9/UVuZzGRXNkozk3NL/yYeO0fEM
vqJtFQyF6YZjKB0aaPTXHQ9ttXR6NRj7zGR0AjKjGgrT74q2OMpZ0AcPALEZ3tfI
2YL/l8W8nig2+pVlUF5AQR0TZi+32MFaFsjgRRv8o9ykJC3VZbaaIUqfu7oMW5/h
6y+gqzg5BdXnTlpP1hIcM9UIZdcB/ldu1frQ7tcTCByp1EnyQ7QehLFfg8aAGZTi
GVUKNbgoYU6DkSOP3nmaU4B2IDXigqc4mTs2YAn05/R/mZOIvZdSYQEloESXxFhV
2xiKapdSKjp5W4BXIL8yKf0FCTCk5pJbV+8Io5wy9WwvBkNj9QOmKTsVnJeetb7F
Izs0JVA8OR/6HT/QVxliBhon4513N/OuRPa/56jM49pXEsTs6tFiv0yPf3a3aSI2
9ysuJzKaNYa6ICJRj6tCXulOER2rzcD3M5E2VzHzvTUH8A0O9GU3rG0Io0uHLlmJ
90K7e/J2p57S6hDWH6gTVPbLglZgkLGd764u2O/tmEsUGpZgHKwCMg2SDyB1pI8n
kxdqf1LMaP2RwY/8RfGUXJ3Pgsy3uJeHk6I+R7KMP/2HUbzoaOgyRVH4gQ4q7Bhg
kofYpQZusv9nRGn3ZkRhbXwL+SL3Z+zniarbn2l7h1gNEHs37H5KhgENJysE+Ssr
54iTQ0Ua+AO7mxsvoaw/DYgaolBWlIbau/t2GFPmnq5+/ppiNAP0MNqAji0vOMGD
JDt8QdChjcH1/F+WFZLesERYYzEtbGC9VZwXQvH1azYGTOmkQOE5cRxSrHXzfMef
mVkRB+fqoVMZ4e+PBIMOBROJoTKOUk8Rexpad+hQoKuQrtZQUiLH/i6aVITniMrk
gqTDl+24G6DndMDHt133eKbRnJcRFlzjCO7dUMzokh6XO1kB0U4OGuFle35xl5f1
2w+y2JOZv5cReoRQSKPSyvyI3VNe1vqdXGIOEnW8R0mvHV6gysY9Y/eO6wDIE8+7
w3UbSKc1a2sRnHixsMIf3VSlm5zX5jhxm9TaGJMYjT4obVIbxXcZb6D52PSNPm1r
wpRJN98LZQXT1HCUpl7djXfHez8EWjsM41z37Lo3WoOx64IsVX6PlRknIBS9QDCJ
XCYKofChMaTJnmNJ1i2WXDgHVCUUhYq+ocUQ4LS4nU3F/APZo6SkjUee6e4WayjE
yzabOiamjuWOZMqkisynnwxm0yfE5uPWZIQX/yxzSCUQ2bOw/57YjcIsKM/95Vzu
VRILJuDCwFcIGG6zagbhUXyl4QkCvktRYxQombP5NYriD5dW9WoSq3vA+dqpiQfU
tMM4LzDnPIaEMBZpwiCQ+KnfEprj+iIbSltKloPtCAhZUH0aBWpRYoxlztgJeW6Y
y4NPPQvt37GJetWALJU3VQvsxtCV0WKkXYCudAiA6Jo07E9eKvgGTNPgA4WXEW1I
mdilndC2dM4YKGx/NCtmEVLTiMLgPrd4e+Mo+t5cR52ARWP6vT6OMvc0gkGJfeDN
uAIJDfQFbBnYP7PqIj5lER1EwsN8XLVVL2LpyBRfEy8fzaoCU98bg36F6LjmYyzU
PAybzWUgQRaLG1rv6ukydvb6K7YPhVgXGWkuwKE7SQZsR1PjZKoJTRayvykbqw1Z
YMZCz8iVAVkPPa514Ah8GsH5ZU5Ynf3L8HQEZZ/IDaQuqPbxOLm02FQGp9wEXNvJ
pudOh4HXORrG1tUEOtOf/J8QT9g7rcRpb5T+MGp3Gm7JciZyZdCCwl47LFIcrZkV
O2GVnC0rXNUTs3aVVg5J6TMkveWo+UMDPVSAmVcWpBTF4kqxY9aGQSS8eYa1LgoB
bUbgaoD0jw6FUbsDc7PLRmErujtRFksLHVvHq3OEPQ5XoBWkrir1CT9GSio/0LwK
zIgodXiZz758ero7r8VEx8ngE98yncQKto7TO3obhf59NxKQdQRH8DvzUcwmVdwY
sCDqUbGv2tRDTa47ckFNCH7owY77G+o1iZbX+LMNMeWwbd6Cn6d93XaDmDuPqncS
gRbEIk+fFg2iSivviZANOwo2DcYHob41o25AXxDWUOrnIszVlKz8qph/TrALSoxb
Bs2qIOFX7e7xM8zEG55ZLmLLrIzKEHK2+I3Yuq1F2ngx3Ub33s8rjMpIpR1GrBW4
Oz7ljSq32KKlz2tUaKHjD3SzYpadrvtOcxjKH/onqgKOIWTwYasT5aHR1K+IEL3S
CiSZxfXnHO/IBxR5zQwUf9OgNMwTaeGPurX1MNBZ4hbJCNeW388Mn2fPFRIfNsPO
BDt6eD9HF0qOXeHtdOiirjlJ4BRtYQguukBUkq8N9aAECJxsPOg6CMNp7aBoMGaE
HpRDWRXMI1clBqpn7LKsM1MEh/9aY6xobWFMAtVQETQPjgUvUUo7ckc6jNgfSlAQ
aM90aNgcvadjFVIY/DzYl3G84AMNvz1iE+Zoz0SYcNdrN/5Ut9QqRWXa9PlyAs3C
0BVBriiTy8+78aEu2isRvlxI3sASl8Dqjmu9GEiZdE5ZCCHWCur8tYtwLoIfhnvx
4QRMvelO7THzGTlEjtvGFF1HxZ3cul1Ix8/705yQm5RVGfvIWxyq/c0oyxr9HzH3
rjU3m49EauwYyaBrb6LqKJtluNHN7TuACFocAhRLZeTZZyTx81cGvhr26+rM8f/3
Mk0XmExu5JnpJPQyDOQ7AyunWRXBb779x6FSoepb6ECouSuhVPS7iagOrHBykxzI
uxHh+fPEhzs2RJOeGC+UyKA6tyFciVMFkNbGf+IeUcdNNB8nKXteXH6VLhWrxAh+
Nirs21T/rRK2tNqtQJphmK8iCHmB0I8C2I9GoPw942Tajyli+CQvHLy2VyXlx8vC
l9f1yzpBu0YYPzAu9AQQT3SNsJCMkl25FizUjuBT3rU0X2N4CeFZvNfHnM/8/wxj
Cr0PCqhod2LMTASCJUttDC7ewcF7/qY9ru5Gl/oMhc8CS1fRdz8qxDO9a4LebTqT
eLlxDnaPjMOK/WGlDUkAyyVlP4c6ER6JoJFq04ArJHKnfwSbxhGGh+KD0lH3N2gC
SyT0LX3bMIyWPVxW63N+hGLKhhlAhUG+GSxjnoOq2OR69R8HOEY442pSPIalRqd5
QA3BBbZV7h7r4v2RPmioXidSHPWZEVy3SM+gGbWaokNWWhFlrbgaWTw8U2l0WCba
nbVZG7U0uCRZbut+78aCcFAkQb4vQzxY/bZNMrofgkK70lYC4I7Eq/5U2u0Nkxt5
cvIqDhVtyZO2sTJx7CRKqeI9tnBuzOVV6HP33th4FjsW87kMc9T10TxztTI/dNwU
Bn+vDS+p7urDh6XOefrjL6adypw6KS4EAAy4x1Xoz6nRKh36Au4SxaCX/xSNCgSQ
/saW6YVHd6AOZUS57fGaRRg5R7BHpLxrt6j+VnYgO8lanDVO+66N01cCumre+3PW
Vz93mct8XTeAX8cxA0mw4xx+f5lxey55Rm6uTIaI6za99s/6saLx3E1j93B2Y8Jt
qpNYxejGBlzKJp57fkUWUK0TOu5DC3Mwl6B1QYwcvLBjuiPkkaB2i6rqiWl4NoZq
uGuTdXSubXL54Od1fAi1TK0tEaoM8SLaUR9E7eKuOswhFg/7Bi8+GJ2qh3G4H6L0
4M9/1oYnYTt1KF1p0FJf9aRmRoErHhqcWfL4JHoLKtJ+LMtHLSwGqqAUzh1agR09
hfNQJ/rT6gR0S5p9ZZjhQsawjpuMH5RYloCbp0y4Z8Wsg04ljsWTKycbP7sl9m2d
jAG1OGVjpGVAmgt7iRa+Tq6pctKPM+gHLwn91yj1d4WW2u4tjRU4DNqVoVLfseFJ
kMvjOw6pIL+/frwfamnc1r1ZfkuD1JmwVqCFpNj7PXx92Jd7AXpLdiioaSKAhZbB
oVmNlSTt7WuPhaGAWaBeKksiFIqiLHIHACiXpdTbLNAFV98wEQ96RcpgvLZmDTMk
vfQHh0ChIInEdhd4YAGDqsTZyoYr8Ki6J8bm/4Mg9jpoySYfkUdpoKsarwNtz+9v
3bzv/GjJm1NXODWxHVstIb+Jz7DL7s+U25Rrh8E4QYOpUsHM+WgFZUp3bRVZWAuF
STYjpQoRsSSYx/vY60Ai4SYwJ4KRppBmcB3wWYGgCHKYaTwefw3SsMzQvC+Hu8q1
Ms2aZkzN6BEudU3J5o2LAY+8NHd9cbczJThFXnlNrU8bFdgY5GA8YGpfNZOdr4MQ
BjIW64ufPUVajc1w4V6Ott4zIY/eTGiRVpfT6wKJZo3/U8l+QotDhuziD8Fb5hwC
3/jPvnM37wchOdWdbbfv48CNB80Q5Pbtl5NULLgizcY=
`pragma protect end_protected
