// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:23 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gVbkLzLpnd/6sQGUbgMDjyIwgQQbvEegjls+0wZlHpCMewBDbW/fKXlQW3iX/xfp
vd82qETa+uRYzN9fdDwKRvECu2Pw6UivICy9TVyEwMa6o4Qs8XcUUCrj0I98HHW/
lWGIaNlWIgGJ9SjPwuKcuzbON8yGcQgEhgt9lqKCcyo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17280)
5JJYJ5samKDaIpJFBGBa8EXpB2Ta0cn6Ev4/KUepKXvI0L2xWPhwj+5EybLBtqrk
IUlGymXgyCd6sXctEhZKLU0vmwnAdPPJVHQqp5Xbvi9k6bITfH27dRSsAUKuikyh
kUAlGx/zLzlyjgkPqwEzZjH0GG47Lj4TqRd0Mxhk/uLLHDp2U2mJKoy3ycL7idwQ
tp9/TV7memN3JHIOfxwHFihZvIzq9da+GYlRXlPpId7sdQsvRpyvZD4odPbJAbOj
BFf+b1qdkfZHJgI/L2W14xFOXyIEbtxjeY/p0zrLwsZcl3DS8FP9hlW6BDb/00eD
tPtytJSbDwM0VN6eCySD/IWoVt4eTzhp92ULutf9Hc6ksq/bBcCa+9TfJ1ZAzfCv
hwqTQNYaDucJyw5hDTYgTM/2Y97zvXy8ovpgGcEsr1xNOPhOm5qfi1hB+X+GDIgj
Zre9rkutj1p6ShRoNy8yfk+CtzzplVQ1ZKisr7X5DnhOUGD90+A3qwJ+v2pEibpB
ycI6Rr3AZXc7NabB6bdvj7sIYi3FuDkcpdGHTMI+IuDALuOTv8cJw67wEyOxtMKa
y8LS6S08qirFw6pIbh1D9KUa3tOjcQp8jvH8qruEjJ9iQ/YV2zwTXbodljMi4YEn
+CKpxYOT805i9uCvFAleR6Z7Y67jtwk62La5IfNkbA9bGcFBp/xTyYggTW33Zmic
Klv00kpFTpOWB9gLnH+zt8BwdjW+VGWE1s0vRonvYPa6rS5Gg/beijJjSgO/fAuA
TVH1KNdLHP7eKg/mLi1qxwx8s7F83UnJUsRC45UyMt/EMTqVTdES4AjVhJBP4UAe
GNeNOFzY7sZ93hCJOk1khh6YYPt0cm7AcS/wDXdlMv9Bg7COz5353DcHvXaZnZZj
AU35h8BAE2m4YB7EUpWwyna7WHDauoxRORz0GS1k9d1jem8Kx2Aqij+8bEsyudnH
1p/7ooWUwtgUuFd5bvirl5YN+H0ZFif+RNYb4TOc+UYMCbR8T4Lc8Aii7IczXVl2
OfGNfh6B67uQLo/AszdU7ppC2DC8I1JE93PnSgXRaeE2OmYrUp8R21mtrjVGt26+
ED59i1+UQkfH7ybXX6HfOCqD8H1EoK7LacWZrm7dslwtegsyFH2tNBGp1r5H9NpX
G77K0TiXRg7YwMiywpAt1j+kMpoF1HqvKK3VfeiTZGOD52PVhE1RKyI5rDvRtT+s
ASTgc+Peq9Xs4FiLl+4Pg18Ssb7zCD07vplLWIlzBKtTrzyWZ3nMZKYZGu/ST0Je
vOqEu8dv2LbWSNr6bHiYC0vRpmD6alOVQ+P7QqGiojLpntPL72NhlLlW42XrzZYw
2KjCZbi+rHYNhGBWwZgCuVto+NbvqZwnprFRyeZEu6YpTeqZOnuHG86fG9nLtSVj
WZnEgS+C10l5eRI9JaxdAez3Z+1fKgDW9z3mG96r+ZofUa2R5PG4XFWvHrNb0RGO
2B+AyBQNJUh6FWaU/1EMu1a2Pb0m1FfEhKqugKHngmedGAS4XQ4GzhKoG2EXzv/F
Goj34KCQvVe7eY9DWhc41SayJcUwGeHv04M2z2PID2P+KrGyh4QVEYq5uYmipGfo
ryYa68IRrRZPJBK0aN3SqbFVlVBwNLlPyAzEMcF1UFcO0lSyZbvXrChrjhtufNPF
1DKQwvqhezLYjkmt8uBDUqUhMaXYmwwp1JviC2/81Ac33smxf0g2kvo/Jsqt7WUy
wh1TYdOZDtiRWP2/B1207jGB05m3W8euTI9RVcwpNnUPDm7G6CQNrwFYG+vKhxEN
KeHVl0gn+YRwB1ryQZeI7uELXtjvkaLy1moW0GVmDuDDArcuGqJm3/M94R1AwtUG
XwaKSSSoLl5MpJTOT3B+aIQa6lsjbbSQUjs3shIw7Vfo/kKW2F/es9ZGmFgllzVN
fqZtO5d1zpF3bwM0XCvSUp/nizcGpmAXaz1uVkEjCOjywT1mX3HoLYEdmjWG7Rgp
VB9YBZ8rE/JWhu+KzEnJW4h+C8G0djhNYkUCQG/amAmrJygMlzNMt79BEImUUNwH
6mgqhbodwF2S7jYl5GZjacBJcBVeWig8iS0X5g04LEe63FevCPe/5cwzVHe4B7iN
alUOiXwxES9SCnXWQItCLoTmBgN/2ocsdp9KeMhHNPzgEaC9C6tP//tYc4HCGXBN
gpV/gEOQJVPVuyHLLEp4rf7KlixDyeiECZu5bvRBMVnC51p8hV2YgIW+Wv0Hr0+W
+dH/MdqJXEXU5av62+cMpUq7EDC+JOaRzhy/hXkzUGEaUUWl3qMAioKfdwhT9ZbY
703qQSeYEkaAEVrGoRpCmnOMn1TMxCu5Z6Ork2IdINE1ajKpBow9OZe1Eu+ON/Ey
4KWl59fE/qa/UXK0aIEYIKXdxXmBj+E3bnkIUalGtDKRZqjluy2PGqj1ak8pT5ju
HUNqdrzuAkT5NP7N3dytcOGypw0aCpT5gVneBUPe0GXfqDpskH/fz9Bi7k344WPx
+BL4NF8oiBK2Ob+i8rCHNlVBnuuD17+xAN9haKe+jh1wwHFc/pp7RQe4MRG85X6j
ITOnY22JxfMK2izc9CUbzqyV0B6qG3p50V1G7Ghv6/yv2daueCRoLcTAwEq7Z9pm
5JmrQ9VVjgRopyIPMl3PnlfE7Bgcu1P+PHkvRicvIw+WwZY3Fx6VTs3513jxAX//
3EgFbp2Cw6DZll4BOJ+4hCFh1A0CXWW6oWYLk0JKH30CQTk1OHG29twRLv7b7wDH
qJqgrkZ5rAYkgeDQRhWQWUdU/dU5JDxMgCBTkQS9JQyAUcKAd1daY7Vl6cnCEmKI
HN25qIFnWKewcqMjLRJn/RzD4mZW3obBF1OUUKHifDkkYdkuvA0vvjGMvLfN+2VG
Rcpil0H9258/ziSV9GHJINn3Dq74lrO6riah9PGvxnI0VJZOhmoLHNUdtoo+t2vk
ha/w2hlV5yZHzm+CXuM5EI1xo8FEmjFmTSAAjmm9vrWnaUInyys1KJjGaiptG+yI
GCSAeRi7uWPJEhH0Zn+/Unq4uhZJiUdeBUpzGo/CFm6tVDpyOX9ZNn/DHNpTnhFh
AWpVtbmiUWG5tV0DmvnUJdYgCCSMen0W8Ym2CN4+xA69WHSMxpXxmwOm4gZePWmK
4okN1Iz8mQKWdcU065y+YSmcLHBUIbPE6cyh/9jE8ZzwRP3hE6Zyiyb18kRa1nHf
jx8NPsxHuNJS60Au7pAoomiNKNsVnThQi6ilFMLezHzBPCItiCmCOCm4kBU/UqhJ
di+bzd5p2zfUe/xrxgHGfhON/oFYMLbxEnWpgCygU5sbbdLwkspdUlW2UDrEt8Eh
muY1Lq5eCfTTMU3c41sRNsHxXCxQfwVHWY703m3wnVYG1gDnMaMVmIIk3N5LH+ln
BbNRGAStzLDgiGKdUpHfQxNbi+U33t+3IE6StcJQ2p7xHVTRE3SmVHgqpIuUagh1
t8St3jwwZvK852UkN3QgjWkRIuwlRml/WOOPBRSfZ7jy/GHRcrdH+gsmUp2HFk89
jNqNRYHEyUCiggTxPWE9s50LVpE5wormpyTHYuAhxkLpiQXPQQcy4Vpe0Gbd/cmN
JpEySr95/LqkpVvUvw6Wqej5h5CNdDkQ9z/rt2scDoWHrkN//uI6Z74tSP970mNm
S8vCtjejKZl8Xn8cIXQPt+onDHHO0WIEv27iWfF1AqbegbVDiJ/tXhQlKani8rfA
Fl5paugE7Jn9HqInVbTyYJLdFAT0xlv3zwhJuSKAbpRishI942DgPwWicd/TUvCD
oS6nRBVH//8WJIYNJVfdRC1axJ5LBKODjKABVv5sZER6xIfJHaxTZiQTRsT88PMw
ooO4WsvK5YkbjBgfknMXaw1ZbQGB/04TXycqQkd6E/JefG3jqtJY+P1pm2UUIo2J
dQjygHmYDVwh/w0yXKjsrT0NX7Y1sIsC8PonhT+q1WEBdKamfxsgqNkDmGthF4iA
4j7MwNj1nhZHNTm+3ldiGNpHJm5huDGaqk9PwCFnY8TGbAM1oJ460f7nQbwgOyEl
zJzORiBF//4xz9L7rpiPwnwYq/V1dbVsWGGkyH3eJCfFxBWlXtlr7TsUq7snN3nO
CL71lErNd+tmYT43JDpQ456n5JbRGf0oypqhnDd4M3bDdS5kK07fU/BAjiwcoVp+
qOcN8P96ngX5+zEYY5lZQY/XUXc4D501hts4mvplhZF+5XqXqYA9mtAh06BBPcFL
zp9o8Ksc5zIZQsXUAWEWSN0rQTAXBpMmaqCgOpIbcijc0YrFOk3/ZudfBbS+fvck
USteWR2qC1ImkJMMkGnLicqpo+YTKYCJQG2qU+ngXGAsGIlMqgcO2Hr8GykoidTB
g6VjFbC7ui0iRJLsrI1YgJ0zausbGjldaYrw5V6xO6AU7RAXq8edkL5MJ9p+GtNp
MXyDcYgegA3rKR8VMDVZ+o8Zl4260drGpO1bL5SCeYXOqitVFzCvvJ+Ih1n6AFjT
hAJQtTKTtJEvMmKngTKLVm/gvlxQJIgDKGKpt/D5eOsrXtB/qpeZjnH/HFNpb9qU
qjRGbHUV+t9UAXcHtuUvOesy9wIBgeiCToji16TSAcRvdbq5Kb3OmmmcNm7uRepA
+MOwRXZTmd2B1NnUH3CK0T9jPT2nt+qDoI7w24Xflfg7Yky0Qct2rP7h7ZEMDud8
CqQGD6V7+IkCEiNkMbW/Z0xZkjDf0fFnsu4swPyduhRbwaZ1CjT+FHXimS5pKmsc
l/gl4rJPLHYtgeZATj5MQ2aZgKA6OHj5OrHc95gs9hgHzFPtU3YM9Jd8D+fdy2uU
hlS+MBsk2jwvTVnuqLBPUhqoml7NX8jIxIdxIzGJMS773MAyR1Gii/shmWP4Jgcz
/34YMn6uE7MYwwE1z++TLyiGM6JbWJcLqn3ASnoeIqVrCCi7c72bTVbMVD0ah2C5
f7Hx5D1oC2HVFHIbSgd5nXVt62UVJc+nW8a8JCQBnJ1WxvpzcTXiElJhHpg2rFkK
29zfnm6+mbDv26DJ5zoGhpj/YYUfVdQl2De5HMfXDch6HbOMx9mHYANA7eBGTL/6
tSD8kAKnwavoIVZ+RBZC8t6R+Qthk6Eq1O3Tv1xmul1/o0W1pQZwk6ju5dZvCXoC
foDUkYca+zCvH04qaVqKvb3iGJAQ80MUfRwGF0kKiFQU8MZJeSzqJLm867Z4cxL7
YCRLG83NbSubh5iiCxSnC4WDO26FykTyN2mCGJ8LwWed3LLu+ll56xghvNbcDECD
z8iozuF5Ef1p26c8rjJXYwpA38f1Xpn4Ox/H0ytV5O31lHwiy6JctMxMAK7oQNOz
ZgP2Q7hSSvpdwdX1tpnDdlPg9tybJePPaohqf/NbJORiKnQP3IEXZVdo1Y7H0r8V
zaFz3vmV+JlOcV+HEgdNle1NDrv3NqUZEcwUIr2cJ2EFpPWHxNsxQ3EgPd5Nmsq8
jbeGRt3ex2SPICszMX8+7aiBKlRchhp8Cy6zVoCF7yDIIAhcBr2ttpDnHx9O2imk
Xs0wMmMPR3pcP5oeWjjzKSzCdi2WOghXlrsJOzMENk1R1wKtSc96jgHuXy6txafi
kGGdj3w+e3EKpNyo3jFZN2shwYvoyZZSFKow7G1wesazRP+uas0PbTuB5EWK6bZv
cKahb0T67wrhSublIwlsEtX59OPCuifI/yOKupjUcw3WnYXf5g94MVjyg8IHLm1i
PAPLOGjBVFEM2G8E/T2AwkPeOtk3SeMPQy+PMIsUR4Gtlj92INjI0hsUp10wc93D
MBCrnacrqGgveXuQM4MIdmKVIA9h9qJl5CEIrGU655zDD8nmmjwIGxjlQiiQDLwN
zfX1JdYDZJW8E8vLwe0a4QV/kySJuaj4OaQYxq6vmxY8Vw7UnY7GdIzy2GwCOWcZ
08AcUnJeOEIB/lE0WGUICXNIa3zaCW4ct6KOVfqBDlrgy1MN8B9aDcDcx50vXiq4
FDRQ4zp5twSfF+KschtDynyeUztnTDAh8ZPBrDU7I/33ihQOw5d4gMfyWv1sgstx
E3rkB+TIetmOsr9HwIGmhMWuQtziPNbAsQ6co3KpnsAORyPxcXAC/Kh8vL4XZ+/z
WgBVVp70R1gU2PPem3PX52IYdKyTGdYU4et+/ppwLWol1houNXVLNdbicYqe9czT
MUIhoONU+emst7CiGL3EkGVLJOA/HjEGlyMOrgBE96QMmQwrsPTtd7hA4uwoW3ud
9QxPK2ocRnc/J7wtGigrOCSQ5wFI8X/6Kul/q+Wccci4VbGF6b2WLU7yXU/v6VxE
HfmLSti4LODXALQPSqnqrWy8jIFXKyD01J21p9GtCIHmeCBXxkGsydfKN9cVTYAe
smvLaKFkO2I5HPbo2Rqd+beG4gdoK/k+c+Gpidl/Q8u1exdByLceOSf1CQNrLVRJ
mDViVB95UeE5bbOzu5WBE02HpuDHDBEZjUSdRknQzY5ySuF0pWRu7H0JouKygHJz
dXkuesCqYw6ZbQEqgmSeFupEcUd4vT8qMfobhPIR0/n7ZrrDtHuKYcmrFv79QV75
4gWJSN651q8Ti+xVH2NYK5L3pqgQya9NF9m3EPjvcj0Q0+hQmGqkEmpxpb5+kwx1
WQK1Dpt0yd36X/Xxyo12M4ewE13PeH407tN3akZ95GMva+lNMl97nI3/H8wl2Tk+
IUXYxCWTw110AzXg193Dc0A2VtuAbDCxppia33q/2TC/QvUB+52K/58oqa+hrEKL
StZYuwzUgZGiDe0+rw7C3ZvLwxSedLAnHwyOGUHS4B5n9Q92O37cim7b15ENp7G3
iNsneX0Ze0pVDZY2PuaXDbRb5LmLiYUiRFhUllfiNcHPaCUDoRmlPdbalkjD2EC9
+kR1hQgJfZ+Nu9Fw+JBP2Q+6iL6tnBZ5/lXA3WBvwT8kCJ97f+lZUZrNfaSjK1mv
ovSdobpuvbhE57hTTZXPCbYWiAp0TxF4Eb+I6+/HWtPivWmEZxAq4WMx6dRFaQ9Q
Gms4yH2sgZaaYdVJn4hCFf/tR/rmO1vdIOcQdHbgx0UxNQiVbBFTicD0UexOwi3e
/qV6hFvYI7+e8D6/1zxhyUQz0/69q26ywjbw6ewK3TNeXYEnhJVEX6w1GVGrXdfN
JpxKeLt1KR8nWOfuhw28rImZIgEH4JJiD5yyrUQlopc+UQbVREZky/9dL0e1xa2s
DrgssVT1jT8Vd+I1rlXSqh00G5qe3tPtYQlv0h0Ci0muWYWgoorb9OgyJ2UzWFdz
WYuVS17zDsg+H3l/D/8+ekOg8697aw/WDgcQj5uTq7uKqW4G/qXLbnE8Xckh3CpW
qacCCxNHIH5kdDJPmqFHb6/8ejJ8+MYUTOwLKtc2WDAN+/pc7Iifxgj32+yXLRZF
QAfniE9DOEZtXM8hRWoAQ0dmE3AGJOMdAXS5w3ZEE+NevhHhGsdvzfcQbbN4tips
LCL4iQcQn03veyfsXr7qexRo8tBJNgUsiaOM8GJm/m8Y1Bx4fSCQz9VZyPRXw1AD
5HJjrHUoHi3ARZdb3vlPsp8MKdo/hNza+12fRYJ7Cq96sSWenmTyjqirbEPXuQ4d
waTNKMUcUZVSZSGRJpd2qK5npqBvM82Tjd2IA30EVMNWSWQKv/CYeo+u9YiFLnIu
OWtqndq93RCs8Ka4aqknBKTwfypLnWzkykchf82MkExPgfDYbmfS8iPyqjQKY20v
0XZAJnirkqyRKcreoNmjr72NCTAs5+PIM+f4cMTUOd4I1jlE+w0d4W2IvZ2Zx5Eh
NUHFMAJpABkmS81svDi1hwddYDTm83h7wrAldXE3olbo18Xo2nmpgBd3Jyh6Uf9D
uGB/mop/yNzbxYNcx2DO/nVEn4HAE8pPGvsutaPLnBg/2alb03ZUI4FeDjQR8qjA
axVgqVtPYGhmiReMlNQF6kuqik2lyN70ex5Ijtod85C7oC/+9uieLSd6KLNSxgWU
fg2yuJc+Uvgnq2gr6/nQYGdcfycz/E0hnPjTu22Taq5UoN9Xjw5u2/ulO8lD2ckr
BFu3dGLTVzbOW2TthZc1IEseIcAfu5qPeM7fWqYkHXfBQG7waBFU717lRuWZXzDR
sg75yGBLUsYAJ24kx08/KERQk1+jfm0D9DBH0Ot1sb9iQ85vZKZ2tZQzcRJ9MnON
eemai7L1yb6rc+yzZ07RcHSW7dTG3fXufGnnhecOsSVx2Kk+2K90NjqK6EopilU+
FM4MqTebMNviZT/vIMjy47l7DpsxHc0ZgDtZW8AWvhuLUbBJTSyT5TpTDCbuwzs3
16+Qki/3yTZrEnIOHEplaED5FpJUL7iKiyBqnQEewSdraN8fakFN7cuXaZ+mAn0V
xuZOA/4V2ASfVrr9VdOBGu+y3rwpeHuBYcpR3nIDHFIvWeBK9gBLsJ/IOWt2ZeLL
/UAXLqndzaVI8/pm4SI2EiGt9rAdyr45l9hm1GnNTE/RIBukkdxAp1e3nqIBmK1B
ZZOGiTpnqW+sKcQLeICnpAl+1qFZp+nHcpSplypIMWTgLybX4bsI9jq1YTXh8pRo
Fl3HZGZKO2JIxm9BDZogS7kswWmA4mcIG0pFx8sLjJvt3B0/Mzz7qpWRFNNTJF4P
l5tTS80tftlZuOaWV+8sQw2sIfl0zmjIHKftXtSw1s01e3BporcLhQjd4hGLyVbI
0WTpwUzWYpXgd9C6xTVbVBrS0+PP667guqtWfam4yi5o2gL2+9RK5RQRelDG0u/q
xv0UJO9EkyS26I7v/U2dVgERveNEYTzaajq2cOA3ThQe1w2xs5+v3Wd6UnTBT0Y5
PsuTQCc7XNygll4+c3ohduxVGcz7CPL4lLIP/20dUakoYV5YsXvvA5P5QAD7rTOQ
hv7aowDKCRVeznfnkmn20MMMJni2cq0j0gIE2JVTTXx6Hm+EaVu3YR5Mup39CJca
+oJ1e5uo+C3F8i6t+kbDUBy/hcXUynpYE6t3ywcjQLh0YaoI7HgTNO2nx8TwEDHw
mFnpOq4zUpT0zZ9RmbhXkbRpWox6d0eb9EytkExn6JOxsrmw1JzsAYtB61O2sfdk
UIVicTqivOfZNEqaneqMtUnamm4rGoYUgcpqZyhOhsQSLAzWts6xpmXWGqXkWClz
zAY6Sbq0Hcn5oa05DSsbretkc53beELdHKxtL2ub2XfJCEkR+Ssg36cMgF+7J3K4
4Yc5cngArCjDRSWQHvh9D1Zoma99RxsuXrV9CgOhzREz/tPLlJWAe4kJ7tHWp3dR
urVmAACSrsZqltL/4BKAfJB47nTjAcjl3qW9Rb7bHGAB0+a/mb2e5UvNHZ3Z8kAb
7cvnFhplBGV/gjavlUuGXb93e1HjdyBYwyyuY+DPDHeSQ/yXcDTgW2Q6MTqI8MGB
R3N15Wdvkbf9mWFQ/FxeCIHYqeaMjzVvaRqrXVK7JtZEDr9CmaXp52kT5en+5zvA
D0FSvwmiGmyQO5F1CrRP11hLTjzqqh0roJuuvrOIne9A6RWbsnLFFJxWWSnobRSH
wnsICbMDU9Bi+5xJIRrmeruYICpYWbSjwhv/iytGnrWveeX8V1XDdq6KAbE2HNz9
qRMRejCfvsdffs0UFf0+wpN37P/mCCOWiuD7BJtUSLkeb0pPB10ULGCm/oi83ImN
ZehAt5fNWOenvpdRuy5zKJJC1jWEhbUquuRHPbZbNvvZ5dBZbS5Rf1GNKYVnKNYv
1nxngoVC6wcvQayWMYm9jJQtiScPT41CNkXJX1c8khi/lVXzKDwT3zJ/a/GiFKEc
Fq3e3XcnHSEUSxEfcFQyXiDnhVY6cGeiePbkLu87o6dJyxqpJP8GQppd4DJIOhxa
31HQ21qKfQU4P8zVCgHyp6QKI6hZ8vibkbfPTEp+92psa9w30FLWrgNYHlPYKkQV
3oDuVY99YuNzt8d/wSi7tsxKrBXBqFSeDK3swiMnN+XEbr+iBJ2Yh91ao0Zx11x/
eF5phTSj2TxuBTxDyF6q9smQ7PmDeVPkk6HnC2inzE1u8lFkipl+Rm7Kdu0yyZBu
jn/o5s5MLaJ0NHg7sOwJEPmygSpd8SU3EPWmrrp1GpWKZvyFxkrKXgT7KcUDnCU9
YpkGYR692HixJJgszrOS0HAGaNubkYq8nSyt0BhjKB0lQJgpmGNnBNhvRZ1KVCZR
o0VdMnRtqH8NEp8AO56+C6AmruMeqIWwdtcqKGYd35vR854cjFF/xZLLN33LL6DQ
T8BPr7fJxzbmM2RMuaGkP2S2tVd2DEXgJBSYFKqGcCTvhLWCL0wyh/yBh1pQGgTn
GR1FnKH9sEJfXFh7Jlf/EO85d3ThZTtCQzMN2POuSvSYlRcLSSNqbpSE6eEd7Tuo
FJMqbw0e+YA3oY4JblutOU2VZ/xkQqxUdspt1uecn7fZwdcOGr0h2zRFwnSOK8op
3NzzoumhmGS59//rcYSyFGW8OnmXRlarg3AflO/tXWluWCF0tCB4lGJH4+xmY16f
InoN2i+Grm7ZLUuH4KOpYuTAYkoihPgfOoCepxyU1ASTRW07+7AyYknGgAvbC+sN
McQx8cBKlGCcoWuLqz/qEFlGdPzatLPylNoUViPINttZ95DwuCtaolE13L+t56Eb
MPzNqBWyHUjOTA6O8UnFDLvkuIwJcSLnpTWg8PHEtlpA9hQRd4giSHlkVBfTtLBV
f+evyp2y02c1gP89l6KTmuX17qNtSKXugCcMz76A0MfivxdZl7mrdLjZsKBDi31C
ZkWY3wcLRWS8AzME1eoIOj14TQ/+UdRn7aGNvjOjTTP7xMcAqPMejC78nnd0xqcd
YqasC3TW5tRqNPRX6D5yQRiXJHo01SYQcXcJeCZOPpyyjWnxCwD1lqgv0ovNWXQM
y5CDMD9kzkR1zRiPVGpW6s12fAX7lIn+cRo1q/vrJ+gE5m+eGsVHsprmFtP8b5QZ
P0Rbd688i+jVt/wspP6kuwNqiEC2uxYNYTls4uHlWzT4wpysBlXfxXJlfKvll5IJ
Nm83nlXQjWlRRnVR0EbofAmw7DRp+Ne/PYml2USN72kkhxfLtCkIMja0Y4Ec5DDY
w2mgeoWwX3l/mCdC51XecowGTpQIN2ENnLejbC1EYUl/hioUDJXJv8IeapYCkA0d
ZVTsuhBwtdi9L6WKXh5+9sONhXJrGd9bQv+tbBz8Ioh2Op4cIY5cEf/DFDerGLLI
FihuZHxHcir/yVg0SZUHjfmqXBtomVLWpZJqQ4IIjDWXmPwDXARNdaGDNcE36/+Q
pp74NxUzUP+GhPy/7ihVtbT60zb4XYcsZo8e+XxdnGEEFk3aOR5yqgGlcseoeKwe
yobaa4iogYA5m6CFI4zHdVXwKJRBghjwj2wRfFFvTV4/vKrsEB/MQxbl/oPIxGZz
vP866+EmLUs9zwGtNvP8qTDjvu7YNE884AaP3ISpmLMPbRS/zE+/HgDetTZ2dzaw
Vn13LOE34MTuo8THZUMqCv/+gj7K7XYUrSsZt3s88P1NZqmrG7kEmBcbmjvfXpnx
dwIeXS7scf73ew1C+0g7yct7wPmlzQMhi/i2EiXc0i5WOzDSfjDdVBOtHg8vmrOC
tHQWOdyGc+1ZKMpNf4b8fbG9dIgzwATKxj8b1GOsQwQvCMsncYcipenGF0mk6jaM
dXzRwABBhR1anCCPGQgdvXSYGuN/uZHdyIZiPBQdQpLaVDDd0KOS5hW0Kp6OfeG6
T01puVEKB2/bTRfgVIqw7qcOetZX68H8R1DU79gBC2ZpHa/uBtBCnH/mNoSNUr0L
HjfU/xT0MdSyQRVuRNGrRGNopQSSg4vEd9rGih+ek3X1W097XmCSsYcjiDTFTiad
iPpoQHEl3klXxJlcFq3h5v29/EpPTvWnB+r486tQveE1O6hHxjzqML5iVXB6Rf6M
nQVa34Ncw3MU5dSjlTr0+sJ62oMjCxCioWj6wd5o/z3wvhYcMYY8nUJ+355jnxpa
HMsA+abr3Kue0325VUJ9Q3hFEegWOcWauGO1wHUiQmkqbt2C/szr1m13tM12lWgb
TOGwI9tGUDLOCniBcwCRyNxT2pRiyo3KPRWsHwl6eFyo9LZBDzS+kgJSA+cn3ck/
VSDkLql/Hh0gQ1jVKWO21T4gnePYrI1myEQlE9CnCR3Jj/m868KO/5E0d9FsK1vP
+28k2L7KyWdG+sdeWBug31RrVVZ+HlxlcputnQF+aJC4Li+YSeoWVjxhuWtMcliP
TjzudFXvQcSEqVUxEYtY0vc0uImPtm5HnTsH+K5CBw3NHaKlwyPeGOYtA78oldPk
T06O82zQP5n/uKZ/7KZIlWp70FCGNBf9c3QMeuxaJH3esDLzBv2RTtFBUiftJ/5M
681PC2dNfJQZ8mdgm2Tk6gN9sVqpUKG6JKsjcGgD3D1Bc/BXzckcX6xlDLsmt9ZF
rg/i8VVTvJQow0qqzpEieTRQ1yEIttQ9sMbRJqm+byyRmHL4f4IYrvaSgyl/IBt7
LUXsBm4yjg1Khu6kkCk4o/naHamtOf1A4WxYKwPKZ12QhdeB3aNCtSwazjadcBf4
vxxIildS9y/IMk1bnFBW+WM7C6gCQbDJ0B0lfbJ3QfxVzN244F22strUKNgY1kuP
Zwa29ZwU8GizvTCjuxo2HJ7Oq9EgIOu0aYtiUjP8jbv8+0BBtMkPKFFXMtbTVfyu
b3cR1MgwVGczX1GAAkh6FOrvfHZaEfVVuSChm36Otf51MitXFcfWFj8ysqV5ZEo7
Zng/AvOFgwpYM5Y6VmoQ3tuLGuCFZFwueuU4MMqzKxDV1K7nfKL/A+9pA856nxXi
uxy38xB/sbpwWnAsNXQZsDuo7m0VOppR1H/0Ms5liOmMuTLzjv5F9mwwL3pDA6uP
T6XG4Lu0y+Pw0NGwX3BRUN7svm1m5ckN1QqRQp8Je9ICDcWU31VKqM4gx3Lorsk4
hSO/bzjUx3b93vvp+1+Es6TIzKiSnFYkOP61BpmGaAn/DzCvBdFMY1lrATMAxCRe
VbX1KpqE1uW/XKrw3qeWK4IgcSfxQg902xdbUuYJC9MFoft9maweCzOwNCmzkEA0
zkILZx2oidLXJFB0aJNpX3qf28ymHV56QN7giMkHyG3gaNul0qsLhGPd4SJgxW39
KWpOBvc1CzYsy1NvEpkiDt3nxQ2NyUSlvcLza4XEgPVtebg6+Y/knuwr0pH7A0CN
BdGsK9g8O2LgnDHcofVev4vDQzocFZYlksXMkZIhatEjhUoocdyrJP97wPIigspx
msddI5ribfLR1TnTlQBcS+QxzyH3A+1N4vRZTOKEwN+fHYZ9QwH3Z8lg5T4ubs2R
GoUdkJcb/84WAfMxFWmgih5IKm8TTsRhD1lhTf1ZtS8Ii1FoLhtHs982Mr4w+466
phLl9Qa5ETto+11X+hD/7ogBdFAxZWiWgb/JsjcuBb8qSRgaeSMwDtQfnySvKKRB
yqzlMBbJ2PEWI7AnAHrJHwcuHE4SI8kHTTFpva16Y9ZSgU0bIbYXQ8lH2SUFrdrF
oqcfWrG/eilKI9Q8+ihBFOBIxzWi5PureOAT93kUkJpv28AEJMtTkRFrXnHHtEBq
qOJuotfkobIM3eqpyjlKNAAUyKlNij4VBs3LmOaKZ/kw630Pet6RMMWP+DzUuwJ9
zd8TnGnSN2YM9HfHVfVdYt5nT0QfWHMy73nZesoH8bUHokwhZkzPeEG1wuPx1DrO
W3KoepmjksQW533AuuHa9Qaqw6ZGvmLbKM5ZU/MW6c59R5WzLYFXzpnIf8cZosv3
Ia8oLmvv2If32H1CemW5jgYPTyOOIfJN1E+QTFSF0jF7w9PKY2VhA0/jCufmX3YR
CdBfVLwafUKVHzx0vNCey+5KX1BJIA5l3As1adXtaeIzQhm+qrYr2zD4yXueFWG7
nx2xN/kpCgghGLcFvKAdZrYQHYMBW87cIqqSu2Bok7tlFomnQThIgcpqZrcv77S9
9LsGBLAzVa97zOn1SijiGZL8b8QENIPD8QXtayqjvKkBqzUQ34jIo+T4+u2DN2LZ
ikuWxe5ievTMFhZ6MA9A+DybxWEBeV3VcDlSlDQCDu127xUKg3GRicQ4PrJmf8a3
iB5Cyg2uZXXVKWBRA/QiItKGDRHlwHcxY15cUh9UjYH1MnK+V2mHyWnlr2JcCivs
JSHKegeAlikcW3lL/11drEIhAAxPs0C+mGoZ0e5xBt/JauE0soBVWyqLPTT4q+Mu
mfvvxe5b2lqV0cS4yZ4q+UkmkRJm4pjTJZ3r+I5DOZDIHp8xkrLGAQBxpeU4hIJZ
ovso9Ltxm2ueBfTWmXR0XXYCw0bp7vy2icHdiMYOv8Odo1ctvjZx7iilPuOmHDWM
3TEyV1QD7wa+VsSs85jqYdiXZiRAEFYwqW3yPsYoPgl4n06pYcU55DLudMRJoRzy
DZRIZnB0xeod6rKI1LOjojq2Yro82SfeOTbkbzJrM8PXpEOLCmfWQp28MVZeNnI3
LcJj+MASEWZ48KWv9HVIkyjGX00ldzl0AOJpHtFYeqZtZGQnoRRFVbeHEl9ReKU2
cxcJkJ1eDRQ3wG+O1Cue/expyr7tbtgdd5jlVokIzDpZFG3FE68nNft4UZZEUtcU
SIjypp8Oo5OvQJuRtJYqmW4nZBgq+EAR2+gTDc8q3LdbFLQp/qinkpZSqsz3bCX+
NlP7yxhyff9AcI0UmxF1x4ERIkpYgSmmmCNpYBHV1JYUpk3q2n1Jf3XwXgTCV1pH
y81h8fZmajg8KkOkhbIETG+sdMdqo9N+X8IVU8rUHMPISH87gDY/D/VKAS83hi/z
R0aHDL8q3rmkTok6KBs6BfLhGUHeTGl5MQdvOmGR5tattP1rXfQ7MveeVcoHvLdr
13rxKzzN53h4UKXGBCXsyCqPm5WxMEWWvDI4U5vNuKtPTbkvCHc42N9VC1sYKG47
BydkkObYGJp1MGRuG5Sq/WTuGbn1OGwhj0a3pB7vXarTnfJ6Swb0W/fQjEPqJHb7
/7+sy+S2rtkLBEecm9lE9A2Lf+wW5MHO9HDXYxOTXA7i+2cqVb4S8Ql/ty96gXBW
P3Z74Ad7V4KI+wkh66ELiEhMc2Zh7Us7hZoefiWnHx/UIyhqHeN/ayZyawE+CRqV
Z0PgOiOlFlVu5kUqXKtJEB+bOHJ96GFQOfCdsujTNO605UUGQg8bf8VAIqQSmVnx
H1NJXA5nTtH0sj3pAxXr9wytwXOswfAvDlfUglnyWVJjosE7LcNrpThJmrdA2JDI
OjSuCcGX5b+QJ+Tb5ghFi2y0zFKeKbwlOl3DbfaYjesNWooGbPUJEe3Bt3Z9vAFp
KKoS+Z5b7lvWhChVrOGhoJSBbc6ZbRbQ5nnDdyRMTCE926JxSQ6rLZmxxU2J5AEv
io+CVu+wvuGQzCDVixnApYY4BdOtiBM9GOVTuAXK+W8HpRdEN4M72qVJ+e7X+I3J
oPv0YCh6YuQXXJ0KlgCXJReLoC2u6Zd9P/aGlNEQkWFnFzcMIndigoTVjYs9gSeD
PT/sB1wB3icV91+vGph/Cib8CBe7UZ9nuDYmKOOB843HjQ9VTsYP6RxcyEFvNlS5
DDrmUU5z3nwF7542OR8LFplaUGZ++aJ9qKJ6h2zb+HR33tVEqPVzuKf1GWg0VIUM
pAtjlb/aBIeHBCc5mqrmy4ASGOFLzGdHk2A/oVU3VsCKlI7uhwc3OjoChr7wVYl8
at6aPR74AYgpeB6AF70y7ij34y/tXuw54xDDBJGqZefYoxRFmVQzmdVOYSxw2LHU
oTfNbA4EXA9P9cWkKnBSjDuF/ilgC4+zpL1g7PO0cc1oWYS01UOqEECaMND2MMY9
xrlDYPqMRGzr0Q9zbIGiFXZCCcSEYXd5nghsGCRIrKyLupRJmIXsDBTFojCef++m
A6cjCaAQv5C5XCzkXoegUXaTIRIVxFVq4bIzaEFej3dCJ8LyVBxdId8NFvOJENsH
d5KJdeDODQ81BsKoEV6oG46eK21/NSIz8O86w3XqP8t9Dpuq50MMEMCRfDs4ENg5
66GZ/bja3MKpql/SzTDlccEi9IZhCHDC/41ZGSxO8yP5PIGkpgzXb+Fgv31rAlpm
03U8RmUqAUKEMbQCELcwOvVAYzIaqtf/iflF/Msnpp+C7p/CItQ04hP/IkOK+icS
BEVng+r+URjbseNzd384pn8VO8p085dA4eGU7tGNP7PqZvuCjafnaNt5n1NKslmv
wknCkOFAYM4eNkw8OZR2hbtKQ9koo1KLfVZMTVpiwMMqGP5tqR1hDWl8Oye/C9M1
evk9SV/Ax44+JIIazK1amOYr73NEoZoJoQ8Ms07nIIKLPMWPYA+fwE4+WIDkyS/U
ue3EoOFQQVEvimudnZZUOMO6hOFizmjSk02YvvdDVUKQx8CK3O+ASSShsZ77YR9y
AuKOvot7FhTeKFoIc8nkCwVEc46aFJAXCfRRstFbs2uhJ3ihkpcb/1cWbsfdcXNc
LJoQ5U53R0EZ4j5FHOldwxR3It78VBYelE2bNe8mj284PLdVsE4kEqwv+gFSvjjx
psaLv1jMLf8TQ6N0IRcEWXnTuGFyPMosRTSRuMbZ4eb5dqlSOc6N3Tfj63v7Usi9
XbP8KHiFhuHSmytJ3gflrv874kQO/uIlS+AKRpXK47mqrOkdPUs69ZmIz6tRev8h
nc1c7PN7mTQmAlYIt+JWsxLix5cRh3/5Y+IAIDJdyHLOiwcQsL+f9CNl1YoMzahc
uhDniJKYhkxl8AMSGfKlvc3WJJJ5lPFkG2ePA+fm377MyoDC/PULCB6KvhChtCou
NHy1oLlKe7V3+MdQ56eYJQxTTWBHBtBHh0cpnXZiwNQKJuXR6Q0BpYl8LbJ3tAF7
cN0LMUWCH1DeDcYwDAeHWnOmTv8xaV7Pnzh9EDJ9vj5L8GKUKsoy6lgxZOGZH5sP
jn1lCzeSHSlWawP9Og5XrAaT495UF1UKo6v/jT/C03opFgDxxzGejXbXqZzepVF9
dPi1X/eeRDGAeS58QS0fl/7ZAKiduuAR6g+h87TnuXqHwJVVqi/obhUePqu5BrbK
7nGKXd+8AKSk1Lpyg9G6fdROuTCqk/1mx+9+MaXIGIA7aJFunHJO011qmbAR2szh
ZYK5KTz8BpkgLS7VnRabY2pJkGt3f3tGr7Ru8szkLs2QDqKWOs6+C0ezJ2UHnynx
YeqqH0FlPrjVch0Mb1e4viOtLx+JcT7wLTsOUka2RQBa2qAb7BgCJkMc19iMI+G+
160PqJ+mwc41bL6PLw8iRU3rB5QXjzWFElEOwvk1fVW16cjG/L4qS2fjwy0prrg4
EIMl82qpUKEB2wmHK6HU1oQmlq5HMN/ThTdMATiCe3ZMV34LxLvDdzbf9cFxrJ+d
pxr043nU/RKQkdDQ7y2gt7i7hmSsfRRw2maI0KmQktKqwvMH1ZQyJI5TAYR+8IOY
vRk7s1PiSJD8hrDhuB6p7NIOdbJyyNQd1dfiCxMFj1l0Wpf/zxuXDtlY0COIwLZN
qoHpXIc7mvosuBEgXGInmUwHqZpsy8tPsmTEmc45rtxK2jkr8HqTivuFcCVhiPTe
01AzDb/9wCQhVIt84q9qXL1kT2C70KXJdZu6oBwScOrJzSvVv3QYa8YVCWt6o6GD
8dwuZN1FbjxdcHEhSIvhUn3lhdaIkCPDX/n6OaEiFHuzVLSfpypwPTochSZcPc/Q
t5Z6POzdXaA663NQp/T+Yd5yJMyJt30EfdIainL+NSLnZfen9+bf0YkvCTONy2Et
rggYk/EfPQiw0KHlutn9hHvI1LxWYZHoKx7uVvOKBePqNYOBUw/PiKp+tz5dJCuP
lFRRfCJZaJxLDevuK9o/3kKRchiHf8wO43UB3x/mDAdcI+Ql3/WycJLHfYpHB1Fd
/YiPX8vtovtLOR5WU9+nGf8M/SMIlL/woC2t45NeKf17tVDRE3nL9ynJIKSEeHdi
4qCKg5qiFgrHuH203n7OvlFkPj7tAzAof7wUsa+4LvO6AF3cZe1+UGCYIEwnTMhf
zjZFiLEVFPkAAbMDF0TzKPOlfq+UCX+yIG2f2ILwjP/H+oNcwRddlBAojLeJCRED
81m1sXxUcdTxGd/KECAZI8DHrb+CnUFlfV7tUZAkyCiJG9Dw9kYK8B9vS05wK8AW
uLlpWzx1LLtcULYfYR6nJMAkPQfsnS2UAj1cfZCXHH+8xzU3yW17Ccb5CFO2CAn0
7TGNrFQDdoMfn/vKWqwxtnnnoWl/w0vALvJWM5adt+zdaRl7kfu/iApMA94Me1L7
LZpKkJTab0iL9H449fKJT9BkseRjAzW5KW5H59qQ4UI/Q31iltntaC6pHchtM6Dw
qgaPWpWSSdDW2TQU4pskJKnzKIfe3t50Q7mnnx1MFKhPivFpiZ2VTI5QHlWw7Ngu
nEDipWiN0jRcqIWUcs0M+085RNXK6vR0uO9+dCxW715/+2vlqV4lJyorCZezaGkX
AOM3cc8MC1L1AHyrZCuiVF+Q3e3v9wUAY696mUTDfbGYM8YJ4ESd2HJbHM1bbYMJ
fLBTWWPuPkJtp1X4FFlyPVjYTwhXPkuOl06CNf4ZPNHiwD9Ypyk+t43gRdWWQwoF
jUqYx254PIJVOU1N6ag+dR57p4jlRXp/g1Vbd/MXL7e1Y+A74/IZB20E1SjdTlXE
5nwf7rZtXLzrkg8crKQtFnyr7YdQxSdl11awGtXlAXZhg5Q1XJBSJQzWts92T9+G
vHFYzxmEkMS3DvNCrRthU/P5piHGKj8d3k4iVqnOzXt59Iad3/7d1VjuFbgmmISq
Va3i/tgnJ5qzb68K1n3IhN2OcIn3PsqFVxFmU5A7vjSK87GHlsBNBIvt7vpv7wgC
p4GKKwXyEJE1/GdN0B1se9IK10CRsXmwsVTCrbGaifQJ/Cw3U1iE6Gd4bAEF14NE
o83Ws+czswdeyPgVs5XIQIGJWX2jp+4MtmgOC4WFFPq6mNP4vkkt5gDCYO339nUT
PEL1eMEjnj5RccJtbgyem7QulvJsRitRNebUuZPWMppM67ft3symrFxzRT/kyb89
EPkJBzi0taQTlGPUrdt/pyD3okOGfiGkcZRuvIMCYP2MvBS9HqNXcGNzUuWOptW+
yQQORateTBBPbp6x8iPwKjbE3J2dRQilcy1laggTTS4CRpcySvEji7rScRwnlHLo
nt+QvI6w4BwaVF6M6FZbRptvTeTiHob1Y1Gi3JPX7OLXhq6SdEoY7O0d8nMd5sRI
Yon/dZ0ZSiSUxw/5w4xMNzxje6txKKTGSZhFfoNxQ9upatZyZALzeCfQo03SUBq+
ufA1UXDz/ErRfypQgFHjNS1co7ngHwRk4cM6A3mjxokqVXUefzHAgZLn+7a35MNd
ekROh1h0fKRzUJ0PJN7ljbjNjQaDBt+vv5dqU34RT78j5Y/SGHVz4ePnvYqYyBjz
lQxj6jAmkEDI7iHxm6KXMDdVXNlVjgJMdhPMoJfDcXGYrLOKOV0hbW8gxfvZxZ4t
mWaxZJAR2hsmHN7a7ndqoSXsROGzA9d/km+shDHQjsUGs0aj4TIfHGdxnkUej6hH
RZT/AB93MzVhxK6v0cSK9IKTWKiTdkeCDOBGa4MSyMcI19R7uVJWO0RGM/c5NjLB
EVBc2gdxTwkWa4oO59Kl4sqDFXExgRZjsWjUvhmEWjBeqzG65DC/sRh1gB02Bvlu
/f8mr6xUhW/NKzvk32+AYwke9J3S+uVyudT2l/47Whrdq5hjanSM8OtFO6/gco79
/RXrmKv6koFq1LScKtC8m/l6biFp0jbYPsMdqb5LczrOSi+LKwben/4IaRQQGRF4
u2c8SaCZ0j8dwiPREDh7NZboa9S0gA8hnTA+YM7FMF+PUiUwqVgpdT1OeRbWsHF3
OaVTJPbzUyBtumAT+bVFPJnS4XjGf/vvfBZ5oocfNtvsu83D4xtH0aD5BtQmIcpm
HaT5sdF4JmXs8JA7RUSeqMC5qXg2ehJPs30Ri6e6B9NFxAIapphCCM1yAYg48NIX
xnwzqyL3mMz2Nm/mjS3vFEER2Vh55WJKXPabsC7KoWpCTipdBaL+vp8iEy2LUvwU
O0g511I4sIbDUZkVb/7Pi4FpvoeR9Ai0WY9FX3ug8mi9MDw93Jzf94atRGNRe+CA
23xcNghwFOOjlgHsPxJ2YuOnS58+wwqFs1n8/8MWjTb5ZXmrz+kDWT9qFel9fFJE
0fJIsWtpo7AmD/XTXaxilpDloKpp6W7IU7MA9ZneuoRUahGG8kQbSjn6HeOAclKX
V2bitxzFW+89WZV0nf4jSJdA7pwQMLu1u3butaP9mcJap9ArPhE5ZJBsEFPjy4kn
LW9Ehg+6PLltSfrsk8aLdzy8BN7xvsPw2TvJDEHd+DtNLxeE3/c1opttEoD0R8h7
s7iNp9haQhNIHB6hiDi2TZFMWnf/kcX2i4G8qw8P66f6ZmdtHcYgMTNEkHMsr2oM
XGJEgZ8i5mn95KMUdwnh0b00kjYzDCsgA1n7KZ2FI1BIH9dmGVEGJd2FWGVksGW8
GlQBIGfXMwKg4pl1FqhQ54kI2rLykGz3Vd3HTGYZEm1e4RZ91PUYsjkJMIhTlKJ9
fZl43n6EysprMmfPxiUSxd69y+wCwHN1OZjg3PbFcSaB8sHBnxq0gbrJeGupAOkg
GXADZYVdHOZoT5n3hYIcVewHCIZ1G3jbH9uhy3nRu5AX5YB2FWgqB+jFrfNyWvxP
r/GEGdfAWCwOORhVf993mPgn5W7kmHykfIfNLpZd8UpJm+kDoq5/JHJCVnsfeTNB
2kbwbLirRIBxx/+9hTvQa2G26ecnCdbNuGcACmU0RxqckCzZwpSfX9RbG65nUY2d
J2hte1p2v+LIAMMWw1huWd9kUTNyWR9l0fWG7MRbLZegWYi0DVG7VSHdmioPuSja
GKrgBwDDyqYPENpYWqF3dDd0HGQLGUDEvSydeDKkFUcxWtt/FFNXqC2qVoTO+xle
Nhbik8AyRKdPzk6q7iA8oDX/q/llrgio6sdcDWPE/nKW+0dtXM+LGeKnaNYIepB+
C/aawQEXLXF1rl8KA06rCT2gsMRvK6j7UTEZJQAlA9q56XJJ9oxdrEU3d8GVdUzq
hHxumpbv86YpW07BknHmigSGjpdxlW+JX/gnAiz7hpcwYfwAKd8/XW6RDTGd5F+/
cUgmeQncRX1MgKxUv6J7JOe4g5GM9Q6eSGGJuHnvnpA5Ec4UhOZ9Oab++eVeYhCe
utGXm21WhupXWuVeVvkzxWtf0HxnsFvYn+ISBszK9Ft/ebcUNrtY3R1dA7mnT2wl
Um4mtAoNmqFheL7kBK3RnqjXLGrB0BY3niJaHPfpaiYMwkLECdPh4FPs3alL/+xD
bRbf7Xqef9hNLaIf4y3aLcNLVPIHiM9sjb8gQjeqMma9O8FWJm0zle5CRaHdxwi/
d/NWnkrx/UCF7jvzmTVFa/BzJj1CK+BCNKe5fvPpbNcLhVcAe6yKpFDJXHYjKDd4
53TXaEK/csJTtPbm5OQodWvDyXW+xCCvanjZfxtsZ3ctv53Zm7y940qFyYJQjm2P
/M1GDPvgai86KSeX25rZKB+A9y+eHbEKIXkVqFJZqR1knInexI/gd74+aZI7RLKU
xCxJcF4FPof7hTFcYjrFDE3zsj7FXwOI04p5kL7bGHDxor8D8c8lAZJ51wtooV/X
ut51K1Lzd3UR5Y3Rk9x66WwZXTxy+ZUlUC4dHTcdtIoE9Mv3Kx24hvZmqqlsHw/z
qw2lsFlGkvG2VhyOs9KB+qW3LFbS+vF1G0FPiiQdMtfWehqmiLozy9q7Z6Hu9o6H
r0XU1b227kA2lbD2jQRsXTtWA/uFKlYgtuOFYwIkka5dbGd12rluQrYapp98KNRn
+E/IQsV5mlNFy/nin/5zWvJreXSWz9ixIUpcI5sss75u4EKJdBWXzCtSka2z9mad
CaVCnp3Ykwxb4ozXO7CJ4EG4ViLiOh2OamcbwmlBIDKpupKA2MmVDL7j29wBJTI+
BmsAwSuao8yWk7S6FRb/KB+LoaW9AVRh4HoNYuWQoGM7MLYcU1IooUu9V5xD1hX6
cA5F3NVa0Zl8iCg5tXfznZgi6jv2urU+0XY2TrFxnmHVTfPF7p3VVurQqEsgUMMD
OTcWFu3DaRAKH9cs0XQJTGmAnQVdeNiFnbx5agx8r/ZRJuJri7QNtHfFv2JZEb3P
v40VhhYNfusYRRrwhtTwUgKsP0WuDv1VhBSZr7xk2WjzH54+fMpU5JjfB6FS+Q5N
OJzo33k5Lls923GnrDxNNNhZ1OtdgBt0ounYkNB3R9xU6xf1uZf0x84lxjXZ4QyY
GifAMu//HLcJ8ir25xI64Xm/mmRSqAmN/YhjWgD5URFdwDJmGpaWNxJTdNE4mcNn
H+sulEhyI/Xq1JvIvWsJUaCXkJ73c5/N4BSy/BSNPlIZkWF0JIoltlRSHYvQsN5v
RfNMwTGG1eWCZehyRWvxqo/xBKAGOxW1LvxfTZrJWTRsB5NumLLO4QibAKorj86Z
CZlIjBaUcczow7ahAMO6NHoA1Z13f1LA2S0dLzKd0MAC3D/8MJsqY/AavXtcurI1
o5Qx4YIINVGcFamdYbh/5bpYqpaheBFupv/bB3DxFHaMjiZ8yK4MS4dls6LxSATD
jx9L5j4cxzZGPG73iO3CiqsS71cgbCWjfiFe/rXDzK/7Nj+hmvBZMe1eB9HAeByJ
qsNGUPHcS+rM32gxvo5ILE3jFJeiFraDvK7XxDMoujKbfCmA9W7Mq0OLImSQO9gU
Lu2n15k1Xb1ozJA0A/mkn/rPRg4P+gbCfAH4Aw5kGkK2lb7cnFkBdqbv2UfsX7dR
0Lqjt6tWtuypMEZz6Ai7LpvlLu9bUSFtZy+9fvKZT2ddjZ7WTIzK+5A2UsyyKZoB
EpLz92IpqtvS/mCMBPuJc11imEW26Ow9861SYbVWt3IYf4nKvgeNsGUeeNWNAo+0
rxoawHBREIpF0fChKNeb2zZmcSP7OC25annGRAuo/t5fq467LsOp27kSIY5xKxnU
TekK+AmzzevbSDEV5t+O4+vFTDPY99JD/KY6HbWZasEia42mv38MNQgo4N4sdOFJ
llz7obePXVRkqF4guJ1BN9sGgmgYVdFqlRjotnBTuzkz1B/j4f87DIPIm4xR7XaY
`pragma protect end_protected
