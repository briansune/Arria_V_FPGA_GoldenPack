// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
J6bsEr3W+rbxHTeubapcNLx6/6MbZ5hdozmWJPvuVZE5BOs9XPdIjKYuUH6IjaXTfW2KjEfJ78A3
aK3FNHMqq04vW71hTi/I5KtJlBbq/RD/vc3Ol1k4kSUq5oa+MuVP3txwJu8uQHfxZELGBp3zUuMx
1o50Y0L5gsLz9HWWyEKHlKDldfTXeJsOW1DQMiStzigfLBFERYRdEeGgV2Lxj3ZrSF9TOqWEOc1P
P4rOOq6Q3CxQug0CHn0BBRwMD6QzwLq1Z5CnvPOWpNo0xszeLN0FuGreDsBcwQuPvNYBCg3+zZp+
pGcPMer0cFbO4Q3bf1sOl2BkgGbc0Fzpu274iQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8880)
WFCg1ZN4+tL4P149r4AFTWe4HsEQyoJzv6p0xN699roE302SSLUio8heLsVVfJhvmMQtUPPJXFfp
0vqxbPU+YRrxldu+UF6yEhoOWUoGTve/2jlCUzrW22XMEHADDJXxUsJ7cNW47Jx0IPkgZPCh3/Zb
bAzaRIV+UnPEnlibmwt/moNyJqZK4x3hheJdmtomRWDFaGzEz7FETV7LL91qJeD4SPdiZh2f3BF/
sO8e2uV34zktS4MiUv6BW8sGlnVaKAE4QEhLj1mNsvaAXdKny126UlHkcoICmCk5s+2dbPMgabNS
NW2DGHKW7HQ1tewTKxw9p4POhXATFQF3ul+kj2C65jJyhD/Mcl2Nyw11opNKUHnQeBJyjUeUw1jx
r7RGvGuH5Nh2wzjulDAPA5OFGMWOoTSucdeNTRClBf/OicWKi+DVulOQ3QRPna9Tu6AAb7AwjfR6
HhGXUNejZ0vH5VReawcnKyvs1kUpGlzb+S/A16VASZ+c9rNFEjPtde2iOmI9lHAT4m4HvCKFFYB3
v0wK6RlAobClHD3OjhnMyriHaf2ljPjqFoe22+4vDHN0KU+FGVSNp5jJa98Sduqf2n1ZRtLajfXQ
MV90vXgZyqvaI/tv/DL76HVB1ffyOq+OlauNWijfM9zzTOAoXQ//y9gjyhJYrhmGYwe08W62XShw
TIyrNMAiS8Z/eQQ/2BTNEKO6/sW0hN1rmldhjAl4DqLgWftSom07v2njNrCytUcJf2/q/KdwEFZc
V3X0myIEWn7DpROvaw/hsupuHC8Z6GLMdKyISiI8XGGs2phFdeO+vpgBqyEDT91LEpZdY2VSwWUY
P+lU9D3+WINIbiLG+5/+LUeuF2SsYVE5EjCutZifQ1R6PiH3KbxADovE745D8j8NKKqjJ2PxMtyi
ces8d8N7ZwaMdqdYvQ74HBtzSe/QSanpXXAa0R3Wfp3lWlE1TiK8sX6GG0MHR8pSdX3cPRkEN6EL
JTQUTlvuxEe7igkweigZdnDNz7V7IoxNqNd7UM41NnScM1h9ISes+8KaLu5/zWgotduRGtPrUJzK
vr6vVUDRgqU9UfYRrLpFc1/inggMbbFPJFtIYW0vz8bsdcbBExYJMKeERxTqlP54C8o6qGvUJ6AW
nN9a2wBrRT/ZY8vQ7zB+h7SUwl7sCXDSWCnkdM7DJHIJbTqpPyunP45G3KyUIM2rCoFhmMVQ+lX0
1s+z6NLnrQFceLkIxr4vpr6HLsIiuZhCYwp07oLevZP+ZqhsBn9ta8Z2/w55CHy6wrUOG2V7J1X8
u6snKPNCb+c9cBNu1CwFx7Ct9HbBycyyqNNU8wsbjNohC+4akh0Ctmfk/MZukU9rVLL87eDAZm0D
tWNRo9vSrKCaxdJZ+IJzOABYKQUT5+VCcJNjsQBNAA3MtV8H/+0Lo+8FqIllb86HYJPMqcprGlgo
EMv/t0QQLchTK81JK5b67y7Gj9W3dPlQ2A/al2hw9K4e7Kl8/Bhf8pcA7FyDvu3QiuuMOq8Yb6ro
BfOFtEp880M3+kBE+gWkeYI+H3XPGj/IEwPyN8EIBYNngLTi7gOD3Ue1W34FNaVaUxN0DFGSzirR
A0TnchvNAMIdgjITPXs1gvcCQ57mbg38+XMaEVk7AlVqv8nEQrwPWzdokFjvWNHIMA1QUd+BqDZy
4KuRwETCBQcC/MRxYYbSQM+UDBLIyCHz4USuQ9IpBGEMClxpMaLDVgX2vZ5da7ICptGyPFA4YtIa
2KDetpzK7Su9VS86eC/J2FFrx4naHtVu5AVgIVSo4bGJ7ydXeUPR/x9WvSXdmMxCRjnMn/vGdA4J
GXqprwBMbJP/Hja4U8avQRzYdcU3tlru3BGBN9x4piVPvxCEjTaGfG+1kiDorRjVn72Phd6oXANy
QLLaFzm9xueeS8zSPZVIyaLjnVUmjjOdklw4Ezmq35i5vEkrMTIwx5EYZAQ5dp9QfLy2h15WAi6v
/JzxAH9wEAw0deyy/uVy+mxtpM3h1cKVKAmaGv2NO8VdmrSaGTEt8y00fF0J5gkWN2mZaOQ3ACl/
IRkwRPk4TT9DPc9XgLsKPt7KJ1AaIECrfRlw77nGsdV3J6YUPKpxARnHj+2hHWlQeBBXP7ByzNl9
An1QRpgFa9Osp7pOKlay5PGEplWp+d2y5RDhumK35DKXpFfO7CXhNhNGv4eIFpAghXZotebc4ly5
SP4i1nc7PaugO7yGX7vfyHoUEO7vZzf8ie2p/U0XF032zAdPLgjGFSIPLKm/7gfMGBFY7Nijv9H2
40VwIi2ZpHjP1r+0R6CloILWV4cdYPpe3BNtQzf/oioiHnU4myu+cReuYEj4PAbsEcEh1utkIXw+
SVE8I/wUm3W5zQ03fE8Y7OtJ+jtzJRRwJBsVl0vrDgkYXFQEFxGXVLBbc0AcU/JHRcXEExMQe/Bl
ATDBHnREPFiOXqwFIVEYQFABQoffkqDUsZDrmb9m6RlPjL4gPL3sCtVtIHm6wxHFXs9iMOEb30oy
No9XdsGZS2hPxreQbnqy1/+chTpASvASotF4vBEauw2sRBa+eTskQuuJVpvVfyyOaf9OOuPwm4Mi
+gUBX913C2z9pU2db+WI+GUAiQph3FuA3d0hOsWX3ifYdl02vDuoVlqPjp09T1/Oy0BtU0bl5zE7
scyaWx/zGOdozfl1uWd2bjpr/aXtLnZWU2hqZpBMG3lL+BF/ALNSOHEvVG+GJgaDD6noXdI/j1es
H/unuZf7Vinc24Bxyo32equPJ1tvGYL6REINOtI4KILuauNRHQQkrvEcHQQG2GxDu7RgHvp7O6X8
gxCZRoa5ZnGPyaOU5mHwKfV0zrktQ+WA1gox1mWYZ25FGdIsinUK92V0oFvJp7AZxURLgx4aXAHz
l9SG4qQCkplUHO0w3qommeg6aghwo/Wqz/xf3xuCGfdm3FwQb4PglHMN/zeW9smQDRFEc0qcisFh
RGd2ZABz4NMXcKtLfKFTlNtFr1Y19dPdsiEvnFE3IDcugrjhkfoqVHfQIHHh2ttUtRtGBoIkOa40
AtKOFZdkH2KuwnhEoHISpdRHOxVrd2YPgBol6p7Kqx1u0qdOMX/otb31FzEeOQiqS2VPk0lh2Y3j
znbpbc/UqAvtg7TBSAkW7kKQWBdeK7gowjsqte13tjebW849hJ/152wlgvkJdZs7HUluvs1P3KbS
wDH9e8uP5ySdY7sXvGukY+KdOXnuw64YgHJn051sNa1mLdsRtPMWNf1oPhqUoCPSVVh3S9jpVat9
cDFKs40y9iCPCOls+LFlHAHiV93e3vwKiw41JgGkXeXacgsVTAva1n0FpcMvhxE3GUja/V4AnKQb
BAIIGr94/7CsW7N3udupWQAj/7uyEgpZSBqo5YIqhgw2Azi5BP33GOd2xyoJfmYxt6v7sw0xZXNo
801BQ7uYcLYkZadX6Qxkzsym/zl/00a58cB58wul8A4g6ilPlzqzAukEmiWO2nw1miN0WCutX5LY
7HefCBoym8S3ATVrVMpqw5itOtWJrvBmifQYjvrPgUlaXfcZIveWKtD4meAdjwkTGSl/ZGjzU1+5
Lz1dFTk3IWiKJtj0Uuf3xqQJE5TFCKL74QiKgC78cRy5EY18Jc7riHj7TOScy2+oyxSrG0wYusEm
lii96NJJjHdzUUBCz5F+OQvgObOh2zLMp1PSp3i6c44Jr4sbTe9JeuEVluBJ6JuHgNsjsUwwjKDn
1zIez6OkPk4OY/vphgDl2rrl94sL5FL3iaJjzSGKO1eUBedUth+6VHvjZZ3+dXAu+koYvpYxMfMY
EGQbgJO0nXQl8cX85gnj8UD7vszjoMd07SKxcG8xDoSFEqrI88aiM8H/2K4dB0BaZlX2D4asBTt6
Bnfv95bvMfAxM0lKwhgzc5ykZuAstddW2l6LEEhi6tZeOFeJP1xOnc+12am+1IJfshL178O5CCAR
ekFcuKS9Ef+QDXZ2i4FNNO5WWgxLE7mUgh37A3lzYoZq9a6j6QgxBq7FKXUh+s8gYWn0eI5TwV9t
WVZ5STo0a6/F0t7+kJkQeuZmOVXPAb6CSafaOc/xpIClDOKEqQ00PzVdLZIXRsYYcQNZZPSTgVOb
FOrsk7QtJsd5vRZLBChmQ9U4oqgFEkBdFZG6auDZHdeeCgppMf6P6swB1JKGWa1XnnMJ+y37ebmL
AB7iYRQoyCSbZ/YEliB0h5BquWu2cl0IW6onjvKaHgiyCKEWk4NJQmF2XNqRlvfliq2NADIgA6ZQ
9BaoR4Ozi0jsyDL8t44i925ei1dmm4Tid7U6TX+tQRkwYjBJqr0fcxDsNaAP6z2ibobuj+aG1SnJ
tlPxpMslQscRqRfcjr7rTo3j6ucNL6jxY37qh/NauGh14NwqiupRRrzoxx0w78+5JQ4iiUcHV6JV
cvio/4lfWaeCICZ5KgXzuenePUQbHS0lQosKKPCkpRhStXyVaNX0SJGuqi9ksmKF9sb63fCC73lA
eKvgPeDdCMAcvg/ROrScXXxeTyJ0ymVCzTDHG0dhann8+BEF6iF1pOqFQyUdDYmgfQ4UN/Bi92Ao
oHDoB+PeFrywQW23hJN1bEIHw+boSTd3lEj6bsT3MA5a21Csqg2psABicCxWE/oFbAFG8hmvnGnD
+VFa6zVDAZDaQ2lhdNv3UGC41Z3QkEUqeVHbzw2d019cEtcXlaPM1W5MEkrBmI/gJhwi/yJIoiND
oyMH82WDy0ZmEawIoE7YwET5R+mELPE0fcTo6yTD9uvy50O6HUGjykZCOlbeGwpqQEfrQyqmWwWZ
y5m6MMPZGnv0QTiljRVSNiQ9qgaozh13r9FWwjZwpTcz4HmwD3gMDyty8DC0xQ6N86Om20OLA06N
E0YzXG+7p0Afw3t83yiFVJeGwVdGcN44OXFH8JGa/WPmW7IrTWIea4RnVf0K2UKi/pI+zTL1ByM3
577Fw4JPv39ddpe5vuEdyEcR3h7P98BvB7ymMVJTosCXPKxEgFVgh3j2lFNAOfeu5FbyvyeS0g2v
g9c6tMXTH1RQ5AZN4hzIkP3lQEA1fhBLKGhX3LODp69rloH5ClGqpr6vhysMlkZAB0Rgsi5tlZMx
PL6jKdpDwCRAJWN/TetHTu9qsKtlNI8vdqPax++cSusvTLB8QeVLxM373fJ6V5S3ZBYoy7CerPJL
JyUvgYnNRz9HrslTt93ywajNvZdaC3zQ4yIH6C6vQNaX+kMgXGzL3vcOImoBgvYXr9dHAxlaX7iF
DYsAPGpHIVhlFnH7F/nlC5WhcJdoweLhafXEQ94qlWcBeTkMBQcPMl58iRsVDpQTfyafd1HBbte8
hnkrNEb1OZ3QCIUBVd9f6/v3yvsH4nobIm27/7WAH3HJ6bmHnDNJ+tYtLnFhuaTIrBexDIHVgaeJ
JBXxDiCEHPCHdfq4Sc/EVcvEvum7KuHVxFXwFjSqM35dHkeySWNH5JhvUxhOxBnCjq9eadSqC0Wj
TSXWpog0lm5w4R15JJJNXzXlW6XeM6XUf+RgJigf/+zb/ZyiyT4JYB/bNJoHnBgxp7WX0MCeB5JU
wjCjA2f+s/Gx+DYfd+62Tj/OE6nGhl8ZcihrQg/907ZWv/zKsWeKCAHWsQ78fVtPGWpiIXACKqev
VxtSLUWeQJ2iW/QdWvFuDdRSCh6HqxT/WyPNa5cEyaEJ5k7D5xy3eMFECl1tLZUSCzimy0Q2RBiK
pTPZpoAvq2PEeVxF0w97VkQk+MbLsZVKCPI5ktJ0vxKCLUL4b/gkSU18YdKk1AlOE1q5LDKX+7sQ
+BZAEzhTm/J8BPrx1j0WzLE5YHBZ2ZEehg1MpMnL/pIDea/wYHsA+aXOAdkDhkwkJSxGEd0yxweK
zW+9DSMVfjhd9ccP/vd1+uEnLwhZyd+Jm9uhwd6imunHnz1XRlhJg9TVQgyDkSUc60DO5t8FHdvt
crhUnJ7eYy+46IefQDiw4xrRnX39WWx1vwz1HzOwuiU4AAoUEAEKjavwoWWh9pnBVGRTO8QBNuHX
ZquIU1gQR4Si1R8fB/0M3dJLGWFRCM+WNLYaC+Vrp8i+4rvTSL61U+TdggWxzhAO4dp9OXJ2mpmt
5WeUWZRccTeF3gL7bSFR7fECjDRnE8pYi1nRHnM5FmskumLhfvs+Ezx+jy+PafiDOwoXeym5JKHz
O+AUZq/erVlSNegPdSt1RzDNkVNgbGWCge4XEM1432Y80GSpBnlVVyYZChqbPqxJi02VyorsScKt
4f0Q5Nl1OBj6xd5RJk0MrtghMs2hT8tAS8I5qTz5ooxLTIVF2arZVejkcYdP3jKVv2qrlPLyQGkR
tYEnliHDdEavJsF1wr/SIQnLhgoyZDL5L4rKKSrSq+Cs7aRMUWWwi/YYqUL+l5Jt6SPLHtmT0j7F
S4zHvOZUPMK6wPDWgKxcdRJeDhSeE94O80CRHqYdb6wdwzoYoJmyr7R+3MJFXVgzQ5fWDRNo1uds
RivTJFAtC1qoSaREq8lo4LEKVsOt2Wc1qMvAN93AYS441XwDsbqJJDyyIhHVYfjMNhySz+SKStEw
tlRsQpHBFBXl3CXqxOY4vcxgTy1nZwIx9fT0IVXpwErLnyP1UtjTUjL+iZU+FEhj10yl49MA5S8P
V5zIu0v6aFxiAHH3U9Vqfifn84lYh8bL9d2jqIC9tlRK6qXXXy5eyyODlyYhXoB6kzFAoCTNQuv0
vjMXh4KFIjlQkbXik2qnJZJ8qmVMhAO1XqITbdfmLZeuae1h2/B2Gn6JOlSFUed+UPbKqbdo0Kun
znxXKBcCnt0GoyeICjKBfV6aUTx1Zj1hCsk9QF+IUloif4bjhLa76WOTCT1Jltd5WhBy8uAIkCS2
mavWQgWr8HCqENdTDaBqSjuNhDcpB0Zoz7fU1kFdssSaVeppikh2TDrgBM5f9Jm8IhyXtBqmblgz
2G/OH6saqjR6m4fhJSCGa4lIjMnZ6PItGfZlgWAzuveZJ5hX9mXTtDhp9O0lTT9pPjrT83Jbrg48
ha10iSzjv0X00cXRTLoWQWBTxf53CM62YNfAds5VehJLm4xHXVzTjTmFiqVRHQtVKKhgMwxd+OdX
5OYNmI+4uCna1wNVNGXFbhlO2tZLHPgGtiaE64y+wx9NPBk/qEgsWX4BWUt7GsUal/vswiaey6eO
tJ5yhn321mSxPbOECUrgn9m3W/w+KKO1IHEFRjlnQgPwZy2G5T3/WqTwKyP6ZW5S+PVbVona2snX
7ZsXck1QUXtDXWeXMYr2STt1rkx6RRlfKqC0dNm3hJrfAbsyqZ2ZtFrtLia6dotC698zWFJHI1zC
ihmVgrLKLNbsxqVaXu/0W7Ep09M+2/BqMyJn96DK0ux/JG/CIwLQp7txjAuP1glBgBkY+PTkphIN
dKXYDstlQTPKpMP/esM2UAea6NXCfzKEzPu/pj9DQQcayljCGn9k1DyDGwCDzSKXxUSTvkYtesEX
gDwmGzR02KT+dr6z/DkA9Bfyjykt0rjfVPlw0FIFMd1tHbs1p9Z1UkyWmTinRuePsjt75fGZoU5x
b7L83pEe+mgco+TA9MqdXTpsg2skGxjAj51WKy78bS1GgSUSvGmXvTq4UoBhjsAzTwo9ihubaM9H
XU1Sw8HuL1G4LcV/5sWheu9ve2EFIol9MS1zUD1yqmkiFM9XyJGPccvK7+yy/XuKYDjmBReuxhA5
oLnwLK/IA+9ZVbvx8DBeybeVW9Whm2H118gV3hIDbXf3Piq7Em59xRlvTX0mUwrIHgCzZNdXwj3R
rzZTtcaSAvYsGBwr7F/JBPwcWIWejLIZ9JVAYgloLQqNPgFNcZSrg/3RFHh7B973qGbvG4jvMUOw
sOgnRmtJRenHvPFAc1bej/248WIA3vvrmEMsk8cfQ322IiZZAJuhC7ygJ22NKtIrBV/BsyHoT2mn
L7gIzDFwp3Afw7asBh67IIa7mNMXpQmgOAjsTedck6xNzeV2n/xJa6m9wTqNovlyt/Y3jffjpOLy
cSRIMKiQGcZSIL4bg0xYq5ljkuAlgRSMvCVcnTFeU50DDFpZzsDZ2AuJRNr6WzjiGqgNDAUrY5Wg
KZZ6LZRWHpdP8mMzTDfpKjPfAxx25rCVroEQDoUB1wf+UmPI/nZ2ffwKwQID1V5YCogoyYt8q1h+
YQAjs5MUyhJRwjMjP+dKKV9t5pA1UEqhi1dIA0k6LLvqwW89VUqc/NKInWCLGvn9P3sNyHKo4gbf
sPWls1lp7/iSKU4q4j4QkvWrsNCs3jY5tu+gbE1Yc9z9lDocbVzpvLMFtwJhjkKq1rZwYmry0lVE
p0USMssMFuExSaOX1EC3ttYqLlTRSRoVb5pPo6uhzQHNf++vIhCfdZR3Ta/xD/eqr+ETBUS7FIuk
trNR+vjvkN3UlCQRHIqGBeZljmR2BPLfrjrGJ/g8EfSKXnpYwQk9CXlPoJJ8QwYzJDx7IK5lvjcX
w2EUPG56RpbukSrCuFV0Kq0c4EQDNM6tKTYJWZEw4IAjvJNZUyJt1arKp0DbRSE8b01Bhgpg7gtM
IbJ4+Xb3F6NvBxKGkjOLf6e3+Fx7SumUqr+Sj6Rw6Pqk4aCx7q6ZITYbrdY5kgWUsllo/GaRRind
q3m4sffRlEmis/HW898ULo+UcOh40sbozjicCXRm0dD44JzEkx3I8z7lUgxzZjT8R4D7rHOlN5dr
5FAOP/RujdlA6tbPlL5fo5fO+t86XMmL0wrC7MYcCTBomwevjcOPJCzAP3uNRKepuUa8fyhLWNE8
2HOKRgGQJabJw7sRevqptCr7ogYuvT01De4Wg+OSqvCTcdXGV81HWixRd4yeKEj8cFkk9viW9MQH
mG5NRMUcwDaladManNdWO0qwB0XydvWwXexmALLp8UefTaVMcpK3fG6OzdNNpe5Zb+Ik8px4YhHp
PWP+t+KM9/D3XfhieZ+vVNOZMfzBc9OIqr81rRah1U2nFVCpzzHK8g8tK5yH97Kt68DLXAX66rxw
CQE0VowcKkI1R8XsgYRSB6W3tHTitZ9ao3PbVrdfIw0bXThM8N829vx2AFd9AwncVcM44JZPOHEV
DePpoQy1XO2iGCRPgr7UYSmGlK0LaAVAi1V5mcw13v2XMcRFbZ9pGnalyNHj82iAEeEJqLCdRGJF
GBdKMZf9hxm/7ImqKB0DVBmvNHHP2qsBmh6jlQIIFaX0G6t51dT5dQBRfIg2obbHPntPOG+Sjyab
clyAVMAtyK3fdWNwGBZt7RepA817OElVb76Fm5fXkZTrgSRTHrFqksQuVxdRaolchW+EMQ4GSOlu
5bV0WJpEtw8vS7nSuDUubcDbvI9a7ERowjk7OHC4WbxC3gFmKFMpZ3Fubw+33/1NnOdjmD3+7gX7
grjjPPh2a04XXje8GLfBzw7tpXoUYH49T5hTOIQpGcGW/oXF4IXBbEHTe1hkeJID0GsOe0nvWV9o
RjP2SssoIbhjYrpD5kNOoJn9T70hHnKdPW0x8Sg+drORBDzQDVcPHamN82qA0dG5Sfsyv0fSyhzx
rywodjvZvm7NlpbJXgWwbebJAa5axwWDALbblsqJ8Ei9AuLLMZTQxRadaujbWgz0dJ3fdvkEXIhc
fBxV1e/bNJ8w8361TWh7Q3x+lOJuN5meP0Sq68XUEcGRh/6859199RZSYwDHb1lNxGY2qxCz6y30
03IrVAyYki6DLadMyXhdW7NYFEuow2YE15jV/g8qyTxtcanI52sW6m2zvU4TWnnELfhufjm7sOno
Ls11SHEgcDTtY5Xgdd0F7W9As0HaJ26gVDBRF1eec7cGYK0HQr5VmrLyH85DChmK2rAP34x7UflE
wTiaBY7xVGHSzRE+iU+UOQFjW+k/CEZzzUhdnNRXmh/l1uU4rA/3yx+mjXkBIbNXkdCtEWY48zq3
tD9vJY27gS9NxApmkRVHLZnyZzms0yQOZWwvF2v0IR6JGATn/hdK1xoJyKo4Qsd3FuCKWUDeeo/C
6H+6rX/zjW6aC5+E/ABmIJQvZ6J+KHf+f2UPZEf+l69JUFc9DgOhbe2ScZawrXaspjIF7YBWhhLV
U3widi5cYV+9ltkfHXgLsQD2wdxn5Xz3IyliPR8/3QHC9OUizamcaYV3wp9KQZ0nkLq/ktbR13Z5
W7DuNkCSYM9Xqzto2tSOJQ65k0i0CjZIc7QK0/jq6eGH00wa6t9ZQ6FDIzDHf+r/WUJyg9edXzsE
Bpr75wmdXUYq0QoE5iRP7qxRHpIHFEyDqoPtQ/847jy5p9qqhUGcOFgZt5/6/9x+lwMpKdawfDOj
1KBFZUNKLD87wRekc5OC3c5I6XR3UBm4ud7PAkZJo1TQdoV98s+K3EqI4NV5/mal1eEjZakJyeE/
j/L3JmzW9T8WMM0p/2LjP/eNTb4iZjbDvjgyFjRQir+3mQHEGHNVrmFA4Lx9Pf6qW8+ULyqYUJ2C
1QWomRnNRGaTvdiuz9GyZAFpZ3ZJK5wBHOm8ghDzMKdkZKZ0hnhp6f2mkVU5y84gbHdwZPQXOQdl
Nl54VVK+vDCNmicM4TS+q67y3TT8e8H3e2S7HskOdJrNPm49xY8zkrQCJKrkk7PyWX8uaB8Ss2Du
BO92lfXCpc5V6V4/FzU6FlrMOCHUrrJ8V2Qlxet79GD4/2oFUkZSfxSd1FgcE0+iqYMylA7DZCjY
6PA2ANYViUCBOMXL83nQqDm1p0A5AMbP34QVwHSxzHduBMPO6I4nw4c/6i/IMEJpns/GaTCJbek0
XPzC475HhDyEHmKkiJk7sVLAR8knP3TTzuPHXf6Hq4SB+CjG2ObsWHC8dPBTx3UUlr/CzJYEXj0Z
vVhsqU+RzKUI9MOK+iAuBWo6YAQWfpY/dK0rEimdlMK2AyHTcEGWnOkbd7+TRQUFVK2WU6aBtOSZ
HrbXJ1d66UjNFbisRl7PGCWFAbVLOWZjLJvl9ZibRbDBkdqxQHzg6HVj5rTOvjEtdVhN+cpw/6MZ
Eq7MjF8QuHibEZc/YNG+RREf6bR5SVKeNCYd87iU4zoW4D2GPHvKt3szlmrGwfO0OAzh0jvTTkrL
aY20QuIXwNvWejWuSH4hacneXSYzeChITUvuZYUcnvLlKATRUBcBtVWGdDp3EBBa0vB1VbpfyfN3
+I2OrVkzFBYvyPctne9v80MXggI+ddf4ve4KVoIhnxgjzODgGAwLx0vae5CqxWSeX0A6Ux9b2XkR
N7TojPaYyCVEmvsjpJEwraZK1HKmtM7D7x7LiQmfbD5sbrwVEkQiPAXCNMxeRlhCcacp9P8UPy62
EzuxNPbDvPQ348qS6lkVPOs61IRG3JJU7BgrAZF9HIs1odcImiE/gLpkTAJLfcQUxJFtl2bDkqNY
vR5jUoCJ+QloWFGBJR2MbcGdvEaULNP1tjkASsXKhGA3bxi/voBl5LU5qJVO/VSDNFKlkk7Tkk0X
64f289w9F48QihlU1PiilgFVP+1ZY+P5mlxfQ50R/5rN9s01otla9OJ0ajvK3Ft8/krrALZ0vWpP
zK4rsaxD3PcFZNun5a3rGUo+h0lqAZdE57n+GmvusSvGqgFsFW/aVM0pXccVM8VcdfboFdw/At27
MD1M3/qFP7Em4w0v7FgLe9b+r4ucV6OFbSnxzKeTb8niQ2bTpd7dFeN+WmRfPyYtK8Wq4y3Qj2ZM
LwtU+DrQ8uI9BXxKBny0Q4f5B17S1xwBAyRkKF7a4XcV11zvfB6utsfzGqydqDgRRPiKRfpBLjx+
Ipg8ZyOx4PQLAs44PDe1I1gYeFPuz3AA1//gpSd93G0p0FldGGPll0ceCfPP4aqUHKYdGWtN4ymr
WVPAN3tdBx3enDXEiah1m+5/YwKRmJZPv+Oan7qNYghmuyjG9J3PRVgCw+kj
`pragma protect end_protected
