// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:27:18 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MH5j97JL9TbUiDEXoEqJRzZDzJ3OicuVVnMLm5tZRaOhoMWY7wh8IQgHHg3UyJl5
O54d0dy2B1FU4BPr+sbrMDAsP/mi/AfipWS9ANClvTNGPYz1livudE3SdFmomMWL
YaMTsk/4CFugWshQc63P/JsVnlCRHbERuxKRMpV1g3k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7744)
E36J0B7JwXxUMVfQBytlK9XR5EI1fR/zHM1f2gQxe/9y0kBiWS53U3HCn9tZKufk
zP1+YzzgC9YuSS7dnwwWY9GngviebO1D0QzdCqRDU+0u6sUiDJMl2f5Aw6FCFT2O
gKCJFcL3CHk2yqXAdqyb3E7e0KCGl9wKN0jYAwooSD89atTXF4taxBMEE1p2Wo18
q4fQ1YQ06NQESSmvYvB4UvGDXI7MCBALjAHRRvoJ0kMnYr7eAMQBENg7WRpqz2eD
GnnbglspsY0rSI2DI22BAqwYaE6lKsutTz2swFHgoEw8mqapAQDnOpR/1VnMRaay
RkFXi8srsd/h9+E19QPOC1MrBDFgi06IVEbA71eSayVTA8p1fJty+6nk6SB4Y40f
xIHHjU1/WmHDslfMTNXYjbHlshpGsMb+MsP3R+dljR/88pR5tYnQIP0TpeUmn/8f
a3n0spcEHlDVOtBOg8Dy1lAx/gPaASlop5EBFjO5LKimFFvesl5KKYqPI0w2RdgQ
HtVih42tttl4irHvIKxz0W5mBVx7EFmYePzS3zvevzRQoZOoJ/irgqCkbyNn6wgI
wKBue4+tjNB94W5pg4SMaoIPGwsvQzdUmtZRm21s4KQsDd7cy6GMFEVBOQ0auF0Y
4blF8Eu/ivdbttDQ80qv+2KruFxUZRtA1U5Lo/NU3O1KaJnKRBDHOsG23zUceJej
5/p0bfjk310G1kzwmMhneSB1MtVfuaAy/geG7YmVAfNkT7oIwW9YLk3E8qjdjdpA
5YzN0kWP3UYNoNndIzjyroePmHDJ1ZV9501Hves6NbiuFlauGuZEZn8attx02aff
AYVEOoMGK5StxJE4bEAHaJGB1mN+PmDwLHiGocBbDWFpGvVJjdMyKmlHC3/YLI8A
J7a8gPIKons45p35tYP3sU8wji1GeYBW99XGb8MK9gqkhsv0tbSLuHwW4QNJbnXG
62KKtgVchSp1+MPf7Eu3socUL5FAbMH/4fSfkGAHtTjXQb2A+r7QoHYdkICrBXq1
0nFlCCDy4c2QYnnF1TPY3snzYiUGioThXjCqFgV/Y/8JPlQHYAKrfpg3iaD9Nsyv
BJ0Z3u/KZ4uCukoXA47OzLhOx6DcMXM767qPYtk8A1GFdmM1wJ5Z831JqQVfMwj2
noGPGE2EnkVMcFPhe4EloU5DZkLSuIwsG7vzqh5A9an+aDrh3pmm6UE5561tEAQ3
Fx0/h1hkTRu2wp0GDHrVwQKulKcnqyFXdunmxqop+ndJBFmI4dw4frBnADdIowGI
nhcFnRNPFNHLf4pwJo8q3DxLDTrA0/Ak/inWfu8Ctyd/geuCwkqn3xw4E8Kenuv6
Jk1zHWE0MJifrOldJH9nnQ7WW9iAAb4q9qlgXFmOeRAvjrrRQNzSV9agtZyAUM9U
xicxRkdNjbJy0BvNd2Z8bfImQgvgh0e9pDCENeN2YkutbAhuyODMjQ4Cz1rTDcXr
f4CTafxUbXUWkDSgH0uSAoWqfIdKZ5U9qNBl3KsVL21ptLhDloidML2+M3o1zeib
dU59nIo3a9ZZk9EyvXy+OhWQGPkT324IyxeHNDNCfjIcRJokxXVvNQs+OBoSXj11
5kZUspLdBtXGm1ZyOZgzlxP5pwhAahdx9reG7KbK62VfDO1lF3ezA98XmEvLzRyO
8ENLVzsljGpkfFD9rvtj030W8T4FnWmggSSFQH1dNDHY17lSCTUNCcH9Inrv1U/I
2PHgpB+FX44/ECDytkRveiPAWHMp3m3EKloNtmS1fXn4ju82W5TMaBYofEZEo199
wco38jmoQFPt6D9siozNzjtDWxTsHmf6VwOM1Dq9dhbirfANLiDHgWnIE7oGaJUl
RQImvtiUa7OV0xsaToldRhfOM/2SqJ4f5MbJfWjbmdUq4f94oanBNXLqdwl/MKxt
Spj+JhypGY+sS25+bBvOlX1KtwWW80sPYqd51hJME3Rltacmqw0xxugzJXcco1nL
kjkoYiFYRpD2n4RJL+58ueGBJc+NnvaGir9L+RJnqHXKErJFGS2/5CIrE+1AUFm0
QOPD//YKKqWioPkAP+IzunU4FKIdbTQV4F5GWoYtB1ywbPwdpvXWryMtz7sPJMte
5ooxaW0wFB05BmEX5+t+5gYsaqihzKEGwv/wX8xQs9rPLzw5BhQyYq15J/4pwNBg
5sJNJEYCh4ri434/5Fyo3MEmcAmgIQwx4oAaW0h1fmr8IVf9m59aJcLuRirJul8t
7Wu/fPff4nJ81XAs+Fz6HQM+wGw40vhvFHtM6A3D76BzGHUAazLBgm3yOBgq4R+1
Ms6UrxeIt+GSJoQNQpNwLOwyuZDvJV94YSrPXmlRak7F9vrOiPdrkJbXITzAGA9j
ouAKKBNCBP5bP6YbGGepEwQUI2eeAB5utVcSJmz3uKcp5mY8J9QJB2vB51ZxZGZ4
/GgX7QCGW/f6Slt+E35kTzLfEKtuyTNLe3qW2/tpHOXyFC+HYPMOPS2LJxER1jeX
Jz0zlFyDyLR1g3raCleGK1KI2JaeEzmbPCCI42doerneVCuteEZrEvgY5xwbGyk/
TeaLNwcxzN+x+Ttu/YMOf73N4LVAsDBVagVjHKO7YwUrz3OwxAYwoBiKhWZycZwK
LZX9g1SP3qrydNAWZvVwOFMjO+6Dgb4ic2CsuNVGP6UgBdeSIsWn5es76Ua1i3vy
hsfxKNovzbB3fzhqj0aO/AhzJydOIJniEdz00tn6OZGhny+Juj8+KD3vkNv8djIM
ET13LIl0xSYY5xbkcBHSdD7CT7Yx5Y3DFlupP9AixyeysHJRNYo6FFPrfVdqnviD
xEAICPZUcmgbx1kqz23+l92YmQN6ppRYCZ9YFNgIL3ZH5Vq9Fnem31oHpPiq+XB/
I23muW7+gcdIpk3iJmhX59i7TJP7vieKeiW3GZthilfErVw1HaZCnussYLUgRS38
AsAxcmJkKnNVi+HUE0nlZiQurURruY/yLw5zYluU+R8+qldVXzfVgegJQQHmKZ48
roDonL5PFpZN1xTdl5y2ZFGo7g5Kmw+Rc326Lcrw8+kPegvPC8c8ggl7ZhetPIkE
ucQboZmQ3iht+edL6NfQEY0lnwdN0nCaUrdI6xaqxqTpQTIUgxizjYYUipPy48Rc
5Tm9tM0vJtwNkQrxvR210VQfTXGS7HNgUf/fWzLAnaCmYY2lfGBW2VVndha9qHL7
uifw1yiZDoGgRuH8rzCnLfLp6WbkVPs2wwD6+RmAFSdDyQQ9nR3fCukVjvcyRMOM
Wv2Yweegei/l37SixFvMDtZfovF3srZFfGlTwYpTSYKF1Pc3LKLS04SWOFbHVIG/
/PSisGYtu7wR1DLnVxnL+85p/UV/2bkxVmbAxiN+Fddl7/W2B/VD9OlyLDcbSAiL
buMewvySSOWsthcGWO9chNTqk24VwezfJDoRY/16N9/6sFZxdP43y1TKTxcqrl72
yuclQU9hbd10qxMKregbGHeY0ceYFIZe1rX2VPvLLfkwd5u7sIsmmPRW47MJ6h27
ZD5VU2UrBRZTN9tgFWGk7KwpjegAE/YDjuBxrAIYIaHHdSTptc/usTVfxpc4GyMN
sFt49f29Mm5IVVMsUPekIMfXNOKNxiFSnx2s3+l8R7u9kYsxWRLfYk+5YMBNQ2Ad
mDnd1UXsa+mBlQ79thk9oV/3vb7cy/UDEKpr8ILTJktvSEuXbrYVVv3tgD6bJXAg
MdFK6bQRIs60pMiudvfmJV7ASv+xh/t/ZUBc/tDLBf1icNPTMJzam+PqbPi2WvHO
3PnFJZbZkbh/7kOXxjmrnkNyeKGNXneKlBm3JqbHdvLfiTqrU1rwqLTTvmIgkE3j
BK2an/MXaU2V/ML8S56EBkivm4aHh+uJYxJEVLvR1PPPKP2webXk/674hRr0t6Kt
k7t5XEoHhhLil1th/wy8UxoRA7W41hkPP6rAxotrG11QUVcvY/7EuCB9ixJD4cCN
uUwbOEp+0TYXt8an8R5pneRB+vpJjKOkZauBfTJyxiw03MnBvAAn81/l8yAl/UeQ
t+ifZKB9ekbqnlX+5n5Norwx3En1MFJ82aTE/FhmfE+hWhJDHugP5ia7xRZX1lRH
by+Pz77BsNWm2pAZv+yX0TM9lG+kr1V7h5+g40F7evI7b16AhAak6rrEXKUBuolD
uRf679N4DTAdqTGZi9IFQlrOFmHjL/546BHI5YmiHCgCMGK/OVA2UOidVNs9DKxw
gQWF0Ns6n/jwPG00obnkZ8lfdZiSNIeC9biJC8mrNcAKPnYbzpEhuI7ERwg74srk
qW3/2iYwIGkOEAgW7atgBB/1kdvpS6QJy+whQZhS9tUaYZh0+A/1eHPm+PoePxoE
uzCgY9fYCyWiMwzOwqIml+2COwe3MRYDww+qNSYPEv+8or8Nl1DG1BB/JwlDVqd+
FmsHWpBNcnTdhG+obO9c+kQ5NZvPCJV/2kVTBqNM/YNy2kqaNkzea8f+77ATcsNW
bsT210Tw/LkhnhPX+KsQT7ENynDv59A97qZplCt6eI8IkON6crO0WPZYyff44lKr
e7+3ZAhPPAHhkeEBLZLYXvibmPju4FiCqSc/+rNuWOVqz6jZkF1f6/iqrRQvsE68
Aq5j1yd0eTBryOR80BB5qpxp4cP+iqrqG/U8X2I9mzaDG3jTq2o0YpuPVsxnF+Yc
ZPjI+lKWHZZX2Z7d6W2qzTwLxZjtwFEqroPz4mA/IQxFe/87/yhLvmgRDQevHPiD
4hirhSlmTUJ5gfWQxP2QUQy/Lpf6PsXzQ39W45CSQ2mSuwKHom60AwrpggLhcwXU
N4GsGOP5n0r2YqMxZhkLTaBXoDFnl0+WZkO/vQIL5nNCLGoPpOVNqrsQHORqU/qN
pCC4DSf997gyMruKu4gCLQSd9AYbzeiVMGtsbYyAwz5V35ySCgsWPZkHVR3r1DQ8
Ip/1KvYcuwrYqpMN0AHoBqzDqbVkoLJ0E8QLki1eBV3eMCSORzJyLvjSYKRZYloK
mYxtf+pIsbJcVe0nrtSfCCyBMPOVnQDB2cK1pMwnpCmdCRfSial/kA85HeAcNtLt
/8QCndIMgH3zu/WyjkcnzJresoBB6pJ5NvHwI808X3sWoOvV0BNLyeEV41e6K2Mg
7xVksuscFU2qy9Z1Uq2eLNvTzg8SCOgOcicMt0YRpmfq6Bx4psMLynuiS+nYrJQq
1uH41XshUH6OQdzxdQUokzevEhgAk7Pj3qDOthE7y7hhJ9n94spWejtLI+Lk/8kv
sF/6KbyLYglTfV5gSHkyPk2irAG51C5fz1Fjp4sc/7txE8qEN98qU9SJG5AwqyU7
g5zhRlM9C/21Wk36ZTUDuBEybZ8ZZ6ibZ96ZEpbXDKyNGSWhAIQ/BkcjumaTJ+w1
gl9VUJVFIkVxVKrCZD9gIrJC5VaKtSVuqZe30W11p4Hx6SOYMUxQCZ9qGvHnxgXv
1ByEd+v44hmG4h+1e8saH4O20yFg5Or6fix5B+/o0PLxJM1aNZag9oUjdnKPKs60
vL86kjjkPUhMQCAzJ/vvGAPZodE68Cxz+4XYyq4aDFkRXaQdIne9FYqkZ3/sJhR0
yM9Y3GOJgLOrHdP5JCgZD+jYf2FpTO3a7XbEwgbFotyaBMw2wKtgw/reQ6NvXOM/
vAx/lzKjYGNp0tMgs7jQHR2epFxKVIt8OmT+M9XfDnP316EPOG0iTN8hjc3PKJSv
+pCU37hu3RlJXQmt/dUVglzrLS4iL8ZyafWBjFFIzZhlwNQg0ZNiIaHM0ge+8WMa
b78GpX7Z9q+uxGiDCZf1EXa9SqI58NvFqeJMw+0vPGLm3zzUWB7cT1jrV/ZIZ68g
ah434JLjfmOHXKx1w0GSPyD300F6fwA3wyN8CyL+mjaQBJckj8VxhUQgxG2Spz4E
lDy9jT/CQuMczKXuPcKK0X9HGPqCWPhxudGvfKQxoQBl0KGh174lTbk79yAXcXsU
AKqZ3UIodE83pt6XJ4olaqNb6J1t+Vcqc0MWsFigII7expHHbJ1kCYaFrmUjaTMG
J9khZreVSDlk0ewyUxzytP+M1ock4fichzgsf9QEMEHz9F4s7re/3E9Pt0f3u3+P
tIAxiTvZSNykuhzagllM4Uj1P9IzisfL4FY7JZCD/q4EWKtaSxBjVXFyX1xOhS9J
rB+nIjVcp48RTOe0HjzEhNDD8yl7lSd2Um90Vs32MKAzwlUzuhuhMroE8UYe762Y
PWhMiUl962WJ4y9Yai8zdAybOjiVvo2vzqiekL5d+E+AGtKdJJj+r4XtF30EmThD
Ev3i1JWF/LRpcdqp3u1WLAXibO9qeE4wNbQH06XjSPDYegWTFBnRJoQI3YhauiWg
jqEekPRgkJd4BJcapGODVzSf8m2by5sAt2WFlNIy4RAhZcuv+yX0v0peQdmRwQSs
XBNGjf6VtDFYClgzUJnpk1NqxF9ExbVQYqT1c9HNWfTzMzcVGod1nYVOGFNKi1ed
nCvgMFtj5kbYeFmcEm6UlG4CcgI6SuVw3gw0H5CrZZtvThAtw3x3n6JR5dQzisGv
CZxKKxypQ1R1M7PM7Tn2kCFjnNv3G2dN22VpJGVDvV6BU2LM83XW5h9Cc/PvLl8K
pL8H9ujVKK2vdrSaIbn62ffbv3Q9TUwOEqbjB3VnGYK6V+AGPASdrpBRv/X1tvY6
ZRndf9oLjIBiNuoOZA2kS5AcjVjRYCU6oVtXhOiroaHhlJ5C7rFKYj6E4aP3v/dU
aadnYbItkWSrALN8UYNDfZ6KD7JikwMIsN3ZofLHmTRNvGd074rnMe9c6QomDBXV
SOALGvJZJ79aEvtPa3On+BhUlgmfykwss3niaZhkKTjvRRGrZgmRcsyLBRO7xHiD
fbblhA0OplRBLJ/TyaMXKLX1qK5P1TP4KK1fdZ8maJk5Z5SlF+JAVx0+jsz3wjNS
k+4bR/nQAU4n0vwJl5emOmkTtpYx3Y2jLjVqcZsfJTsrDk5WJuMvYJTy4M7Y3Usl
C6aTD+ft3Y6/97krEOdwbI0IA/Dmlpzfx+43nCEx+9LEcqlFwiAe9OP82AM+8Iud
wka0hKh7mmI6+6d90PNmJLAlbUQJWQfrDpxhMH8M/FJmaFu8Nap5G7BKg+dQ5XYx
DqEWZQ2LbLEtHA1Syb6XG4hkeZC9Y4uWQTnVqwbtKxZq6fqUIn3PsDMu0SmfspLV
kE8FSpuY5GyqTG7qH3R1dzGzC8KVFjMaaz1VQoUFQs/ANf01VIdxH+OyXRcCwkzJ
3MSHpPtHoLYZ0VdLq3EnRs3qZ9EBya3FC1pEQDGfnADUfMqoPfWXEHgQps1s1Kvf
ju5qW1ELgc8qjP1thK4mKvptOI4ESzXfkgsvkAsqTq/o4VPAxdftoi5mNg7wniSr
GvvLNkxiq1Rt6wT9E+ZIsyRAHmfQV8q+cgmrTkSYC0gz+4f085zLE3K/lG45nAip
MbQq7JZMAunr0qCoNK7s2/h+Wkan28k+QVxwOcDy0cymn97iAMqwICdEjMVIYvh9
rFiJUqa7gqYFc8b1qri9V7WivwRjYnOaCzOVT3k1TufGS9xKUciT06mAFAItfz9F
fCR4koXkBr/BIdF458c6ib6Yss68pE1qFmizr8yoq7RID+Ex5uZtl0LAgFZX3gEk
qpFmKBotcM1q/Igj8JG8MzH5HkHwf05HHjwy+TOiYaCOiQoNC9RBrwkxQsL0J6gV
U0c6h6oLMJR38X2fnIfj4pWZh6T27nsF20tf3ojO2QAKVuyDllEUl8B7H39qXLOh
BJtmsQCwT9FQY34c9cRJirat8sVHmdiqSBt4yj0SV+epcD9jRZ4quWldpbbTCjEK
ZqZs8xPixwcLP12M7q4AXXaKntgKAZHT7KP5XvqOYeCKvqNif6WCXjtXroIoaH/G
TaWiROECJ1wpoD0iuIqfQPcn1pjKYoxNOtOfsYwxbTw5PHFC3xUTg406tsKhaExV
//zZSVV7xBjd5r+oc0L6XsujnqK5c/RakR0uPmbSO9Nv2FoXh5qYTvNHk4GCZOS1
iqHp5/lZFPMQ+rCZRWx/gdZTWRivTngqgmxTVHxewE0FUMdmEERuVnfM5bZ6Om7O
Zr5YH8jz7rJENV+l8ZQtzS0KHzD+M1cTiKzDv4bGXeLn+/91kiPXAlxAhrelIFcg
PqN2IJj1xFc9a4t40OLB/7kkhiuwIyc+kdrxA9kCR9d34wMM/8Mk4PkPjU5i63v/
e1JLeegulHqfz53EazT+lK07ocWPPmfpYqKk3OgU2zscKuTRbdRnHrUb2EKjmH+v
1xUyHC6atQHeEolew0B3IgksQg2BjdmVYoPS0G4gtw6ynOE3sOy7HrV2OZrF6bmS
qgkAKUX3g9SK9js6Hre+ZVsGaOoOSyUffmJLm6s/3rPb5pihcD5Or+IvUChgG93Q
Bi2m3EnLs76s5rLsZ7VcDFRszFvxA+LwKBwwYpIojf1H1go5uXLjnUOxtKDKXIa4
m/vqZMCzscfSFhPVxBNl4X0z5rTH22sd9Ok5Ad8nmYHG1gH3fJs32HmGsgyt1rRt
Z6Zb9HU75heqdrQTYjCWCsr1B9a1c6W+uPUWTs/LwhBGAU5U759LEFXjGQCJ4YQ7
MS65VFVbWM0w2goiVP7qantyr+vWbAWRCtamH/e28OLyMBsRkm+h4uBs2ctR8zCQ
zWru4hUow6vckouzmpHV73oFq0qyFMr0tkqXiVo9Yy21SjgSn6+jv7ydvOiyH4Sa
9XvSECGwaqesrFN3jNgf3BzDoSwJ1xZD/C55m0YL/EYYSKWuw3ppZETa1ItB7SOH
w0AHfHNRF5ucs2YWFrUAokipQmv5ImhnUH4zFp1c7CVUfX81cKny/FaO+i6kzjOD
4XCnBbI5PEtsJJWNfAQB367Rpz5i1oc0Rpinv0SSEBLs/zApU6rhPtzWf8GIFVfA
27Qax3WZzbAvbQQXvNPdRItePDbfddnunWe4gAODomABTjycI1Rn78gIHnNJ32br
gVeZ1/eIz3Z2XpANZ+Dx2xi0ddiiUIAPEo79lgkHRwlFoO9gL9Vp4l/ArKGBIerF
EUjqgvzJiPvyKQmieS7ARyOh/OIGgADO5TkusW/TBga6L5d4ZC2RaPaTEKeWQwXd
n6nOPfvl8TkYK6O9HlPSuJbKNMF8kXBSwBKDDgMlAV66+N4J9Olccp/VuhAOxCnV
b26uBK9PrR+5e10PzsVjgXIpiwx1PQry9weDDEVOK9AYIUkTQSYISG1usNFOr1O+
nuqYFYSbocH8Sf/nBBsBn+iW3qiI8/seOmsF4mYLrbrGCKIiRJtkI56zAdnXdzRa
vmD4I3GR8EKZ3yPsb+3OPr8QKS/u0OxdTg2J+Qi8Rv3UBr27JSy4w4+fEqgeyzGK
EKd2r3BoZR2GFTPWLt0p6EQkv7GtAHkPNf0iwPaxL3n6Jk7iwN2bmMrbnxuJcyBA
yxkCJ3pRK4DpVYJuOSLemR2/coPa67auYRzysfbyilFS/dpQeoLkwR3XL0a6zrC+
V61kCBpoKEu8ZBffjE4oHvoUZlJ+Dpj+tScvtXyqIhmwLXBtQRDpsldp96XK9XXx
JKJq5Ai4X6Tn/UNnvAOfXG7+Xbkku+C7NtDWM7wUSRsptRXoUYdBQutpAKYaBfol
ZR6t35NDaQYG4nx8VHmrk1usIK3MQIRrF9SbSJPtk+DNcT3n1Ko8tWoP5NGgzUhq
Sj4m8XL3kwew5FWql1xTaTITvCG1dQ9ioBrQVVlXxAc8Ga93FTwYMUpBxddxtOIM
nrgF25vFKFLFRjtLKMqXyJxA9q4wtZNRhA1lOCkrSlQYie9UQP3zyz5+ZC+QsaZS
bm7eIs1iX5ImPBWJZnXRxB0mtG+JB7s8ONYQBgkJeXHOAMx7ksY2U5gvhKHlhq0N
E2JSgKDGuIHhNeVLOiQ4Md0lFOgEOQWPlH5pnn4IPlcPQ0ANMvVyw1b8TTYLnS3y
4WsQJgBQPbT13R4r8dfEc8rWlD3m1bogywrzJBW/O7IK6xxfDEedz3by2QSB6giB
197JQCzgYhlmxf20OWiOC9LxslqPsVNDoqMwbCig95C2YZw7aPGTudmTqrfd/Sr4
shbQGZWnPONfemmfIsud3q1imKQuDCCeF5NDkdrWBJhxjo4KHcxaOSTbak2cYN6s
vfNpSorJrCfz9qw2ruSbrx5Qjlqjp5x5yFYGa9ble4RDnko336avFS9RqcTHdtVi
eElikhH+VXaJQoEyKFNI2y5EWGPp+gShKuYqmFxiqFu1viqtmyzriJhgI4RY2Pwu
hFHKfH38XoP4t9UtC0URSnDpD6/y5YwL3KaGTH5yKvtQSRvqvb8NHsccAY/LyqPb
3ydSAe/4Of7FGCfr/Rn8PQ==
`pragma protect end_protected
