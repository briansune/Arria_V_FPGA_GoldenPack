// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:21:08 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FwQBx71AzshyNckWKV/oA7bGqWBl/NquYmc1RCTCZxUK6rAPQay9yfafgBLYpiDg
MwwSpn812ZzSCmEnWiI2Wg6eNt5G1Rcx3Vh5Ffqmg/b8wLE1l6bdIi6SLYXKI5rV
9QoDGOSBQBqgT9jsZVUkdiCOK7apKeLjpsBD8OQAL1c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28384)
Z84RsJO0Rl33xUX61wPoThlhrZjdXB7VKI+OpWGdJEMFPnuYiKjVPWhC32kRPaPG
620Ry31DKvAMArsAqlXdbkXjSOWS495luz6R3FliRg7nvojstJb8VRlxZ2TF41ys
xb+JBU/0fMcJVExq5v6CZnxsKI+MqZ8Kxww6NF/qBpNAiYhAXDu37O7179fykNAV
DgUgaO2An43jBuF+rshjuLHB0r1AC/FNSLvtjWnioV795n7U4RUYhIyXxPYx4Z/d
E+lpyMOEJ7E5qK6m27pS8CkWJuGGF+/aM8/J8atcnHYT1JhxaFG1VC03MIS9Uqcs
+oc8IRqEOm3Ys6Mt44iyfn/1WOjGXLzB/rPMyEjxCew7s32ppjkfmheiUyhijOVl
9eUHk7OvhaXgx6PMYSIwL+E909PErDfCjv8HKZIZJQhESG/wSD0JCOeltR+OPl/v
iPzFXXrtloozdYab5iukd310X2DoM1GKDyE1qWE1ZsBaonGi+8OX5Ln2JfwIaxI6
jwnktFqUAnnvTswaO7nSSfbzABfQoKLuUvQBVWHTF3Py337+CnGL+FTZ2VKeq0PT
hTI0QNFujmgXLQSIr6+Uw1blvnwyjKYUUH7r89H90k5vgfqrehSm5zUR7sYdR6jU
yfDnTJ54meElUWWVAxqwLKZVrMB6xpxb4twzRvXEpz1bfMvDQbVejNkIH6cuDVvx
y0o86CoBmZsL519wO9sufJBKvDK2Vrgvl+tH33WVFRY8lMBZFpZAVcVun6BBquPT
xHlAOsm3OT00xAPmOgbhObqkK7FnAHscsCb/sLPbDuXkNBib8fmBIkpaQS8M7Dit
TR9d5D/Su1TbbE9onB635ZvSP/CHKGi9mYk7xsgMBbqGDS0z/GftyVOrZ7SkUE0r
dyosNzSfSUqFIf4LRDKZu4Ws6cxBmk1kL6surbqB8HEunvCrg14htv6SGEdFr46G
s0w9alHue354mFU+BCgsVceu3CjYfgu7oFfbm35EBd2zvCXqhITNeLNCv/+wNB4V
jjB0kmCFH6+zzM9gBjov8WeLLaacXsI63mMZM6xh3WuRgnLnpzFz6nlPf1iIyXm1
JEP3ItUp3kDi39bqZM2gm3OCnzPeEN39B5S8DJbgDMfiS4RnJfAZhA2vifQVi9u4
rFLgOS11yt4IH4ii9EpQzUs3PiQXGJ7V1W421uozoHP8lJJCgfXCFehT/QzRYq1p
Vg/IQkg5rpMsxWIV6xzNxkzW7TeN2faty+h4kUKZDJ0lgFp+l3PkKgKE6p7wZkRt
ghuQovK2pYAlsn2khf0viqrO5rCE3P5zNmb37cLMgQnNO+4vaytNYMMA4XfhDGxZ
AjlwQ7qu8pSRuQ1fNcaUfpBYwwAZvRb08uWptgKGcadP2LvzY2YF2GMn2YYHUKXc
AK66owDDzgX/dkieWrXxDsFZKAX5o0KNMPr6eFYgO3ArJ1shdxSkB2Mdgr/5ERVI
VKNTbGSK07klwFzNc2OYaKifNkKy5hSJGtIgclwfeZucyxxaUi7lahXedqYG1l9V
jn8/x0fBXX9kpQwBIeVSikd6T3Zb8CtFr64kJEqm35wS3ikeH4vRfKWh07iKJMGu
lgNeAW8nmdCPZ+hc/60xBJHPXd2hGAQpq/02icKlcK4SpplX37TUOSECLzOMS6u8
p8KDsZJCF1+uAn71SacJgsUN41GV+LaBSznfUC5YnG92CslUVX1WAH7Jb2lRA0df
ts/sArb0oAztRRa1++1qdU6/cPI1mKdMWp4SGmxI0BsXN68W3+d6gCpKYvz9CvKC
vWQehspJkpe9GCai7X5eHlHbeFUE0y8qcKMtY+7+iZX2gQ8KxJu5rpPPDThwh+LN
s0qqYYcASo8lAUBOKJG+TGAXY/Pgf66Fejxki3HgFCH5kPqbcFn3hmL38RU9Kisb
ae0CqWUQri+OGE8n23uLhz7XJyiio7N8CeSEGZcZ0afMZQC/WqY6N0E+QD4MNywq
p/8qNyYj7FANS0iN80VUfP5nfG4Nq99r0fkG9KOr/4SGQoB81/L5MxFxN5RWaVd6
2aKW01fl63ySbM1qryNUHXWw1XWInyJielhlja8AmNZq3aMJnxKrzbLiM5Ojz0HX
OUYTdJoaAKflNYe8p8tQo+FJhaj+j9ljmb8t24zRSPhSonDfuRftWiO0wOsfYZWp
PXH148ObiPzi+n3DaTsUrlLlrIBXr6vcrSrSN56I/U2fN6DfWuVoM0vYdeILhKyj
RknVh+ptxqBDKCrUeUo6SQZzUFEuuRrog7MWZ8mdLJ6QvtMyhV8rr8Lgg+HMByW5
zXb8+5WXAD1M4ozZ43wZibuvTdjMMFZ19YTIW3X6AXmh5cozGxs/9QhkdMHplbtO
h9tL5JsvGV05h8ixGjnw1xJGAln7bY83/2L9GgZCf/ZwlsiGc0KP5MwL/sahEU5G
+zjDByOkr9s1Uufmwpy6vbYqbcz4zJOz2z81x/UHxfk6lOt2+RKBEGVbaSXJMBvL
blT98e1cwiYk5ucqfDgx0TKIzUmg652EW/vTBIJnDfGExVy+YO1miJT5Mk3NucJc
n+DviB757ab88O++HgJ1hCes3vkErWSRy+NlQ2aoc4RL+g2YyKQXi1rXuJ918XTn
pX6AKe0KHsg97m0QDvJFGB+ez+23Nr0+fecdMVvjBZEOd0MM84Ebjws6PYjLCOLP
LukCcUKaj7jSI96OczLVgMkTRxilm0kTkittxtGNOCBU+f/+a10OQKsuQC4famM/
mcrIrJV4vLrUmCbPQNub1MBG8eK+f7iSin7p2KR5Ijk/jR1Q+ZHsjUAm4qYmTg+o
ICdyv0UPHAG+0oP75saLHZlXoDWSz31V253w99u5Kb7tMvm2hzUB6W/pGUj3p/ZL
bQtUAN7fy9F+lQ7B6HLjDQRAN0QHwaGO5K8FH4maoaHlVLsS7L/icae32CMeval+
Ioc5zeSBAy0uo4Cc2kODREGZKGS87iQrKAThqVzjqFWm7q+x/pilW0qRwM3C1WkN
CDKkakorC9bnx8u58S+kXC24yoGAAELVs6+RHw+PxNjR1ZYubmjxD3WNRCXx876+
Xp4yS5RTbZ7LxqendQbs0PSG1xp0dvoUxmQ0j32j5PvsgOZZNuOaUj6OrIaCsmnp
Xgo1XevdtqTY15mgSVVfDIM4+7xp30LCxooL/3nBye5x+/J7xyy8jkZ9i6fOT4Sz
boQBnYk0w+/LAh6vjAK9JwKJarX0xOvCDrJu/AkbxS86x8hc8dPWJNQQNR58TeLf
V+r3pqTt/0RKc2fx4M3z1PaVB6Objq1onaEXUfnH2kIIpfuF9x9T3c7TOWL+DQVm
40K1teyfqx0JMUnHeM1nViAAPmYF/vsIvWCiYp9eJTpqjWDkdykldQWLu4S5w1sz
B3IrwIfNWc69AmmKvXtrPTitr3tbJMyk09C8ErwDu8nc0N9dIdzMxkeItZsoiFXF
Tr5fEYi/QBl1le7vJ1vobYBXGonrePklGfaWyc2aoR73lSMNMyEpUxUa/1Utxtn/
KvbO1jCAX8+yBYu78yS4PqMF6QbyNcjUn2SWW7hSkdf1BsEwkWM2dfDumsbp/GSQ
0izhXymBNlKdwLl0weImwvDYr21fs9bf8hW+1L7rOn2gd38vFE3ws4hiJwNGS/yQ
Ji6A86P1+Q12AiSa9cUcxonMqtvB1UhXALwCI9OngnLXQF3mhFNbalsHruVLvUim
ZLxiil9esuSpQSSRAkRc3CGzlgBBuQX52nyMNZkPJ7b0jc1oeTNWS/5TxIdF/KVH
nnYPwlwBO9bTbLIe65wqnTtudYbvnF2dPQc6du7BL6vDRxBejh499XpTmVOZ4Lbz
sG/XWfnkWVB3RQWYTXebuad2Y1I0cIMkPfLf0p5cP6DFylNlfaG+D7tD3kwx17qQ
20BP2pMKjn+gtPAxXs2jsud4q856n2/5L38jGbGiSIYidtnb9+McZzeksF+IDksW
OtCw6K7yZhAM3VY/VqAezySNR1xEsoqWtMLJDBmVf9rt/WnYag9i6Z1Mg2iw/p8+
YYQ2KcBYYL/1XBBV9avuG8q7tIqjsHfYErIlqi2+xWMiK/Nha1G/a498p3UMTYHW
PFoaT7COdl78w9kORfOITTWPYuJ6198xSmu1tTVsINAv3se2n+JFN/7S0DZmmXa/
8IvIxuhw5IRDp6J2T23XvAoIKbaOqKT9FI7dkJVat5XYMeGv/nF1kGSxSlEQXnMu
ElewsGdkRw+q5zjEaHX5gWm31k6mTB/CUMFPXtebZJ2+5IE8e7Zk7EV53oTGuKFr
J004tAGJKVRScy5JMMhXUNEbkXQ/KOn3v/dqzEx2hNrPNn9Cxa9p4HLsrTkfIppF
eaBttBnYqsG01zlK/WNUobvJR8FrZkRxk9aiGCBIHQMpI7xumuX6bPjIDcAHZuR9
Obd5KnhqFNoYu6Ei0sDExDRheXo2xNiSrRU+vB2F5QbuauW41HJGNEZJfwr4klaZ
WXLWGyVgplIJbTwabfoi3ww7Jxkq1jfM02m++sNz5CZOBKMm1+3zQbk8e3gaMI2q
5373zAY7+pF7w1QJtAhkXlQwYZSEztSn5OonDWiEzhtp/HC7UETbs7Q5Eh0H3043
iLtRG+hPMnfFkwzGxvegX7pcVgyLMNJrpC+uU81Btccs2TAtqOl5Qr18x+vhUu6S
MvBhmGkeAtcyYlbzwaz3XmsTF4nt9O1BRNPEj32Wn3XdugtzHZ3pdTcTUIZ7euSR
v/qE/k0UwxuHwns3/XWLipR/cE7cMvQAMz0i8ZGi4lP3HNoivqTiQRzJHEBwi6Ii
NWXTRlv62fSTzWyN2lUZFftJ1AEbKCpvIIgmeSQpwqHAg95ezQ09kZnKjeK0gX03
gukroQCmS6aV2ifo1I7a+CQmYyWjU2uvovMmUhk1xGl7Z8ZMtrZHCAZIrOPWZIpJ
R0QeDltDG03AO9AQjLQqspeL1YtN/kwMhdmSpSlDKttPzM/U6pHa/IzkrO+9tNhm
Yu2rZuY/NIoRBte4RV0cBMP6jiS0Jdf/saYftv8ruUIM+imuFHQzPGPVI+2+wwqZ
m4z2+F/Pb1sCaDAmc19BOEz00vE9LCNONi/YCRFVcplJzRYFpv3PLGawSbAZrhus
C1aOx6/IZlEqldEe/U9QIoKBOEf6hWPi5Lyu0uVsy/eLUlZeyWOCzYf5iV/Pknoq
C7OwcJsJ1krL8I1aPwxUGuEpT7vq7vbbT7zHsMEMGIhOs+YJ3uLNFMV/GR7CkZC+
mNVlGgIiUMWNO3V4SmdjuKOeoHWYLC/M+Jdlvsl7n6lDIy5+EBW9LFZg4Dcachit
Wc5Arwp/xnyQMNwQBqFSfBEh235O39tJsZPJ/QhwTeMlHyTlykIeSgBAFP0eGYbl
qudFh+mGeAqRNiO8FciXvtPooIRnD3qTLOR1bjFjCukEHCjHzvhKkgmebQY5lkRH
3h3JG9oJEfiOJDaBK4L5xNPjuhTWT0O493c3sGcSB8S+ciWcNVZlwJSTpCq04yNi
MhyF6f8G6ZOZ/5IMqOBQTzDM+WKqgH5tUV/CmctCcwhBbyCqm9ztZrFCZuIchT/E
Ls+cixDYTnto9tzq5ewQuuktgBawdUw1Lk45fG5y5m89MA42hb96F+5QlhvEBMUw
ebM+w7nKMXR/b+n1BJ20yAubNfhtJSsS6+mFivEQ8dwQM+QMp4qcUxFJryylLSub
TTasc+XYTr1piai+C8rPYVhKdn2RVC2g17i9IQvW5EBfr1RmyzG3Ohpd9gGU5jLt
3o/nQvxkd5om5UC6mxNEMrKimLaJrlhw3Wb80R3R9PR8ybrckF3ohH+15oYC4yvn
0Dgd6shGFEfxc6efEHk+Bv8/QX438K91GKYh5BD/Ot/i/LDD6nQcfUoVsYlKS3CX
TUL6EsZSEbph+7Q4nr1v63b4voPUTEQYBPx7m4lQ/y3iOg0PzfKR0Hn0Q+sqZGEh
lowK8W5y4eAGuY0FgyqKqXbo2WUAhREXrs1NWrOR+L3IevxxdAL6YORvDYMS7n5a
Cyt0cVg2gMwq8OGqQO2qPWYijT6PV1Q/GeJh54Lj8qcSLfUGsn4Cw5Ooy3tK/Hzv
gbP7H+xNpglmxPWXeKci0d5SJu/tHsYYZhvspdLytXxHqBGXV/1PnQKZWc0ZH+p8
Nino4w67AgEBjdjTOSAi3xbuxJIzGBgvqoJioQ5Ogk3FX+wbPS3QYYTLZhOY2Z7v
rVLK7Q8dMw+ttmOBday+KDxtZ3lDNLdKs3lCBORxQehX+iFVMrJBLtQPwPjUX/k4
UDNl1Clz0rQJfSX7llKZD1js7fdKbO+0wgEmLnVJUUbeZ2bIScSmgbQDIYR+0Fd7
rnkcFsjipB0gXl52EmoPVDT5KPPM+s5wX+Wgr5DT4XthczwzpBfGV1ocRln8P4ol
oS1R29CqqeJtg7uJLpnowxPOnlgaE69uro2lJX3ScJJ9HhKEHSuqWmLT/mTkdVj2
IqyUt49/yOGbIkzuOztM13Qf/zfQiuKliBqTWLVxeLiRU/DhIg6aAbej5KBM7sqj
kyAfSsP1ro6QR8E+XuL5V6W9b2q8D1wXppP1ude6OR2+D4eGtWVidNyWMCUt4D8o
wWQLy43rHVkrHyPZKEJJU6pUsmMkAfpocjy2C16DiIWL0Wb0CgM8/NfwpgoJU3dN
MknyQyLlCkujHIrHvR8ut510HRsyyIuSscsNs6GnQfxm3NoSA28J+QwzWJSeszbJ
KasPCrv+rg7UrqIUbbFJKOsIRUF0BZ/c7X9whQsV5c5NMc9G3cvdARuawHzlJKYk
J30z5PjIwWdVZmFEYXyv8HBNsICcVHyoc/sexrbHUBkzgpbbiPyp70rOcxKA2ZGf
+4BnMHUKqIzxh9xXf7jHhzt8Nl3RQllbmV8iMjISd4wEOVmEJNe2LyxVyz9jDyoF
xBCzIj03lbAtZyfJUTG4GP9xUdQkd7r8cfbTh+7C/BFKLGEOe7VzdSUtHcgUt1rl
knDqc4KxH/RoFVnRxUyzPSK32OGSKten75YdyUY8/Q72ec9ehL9ASOEs+4Zs81JY
kVW3e+hG/jtHbXawl8U7JXDUsq+O4JcxiSwF01ze38kNlHLMZg0Z7QIqNURGSua0
TygPfwmSavMouro8l/8tFeAFSKhi+Y0DQQoF3g00MIKfFMGpzm9rEW5F2Rk7lSN3
GK24IehjSUs3zsWSMaFs7wWY3LoffTAG7AaM/UOKgdYN0+ch97fk6hyv8SqLs0N2
LnTq67q0+PAFyTOHsTQcmxiSp88u1mzlV26OJbSqaSk/mdCkd5qimYP1LSG/ivgH
tvaUWx0tIzWnCNjL4Rs7dJ7JYIujvfaDjsnfIyJ+3QD0ooe+/bvsEPeUR+mtIIx4
RRO1SDX4sgSWEDhMuSO3g2iI0KMPuRqzRFM7XuxWpBBYxsNj9A2RRTgzwrtxB3/Z
coGKzSzDDAHx7fhuJYThGJ5m0+RJzrN+MuHjMv22r1S73FtHxZub5EXcBjE2ctWC
WHNyGnY/D662dceF73L1xTP7oiHw49sBePgSn709zuEWj3kDO1NyPbRM9W2TpW+M
9bp2PR/tsfMlrrrO6DXhqXD0x86LH0k3EpS8kbWV2slXl8cfgLt1rtKXnyr9sJ4w
6XZ+LKW27+i4LT0Y7N6W5UJ5RSmjgJh3e92EPf7Wkf2Wzkueu4kAlRkmUyFLlWkT
E9eHT6s7FNEQskHjfRBxdWqrifjNpeoqA1+W6tkd0xRnXq2vVSuo+uAfneMe7Hwv
kcE2KbdDVf/TlkbII+Tv8kKbuKJLVvyvcCUerK2uX/k4Xa3W4ESIFYopEq7TkVW8
dugKX2pFP4gOAXHL8Hmc2zDiEazHXbrIDOJ+XcYKKayZsjGYTEe8qxaONKNNLrfd
EKb9DtfIBhYfMBsc17OUE1s8q6FIQGJ4U2/0+jIFSlIxW+GFYPEZKjiCAWaKxhGD
r+8obS26QoPOpaRQeDzE4O78L5DnZYQqaqvVkfMR6AHam+ZNU9n9pBJqEJiabRZJ
1qSm5NlDxllTd//tZ8aA25j/PiLL+ssWl/yxbgKhBg3f6+1eVzowUn6Klvk2m0+g
LYceDLiH/MzIayJA5XQYjcA2T2FgJhkUk3upmqLBftztywosLKt28/RVAQWE1nB0
sNwRPMXVuwTCKdzSSLVagu8WT4ZepWTyyvt6CYGiKUEi7HSqREHidxbKFNTGFb1v
rKPcShVVCzXSz6xhg7mCXGulY1+0bF/NWqVSBywux5DBHTdYzE7UpruDiVs2Wb7M
qBtQ00uhXWKoj/ruszVgxRSQs7lz1xd0JE/6ZqCIS20mXp3VjCfEc9naT+jFKFxc
tMCfBud6V4B6bKSn1z979rpUE8ptSBJmqysQ/kQaF3ZCFbQgFMccS8rMqbXvcjPK
YaEkv31fUEH3AIYF1UhXQs2zmDuxDEOIF57ofYwPhOk+/tQG+F1cuqm2J42aXBx7
5vs63PvsHrfNV1qwVEazFwB+Yw8tmN+dgpxSwumM8CvG9o+cHC47uVguUbyvsERJ
O4YFt2IsWcPUPhpQovfIY2mff1V8VfjfrDkxh2QkPfdNvHQxx7i8bve0ZdTdATYV
mZkzv8TzwSYfEeXTnh7LW37awp8sLsPetgZsdemavcyKhyufItyCtQG2Sg7fQLz9
eBiiBegEm0AaBkUa3GZr/eO/kMaQg2N5dHs4T+yqrYDr7yScAjcS8Bkmt82g3Mkq
6b5dhCcfjHUGYkeOy7iFqbYZ5mdUblslOMnmHr+iW9ntjCsrp561tbGFP9rxTGgz
QYwiDnPq/xVH6646ml2VuHs0P3NkKxNIkGRIXGbBTX16k6VeD/87gxvjkkLv1Gjn
zVXzUpLiiMDAS2KKYf0UnyVeucwXyldOsOsI90GigMiBuYGsFr0yx5IpyEB14a4j
EJZXZHWTi3ti5+dBBDG7panq7xmHx871BZ0ICp8jVVbcM4cXdHoVkqBHczbKDh7R
SGiYSUky76b/dRW/L36nbmNGCkdaahVkhjcuhkQHCwchqKYCqxxVWA/hDUPLw/yx
htMWQKbJ3GAdnza9rPBKSu8s3Lc8o4Vz45Vyfdc0e6H0+HjufyY9bjHQzDYHiGbH
eq6/3lJ35x4MA4i4mbtb+/i2N5VDHkQIifMej7563DOKKkn/wBhT0l6AfZKc8KE8
ntGnjS8YBms9qovK737nHTaXHdsU8MGxH5zMI3uUeW4M4a5fwSuTr2NMJB/3/la2
2IqRUXjvkaebMS/lA9hDeo24p0YRjEELZ63qM/FBUewFyp3WgIyEMCpqeyBqsrX7
kHrxWP6Ta7wIXYuLuHeyZQRIWxWI9wOlubt8Ito4UxMliAEx0E6z+w+6ER8oS7Uk
OIJsx9hhWgGiBzo3wJHLhMMBfgTGqcH6tjA7p5/OouYG6pGe+cYUnJ5b5zptnSUO
ICUU0SESVIM6ZytNqTyIq1r/RBqgZNJN7XJkjRp5Zyl2/1acBQ8d0hiXX1HJvV1R
Euaa688++oWZtj8d7Mnm+Ctpj2clwh0Lqnhg+Zt26hMXlrnsBx+lej+1DUmsEinj
qJA62TLtWIIuI1lj4kJb1mwjktBJj6wXkxydSaKzy9Y2nY0anM41GRwleKHB7JgX
Fy+nNTfh8DOuNyoF2g3w1rET0t6mrBNOwZHcGPQS4IhhstUw3kr2cgYbIrJoLS3/
W0ndfHOicK9oh46Hn1QcwJhm90qBy9gnYOqd5VXsNAUag5Dtr2/+drhphNVHa+WA
jWFDIX4SU9X/cimP8gzlJ6P67qWzGicbzR0XcVImUQB3Cp2TNDAgwpii7y6y3A7z
xaurV0ZvxZ9tSoruwvPkdwCNP9V95ylLeQ0MEXMayafDNaCmFke7XHwkjsQzQE8T
93eVIKx6HsSAWtvTW895GQeOpLqHlp5AW612ri3o0/PLRvnxgJPemJ5sJtxx9Vns
YNJDdaCs1is161Hkw89S39g3nTq60YjhwYeLVFA60B+stqwJN2iBEeKGn+N1BiUA
jDPrpoj2lZzEckGnp+YJVk81FqxC31wb5lqVnTB2jk6DAwgZVHD3ud5y57lDS0Sh
Bf7oGJ8DnHsiJiUgx2fj4EiQf1zQW8CZ85xz1FRR42FvHTFaOpuG9e6UKRTRnymV
tVIDMzDgBgbQ+qlWmp88L6TCVTPOyYg8sNtANbyHKm+jWlF0wAWl0CPleebNQYYh
Z27txwRJY1dnLEHqBWN1qxkhLEV2y5Tr4Kkh0z2V27P7tkFM6IP1WREuRz/5jocD
wAoX1acqPZC6FMNpp5G72Rm/Y14RpWUUUFXD8ZcUnmFEsqBHg88YrbMCM33MHDcl
fIvJv57RsLkfIEQC0wMInVxGl5d3pNVRJatrcnGJnl86st4krDQJCusi2LmryWzg
WyTkw4qYmm6/2gDxJr/dzdfcgX0hxsJUgwdHzHMw5BNWv2GkW5ZnxW5QnJ9H4EDy
irRyengtyQB+VF0mNfKzduI0FXPila6Oah3FHamPJo2yfGQcT5e+24ZhdmIGXd9q
k+ravAwU06h1VovD/6Vm8door/oN4YUqUvk6yNKJPTt9iDbnsJAOt0hCU6qDA1MI
1P661371nw4y/ji3xZ40PrtAVNX073dKGfNQWtWEldNNFaPPYU1eOI2e9uBcfIO9
v87rF34JYJ/WKYD9HYSG+9xir7R+10zyjiV0eJc+V0Vg45XNs/EOLg1RDXNTCeys
aIKMArl0W2YyKxsWnstTuTxEz5QRiZ5CsrXCx3wI1V/SHZwd8jR0HzRXB/80d1H5
OODEUnCkvZ72VJIkv0pPkFmtNe5YeinhKn5SqDG2t/oLeFoCpvraNTFtkNwq6JfT
hU7slledVkQyiqK9pW8alIHUUfJ6F0RAA3a/4MhhXqrxQ148FwW9IYPwvbD5Fv+u
W21AGxu3ZJBroiaA9x7zRg2wiurX3tEAvnD2kunn43IjhQn6Roq1vU4JOzyfB75u
O/9NH/6lABEJdUC5S5rCVbQe4BekhHeFP/86BCc6pfklaVdIABcPncUH2ZKPWL99
6UXmPD4NTPczYHEHkffbxRX4U+clvik008XawDaApjv1RtQYEj5hfOTf4x/de1SX
OdZUJ3nQEvOBc1Di3PgtHlv+gGsINWQdithKP2khlKUfTsMvwfzOdqhXY4Dnk7lb
y5w20Qh/hoHeLqo24BaW5lGpA7kbHQqJPUabVcIBawao59VQStYl80XvLxzlAsZF
IwivVEzrzrZ0vZMIrTHwU1J1yihH9OUyFEZK9+jlAwqp502pxUyGl5ZSTLpb9Z1G
y35eFrvDKPT/jC2fDJBSYFpTtT81fd+WVtnbowM6daHMBiC7XOJV7QuNNIBiKa7u
N9ChdBEYiAXDfaxI6uoGiVJiMbuoteRB1v3qN/j1BLqL1lRCWPEQeEXjnygTrI3A
j0G15/mmQk43PJAI4DzBpPW7HcAa9q/0MvEgZTzWI+Off+eZb/6U79AnFFMXJ51W
pT/UjZrOFAf1FMw7pDG3MewKCpatX/I3w5QxiZDiOz8k1Qz1JE8qHGOuMgCN40r0
hz7UiHvdEbpAjCv9II9Cv2mNjs/fAIC0NVCi7xN1LBR8dsfXYuYiMRhMZWw6MrM3
3XdQMPTyIg7cEWhdy3BbMtGHUx4jh2EBj/bVWWHPqh06VyWnuE5nxO0/ryqissLg
vH7r443lEG/TIdjMXZWkzutrT+mkRhLH469+VK8YsJjl6gNbgT30g1SwYbKZqgG9
8sgRT4aRJVKLMSehv6W5oAVpSLYx2dUbtjXGuVOfJdZ3ro2Zweatl8GpmFnxXBiI
NM6hVEQXGXYX7zlLZ2UuA+9GjSpYowzJSH+MqGNSOMfyzJT3e8q9x25SoGlJIrAq
MCgwe0o8gVDxS7q7Zvq6LB/I9wOuPkfp/dxM0zQ8Tf3nZgFrNujvqXjoIJNo/LOI
aski3NQ5W41JMdaGYP5a5/X4kdinB2u2z0NrFt905INZSBF/4UtZS9XXdoSK2jHK
w39Juw/Bwm3jB8Im9ihUjrSAO3El6cfQ9l8KoEy7Vj2XgBoHTBDq1rnLvhH4Bc27
x8Uv6he1YNkNKtnLdL7YnelwyNcAzj/ElojXXc6B97j9nIysTyYCtqUohf7LQBJ4
7nUZfLV+r4Xp3aU/HSMBr7SkZUV75pMiAhWDkW4EGcn2QZ8b0pA8FzCWs0tQSQk+
xw7JfHH7l+1EMnTs/EONzK4btzU3gFOZSTV8GQg1l3ms8ZSLEWnkadSqnIqRaipA
fEfggYkfM+By5GXwzbWdpR5DWM3kPFPgKgfaAApJsFdOBSAJcvzUG2u+AmXydc9s
XzyWMzECmBdG2APlAp6xnZEVpyBPkZA9RljPNwvta1eQ71M3rvD7ITk7HRhsfjTu
HjPKxu0Iv7YDLP9FY/QZ8wlUgXHU8qFI+o+bt7IIzULc6gK86Jdowg9/ZiXJ9yHK
zYbk7Ad7zaOGBiIb8FcLKyNy/v8HBLVNcY7EuSafLld/hVJxbU9rjH6uZFTbCRFy
WGGbGrMyk1lcN+ggk7nuoOE3Ax3DZDLWaZgA/4FL0IfxOH79VF8MkgwWyfOTw84w
WVkO7zgDMUFtkVdqtcoUU5wFsS42h2Y7kTG3p1Qz7jkFtGmCikCQcenQixvKgqQ6
39IWZIFp/IDaCXnci5M58WDGqzn5OkSOBdEdXSKwXsokGfs21EwX8c99Z+/RHQX6
fJpjxbUF6Kmfux6PuNv2AcWfjK/+Q+c3aT3eWvXzaaiGjAiwqXYXheeBpAySmiW2
5O7notgemGByzbgf8waimiCPqqfMJu4RXwQly51DFF48MZX2Fso0bNmd0X0ouJwo
kMQ3dm9UfaQNL5gbhw/BWVNfCIokFkJwEcFmRfHrbIr5fzPixhkHK4esWZfw32Wv
dYnEiEL7SJf/RUh7RAKeq5eFZLxVta6AhL1rEocpbbh3eZwHkoXeQB4w/XxHpW1G
LkgjuT9oycB+cxPciboywRjY5lV5ixgptlEww1RqhuVvHOcw78YfhIMIB4EKF7sb
wZ0tkUElhUw8eFaDUmeh1pKXYkl3sE5Peks2X7IFTQbsYYKROjyJiDoTVYPPeWA3
HF79anXjsMuaRwE4nQywXhsCVZDUcIt5ZVgMtFOQSsEF+ajYhvOd4r+F47hFxBSc
RmhiSV/Ma21MBZZ/TSGMTTrokzJgSp123JUfSolxKvM5zDV2hUnXEX2sm4qh+rWt
Mg7Qa2Fuv9T9Y3OBoDMeKOZs52nlqnP7FKXaQWmMK3pKPNP2TiSLkecaNH2jjmVt
7sz7PxfzPN+NqGbf6xla5e3+AJu4x7T8hfU/IFKBK8riCIJ2WLQM+svlwuZLWWHc
T50hI2FMJHVJGL/RFjJUqeA7uvAKZV+gyESGJEt3ReElIflBVBZ+Uj1PqUkFRC+7
bsLZx7XbwwnxoUEe46C/Efh36jbVU5fXiBzNR8BE3wrWrm3XJRwK++6M6QwE5Vd7
rAldJf+QG/7U53W57aeYAqYN50jcsQC4d5XQOal/dBDXKOs5ejqZMIhAZ7wlatNL
NoRdHi1N3MzJCQH1IkQhS5yTwxw5JlbUZ1Z2updqXHr4MSJxtwUYlmX/m7FbUN4a
JeDZCNIMsjLOKPq/35bUNuGnSHMrR20zAUmkU+rbtaOfdZYqPvz7Uv2VgDu5QC+8
CFIrY7OSfOaHWJsh9opFBF8J40bO5Cfd+cF4ha1jgq8mLwYmnLU98xDf6WDeNLz7
r5suVBWXiuUruihU3m1IY3/7cqDr1NDDSEq7gXN9HqjithduHuDwK8UMdsAYcxaw
h0nHVTnfotZsHSzvLoZWa/vJHK0MBOrvQ9ivXkxlTZzqwmyyExLpgGy6uqaEeeEQ
lmJZOYxm44+RvZVj9UO0VOPVCcT2nCmP/shkni4TnPFXUaSMGdO9iIYHV6pBx+zR
yLZk8IoXlMYgvpuMv9/IseSI2gGGgaLrPIKBtv72Ub6hHxPwLhJCohfkwAfBDid1
ny+RnjVvtcXH8DFJYNJNK2n0D9Dt8UcDxw/fXWdmQvQwjvDQ8E9AVqwBi9zZ08tW
ggAjateAufmwmXIpT//lILiqQG//IFVnUl7hr6aIPHv0CNMOnj6ZwONvjrrMBtdX
aFJSDy68ByYUt/IpXanAmMzPbFfbZ0Sg+NpJhRBi05PEwnFU0rQd18k6jYk064l4
qe1mh85/HMqs3N6AJm15SjdqQerfuKL/L8rtjr9ZBAHdCU/v+c7GqxlYw2o90e/7
qU34hwYFS8ak4eS+75K0ZzrxB5JiOIikZlqn5tlt9yV/oigtl7lq4ouCqqjE440B
IppvDtdXcaN3AlVTzKBlDVIjJdNMGThef/xFt9M4InFDmgF7X8E4fh07BPXbEBGc
aB9wvmPM3LCz8TWS+wBKUXxQs7d4B3fb+zIKHeR0csoNp4b3j+ztqw7ABFakNKnB
l4gEPB4kHv//IABODOPoc0veckB0sKQzCFUJTPocyjVEidp71o5oXRljWfMDq1tx
CW9RJFYo6iyIxFrwQNHCPESG6pqWWpDF6fnKoePJhmmgiHkQGRC1jJR1h4g/K+7K
k+CVWc/5fCz22kywjouHg3M6g9Ap0Lr+pWomX32ZA49Nkm7kq/aBoXIIGNYiqDWW
6C48uBlxSz4qveKz0rY2FnK/JIieYrhEGxOBOmRI97Mt3R8oP+d0tqTPctMqEKnV
I82FBKHlfnVNsBxaRtDyCBQ0e3xSVKCOBvTB4kWgQkG1qud22jAz5q6g9t1FkQ56
FWyjO7bdviezwz29tNTzxpxmUcmUQfyQ5wmZ9BsnPiyDODvofKhGpSyI1Dj1U2p2
l7kbAlXmjV+aqbYF9mBT5Gt919Iz1jXiEJFxPLdgdcJv5RpfDjv5orEC12mOgLs+
d9pve/jtFVFKIE1nWVE/1OmCTau38L0FVt65rAiI5N3webU9WfLGAyWablsJs+ja
hwIJNK/pCpvI4UcuN6DNMmL98l92Lso+mB3wz04W5mNsPXPLg5cbDC6yVD4EkQO9
SN75K4GQGStG7zt8Q/vJEz6P/x5eYYYz4ZkZr+3mzaZFZ4nWYXE61OLOr5RFOhTy
fP2THrGY1LBdvn4ox/nmVj7LmLdf33HHGCXjViGAXVNvLjW/qNs/Vl0Ee/y2gH8V
IHlItAuzaCtRc67jPVPeQGRgq30aRp1jfzQ5x/8wkU9TSW/seZ0Z3JrRbOElyaVl
6DU3rprV97kakNkSzh63vfP/FN08tw1S2aVI1bLPmrBv+KcggtQbj37YJSiSM7LE
zPtNtvCWRQI3EJ/gHbc3Or2svavQcQRGFs7wJX5Zy1+pb5h7WlW/pvEpVjcfrg34
s19rRL7j32i9bPKgTpkEVR6uqKYyFUAPqUXsdhMRFUMQEi681sPUwMiu+ubXK7uH
vC/C0hCNpBP3jIw72nn+GXmvXVGU0oGpVHYLY3JhhF8uz+61EgVH+1QTrbn8Y3t7
5gjoR248ykI2hHagZN+vMQXNpA9LqmKDfNAmyswJCCK+1ttI3V0Y1BZTkgjF/rFJ
L+7ChbnWU842ce8UmdMG3njDle4e9X9sB/jqffu/MAJ+FRe1hWsyPrEGfXe4ReG7
QpkGJN88f3vkxzVmX37NPpxK1HTkhs0oAPo1QN4qobaBFOKv0p+y7YLaaxuzqteU
PK0YTSY+cXXm7m+pRawUgGWwB64mUS1Yli0qVCQvd98pA9hrfuh2sZbr1Sgi+bFB
0dNuE+CgGVjH4pzS7W2sG2NoAHzx1Pwnj1aJKndvaRedqHXf+gYNNYOxBeFF36NY
LMAH/fA6kte0IUdWZ+gvUc5y8oY4hfs8arVrtKqqP1YyNctRSVavRlO+YCIz8Hcc
BbVoV5QOuUzCpHchqfwwVKxcaRy4p8zvZVuOuhdmRSTiOacjE1RSO1w51HgZyqbv
pBubMnFkrLjB1doE0XpXkoM8PUyUdxZl9eSRQ3WTMrAsoDUTZDb3km7RkX3toWay
cLEY1bEsPrz9LqqBJOTobCXd1C92loo5XWayJnI4w6lHL0TFrAC7BYuColaoyZDS
3UPvK3QANYMc1Az9zmJuhOFL6LAUx45di7GYimQ9NZIdELP9XAa0aO9hQu/RWt6/
Hmb62PoosQzP1Ed+Ar8xKI8M0U4a4YOZ7ZjhwS3YePQAnXF9b6HDuyGozCTRDDn4
qPPpPCO5X/JL9Dn3NGauqtPSY4uL2wpccc5i9cIR1ZuffWfbwrTW8E1LWR5mkyaF
8Uxa9PdWsWMtqrf7QyJ8kERF34nIXhoDpu0O+XKhs3PI0mTOLsUs/NQC8ss13JeH
/zI90jLXy4ICfYXcYW4qq2LxCRJ/IwoNnzVPwWQY7thbrFGgszJIztHm/nIV7oEp
s9FJZGp3d0MKFUE6LM7aR53qftQaSZSbAjP1sSUdH4VXFSnCjnqzD4c6Hx2vxYKu
JSNNkZup+b3FKDCq/+mY2VgCGtYG+sYqt6sRY7kbc9mK5DwTdrntiV/lKO1TVSMm
RfxzaTB50mYLIzHwVSX/jHDBkDpb6NknOZiAUHjC+dOCg4M2Vi2aBZa5EKYI6c5K
NSA34xuVU6vMPbyM23yRsqM+QVeaUEM8p+/KZkIn6mz7UhFJaZKbq77ZiCYgAN8J
PPLJl3F1MXLEyUNvFnyj2BkNnldtg3x1T7qM7X+aoc3D14Ep90jMkHbIDCV1dlqv
MLhInX2a3Qyz78nTSoYR+fGDNtcWaN2SJHZ17Qr8+LL6XLG+qaBN+z0MoORLSHxb
uzazYcdrjoQXWmunqSu1GPihRE1A3DaVhbmwpjJ/syCaxy2exEWLmT1Rjm3vTSkO
Ccxoi6ON8bkYtAC85BYamYPyf3W07hj9ZzrlQPuK+tGOO150T4EbGQ6nQKv9t/GW
PxwNkYElId3h3w3C0SSXwAgh22otLa2wXYS7Sj86wrNRMwePMpHIB+h77vamtaFf
oL4m3GCGu43W+JD4x5ynaw2RKsEYfbGOsyAXuGSps6bWy5AUgO8eWWedXPfsBDyH
nbh4sb4oe5VRZZw4cp+AT4DAUztIbsheNlb7hiETFaak1weosP1DKiZLUnyizu/l
8EFl1sH8rk7tfq/Un12QZ8bU1K8yLmHYpui6BkSXcOVk9zIRyCgVylQ7YKdXBceu
gAvsmIZ9e+erIkUoL3oL8kfECZRLmizdKL+mt3FPjaR4AzsvC3MPBEF7qb3OYsXA
WBrTtGTU0UEFpTsBbiM51RgS0MN3Auwt5Jh+9HGpm/DjPkJD08KCOdgpzigtMqwg
D7vYveP525YOv9xcKSDYwdTUMt3If6dBYmMLV3WfKUdioWVXa7TAqHN7Yz4DlmRB
NebDZQBaKp2gfRydTLoBmdY1XoNlE0ht1eplVCAbdnKNSKENfWR5jc6jQvH11P8w
1CZ9EeGLADZnSN4b3uTWUTyI7+ZHaSwNee+xVteaYi+ilGXLpq8KWeyPL/FaS2nj
Uhox7/jm3Y1LOB+2YFipKksPsVQ9dL3tt3rqIQ9tTzCl50x/7SHHuRc/pqZHrv+f
gbjy/w/aQCtHu8HedXvy5nswEqNYmEAd/+bwzrhGFpTFkN+n2I7Hiif6fQm8zmYs
W7u7snCfwp7Www2mYzRV1qxUS8F6H0LnmCgSiZZEAm6zB8D6B85U7WrkLXIr54Lg
nJKLKvZK87UdRX83o3GA4X8Q1sdNkvJatC7NOd4ChIpihWzrYXX6qYmJKT/NX8Cv
UZ9voi5osZR6C66JhY+A0py0VU6zydGeWdw+tfGJMAXYvQo6UvWvktkuhqupEmei
oSz3lQd55jjOC/S1+E3kkMjg8dXiGzxHwqOf2OdE70qR/ejUcbYev1HLthU3gImk
9JWlVlRjHMSqIYwmhTly0yj9dfZ2OXkd/ZYMe/exUIQb1zbMA2QUKZsiDHCMl7pX
g4LnASBJKC7aqddrO+bNlSO5u5Cz2FO8/WtBdomaWpLgNKtAn8uWQXOnguKp3J3M
TwrbrfI183ybLqHWySoTnQ3Xq6kMN1e06FwQMhqzi4yTKuXjEoQAYKIHRLEjX/nt
amC3y/qTPlaXX3dYCbHVCN+DbNopzy2Ao0mfnDyGOP76ckWL82/QkQOYJpoVkpwc
ZJE5Y6XSnfAkKBm264dLBXlStM5FpkI1zBbZz45pfa0QHoj4qH3+KuGWvVFeXKay
RoGA0Z6M2yCysxJd+NrwtAh64rLLmBJAkci0fpQse+7/TxZSaqRGLBVwCGhwGo8W
U/I/AO+tcyDlHhJEPv3mfmD8LAGqowaCaImJr51/b94T1ykZ0qD3SvqyNN7gJnNf
+jHpGG9tGIGl8MAm09aYTPq3hjKGYtmv0cVWCxU0yATu85Y4lXEZHyAN7Fjn34pG
5YZS/VE+kUqz+yCDjUxppmFjrwlwOnICh1OfVmhB8YbKrMa3RWme8T+CG5RgwfCR
SQhtavItvctqIRnxJDwLSzSKiTjFbUJ8bXmxdu8TSV/YjNKLfx7SJ+tUV1CO7tuI
FDyIk8+ZoT0vpdClehMcDdPMW2IXlbiGgFm3rR/JTD4tq4sNO09vuDn1R3Ln4KDB
D3qxFarObfXDOBJhL5gbSjclrvT2JByg0bNSIHPGYuGAszP2allDbHjjyzu5jHIV
CmXNmmV+MV48RI4/87ftx8IyTU3+47rl5KYxWNFft9x3JpUc9kRMAu5onOdHSs9L
lWeN0KuVz8FGgRZQQAAkdNR98KD860OsMX8lYjz3ad9IDL33asnhQrN8LQ+7fr9C
2xSJ0Yz/tzViYQvl4meD6nyU/L5El8iIv6MH3465cZc+XiDmSrqvYQPNw5j1QFgJ
kaPbfjxyqdTZ98RNd500V9JgA6in0p6hw1TWAbKaWlys0tW6EoQNx0VAmvv0irQX
++0n7W3hl/PpxsGXXLk3MyyOngV3NAYsa6UpI4q9LAmR5AlbZkKFjY0Rto1tpHfO
fxCiPxdnQetIi5tN2BBy06IL8D9Kqn/NfumlA09tjypumZsHMN5y366B96ywv5wh
TKDNFlx/hjAzFudnHiOKVyDyIRT0tVCwc4LjCLNqWpcUE4KzdBeUsEQ5SmqijiZH
TscvQbaUg3SHB2Ag3uNQG1h4QUerfRg65Hf/XWhybiRPHKCB/SYt1edSMTApzBw/
QI6uXFMZ91oR+U0Lp4WaYmsREBzpsUHNQJwp+fhX8zyHxe5qNTg0t6pWVIgU+DjO
a0Vu9bd9WAFmVm63dmQFZz7KAOch4k2hrlRPtk3gNFqGi6omBQlXbW7wXfQsLrd2
qiaZeh16l/rV+wzGy3NxCJsMGsPH3YRj57urFzPgKQpbu7dG6/lkh3BNeUlUPlEq
0WYnI8VQ/iTlrkNbTbRAkegEJZF4rKV6tVLpbClvgVWirNWLSWcmkLYf6gd9eYb2
Gy9Ald9INz2HscCkqbF1/YTkxGbFO3qUF2mbaUhdvGuttcTZPD7hCW7uJVI2/dum
y7ghl5VhNA/mocv4p6xK4BhIXz0avEmZ9TUxuqFILwMmeHuOOC3W8rQSXkkljLDR
7d+XkopSUEeLBVDY/1gysCylZCa4TYqZ7/aULjlK713vjtjynmPf+tAegOFdxDeE
KGBi25AOQLAPLjSiTWVvmHywmX7TmGTUIlWDrg+9mMF7nl5g2qo2/mgTZBLvpP3W
SrTh6iXlkEeMHNnhNXiMB+Z73TaTxFQG8KOLkxunMpMMTUj7DU5dlRoOXTvYYpev
bPIa23545/2mR0IWk5eVc4Aa5RwzYI8nYOUzajo4dkOa7NUao+e6U4vjF+HFnG9q
aQyMMJ/2X1IlCFzxwFM6UFbEkNd10XpoSmvS8Siq7z+tg21i0hAa/tKiI1smrqk2
8tVmMBLe4M/dIgZZWnxyaAvZMrL88BAGKc81/XJBhIFUDuPCrHMt/IZKOBZUTB0u
U4ATX8r4U0c5AmFu/CyYnnJckQOHgNpDp82TW+tob5swgHK/Evy2SRIbi510LDE6
gjPcgMpvhGG806s5lLV4rhkv428zno+H35wDJoq4oZw3LkV/29ZjUaDax90QGGcV
gGWkXKNv0I55PLtCggieTnpQTmMq3W6m/qHPtS2aYl2RD6VayIPXlS59LgggaIV0
0WWo7uLMwLZLCR0vqSGbTglqa6jebnpr0WUarl00vcVIr4QHjVKU66L3oBr2umDT
P57Mg0rh738irDW27ErC2jwqLY4ss4s+65UOvhY0XkEWTzq3DlxqBUSYthWocypX
7L46pFYU19jf4bbFvetnMEbUaemRQMY2CT62nDnQlgskxx6gDukdnEUrQbAaxRVe
K5rfsEeH15CvZPVnzL3GU2Aj/v1nKfjyfh0acAelyBoer3qRUT55a289bZv/Iap2
VgwBEJzaBf/nPo0NyrGk0mFSMb+0/rb6fq7mIpbitoGADkry8Ed9BJcUbQ8tITdk
pmwxuHImobRzAqBc3MrXoEgzBe10cQIBLIBQCvpBdiXgoZy9GKyin3S+6+94KFX8
00uRVqXvvHi1ToeZnrhzTNP4Bvv7AKj2op/KMFuJpmmVoytGtCdTjVCFx4IGsLCx
iRhe/eUUYkKbDMHDtEQb8mIisqpJFQNGFOSHJw5kKxh7PREqFmf23skTZi0lV9Mu
V3yB4f6a+0V4NiA9KzREzDnt5MSjKkmXAw0WtoLQmu36b4yRR+Vz5k5FrKuW8qrp
iuHqpROp273JWYY6Me67mUIu6BEA3HUqkU2n/Djn5LGA2LNgXjUbMGjaBS6B5+l6
bmrOHdGDpbA6QFbqT961gZ+yV7TjdkDU3JCS+NUXxM787ORkQ/pa/VLGy6C2dmUi
AFbfD29t6H2u7R7Agd/2NpIcZxvInCSVG3gfeynSyB85HLbctWfc7Hd5/Jh7DdZM
HNPnKWHQUTR/ZTZsentRI3h6DrA22G3jNKYXTDnuGlCBopTaus8YZOH5EjI94ezG
9sziuOFOpXRg76RhxjvKdECf2HQflWWZF0bAq/WT8lOFATmbYvvT1oEOp0SbBdi7
EOMHu6KvmzVJFDu9oitNCbEXvspv67qiAYUH15iOXCTXwdmghfQZx21qfuQ2vozd
PbcFYSrPAvs8QWyqNzDI5FpAyS9yoPqaD1dSMzveDjXGdyw0+yFkhJPFVBF31+aA
mm10UPBeYNCdL051PdcSdAEZ8BeIusvPjzY8AKxRqZREDQQgAS5RLPWJse7wQ137
8WnlwtXG34iaCjZevkfd4UyIf60gdrwNfld7BLqt2YyWSyHt3yfkxmvdqwPaCqEF
d0Bd5YjpERLoMSUYMh4B0jCj57IhOhuGcedbjggXArKzi0cppADAGzVDAnqTC73X
1+vNRaCZm5SiQSiNKBImqqrAm866nmhMMkimXEYBFmOMysnwYZjgX21xuduhBdg8
p26uKXcqjO0ttgsp51iZ/gO36wRk2FkMQm5RFm8fclUMUPhaFqu7m/mU5N3ACQsr
U+KoO7IbnPHQNjF4AtD0UzhkcOICGyMIBi5Vm1U6QcFVlbyOEBuBd2+I3/IsiRW4
T6beh3KVKFHOmsQUJ9nVFVjZ3Fcu+PEHeqyeRP9BgsG/ZMID6AQP3G3XHPvxICxZ
PPAYtQIREuxLuInxuK/HHJ4BMiUypt+sYnr162Xu/wtNOJuNmlB/1nGOgY8ZZks7
LgNa9gDpbKhhzXn8Lyt/XNCuZOdUIJ1cqcelqnRSIUl96dv4jbtEi+Omb+P93TOG
wEPQCDObsBBnoEaj5gCRU7GUv7Unr5lHMavANxficBzfVfwqcDBOxKVnf4DiFKHO
VYVW3IcQnzk5lR8+XDveq9dWXyCDsdJHtVz0sDUblD8HKDG1uNOOGQN5zZlNO0i/
JDTptdb4SM1YKF5SP6aECL96DnZUJLrrIxk0+vyPBWLspEPw+m+g6GD93wRAcPpE
l7/GIaw27vN1EwaMg5dpZMbnmQYSZ2Ata+34gTVd+McdmnsG3zWqfT31cls00ayw
M/Qa2d4SDlMRA/y4F5sw1N+vilSUEcrk1HxOq4qDF88AEwGvLWy7U1hjIbGD+A07
7vAMY1aZLf8RXVkmxIC67EEJm9J1MNAbSpdamS0iac+0/vZrWC731X6G5LIGgBTQ
FwBCx4fx7r9v51luV70spfSHvcJa2ZHKgu6lYs7aIXcwNmuRXkYgYF2CKKNohwA1
K2/H091cqOedpfxgmZWQgNAifHeTKbYVMCzUhqkbcSuE56CkdHCgtnrOU9BkWHU/
HXFjj5BzeGW4D+cTp5vaNH3+W7sfVBR1exHjAGcFzdAF/H/V9ro+eTIwCjsQN/iU
iDaemdEjwy1zd0w2vmmWVk7IH4ZRJBlQVfFZ1QvWPlztvS/Oo0dhb+F62AYiHeAr
ChZAxEXcw4erZu6tUesXdGcKwEGiCBHev2pfcyttvjblNk4zs1UXQ94Jq0mnqeMi
NbljodS187iNI4p+/6rZqL4LD/rnOuKdVnt2UpBXVBUfFDY452tgwggvhmxrr72i
Q7AhMq67aEvN6ElkSUpi3PnvCSLTjmPJsoum+sImXkRUOBqfMmiXS8QKSs3TtjGR
dAirtS+M2rVI6hJ3SLcemPdn6IpK3vT+aey6zdBNDuQ9fWgBQiS+PaeQHOXUK2xl
LnRpMhpc2qgFhGbBRWjZt463gCx2ASK+L8d7gUZKAe8s8cav/BLSQXQBfsyEQ4vN
nhKoweVZ3ZHIFgLAKxkLcj5CeXj72q/30lmJwdq/fKNVxEyJwbJCtPdnabfX+JIK
sA0Da2dCWeTtGaEM9fbUZt71Uu3UW6cw9519wXYhyq1gDIa7zZxC/qzlJ2zrOLFS
taeqWwxERj9qXflVQN/g6QxDV5i1fXxzdHItZOE/ipkRDcmE12uQ9oSz48AgNnp7
c9LFZox+VnZn0mhhpwKUGpYzikdPKbQsXy02yxUsxu+OV5fVwb54wI1V8rF8kdso
dHMNTAeHrC2LwL7AZBrkUa2L5PkLCaeeCIqw81RSeCgp8PUou4Hq2SVOwKCwaMmp
DB/V3nGU3g19Es5jSOwpI7Mx2cLEQLQMF+HuTCNJrY7nJZBCwjTN86WJidHct+FP
DvwoajICAOgS2C1tLG1bOveXdosCUm3gXgdkDk2i9K8UkCz5rDIGFbKJpGuxD8M5
D1bqKj6mug+dC3onCK7bCWEhMkcmw1SGVsvUg3thT0w703h4RVKPC5s8rwlfrZl4
HG0I+MtSQXuQEvedUWBeX9il25EYraKjkXZOwQU5YtW3xEZSOLCXVa5n9e69ltfc
w/H7b7bgcOJtG8OCkRkJ0qKu6yMd7dgSaEnjvQNuDOiKgEPuSqrT1mhgV7m0xXM8
sEMOQUqH4EuoalrQ6LekFscYaq3magaAMxO+gi7xpfDf92fKclu55I5GkVhEImv3
ryu+DkmKd/+BP8bFpCAMMSTc6nKatrRsppOqoTcqeWRMwnZo8xZ/CtIhkcymJgAf
o71062D44OoMloVFCJND3n+Mqi/D/A8JyIQzz5b55kNGyNaxl51ncFNZ7cOF8pV4
uZxsE5eyAkyOVdKsUKazEPpfrbkYvXCJG7VOjWT++Hplzose4/MyNbe1BsHxBjKB
86e694uaZxTCiMwKAXJDRDW96Pul1CMPuazFW9uYaHdIx37yLbRLIQJkhAl6PuTd
ArvNsKrTz7U7TOog7NlhT5pEc3eBCwj00H0S0p403uoISWbBVz3Fd/sE5y70sIG6
a10k7UMfztyq+Gem+aVI5+NmWbPxGBPNbbQzqBT7xgh37OGOv3ALh1FsNTdJ7/zi
Y6gacymZa7OowVIFJyBKI4sey0mKLgVCYZeqhb6rQduXzs1v5mbudQfLquOLHHC1
FQW7N1Hdj+IAaleLQwUpNARp0wmtqaekjropqZsq2LlaL7IQj0+GTXtDI9wKfGB+
FivBvDDbQrM/gxqzQjP3yjB207vy8rwGJVTx2WqhX6PDsOcWeOPYzTYGmZ4HB94G
9GFMkT80p+EVl7Dkt8lIRYP+PYymERSBKCwsgu0+jb8xAUAydU7RTF6sWhS1SI9d
S3vdOEL16//zvLUp3cbriFxqU9hYUF8PCvE6HWB6CFAC1fE/+tuzYTS3Wu//HM7C
Iu9NtNpXz6ekeewAWIPKIHdqbvgpljduVsp+ohcJiA+snRA0neHCOAB9N8O706O8
gXqH+Q03paUG86TfZtA73Q+tRr6F3S9E0WNKRjC20snmer1wwhiFXf93dgeZ6Kbx
RheR00Z49NLIfG0TPw+pXoRvvowzRn3gaUB6M7r9t+9DSrlEgcGSDViAp7jy4lxC
LBJr6eCL8ALkpZ4X1qLzRLvG+Lv6RB/8kHzkZk4HESAlkx0DhWrm5b4QWtCj+hXk
Roq5Lf2HqSTLB9X5EItclgUYcpq3hbLTecXOnvsOEfhKntKycbnDyJ7f4EKkQW6v
99njZx0cQbR6JuzxP1neTadHI7OBTV0vD2niZJ+UUlwWmQCC3yCMJTF4DI14C4q3
YUtHIYSvHswNZIYsTOeSjNVidGif0pKLiRmBXB5ewlcE4/aeDNNmxAaFpyJGspjW
ys7Asai28EKPG1neFhuvf/snAsjG59ql07ADeCfnRBVcSk57fJeXjGjkZDUcglf9
GmJwzNyebuExTQllZDPF0eGf0Kt5j9PZhqKRfnkz1skwG7e/1pvEBoRcTDO3xoPi
gPr4oUvP8dV0J9hqq7XH8xbuJzQPfyy0EQfNZEeN6NbUyUB+9ZorEaF1v/sGWzx1
+NdM5rxqEoWaNGyID4qRQDw6oaV7zKJm/tstifKrD1OHo/6Mzs82n2kRhi+EUY2c
Z4ef0EQwB4sjEiHzPgBQ2832eNhQ5Qi1qHLvJbdWI5ljM/x+NrQHheecIGNZs5bd
YChmtiefdVBgp/2yOf6QK5FU+kizoPsPwaVsn+DpfJVFLnXClIS3a0D2lWYCUa84
Ra6d1IYCsdtaS3tTLDQ09xQpR5U8a3pyMI5I04Nc0DF3gKNz6X7K1ECY5jLe5QcV
NIZg+EyArqhusVymNea/sH+0LusQBVeAM3jT+8ZL3WoqpEeka0X2uIvKGMNDG5Zw
9ZZaYsQLviE0f+5jiaEytySEolidei25DLmyU1E4ipg7x1iYNcQi4CIaAazS1ly+
Bvhysq7ZPwXzGyqy/rhL5ewSNyNJZrGL3xqN6qX5D7s2Dfh3LcUh/OewzaM7XBnf
e/SCtsFk8TIqRVJQTA0Q6C3ahgofMTXgKzBirewaEHrnTyNNg+EPZ20xhmBEaBpV
XsFuFBcJ9ZxqznDh3KvfdGbNohDSj1ZNHtjnppqdXevDGL8wPXZp04HjcCsZvI+P
kDSP0Q68S2yCDIA08Ek5L4Zlv3YwIxSOYI7CXyqTDoBwx5e0jomy1SQs2n7U7q1L
IJyJj7SxEUN12Q42b1s3WeoVNJize/G5O5+fn3+pKjlq1eHnqbL+zvk6syHC2yjf
jy79lI6q9XCHQtnXPmCO3vgrAYZc1ek5a0QgaeYyu+2MhwHIKOFPGCDTIgn4Hxnw
dQMxUYTc2hodCmw6OYHyK++c2cBYzUMEXJiQ7hSDacH0aeuxMcVg5vdolrHybTiy
XfmynmQ06rnS3BpaayYowO9SgxYFdBgTm6B3NF+Er0k4hes3jWBDk7RX/Q2cgKOu
n4nHjQXMHdY0AQw3wcxCAShX7bGJqI8fv0/2PgvZGRxrFXbd8Uh3PNO3aEfTaJjY
gstBbFgtUYMDVXp5/N3xu0jTgGf0gF96BDbfPAaglSGr+ZBEWxGz/A4/WbZemYFG
/WTBB2HnTABcSlbcazShiEhWBjbsfZcBQ92zlLZRs4tny/ERgKnCA6/ZsbZqY3ut
Q4xHpcCS1BQS+yg+5e52TH6sW18dO+ArwB4UhhVuJlc1Lzw/iukJ0Ab/8rlEOOOV
4h7gpvqcq3YME8MDFc9765SYBFUpxVHOQG5jsRHm3WauDjGZLXbKCz9bFo/9a9PB
1Fvw4CxZua28wAGQh/tT6HzZa4AxdJMb0GUHsig0Wzg2yOp8uMLmC9mkUFXLpAEx
c6sODgaTppW/A1JJw0PwkfccEQCO28DZuYTV2aBtpZ4kckDG2y8m10bqk2WDgHcw
mQFIM/mNbZU4FJ7JRyiu8m548ql1Ypx1JdgofaOcE5ww2m5IpVHxvBju+DOuVi9O
+P0twD3YvW6aOxsOPp15CTOosMmdnrMlP46XRC92gDS/iIr+oKi6XKn8aD1uOY3H
Ze0lLmQrhGFVcrMxy7obwgWDguX3j/f2y1f/JmEB9pLxFAMMDuNRdu2Hidl3pqIS
xcUUveLgcEsGqeWGrmWqGxoH7PDYqM6cou2MV9QzQkGkmjq+9Np7Lvbt1EYtHecn
S8/UfNngs3SlrzvUIoWLQ5ikZDiWYwFU10hQnr2+TkFXCPaE2ZU1wc3HfW4cxNv+
3cmA0EC3F7jacSoDOV7hbrZ7nHMCfLp7mMH7Wm6fjcopXZ7MlQ6VWPikN6BYzgxL
qYSLm4XoMpBM7ZeIjCjvgK8gMg6IpVbJQKq8YuCv50JIYUZMP4Ee3vKQgkDC8nTL
NT6EsPDTtWOteQ6zCxsrMootJOmB8OKJpWtHqVwnQbmnA5++mCJnPnwQU5hDbEqz
jxZ1IDIiLaPlXpg1cTsWLtKBeOtnaHbd6id2wvEZrNRgW0Wzoa7Vpu3o/oM8J+an
im8bpRXYnQUrn+BLNqunPMVM0jpdscBEpwFlJMDsdd88ILhrYWxQ8Th2WxiImDPA
i8CaWWuqhdLDThyhY+diom+p6F6xqn1ngHsOEC6IwSKZFVKMSkgGT+qOEXTkDjfL
DBjpj/dCJ+5C/6plSYgPUeQ9lkpjQC4eZUDj0jLJ+72tueliJUl3590FBMoaQ514
6uql1SxxCdk3qtyhmoyzJOPpjDwAbqG3BttVDl2+7e2efB+KvCfxPbQBqtxYcAK9
8ZwKlGKoDwaLAlCWOuLiOu8aeIv4QnKAoxKmcvQwj8nHKh8WFGCSbgWOdGJwz8O+
jbGSNc0xcM7MRUUG9CoOCmM1Of+L6n40DN60+UHpcXZqJPwjKaCUCj1tdETaMstG
SClPa7Eko0X5FR+28e2NT2ktFxNAiEc30YvPc5H3047OuGBUFWwovj3a0Ny9u2lR
xd14C9wPNhPmeHZDN0Ffoevu9WJxPR6NL1DOCZzKQ4fJeUmZYYZFd3mX4nblYuqk
f1+Ep4lBcoT1eUkvP/H9DOLjwC25PMtCXrS3TJ8W3vNJEVgF/oebb/wtLMmyR+vG
qjh3vqt7dn92HzWstFBrAXPiNEd+30jS5CQX0vruVluqi1vPztSaf4wr39ySC0Ss
u2VTtRmKitPaN6HXFHhz4c5M3l+MTjVCqlMFTUAyGBCiCKQWvxczjghM46wpR6y1
eSwc+yiL3NptKs9yYyuNKOsIq260RApGSBjU5qRbyLd3Lh9ak3Hlw30JGwc+zLMU
oRAtJVJcMpgV4k7StC/V6cFPppFjhQ1QmEH2G3nFmHQgcFN0dRRJ31llgw+pIkRY
E1U4cLKrwbTMEL2X3s7kXId77kkMJBMRMnVBCtgEP3q98cC/3G9mWhoCzWrEwqps
E3RFcr1+IBkYMuoWH5V3tcMrXxHHXpCAPVYjvGYo9eK0M2DkVnt2E6+q5/V3/XOs
Puaf8OWbT+BElFtf9M45jRB+5X4PijjGOdutsAxUfBiVSBXNVaL5bOghP4WtHLzV
IwQO0ptbg4gDIEXdvxOBqXoAPJ5ZOpzcO7UFaLg4yvsiQKgfd7S7YRlOLpsBkPVJ
MbpVnSJeTvgxM6hWPXIA7Ecq1JjhTVzFmsSR07Dl3EQ+9AmLROJrnn8aIMtTGMUX
qVLozC0z8Gt4qet0foXj4lHkQPU+LjSGFLOtvab64y/Yo3cd17KPrE05yrlEJDqH
mHfgKaPqm6k0Aj+GWqDH0eHqqj2ZHTQq+KRn18b3sx1WhGGE0zZsgeZ0eqyRvsJu
z2gfj74ry2TymmBvHF90b3hxycZ93/PGnR3bWQ2TNkr1y8WpigId+fMYbOyg7gm5
Rz33bpLt22WDasNLwDqlAcmi6jGnnFb1XoZbjPLXYTqNiK4M6lvn6BQgbW7gmuNZ
bJe1cC0EeTMAW57oijsZDu4Hy9MmfB4ma2SKi7hiKiaEcFh9taAMcj9wujY+k+IC
1SS6KwOJ4PFrca++NmtoUDp0x4x9YniNUlPIlWddY8bgEG5yAtM8WpcpAXcUFdCU
YnDEZvo6ns4kvsd33HQaX2o6iTUPZp5SG0R3phj5TNbaQXu1XSaW1wlFp6nbghPq
+7AnqhnI9Wnt9FKwliGeo4J//PcW+IgAyrxMaHqQ1nUY1VAPDOW1x4UCDMEIO3xw
LSvxUbkSeI46gW6NvjHHF/gfuZ8umAHPNLHFqSh3TOEVfboGykoUQy4Jc/vkk/Ny
zjSPTIqqQ9tHZ4Gh4wwZU+l2897DuCboQOcIBo9vD6nQ7le+fTpXgvRp7Zi246IA
ZbDtc7hVRa6v2T9qWZkvTUyKB2pggkOZ+mXthhUDSJ5zJ/XFvE1MRVgCxDIQWdj7
L6mL70vQwsbZI1CU3lhvR2COfoRpMae30p9EqPDNHUpD40NL0yOlXIiy/3Hszo2s
h7maKvK3t79314PQvg9gJukooVX+tsBH+yhFW59o/DIeZ72u/wsZUA29teEY+N8g
z9XpKLyzF6vQ+K914NcySQnmGksar5r/gyVYRDe6mltHjxlxuS+xfZzmC2i9LOhk
tzLJy71zpitzHK0xgmifGcoNjH2LvkbneayAs0IMMMwJnC/4z04MkTz6rslOGhW3
FRwQ9KLVdnbue6ooPBBehTBRjYpIX8GOrv11lEEcEItr/XBWuQVu80HhtqpNooNK
HOW7VEfyiSfVvvm+RPj2mpFj8LYEKDajzrdr0iX7+QAnZMhi8AvnxPUf4K8E2CE5
vVXjLK7Buy5Sfra3UOWmFiQ/YJgIf8yA5zqQ8nagjqcuQqfZycwUaKLzPlZ2Ujhx
9yJrk4ArbSu1Xl9mqInoy83ojXu03C2deYV3mFx2tTMG53nVtKKNzMa3DgDctxGb
1y6uFCq0u62vIL22e7hmsrwdP4yfv48Uom2k9WXcXJGMoQUorORkEjbaTVPpdYBd
IYOmaxk5w8CcQDsY9Ma4++VeJeNmYKUM45h12Au6Xa7KI+R8hA7gnZpiUVuaXpDj
ggxb4Y/WNpgUaPXn86CodZWXWZrWq+UEHjETFfJ3pLdKuN/d4q4E9EB51qVooAVI
fFqLyxLHMFKf7FcHPwBRFCRoM/GJelrbXQpAVxaZHOZ/hLWv6jy1O1A/gv70BQBw
0JjPBtwQB3d6nxOOjlLaSBJZzokchzA923Tw1WVLx17XZiZ6nbIanBA2Nco1yGfu
S7sYVjW3nZ/STEe2Qd3G6E5axid3UeqZccKosfVw5g8XwjcORyrXPzX9lGwDR6gV
ql6Ln0RSqrgBlUcfeOar8NEJLccVDBmjU2ansWg50tT4BJ46fneQKMePMXltkeyx
NghlvLyArZDe+WdqM7BqnudfOjyFCpsks0UTklAc3vkTZHPR0ypihD4HIEvl1tck
PzrKBpokDL3uxQjjifRuHpyJLQZP0lMyWD6iPSLS5aGAleSjBTuB5jj8V01wWtAg
ILmnymmmAbBEYw1XzSX9XH1qz+cecgyeH2JZodr4rygNm88Y+EpIIsD5uX//jkO4
oEWF35KB19SgzIRxJaeQtXqL/qDpUG0vsBF2sM4k4qEViZdPAd8VAzv8z+g3J9UD
R/JGbNDqwOE+Pz6UbAmUQFK0jD33aBVdvkkJT03FgbY2jjkOLp5Z3djCHooRRmBZ
12LWY1Q/ClwcdE8x3BeXNVYRe6HhE3YvSDERYdgN7jwfRX0X+WNlHXoJXYyep9t0
Zh6JAEXqNhlisF3V0Vlz4zU4H13th32/GUdN4muEILKbCW+L/mLD67FHwWP281JK
JKEQ31cZgr/7jyLYLv5bYPj/Uw+lkQWgMx1m7+FimZvqiu1ycnZQMlsLbvl0WpaY
KVkzx5Ox6chhLJF/HRIn3AloAbAHFmS3HaihErudbjyESH1vF760m9Qc/KxJKZEV
Zgb7FLDUI6ViUagrAjVnJCENdMiUd4v5zm5kIfh1ADV3Vo8WAVO3LEr6XvfxCPYw
ZsWApKPz5vBfy8LDdU8Apx2klQmxuvcYNHZVq4TgPlfAjMFBpSHP1zITgPtxZ9N+
yhYGal1JuT1oGwOHFiZXsOJBIYD7DlupU8VjTC64QgYJvaSn4u2mx1K1W+Rq/KsT
9C5GL+uMTWDu70RKJkq3olo7VfX37AmIHEzDA083rF0V6BD0KCzyewCNQz/HDPI9
pnKg/tUaMacFGTVcum6YlH+ijr3vUBuK/4li7ABMIrl8+FVGPVfatrQG0ER0tiN/
UoWlMmx1JzfSV6uHrsIL57JbDzcfAA0wHd23lKcui5Zg5W/rHVBJD/g2qE5EIp1B
gaq5gWks+HgbmA+qXfozY9IXzy+SU7nqyfpJaYt5epFqukAsDZWd1aEfA86Gyk11
ruHmZ99WBzvDVgvWsN12r+RBbhX2WW3pfyAliqzQrB8hUT8hELiTJ4/AZu+DfIeD
tKhMFF2dTZkhzPaUkzHCShEgXiQ1JvCktTybI2t+CjTqtZs4S0qHBQXAzq1+LZgs
ZAYy3BCJeKXarXs1I3dolSlSJqusJrg7x6gzRPILAntRRrSpuv4XnBdK0vM3dHga
hS1grZUkoHMbBjtw3oWiwf4J0eBYaQ76C2BqudoBAFMXSe830FK9SRhufK2pg4mD
7NjJPPSy0NeNgWZM0VtYnqyR2kkjrfLHtOK29pjBc8MrSBkjILeHghYFOCj+BBft
p9UoyK1Cu9jwoP7oO2o2NYPuc9XGGeZ1JmE9eSAgXfxXf3xi/fD7QuAwVDKHbFZt
YmITZUyshsuO56Q9S5IrM4EXE9o/uewhlEptey1nokVMdvg2NnLUTIdUUoBhgV9l
ya4KZ61lS8d0N47OrDW59kAWmdDuvBkj5vJwbQ20dwQEnfPMEHBLkmz9HIzEMqI0
d54ORAKpMqi3fP3Imx34PukuLdYfBJzVUJJwoZ9/Kp8A1WaDMSpKuFqhQz2fFiNp
XdfsuDGKOC/9vulY8q3e8DaJQpGlFzO9l8/iXdet2JhU7NodDun38B0+/S0ZfBbm
e436CS7HO8rfDrmInE5xbe8utJ7ncegWeJlkZXOkt+JctJ6IN/4wXyjALzcZIuaS
05IAdN0KluPAIcMbXOAnc9dWTaQqbsJARdxumT24erEsNsjkaeY5NdFsDoBUYuF2
RK1eG2Q7M2TneGR9B2pcrPDTM/aZHZ30XXp12HGEMB8fIT3om2jKXwTmpn1VyR9l
ZrSZOSkGb84oyuGKjJBWJqmiVOkYbh+MASal/5wTPF4m3whjaWrb4CcicAI7uVPh
eSzlfwQw8j7x0JfuukQ05vt4CbxZ3Bx1nRfAAhu01jXQTd2woJKDDea4GVnq6oRA
XMBm7pwdlnMOtYAJTvDW/LVNcjj12PKUTRr2J4Duc73DkB9V4jXg8DR3/hJWMUMJ
YivH5/nc9d5xLSXNQ6+7fV1yyY7dMI+1xOweirAseL00GHjP9tvxEpVb8GnId9EJ
BMswj86lnpQTG8vTVS15jY5T85VJsCtl/qiAA3yciPRodS4qi8WA/sW9STzl/WcY
L5zE8qUQr4uj8tv8h6NI/p4/8Zq8rFCIqNQXXF4t3SSe3ejbVd4F7lu5wxnenJ0e
/BSN+GbrTmbETgqKv1WmNoTH+DI7tJIn+u/gztdDVvLb1nd2XcuCwq1JWnp9EsCG
LJNLhKdFJBDloxRfqQuZQAsKkt9qCg5/uNUFqPEIMeruiYyrw8svBXlHlM0wFkxw
c7/sK2U+bXV7una95NyhfXrQEL4dc+SOpbSZFpDdM4BH+IhvNybF7XA6MxWwkQOH
EexPO3EHKx46cSxyRFJYHHng+nf20oDDeBPqEKDsE+Pu9N6fTpfRGap0RpFE54J6
Vr6meGPN8MkCBYyrG4tyU3FYlJrcIElfldl/BMeVNfAbJ9s5u2ozlf0Q5b/MXwen
8NbWISVy77EhQpO1+CEHDeIW378f0qFH9EkY3Ime5HSvA+dGjb/S4jFTnUooqF01
wE48qehQIxQ5jPu4AyPxkGDk8lg7zklm+3dHZnh1lR5tnWcSjEwGPqo0IyVAmSDK
QBVNZ+n904Sq0Z8D/FOUHPGP8SoiJqoUBLGp6VYsWyQXnxvuu1qLCU/FJ33FKLfo
Z+NiymEjg2LMl/pd2DNPcNDdMyRASYbXyTMYLobIAeG8XgO1Ip3a1xff98HDPXtf
l5lJyjRo059HxH1Emc5O2RzxlG7gtJLMq0by2EUlDYSfMVJAhBeDJQYWQkd1s7r8
Z00tR2bAewm4OgLydUAQvWzkrVSk7NTibXXeNaGvkYbVe7dySKT4Z4UWtcGRrl+W
IpF1wZ2qKtl1uKJCXj+v598K16bWzpJFHjWSGibyFa/YdGBRD82pu7gjFjglsrd/
+4cIdac72GFhNbIGyawOnJ79elkp+uMtmagjyeDShXubdWdoGD/Jixauwm9tAmuM
h3iEkq6N4FQKWE4qXgqAIkY5n6OGrHaAPGh/n/db4J0HiG8R3OE+6jdKGrxSUiLH
/0ULWAbY0+I9Yk/Iu3zVruS2c8NOeB+vYUHxFWBxnMZZXuDev7EOeQ3GgSJ7JUpb
mNmLgLkG3drGFrrHb2DmBaICkGZ7zrzCbpLiy1M7d9q2BpjtQu1r5k1c+yxvAU3+
L+ksqzrQuew1oKWDRVEa9cMl0uebbuEcBXVe/xhNNNytvBAwOdrnBWhMYD8N+STF
qFI4LNfdPTAxOj8ORzeWQtlRRtHz6uer1ntGwyrJSAodIb1P9Ofm6t/67Aj6SEtn
Ssc0viMCV8yeNpRFJ/1nVb6P0dHqWUuD2V+aDnMyjyjtr3b4TYQnenT5qpj3D0p2
KmnofYWx/YNNexruLO5pjXN2wLgSF7ykYbA395gAfPxmfh6zKEnkxRXbUE1PXtdG
9XSaJ5Tfu8GHcZScrPaDn9uyjdQhD9RCO+dnE1Aue7EICBXxO8pbmL+xBAEIphyn
3t5ao0DaeJiAKd+OLsYvGIzaQZUjlcvClFxhlteLgFe59ou9REJB2ymKU6czg1cm
L2Izb5bZT+bsZUn5edLMgUr/VDINBAHw0i5Fs/DGb1CqnGqEB3DnwF/mFQEcyCRd
j6UfOyv9KPlDDixa+arDDtkT5JeV4k2T57S2IAI5g44IPHfZK/B79q7jbb1glujC
NQZ2tqMpB7/+t7GqJxsTfQEmJJqT8eZaCsrf7VQmGOAbhGz3G6fCpd95tZyb7/+D
lK5NSXz69Rki31COMCldwDSMAnLt6CQ2JEDnsTlwg3xvF73ikvGkKx4gxyTgTDGb
7bMIrHETHbIcej2vEG13hjYf9xBBwsAYTzjZpZD9GC4DN2mtzz9P99ONRW12Gm85
SgelDM6QenvuoMLipqcydnn4ybroTs2DIQrv94iv35tOZn8H4LWMpau2N0QKKgCQ
oOQoxk/YFzNiRtXlFzPjIUgsdyWuSKEIKtVGA3yZ4SIqJj6+UtIx5KAeC2Aa1bPp
7m12KlnofSLBmAFMIDLagxOG7Wd6oZyBkc+XYr4G4NkuS162uGippDxi3P/V0pWH
tmP6Aq977aFfEtBpQlEyUqFsafPj9vsUFidmpdj1YJCYOfqgl7guNth8tX0iKm61
u5ppDDcuZvth5w8ZLgSKJUmEh4Ri+oAGbRs5+oeo4o9d3pRV5qwnN24FORntLh11
8pwT6Nm4z3hMhLuCK99cs4+yg5JIVBYD/7hyI9+MYbBk/QTTaHem6Qg6KOSQLSuj
oVPHUKAPjeq3cPVU0/BSp3K1zrLbX4vHpvPXSDNf9RssNf7mcx01iCmMztpAQwjU
jJarj5P9q4SX+EStlSd15SCHRD71OvSdKbO4vvFtPrMV5dXVNrfjoeIgymPzFq2B
P8RWE/4i9ub1WGgr+RFInxSa18KD895evNKsrCYce31YuWDdz+sxAhb7HycmJYS9
lTrNgo2ODImJZo6hq2hIbpnH7YrgxIlXAMOvEu/iGTsRd9uhKskLROcm/RUMgVV9
Si17MZSVlTQBCQd0r0fPicXsxR5ehblXvgizyX9/E0qL6D+dDF16bx53xViglD7g
bOMhY7PsTxvikV5tBBCccfkEOqV+KNKv8pL5rlHIbA4+XSQn7HjwANwKhjKHA8Nu
vauVXY39AXNASQcUPoEUR5y58cOqM5YPptJrGGh5iZbOYEs5sjOF6ERJNHSqnCOH
cCQv9z9RqETxGvkV5nWZf6BHeyselSixwyTobsxlHoZNpsfnl2rJhpCc3P5saLgb
fp3qSjawZSBPj40lfXZEONdPPf13Bj4K20bOfQwIHEaBm2osuCMq8V2Iunz/6Vmk
mlFXUS0ctRPDZwi4j5DBAqeZ8RriHSN9UYW0NhSR37ZzZRPygME6DiXsm+wYz5ca
m5/gXrn1KSJehN3tW88+lq2QeY9q85YVtZ+Tc8j3X9vWypukGgO5bN8wrDZSA5DJ
IoZOlxvSu/aVzZH44XYTUGYGj5kK3ZwFEr+IRzfgXldgBpF3D9O+La3/QqKewua3
7t24bL1KOb3pv8sfwnZAQa8ewxZUOS9tAXUn8VgSMs+g4RP7uf1aCvk3J2I4H82Q
Oji4iF2Zu5uhQ9tL4AkbZAWnm2ef6MgtyiLv+v0r0e9e9iMNaDlX9wsqhmjkkhZZ
Bn3pQcpWb8zkH7rsyPOxpLp0wCTdirWAt3PsoqnfGCAhtDJIREALlJ8dHz2EsgNm
NPeP+PoCNPzECm0RsWNn2akgcFdh7GoM7YePtALAmiv0p+Z2bHfilRLsG2r4Zv4b
szjBZljEB+L7qTQYxryrUciXGzYKH9H/822hgiwdvxCAmCYuQW7xmmlGVm2sWAjj
HJNg01tud57NxF5h25/i4huFQQTMrYf+X69/huYnxoQIptn7KvtIN6GwH3qqNnQe
tG+4KNM3F+lhiD3AuSXJDy9X+6oEsvnfOTL3ljbfLeAoIkBzjRz5zZ9KLZ7pnzAk
lOSg64dpmcSOviYTL424OmMESHQPWkucAEeONgctunHKyCfuBi2I8vjkm0lZUX05
fWovYtqzkHWz4KW3C25PKth/B9s4Zp83my0dH0AxrlU07uxM4vCdyPmkoZktYlN0
FyfTfZWMtKSF9mxi34CFmEuTRM26aG2L+EDrVM2J7BtKtlL0YcXJLiKDi4FYnp14
lrx+PeY39dZMBtCGVPENqxuPyCyJRAi/67Afc2CzYs5kznn3mLl8REDWZZtLMyAk
bGCGHAW7mNiE/q3ylXvHct7HvKwrGF4vCoFLunCXgY/mZLzlD+byrtnWYOl69Fxe
B3XWzPUxQNm8vMjPrF/8s2gfyDn/fm5eHvCYNf6G76kbsX0iNwUUGwU7aWW9m+X9
XpV9+3TX5PqwA9uflJ8sF7O6mtOvDMb9TSozOqcoYzdDG8tTG+7za3yKNm6B4dYU
57/pQ1//8m22AQWGw0a0DNTwz7sFiBmuMcnG1GvzPYTBvryY3QImJinEh7oVB3Qz
XdP+w3611A/+bj2+bnIaxCfqPtJ/GD6Y3jmEijfMKXOLgmaAfq5mIwj6czthM1/g
sIpeKp7COdtz+xPBAbrH+3IpMWj37LKWqLL0cBvIEpgqF7TMTVIeRe44dJ6ex+Kc
SzRturO02JBOKScGiUeKSah6Xw/wngR+OHerpDFSbl9TxotBZikXwcUk8PrwXezu
P+SPw+5h1vyPumS7KSO+wFTcbTtJYiLXKGTcBgqCKgCfO9RyxblymcnCAiA7vCgx
JhnNPngaTezgbVhBDTDGuqBnRgcMe5ypxHrzKqQqwdDenVo+35UMoTYb32WhMEfh
RLDLvgbbDM5vXRTGo6eacX99R/jzeWlTuSJnVa9PVXpCJnhy/KdeJHf7Z2vSX6ak
ndG9fETz94sM3sO5KQvCfy+lSggEgRGFfH07X9z6/AYgZr/A81u41+YW73LGIFoG
AxkiX9VpEqKvqMK1OBObF/+jruuCt189rqmErLNEpCdDDr23Ga980lXyzKx5DUcb
J/0CspKLlyhxvKFSnasHfVLsi3wybmn+83wVjGQ0uDoGHSRruz7bq0ChsVFV5PRO
C2jDBVDCgrfWiG1lAm4VCQrEmrKRNuW1SaqttiX0uZMRpJB+5EuQgLbsBI+yhZ/d
PC73M0RY74JYM0FcrN8k1n44UvYhCrLHJwYDxofx5TtLgoeT+srwNgLR2RHtVcaC
mhtYdY6NKuCpkwe4GCJp/U7BSGjpJm+W2aZuMAHoxrURAjTRqHHqh8GO7B76MfQ5
W9GAFjkIkgkJEBcmpkI6v66WEZnIEWRSz4ljxm9qSPn439bCUC7+isDSslPsoVfA
FQ2r3gDQGnLQYp+EPAR5/Yu/Gn+kZ2Y8mRQ2gEhmyU0gSMRZyafLiVmPRXalQrn4
XF16iy4cjvt+zbnarlFweJb/tLoxf0KJkh0xQJi/Js4rMdCu1tZrlbwmT7ft7TM2
Brm+sZyYC7LGtFU4/2fUGdpIGzJI4O406poq1Fk4WoH1mpOD4qRMFTRxNjzHFY68
mpkbZgpv8rux9d7Knf1F66+oVJ/Qe5L9qqJecaJLkc1XYwzfgicyi80I80uyc48x
oQDmTz3OGgwiiX4CQuvBRvJpUbB4Hnuj/v7ZYdKJn+FoGfr5s0Ka9E/FQkvOudE7
pauQYIdFh9Eol0rwyB/qF0azvGghSrCx0vzMEyPW8NmG485Ld6W0DLmwdfVWXCQJ
YA33pnNDPAgaGryk405ICsoDLKlDxeGWYw3jNIF8TDpF7k58jEcNOMOFC3MGB7Iw
UNACxGQnjetMoyk8+hCe49TqzMbI1EXUQ83Xpiq4SmyQML+9idAh1uUm7rETNsmO
T9H+k/iRAWYQEvQjXzNocAPJxxXPjB1g0bSZ2a5+4UAby+PlLgft7m53de0fIQqJ
/lrxzWP4uJcRdkDQFGTcHnu+YgHodglRtSUiuRzsJnwcyWSeifd7aEeypzTR+I30
Pv+xFcpme9Cb2ECZPGGUDKTXKwkccarJcKpkbH7BAxCtKbAopf0IAdQYotLHeMf7
MZc1GbFPFH/P0zPleXrdJk7MCHkv9z2ZLRgmkehyQoA5I6O3Bix3PB++eFWYFEoy
uM4QetUlT2QylJmkkIvpYSEyj/wd4Yn8/Kv9sggaPQVDKmuoDv5XGFc6zBQJWiLh
jtXI70YQ7naqXbohOPtYaBFZORiQGgDu1HMjpp+xL7F4bImx6NFirVR9UxGUTRUz
zCY9VgJaZeuQhOqxVWo6oC1tT8+OTW+c4S/ou5KWwVH6nVIyCZv0xOPKN4DscPwT
7dpmZz6+pMXIDBy4Pxzmf0Cpq7ewgR94BY31uaRsT3FPXsaNws9AUI/reAfh1CR1
15LAKRJxeNGAm5xmmYr99LO5hFWwpOdL8bCa/bVe8ZtQzFPsMUHfB4h2qnTHH6iJ
qOPpdm2XBn1pY9fxfuJ0weqlFtAQVY+ucm3Uy53yRgAwRwbC3A8AHbOEWP/eypLZ
6HLwPeUc/qrpMqJZf6Xs0JKMPEfrAsS5/l7cNbin333QjE24wMzuHzgCmivenVQ8
v4SAz/eOQSNXQHU1yHQgcb+p/CD8hMr0uiD6F4g0neQSzzaa7LkRRoJo9olppAIj
dEITHRzMO502JFeHaebHRSaiHLKlJz0VliqgiTh/UnGQrqYSAZkJ9b28/2XThy28
EdxFq/5Mvb0VhE8xvXgAKQNXIcNj7xHHtPNiNHbWi4CJm3zRy13dmwyjG4Ll99fe
7Ul6tqo2Q+l8/SEGn37ZxqkOXX8dXj9CdFu+T1WhMIYCYpNsY1bzlwb0KbOXHehi
ImTp+Kaq2X+Mu3HBfwZarnJiCBRilFZbNfkazMYt7CGZ+Z+4ejqHk0kptYTkDBNa
EPxmMP+YUNIqsDqN6dxIdg==
`pragma protect end_protected
