// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
AgYgjayJrSkZtKrYQ7nLwVeKIZokg/fYzMxAtW7yEZn7QCJnz1L8Tew5jgZvRkPePLjHVUXafTEt
KPgPqZt7AWGy86ZDG9ounOa/MyubyF7nmhBmr1Xr6YQULYxY0a5xgbjEM/tg8ikG41jlHt8NBluC
eeKzOYGhRzhnBHB6nzMtFD5X3WNSauP4uYJJmfGMpcatkm6eCB6H1MGM0beETBgJBLiNqQqneOvW
lGOeVZ7CRdA0Rzfhbu8ru5GggF9rF38TBn5ab7Xw0oOobUVpyBrudqjQPOH0fx3FmafpsmQmWYUP
NvlDo6CZQA69A+NW7L+rvbVP5mfEXLSMH1VSEQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7664)
c0PaEvf5G+aOR76NSuhhNJDpbmQBNVKQn2aKPjG9P/Xx7CyobPJYJ6S68DDRgb6MUGzvazCUaxcm
5s16BjB9QxW+ZNVIPKPUgQZPOzZB+sAfMBZbhIAWZFzH5kirLe2fwl1swv2ZuSZ7cXms4/haZVSK
fh8aRhJRmHTp66uN/R+PjS6jT6waxmqwS9rnSdP9byPZRznOGxc2IlCpWu9xkyN3rw8korV2YUGz
01XXsTycZ1YT/axsOAazSy+8yE1rO/8VcnDOhIvUOAoiOyMlbUu0U7I9SuUv0+flc8YZ4Tq+Y11R
C7jtmdqbBoSpPAgjdkCB9DoNjH4/Fa7IRE8XF8/DckdbXhnLG1yLarbiCf4omnUWISwZUwFkOROR
rHIm30QRTeuwyp32eda/2SO3aqHTVT/QD1RhLqJmjS9SxKf5Zllj3NMI+KlADGrTj1v9pdRs+ZXh
Z6QLafFGnhLknlHRMaBLLy2Hi9RB8MpR45pr//r3ztj6TaDXSF3kWcNyOMOfSXBMrn81Hyn3bZok
5HorIi7qeyC/19vNqCFt7DxNxsO0IyACa9wOaBOPeDP7BvaQu0ro6h6ZN/9RaDKQj/bw9/p1Vc7p
5CFEdkJX8T9zlv1a9emQwLsS3kqYAhXWIEcfJLj3kjYVsP7RsS/ZKWu9ILeSKhNnpJ3bmE7/Urbm
gAOmEuaN5RKkWXbT8mp4zGus9hJk7f53JqJ7PvIH4iGvl8RG9TOyT9Vo4wonUbao14rDzW8MtcIR
KHpKNc0nFovXEoyU1KOQE4dGXm7Z3TYfTXTKWQzQz1KpobDEqR8Gmj2eJnoMiSD6BA2vxDnje93i
6gQLFmzC0rexQPSXjujWgnyo4RSe9j87Yh+AMfELOlLfJdmlJaRskPub728GZ7Wsw4adlNeQhp/j
SY7M8dwHMlbgdRcWOD1GA+7HkNgYwmUJEtE0942umLNXENZsj/cGiude8PpCkgbHoi1xMb5JJZ3/
/mmlwqE9qVk+9lNoKpl0NCj8GQkkBxWuZs0BYFFe015mYCNapUhfJNn2ESY8R2/oAM/hEUPmrB3T
PpXzoH59G3JZK3EWCIfjm9zC5cWPp0SswxcO26Xv6I8uvd39yLv5SF5jW9m5EBUrIUTpdz1I61qO
+PJrWVVqEscYF8lMd2n3lV2G8mAGo5WOUfVj+IT2Vg/GCUPKlz3GXQLBqfsYPM6KxDwV5AsfRXsP
PW5zH2bwV3tBd6UpHnUq3l36AoqYar1ewJaS14U2Yb4wF/M0rteEERMGCSZgUUivrVd5NN4++cKC
T/W4ilsxet7+kjX/7vLVZ2E1dCX61VMHBd9Eu0Yqv4i0Z4/tK0HXqc8/3jTV+VzrZ5dedi2JhvKH
1SHcPh+AAzZPBCWfQgKFsdbj2jxZd7HbXE0T/BAZL5PuT1eTutzeZFTxu20KvE9wAhSWZJ7AkyV6
hxbagASJuLQpyZUD7filZ2o6t3OBbXvliEwxqqStDcnqokBPjrgpCVUSM2UkxWz9GV4+1NcPAtt7
atRirZQ2DZvcLHamm/ZGPITELYT/V4F3dzdHQThBEEJAcb1O+tX7kICxf6Slqi010GaKUmvzouFg
sJGKXWXmbYHvg2Xzb2/tdrezyNy2ckrUNfIJIOAEBQUgQ6DiYaJe81mZXMAMn/7Y3o+iC8iZooBG
dsTNlASjaYpVSASrjfIFGUX48CDHOGu+teCqmYm7xu5wAi0YTnPUnkkvQp9YajeX3OYHOD5KUqHA
8gWHUYG28Pp0ZZPYc7CwcsyAQ51eyhbg/dsayLuZmeUG9YupFEO6sCxzC0W0kXXomDHCCqfHml3q
MLA/L/5BVsACCH1xWT9S8zh+0Vtop/ywjrRpdBUKTI0b/FOtN0rU3tI7MpaD/yaouJdlPlZPXM7X
oM10sY+y8Cc5kzfidcDQ8b7T8b9sQ+XcJ2A17GLi9oQ3i0URo1O8ZKi9yJbN1aAbkB5vCXIP4Ya2
q24vceLz7luWceG4CLyeKZlsbKbTmm3+iDjPBMUvAEIDHT2X8FtZPbJi6JOBLj/PaECc9152zXtQ
wDa6tbZ35no2gJAy0zR1tRxqtI4tdu1ZUv0Np/5lwoRrR12PA9L7Yec6NnHM/m8UBmmkw23r9sBb
sBdXqffdX+i79bSz5bK9Z/M8qQFdCPhNPRqLWSs/MUMN0IPWz+CWIWqL8uRxhTAUiodmFM211f4W
wJ+HWYnfwaAs15hF9bgCHRXSf8L2V0oyc6qQHDLcMc++coCKV84AgnR0oRrGcfI0DzvvS8X8fO9/
q6+GQ70oGP541zKxfrIgtOy7fIlw1A12rYgow18Bbts3g19PuRMdH5V44RTCMe8aea28JTNm9iIo
V9GfWkq/SveJFG1CR72haapnxX+4w0e1xCIETcmmv3aKfZKJN8HqDQDg571bEz5XJkGSRodw4nI7
XA122p++FpMIxYVL2iOGGlFsvtZ0H9Uhg9/QQWlAOhcCCYnRwNOhTWixabqT33g80hHbMZLBxR6G
L3KlrfmrIqgBMsOUze2hd4e069vpPSQGgjdRMSgLmrVW5UAUQZ1BlcgSJyrTy4EEd5zL3bnKcPDz
HO1ui/5TJO51k4Hg/Q8Li84VFqdatDZIGta0Uxqt69BALDxlAedgEsIp+abXvD+3J8vj5tJi9qhG
dSlnwTcjdIOii4wqCZfVzLByOmaKC+X/n+yWg0lduLo7osieuRR/o2QE9WaXXia1Xbef/hrAK4ys
/1ev53rwFJsyDxlrWoRwEWk80I0h4dpfUfBRl9jcb7MmBSFThTbv1U64W3KBswMMk55/jHLRk0a5
VU9hOkxQcCn1urQvqnlcF/mAl7OBEozCrMWeVm9WNky9Db0RhAjuHhR10FHqAC2kZkdEw/9nCKgr
v3v6Bqo31FMJGoJmbc/ueEhVtl4wZ1UhxeLQfEQ60XEX+t7q8bHFs1Q/NnVezlpJdfAqSfnU7U9k
72ftVjmnOK+vYlmO/D3m9AQzPB3c3Zqc3I35joZ+5j+Ras2RmkxtwNEFxbX6m071DohF1Vln7zVF
/fClMy+nS4o0TpEX9ZnG689CcBGwsWPEmU/0vSlhOWlf8YYyzzOsVn1KKS1wD/9FNzxhzWmNO0F0
/TZYGiviiRoLrA4qFfEmP5CJ/GKCL9MqLu9Sx/v6GBfQ5iyJP1wwRRflAWYTzfToD3lIgNukZAxw
AiMxENt7ObTIHY6bAv3/OW3nBQDNGiubKsYKAMCxUioCEHXvEzNTSBwU5svR5PhjSydy6iwWeOlQ
W12J8zZ+3w/7xe99JaDQ9fszAgU8TS3DgL2b+88fZSSCKpX1L69oVJhHhfAJo+iHE17PrIiARph3
GoAHOFs9jpLaKa8a+DRtGQi89NRzkies3aPCjUovTcUmwT2u5RyPvSbx7Sqr3NYwpetbO5Log+ex
t3K6BqdCz/Ny+P3c2G83mERIei3mBr9LRKPYJcmL865YVBVJuUwFgTcfPuACSexIgEbJSoDkDAdC
LdvUF7lSLMFO0Qtm3ehYhf6NGcAi60I9CVZe7e8R7TXtg0SAAPpq/u3ulfQvn4EUQ7pdDMPl4AVN
qIhsXrT/+i58o+ntyHbCkapA+Fwo3N5s8V2T6GfNUhLb6zoZVkun+vvVLaARvVxsC0dZznpYUwzv
bTC8IvbgoMj6jv5dkfHHoNyiRJC9FixybfTw3M+/xvz7L9q/A7d1EWt5r9E930O0tgkzbRGMQttB
PUl7rFdgYIed1wZd3a2+g6Oedr+pJJT4BAPHkM/c2W+UMvobqacwT/GXw/HataHzOvpdwuxreHEM
GUQqjMIdex/96kqAcQxpadkO1TNTZ46q0mNlfYawvbYJu34yoQHsiNsZVInFd9/yScUkGLTzgUjk
xT0QaqiMSH17nQV3fXSrxabtDNCOtjmMmSh3Wn93UoFWbuDkuBzhgnHLjJyM02lUeKD/l3XLeKe5
zSXz2R4LHS8ESeljVL7XYW+qEjeGQqDS6ys5FAONWnjLL/oirX6rzLcg8f1Y7mr13f4unHJpPRz8
reNiHyketqi8wBU3AMZdhsumpcBBPF/Alrgac56BvmGidZ3KY1S5DcObqGMdUvtnR3N3aUPr7aaN
RxnscM7qRYGjEq8qUUvk8QIxB44Y1PT8D8OKbl/Ik+X/qLxJaUbhhFqJLWb4jkJZp6lyErae4Xzh
605IrhKpcBfDs8bv/zvsxuvoxJug4ueetX1qtY5B2xqWG1MwVd84Jmc6NJSiBqJNFfcdmHlItCoa
UoSzN9CjlGtv78BV/VWa5coxfHnccG+y/YUJPQrhTePcxZcRv9BF1zBTAiyfrFoz1J9xehBg30xr
tdOS6aE1sl2ZdM+KlwNCVr9vbfSkFfP+/imBclRWgfrOrchcC9TgHhgrJtZ1uFi3X00FUjpsauN+
a9kSe7Qpw0CeBwhBcSYA4m6CpVH6CM+x7nWXCrllj0dnvPn5rfKZDFwFDh5T/zxQxTB7ab/dq8d+
+b8pMhLFEY6rE6JOjKKJ17PVSv6SpfkU9Gybx95KSGgqA0o/f6xDKTp5rYRwFkL29rXgHQ8KCdD+
0S7jN17k/aobTuDI9F03OJO8/GP+7bdx9Y8yQBisMIE1qHPX+CJrfNduDKSoMe8eK3txEKIn4AvF
QyTHk/Do9mk76tCvDXwsi3lD6IyJirraZujzN6+myVRz6vZmcxfBvz/o/06MV0T68/JwxB34ReOX
MzBTF3qdubfjpF6GCAoep+gcV3dE+cdTnKQe2kvjzj6pjRI1uNAx9pt3rEp0ek8KXEkylbDo/IJw
J/3Zx/CiljzMt/mRa/K93I4mvGWxNxmHRqhJ4C22d1+zqtHmP9lLCvikyvQeAjBWO37tksYmFDDp
VXGJpqQ4S7NLRhIYxjElIE7F7U7r701w0DYwTWlzFLzqfDyi/Xav5L8fAoz+4PPkYaTCqNDuSkvU
JJQ5Hft30bRaRO+GRd6aeYyTOwLZBnWX9b6kniAP466XSE5It7UyB821cp4VX0g1EXQizXq3BlvW
6SVeiyF4Egs6nkbby7f5cla+mFOclxRfbl4ZGxZNhCSRm/WHBkXPU0YX0+ZoL0p/xGRQMihCTdGk
1WpB8sOJyXKetswMhLoKYNzr2uR39a4OnA0CaORtR9nrHkHX+LcCrgaryK6SbL9iKKVWVuLubUXZ
IZVPG+0FK+VcQATjwP0L+TzcC4nj/3+RSCu07C6goXCR9FUFXhTk8tC1UD96zIm35PVOOinGmzfZ
FXgqnK4o7GoC2TAZ5Jm2RaUWLpX9IZ5EKh/Bmr47ZyO0Szb6t4TaZjDDp7HPjQ/rMnYsdel7M2i+
7D9NVMk7wmOFBriIyU1edPdPOrdeKPDx8BwrRN9WY/tUxwAdKxRDDo+Bz6mfQBTbXfVakOCjCviC
iZKgV0e3xWq7vXbqydAIcUNFVbdX9IC0sMEjP8C/sqNibfvyvAImkJqxtcvhNmSwbhyysg+rV7L8
ASiIXJWJWSQ4Rem+HmDMRo/Low6z8DDTJhuyjPqCPzwvZ2hUu7vwPrn4yOb+U/aSpr5nMVL2Nmw4
YtzCHuklc6x9HA9WCqMVPPSk/cxmcnSr7DjeOUOIdF1EYnlta3tv2dL/NYKSGmUbUDkbJ+TldBVT
z17JRN5LijCkp9PaD2LgUfWYWGs/s4qmlUWcI2USYcpxo7f4kx5g3vf0fu8eJ1i+UQ2UlDQd/uvF
oTb+w/vjfBW5kLHdAuSFMSLFISYi+RJtOJET06aToRMM1E5gtBiWz924GtfBpTwTVxGHBavTDLaH
9hy17Gf9xhxwUiqYYL3qzVBXLSWQzpyvbWDo27OELAGzJCr/5sGd9k9qw5g9knbnToBTe5ne0G/H
zeZ3axnzNZnTTmCoKY6pRE2mUafSXykql/fdqkkgJuoJXuTs4UY7Jf725KgjHqqteKSSCRHMSJlj
yju1AMVlUqj5mNFv5H6s2FlHfMmXSVHA4Q6YU0Y1pO+alQdvEFUSB3XoWEU6C3TntDvDT+MJl5Ov
uqCsoa3NPpBZY3kaBfqG6FRgkGA9CwMiE6k4gsUmOdHBLan5cDASJcQsvRXQakF/lZMgnohRDT3D
gQYgwfpIk4lSgWQde8qTcSfIUtsPjIs+7nSnx86yxUjKqK83v+v4hQdOiBN0Hg79Jbzo7aXk+Xky
VEjRSL60MYFlxtKEskyeUUXdLeTsToW/KHuZCxyiz9RmQxdxg7vmY/2iaZtHg562JFNllIIIe5IE
r8lzORRNhb7TcKk7tddLB9r6saAnaHMoFy/teMrc0RkhmmpJnzTUfeOHTOPDSN4btEKmt8HEC5QB
hJTCWwavTgBqxHGJ0Qhf3tpAMuLpulOB/44R/5knxAQxHKyPFfYgFTbV3gKitorCTXFNPRURWDHL
b21R4VeBBfr7qC40RwgbgjNr5YsQezwQC+D9gO5ZJ//T9YVPaLTq1WV8XZ2mw3XaRi6x50sRO+sE
mk4aLnwLGsbwCdCrA9KINM2lppzKLxTEDMX9yq1Q0pjWqGD9LWXazB6TTtGE66ED8ok/rXpB5MS7
2BQc3J0pG/nZh1hGK2bu+uc8J3Iv4O4pu4shjoy1c2ng0q9eEWvcD/HljqeORUMycPqB5aQoxmDo
EYaVQCFNZsFJ5k22gpdr9qTqOol7jdJO1ZFrGQbT0WOq6JKxT5/+eg8cHPLqnycJH78AEVbFNRI/
8IE+iO4ghqGN++mhIHkVGbc43zxz1U/x3k8YYNiJUEfngU0ull+a4Wpu4G1uysHG2ajUljy0y1CW
HqSy3HuCcxiGkEwC55ItsjUD18N+mqP867lTt89B3AWSvoDqV34hmzPm+YwzxoMMcXdPW3pqu3ku
WFpjRVqSiKP3DXqwae4TMv0vqKgrlmvRfjhP1VYr6a6W0dvBOhJ5s7hlhmbMLHc8NXrkvkGuRGPa
sYiud8yx3SXxa1ROL4JcGM5x5Opezym/JdJEtCdBlJJ45fYJcKKr4wrT2VHKyMN9TSamqnsuwSzw
J0HqRrOsGcGqTx1bD4AIH1A9z2MCve2EooqSDW/Rp37z6w6pvsBzrvv3wQfgzTYutWlPztXqwZjT
P/Ev7Ycz+0iTQvgsHBm2sOkXTvI8t0uOgSJ2irvZFageClKSsaba3xIOl6mqdVn+JA8eHauz7zmK
uLmMWIENexGkni+WtjzVq1mjyQNWdI3HLyHfX0c0Rwy7/nK30K+W23U/2ftQO+aCbd+LuEAtbSha
i9BX38YPAnxQi+Lxk8K9Kk1X/UARHbnMOyh8fZmCE2tlQefu8Ax8TFhA0LUGNHXE2BVlEZ8xaQ7X
hEoZ8hlzll+DIwKW+ORKgJzhbhv23UZkG2p0lCgCCC8FEQAbyQ/vfLTZZu3XExC+ePaRIIG2YEeI
qwTKnj0dr2vgqNmYbuEuV1p2dLQSscqypQ+l7DU13C3gfJjD9wO5L9G4tVgFJx1UZLrz7MJq+LL5
8tBNIz0snHBgHrjqIUT2VnCdJhm1M9Lhvir/RaREDegWwxrcv+g5uNFVa9TyHs+ig25oBQ1J97K3
wL5F6a6qKHkyWIA0+DcLYpVSk7lEARB0XcaAQJAFpZwOeFjMoDU7Hv1idddWEITyskQb+LqOYlXP
HGSQ1gwtgKBpZdrnmMvZoVVCxpE+GV/VKHGJR9vGjwmliNBG8NdvJBCcgRXQlZaKXibnH5CWuXYg
67PkYNgLAqQPjbMQMTdaTr0/R3TItIWuau+W8WC5quoEyXzBv36JnfsFCAMjsuy4o6Pq6bpqxqNV
5b0m9SkQJqPlRiN5wHz5G3GTjHXBZ+1ZqY+ohhwBDe/P2pYMY5IrU5pTQUlxads92B5dySZShHGR
Xz2mHr0gVBuFyyy5mc0hREj3+0ljqdXoQyFD23pYY23vVdHSWE9qWksx2UP38ugy3VIwt5VnT2JL
TiarMDpTDJO4RIx8wBWerVM9gClmRY4mB1zDNkucSr664MCSzyGMk8d3tfUdrIOhCoCHm4heOPEI
942ENf9iRfRDl3T/YOiYtsAKKnhOH1H2Loc9sD3gKqZeg5pCtD/xQWwc3gm9J6ywWuGDAR7bWFW1
UMeQwWIjuKUy1utvFC+Aq7+B6m5rFrrC25ea/5+XTpp5grrhMRD1PQNhRiEnd7zoNJeYU+fEOSzm
cdFUkambW1LsSDJCOr+H/oEgAD3ssbq6XpvP7+k3QZIR13p1ZN/kLRyA/eL5+B40GtGmRtB3P4Va
aJRA/hqVI48k6EYLAjVC5QhgMnbcAKHv/FiQlqPQ6QLKby0fSbPBhiTnWsrry0Fq4j1LZ1RwJvzu
QgmiO5M5MLmzKldWllWscUWcr88XHkE30Vmb7gaM2CfszJWYF7udtMAYL/2V4b6T5uYAq4lX0/kx
O/U+eQd95EipyS5jJpw0BbPhkDWhAIkAPVsTBo8Q7ziCL2hKanPnS0T/wU6xAcgzSWUj6Z2n+jQZ
w+ea6MGFZDdSdi9BOvvEIOBynQfPmE8TMKgCvtI8yL58CNn1Uv68PMyNsfupMRKtO/K2xC2UXQlm
u+SKHY19V3zp3IvHnaTZ9HR9pSpumIw+0LFFCpbGRnyHsKeVxfkp3xCVpoheBdz6ONJTaaainnIp
ELXypPe7DbVMQn6qQ07qYbBJ+OLT4OItXIUOb4y8CBmqlj7aOgsQx5Dw4O0fCoJ/BMCT1a5yVOXr
tEcbPx68AEBPzMmj+eGKg7sGFqLjpSOWdQNoRz3+7SmEK8MtveI9rrioEULApPvzklqOR4EbkgQW
wyDFKraMpas+FbnZhBb4n/bCeL08SM5KbktnQM2E08biIM9NdG2CQRcCI3JIbJY7J08Qzw5/7wG+
1EbrF+OUqdYeiQwJPmByvMSeYYvbqMZTDiFxx+O73ya2sOVvxD43MGd+vn0nN3ECXF1MfXv0A9rY
p9kRVVVjAjr0c75obfXg7LGws75XA8csnjJn8NIeSkuc+2czP9kHKwnHVE69pAgXJZ4Xby7MAwdb
01KCSECLNpE7zl6Ab6CogB9ntj9tqKKLOi3NFc4VR6NQAYiIK0mL6Lqi3NxBRKmN1lRefYyujs7x
k7rFYgR7jDryz/Z4sCWWf/sjrvbcX3tR5Zqok2jJmihGBgNPhNGutZrQDpqQ+PAc63Y0PA7DtXt2
pFyg9Xkvl7Xj54OlJ6+Ab0xLwRPHRgk3+8/AiRFgYArtn2E+M42PCsIIWLph9wnGh2gfyLKkNzzh
elqWOlO2fcSlkhM79Gs7b25qeu51P69Uf/z6UZPTn2A/VBg0pTeiMDCBK3ufs7cP1Ze9yN0TDDhC
fOWaHL596Xc9ZJJ/v2pUWgTgtTybP1wGOSCYVGNRIGtSYNPId74ihzy2m1LLXdRMAvUOYIVBZ+fE
TvKKwl3tkx92XHNGyvSJwv/jWpsCu3J5XJ5veiSlc9Q6AC/gg4kc0oy/LS04ARh8IXxxg9mMc5Sk
vrPip5MhEthiYyqBUuMFERjp9YwzW2cXx4E/TpbYxeYoWqsUehpuOp/8Okb8gENmuXMYdBT00lQf
jm5Jq11LB+8mvFDK1tPF9sIk5DF+o0iel29s8iKA+seTuz/LRD/y2VMunSysyk8K1uEK4voDfaEh
XMyBVjNP2ZgncRg0ctPFS3/pCQ+YcjeeZcm6DC9EDkDl9M/YpHrhjBwxYdHBdpTYmnU4Jg8mBSSH
Hx7uYESUc6TDjY1i7nvSTxEaJXP3dSKMR4qF7V3KApQm5r8NBTEm4O7yfdvQXzcbLPksytdUCvX7
CjgEP2k28FhNaDi47BMQxygLScRmeEPAzcMgev/OBUYcj90RkSVicSFsmW2/81juqSmL6L5gAXqs
HuEeLprkMDD1WDzh3RBjsFVDU0dxW+yOHhvktcDnnz3853mVw6FzBQoDy5f1OAiI6X2Rxnlg7QcR
3WZEUim2hZU88EkOMkFS+ZU3TDBoE10+WtvFA4zkz/dRjfBtI/r239UA1SAX3e6rmSkQBdBAqZZT
+BSUPtWPU8giSR5A6b0iVnLNyXbkw6LETWc7mi8dtpT+yKbUonbzv9IpENbuZS4rTOlTOG5RV9zx
0rXFdBDAiFNmnzqGyrTksFYaEKBVwPSoT+Zj038pMKx23cZujROf/RMAVHd3KjfI0XRa9xhZ0mG7
d1vrqyK1FphuL85Tvc4p+J/vmDBWvCNZwXknHaXSWK8AjO09iUWbu3DpTa6wRFn7flxYaWGforbu
wPFFaBja/2f3JsXcYc2Ymd4PlP1ZqvGc11A=
`pragma protect end_protected
