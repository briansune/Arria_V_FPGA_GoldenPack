// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:18 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VIK1UxbOcd0QwVulNZx7pD7m8TsvoW0uG/uaRcDcT9u5YYW00V+I0UYu1HTpZSEh
YGfD8BQdzCWEFjbaxkbOpGk6BlNtXSfyAOLfqMc0OiJCdq4hAEEhEIk3GLX1MBq2
ifO5F+CkWyqlHz/3mcLUG3/5/HnWm69rCti85w32Qlg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176768)
bCrfMQ+RDOnef6C06Bg7FINYu5zL0nWm+E9E5uusMcVypBjqSvWT6DpGZGy3Lo8H
tGyEeBi1G2KjgndsazMqJ1eFLKK2cFQjTo6+TPf0u9qzR+TAzwkxJKX3u6UkLOMH
9ZcWigM391p6mpfF72217R1irVp6UsO7L/aFIlJ6+cL+CErKzCQ8RYvziImuF1eA
g9SiGHtEbCgk1AUaS8vaCAEG2A56VV0kbk2OwEQu4h0iiOxutTtDsYyQ55RylDT3
JGgRIgPb14n2SKNLm8ufWnbbopHBstU6zJvpLcYKO1bp8F/rV25jU38fiOBw0rt3
VTwUmcH3dF4oKJMbSTIVRTCFsMc8rejdz14nh6LVzwBzQmbz5XzrNUqrzpPxXZfV
G7/RcuTRFa0OY8935LTPo1h57oqLxGvAn57wEQjtpUbes1b0TYUGLi9FU6lRVtPF
tf2zHzGx7qVOKPEaGaubQW0zcUSSQBqFn21ToFF6vnJbwGozUE76i9/kTuihzoAb
g9X8ihrKG6ADEnN7Ib+z7cSIjsPVvxIeFXEpxqvoYd0QjCrzKnIVtigPdHhwdasw
4/hFoCia+isSlJqlf3ZXWbXTXHQUc1IPKPrCW8xgNGyVeCjO1w1Y84zbNyu1XdGV
8OLYHv5yK9FBEeU+y4TaSmnmbcUAkKLMRP5XaBJuQ0tOsKAUYUKxV5S/dmApFUxH
n97mmDpgmsGzuNQKl05alEFJCTODCHGkvdlQ/CXqJ/c4Hhaycp937GW2Pgh2YaHP
WbaucMi4KJSm9OtpYaZhfFpfkwpx+l1AH2IB9NTEfg6f0cZWk8ZoHkhs0v9UB/F9
r34FU0Yn1XCQHOxLzX1S+GXe+9VGeWMZD0leQ2H7/c3h5ONeJQWF5+8B2vVnnmh3
wm6bFKMj9AeRwLZlkVKInPeP+s7xpnRu7KvMrfAjrBc/3ieueWoW45CcSFgIKEwK
632PttFGgKY5OC+9E1u/7InT6m3CEo+6u949qY5zDbV6255DBEmx03GgXISaI3er
9fhiUySRLFG8uJ1eQtx8mXZs2j1/b9w92zYM4/g7Ifbf2NA6o3FElRXUMrmHd3aR
EgRzSbKnkNoukfetpbHHi5rRHBVyPngKXwOBmzgCYG2kpwCgMMz3xTj+zI9utD30
IeJ56jR2rNpHYetQUClZ5Yo1RudIbEHltaF4GLgaj+LI1OQJK9mZ2VQoBfwdJyrf
zVcBmXFIbkJiScPKyBids0TPTplxGQX1BK24QUpS7jIUbQYX9U///a7HbqvCCnME
+CCwaipd08ArtwQEVJy0mDVCgwkYP6T3VhwZUUi7HNb6QGf6fa2WDWl6p5LtmhNt
cVtK5rsJw6HAk6hk04RX2YdEdYGTL4/W7/7Sf2Sn9eJQBWxxTqmXEqnVGRULLkXB
jFxtk41RYQgiRFRJCfqcRRQROnwiQUl5iBLHAXumdAHLIqj1fwbgq7vsmUqqbzbW
ZBiMgl4ZBCeIvFFBnHh83CZixKQ0TudKL2vkVLl0I8yqRQCK9tihI9fmyxRACrKa
eJ+bLff8mBTI3Aw43hDPiPTCQ4D1qdw//lAUOEE6qGos/BqsGllFpmcMHcvs210J
YgHWkEcPXm31fqeOAMluRDkZ3Ddi2G8pF+FQ3mBCIhNRn9d8hMbxZ8f+jjukupsH
iLaJDI4oqW2mHagpfIKTrL8eCRoaLu9jv4v/aB+7Gz9bKbYl2nJpYl625lKa3ZJw
Y/ESB0pRI+AVvap/lMQFXY35q0uO8g/8BEcLusMRdu4GL4s5YGYh2u7ppH0tFm2p
TGF2nAZfjkMNvRR98UEBd0Bl1ncORCAmuv2ma7PZDnE8P8aBn4dVm18Dx7fgMn5t
C36hJNSTYezoMA4UpNjceFZ/qzjgPy8INwCjOnjmsQdirKzYPJN0xcWQDkMT9W/X
MmTKRzN+xpEdamf83zdOVg+rJ3EgJHiKCQQ8JHQcqBawKGiOJt65fd7HzWkxqYkX
vXRw8GGWWvMtL0AAlrWjbCXwQuekwFjfzFXskNCqLPYyvNKhDM4jH2OCbhsXzY8p
ypz1iA/jF+mGkNd0xLRVOzUaekVdA86v3vb0K2ofhsJK6/CbeA/HcoXGy04B+oju
ohjP0YCivK5f4d2z7v3Dmdb7gMeF8q5Vwd8ey4xLrB2dkbaU1vr1Ooj6JBTOmxJj
+wLfCQ5rA6XvqavfSlMrRKsmbuBMetccmVZqOU6sJ3gV2C+IZoIp+XTSNYVQ0gXJ
3p2ZgO/nl2DSuIqLI2wO2INBI8vdfJXZobO+GVjH1QIXr5jFkBt32AG+BP3FNRer
udKYHSH8VrVbIhHwYLJ5mDZbdf2ngei4/O5kNqsK/A3lY5IKcOlPKVmrjhdtroV8
oeTdjuD9xwPOkjhb3/O67/9Ix6PVbjst3vIFVAg8G6wVdrzWOsGcER/RNy5C4w20
L6XBSaVEAshOV/4dM5rPRuD1QzWtCyoxjkk+Ua+jd0+3PbHnykvFfaEnf2Hp+wwU
BLoXOB09hGn+iG95yycFsbzsPpAUXnBNWUzFBbDVBAKSoFt2eAzBLa7st/57qI+K
LVUaVXWAesbtud6pOYyjTYfd/c3Z3TdCOn/ZsBTv8uX8xejuMbYdJYvc4GD0G6HD
jTgm05jicdhJGHVwCB4XnK/X1dUbReFR8V25xf6TWXzJQUYxtwXKB9idBeLel8Py
1oFrK7kvGdX922ZyNsP9iqgD3Vj5nRaj1gnumTfuEMvsgKG+o74MFs0Ytbrru8DA
ktl6eTAAE20Pj0nkNKjsRFKTqwpKryh/NY+TuK33+cdbN5We4xn1wXbtX6fXaUHl
J7PsvWD3gxaos785dnKsUMeJY1ZzLZOoJoTtKHQxlHmwWozzmOAd2sacTJXIvG8S
37eNSnbaW4Hl5wBAzdAhWPAugFOvA/JIKSQe5n76iGINCp3krOJUx4MBLKXLIACU
JDvKRdWKEXqm5do52Qd0/nPfbEE+g5fbIRpfT5EZYzZdwd8OT+F1m9ygiT9JgRtJ
K0LHLa1gJriwInyLmUDWMw7RuICcPPdYh5rb/d2lJWhRoAZG7Ur5aUw+J9SJVix9
kC/kN9NATBjiCd/MdR5qEDByG2K1g9mL+gjQEf5yYj6d1hIDX8YZ/lCuhzWjfF31
eLIzZMZmwfl45ozAQeiO4B0Wy4j0O+l08HRRcevZvxKhdroXykoyB0SFw41pnaxR
ggg8SvDO/3Cokmjaf3p+2h2Vef/Edwp0FtMzhmME1EPSjnrZGPrrllfW3JHJM5WB
aqfXeKaRcw6fZLqZsb4k8IXm2B9jFFLBVzNw7se0y3bVWttz7U3KmTZEIcr+BLrf
lPSk+xVpFAq9hteuTD5R3C2W9IOcAlbInZ8oqmPiawss0CLHih2YsW9Ze0OAMbw2
QFv/1OmXvZXoW4UZ4Ej8O191uzKWZ4sB3bc8jMgvQtfvAM2kAhE0eXr+qwxAPd3X
4TZ9+GtRm69+IcBIQPxFLI13qtNSQHwatv80rsEtYdsPQmA2wmSs7X1u5kMn9p8O
NZpYEGFtV2Yo+w+q9KMtTZGbZKXgKoPCufBnyY0FWfdVYu2nHEBD4BXwj0JWifig
lg9PsZ4ULWcp+YCyRSp5YgvwgxDRYJEHGqFTHBjLjq9Sw2GDsQIvbhFFGT2ei0vO
RoNsHdwtFJrHewrPwK9tle4SXaUem1BP4J/HKim+h6sMZIMARKaGgUQdeG62Cgum
UmAL4RxG6n/Izp/YWzIlKJ5xAI5/UXdsUwR3SVL1sKCfJDHb80SFabZEFVsGmfDy
deqW5HEVqm4jLALNONsVx/W1TDNW0d8q9SlJqnJxrx+oDd6Jzo2V/ytqlehkL5eV
dVBj9RfYaMKVU2EY3t8DWYb+kiYkSiiuxp69+WKwO7Uz4dN/2DvbOzJou61NO6v1
e2Awq4COFi/Fx9NrLpvltDhlvduHkkSQ48M+R3lpM+iQj0qxxfdd9MHVvj6cCxiw
v+yCVkQg/tGaN0y/IRX/bW+U7HvzLgaL+aMSpe6yUypSfmjMw8ddbtDQ1zjnvKWT
rLOzh4ZbOFVLwhfseWSkgbn3Dtgu3RjkyxzAjyX9HkD41nxZmYfYpv9rqHi9wBNp
Ts2w0rVGzy6FfqfncG9iM+b8KQsipeL708GGZ8tE/INmUs7fVsJC2d7bEzH04Gry
XFEYG9AEJuTenRMXMtD60lSSQ62WWByEa+/fPYldOi4s8Wa8h81VkusK3zR3PelT
Ugi2LyKPgSkbgSMXqH5v77PsYtPSi+ngjKBwuwzcAZn9xhcfzWREp6IsCtx0LT4E
dj4uhfqIl/EGm4osXys0t7dOAJUo4LRtt+MJt1pB1e1e1QXK2WiHhJELAZ+oKDtU
vIiB49pcXKzh99rlXbZw0/XwhZkdSpc5RwUCScIfQ/Iaeig1b18rr5YqTAA4FaGu
rNzSlK5Mg5udj+HpAO88Fc6+clsKckE5hq5jQjwrGcXL59/CHsV78Fe5mWH/FliM
GKWC3TrXDsbqelmL71sFm91musc/Pc3K6iFxO2hAmGw9SLecN9bW34EDMeLovN9l
pw1ydTkXMHKzjsZ+CamRke7Wzcp0Yy2W8StNEUv4gyKgjKAieH9zvmmmwYGJomFt
tT/Aif/xTBW0wvZYrIkCf4pQB/oWrchxd5xTNHbBWVZAMfF2T/7945HVAhu7l+Un
psouqcBeGy9839wNMbbrmDCPh3/LJ1J49WCoMjV6ISuSiSNt4MiFTf+YTB23Hz1t
s4RRAYAv09EQBDoYu9KKgvcgy/2lBOEIabG9QcsFQTW69XfRJRXIIXMpTA0NO4YO
56XtrQiZ9ksGTvr2WE54McHBno9eiapiSQ6F/Qh3AmTYX71ITuWIxKfLuHatp6RA
XxpDAC0uchHGIxrGYjNM7VswS6pinFFaf/AwIqPaB+dGMdguUi6rTtdy8QGwmiwi
CbI8jANc/bbdtir0dlTXLEZL6dGk84cBmsq5nc72skRDy7UhXdwGG8Te+ReU08ca
3bIUmzn2qCJP4mp8Ad4WIWhQ2r7qEyzd/KxmUaJtHiun2KCvy9DoFZORSem4qJRx
QA+lB6PPVt56ev3yEUWMI74Y9UYrqxkznotJzI3W2mQjifJFliK4tCYnlv3I2WLG
ke+K23VW1u7aWGC1X9VEEWRAQjCxgUqQKw6CqLg66rJMRIdxFJ4ffVmxH/Gno61n
zh6vCOcy7vaNVKfenbyI7Ay1I7VszcVTbQ/fJm/1DEwbcrIJ2/rlWaRaIoZ/ScyL
tVdw9/0RcZYreOcLlLhy6Vn0L+I1RJTYiYVzFlJ43wKEebipLzSPSezvuCu2R4Lt
rE2L9RvoFy/G1/sGjRqd63lkgVTugU8etDo5P2/jKDTwrPt8+i1hQkaLJqIk3rVJ
qLOphWYlq1Scg+A171ybMR93FBXZ+tLXGl5PxSnoYarjtyYKlEQoDPmnQybxhY9A
wZZHLtQr5+Cxz7Rg+Q9EAMyhTsEVYmfDO8Aqpa9zE303Yjpc7aQcIYZiNPZMdGxk
ITlGonfOnZLP+Hd2/rugwCY+o/NwRPHK5/FjLnQlhLkeuN8PtqGAbjzImt6a6Nto
4Pf//ynhND47Z7cqP5gJtYQiLOaIXsctrOQ9S2O+f/xhTeLV2Lf/3oVP1USj6sG8
S7Ija+I1Z4DXGNoRCm+rVQY/19Zsq8zS1/fvIPv/aJ/6gtRBjjid14fZz9hzfn82
DvUuup3XMYdMeCtF4Ph5lXHqIn0EnwZs/LQkv+M6VfpAa1VZaLKr3iE8CWlv7A2j
V8VoqxScDMcfuHkJTZSL63f3PL07Lm6I1j54PHIljnOVOwI4WWrrmel7I9DKCqXu
73zS5DtCjJ2VNlgyrwgxE7Cut0w05zPYGOdEnMltgcyJGa+vBAHIw0f1n8qncSHz
FLI0E6SzTqcNJ5zqKa6sngEougLgQlK5SW+koa7GeANML5sbfSU4qaxqtgmk7Fv1
h5cBaYn+aRYBAT1RQSVIRy4ZGceOhjOljcWaFQxjBU3t2DhRhSGcxSsa4lkj9ZdN
yvZMEsubLaYgCrIZRP51oO2IhZ63XtEhlG4iUpbcgMMhZ1ESa0BwVYnwt08ICJs7
dVeDafTEVSp5+cMxAJdyWm2B4lJwEMPPhhZoxtyP8V1aoGQ/aEdVfQDPjPlsOfNM
mUZSfm28/mS6Al/Oj8RuOQm8RXvasQB4XPv2WCtW4tIBwf2SEfXr0+ueZM1gp1Q0
ds6TKxcw8InGAWIN/Ckncjnf0haW7RLLmQX1aBqmH5PI9nqA4hATMz8u+/jJjcGV
5tKK4nVbV7VApcVT9YYt2PCGtWSw9ZhXdfoPpGNaG9oWUiDFhMcJrOTLe3Keyi4k
kkUBVgS8R7PTg7ABg/C1y/A53Wex/4F1hViCWHTsbCAZqJGbvrdnwCcRZQs6zU+0
E5woDrpsdzDHxjKoDWd+kBRo6bms8oZlzScIheSrbDwuiXmdIXTj2+po1PSynpHy
KnfstF5rzGXy5ncaMyKYycsIanjsDO4rNXaJ9EOHEllMgIKPcVJNZPnqYzsJnCaF
uadfSBBjfBZzu1IEY5uGZ9E1m8ANmSC73jf7/D/eRkdypCdivtTODUzPgp5i6HWo
QclsaGNYu4FhUt7P38EXypEt1jxyM3C9FBluypNzAE72lpfX7aU5nv/451RtINqe
3JacC8a3J47c4wzjGMX7TaQgot3vB34KuTOWpDPo0WSWwoQoKgqtojIb1hoWH+xt
CPvkGZyd3xNR3lJ2oq2DkwSwuCbYth3gtYuE6sibmgwEB9AyWqQZE0J/BARJrm6T
+pPMjTGF6CFksFZ7tRYFModJwrsjvnysdBElhOHCSdUJO7XxFtDZx/XycqlmM7D7
dpVigMPiSsLtd2g/eEir+zgq4BJwIiahFvuQb2Id47yinK1YNqhJNoZTQpBLnvzQ
phTz84oOqTYltYvTZEAr9TCq+2iwmcok3J01L20qvfvYLVA8pqigDBjvN7MLO0c3
9iGFdyAFDeqbLKffgGiigeIlV/H3hHb7AUGmmXqjsvLK0r1XDacajEo1RJPgUpyy
WJ+7/V6wxwARazXjfw+VGZDYUJg2tXV7flx/gqqe5dnEZmErSUwbfo++eeXjZgBU
py4BxAp2DnvrY1SQG/w5k/ErZ7Ml1lSd3PNaF6Jsd7FIMegG55m2xjhuaiQZqM++
szVbiLFOsOSc8NNzohKP3874EDqkUMjlEDrxuS2wvjyn8KL2e2CKYjX/rLBD4wM3
1Hq1sZrNjrYauEirgkuYSBF0FKYM3KIcVd8/9QJyxVCtncpSHh+LYtXdCMuvvXb0
KOwW9n2Ujf9BGzdRnxbgkbmz5scGtbHw6OlU1GnDWaMYZh5JuCnjT4KWJq1ub3UH
6E25smf0m79t7xb12DHzl8LVVC977LX0ZHyvvkWw4JuZrAzRqF2ywiVw1rihMHsz
h2rkIsWQnbqyFelBShz1AdeGDoRZ6PXn5GXhD8IxNf4WOFX/KJnR6ztAGUipQeNk
8gTrJPwtXQau+UC4bsVaduwGeqBXh6dcvh+VIrg84G2OB2nTouR1ZDv7zie8loTY
REFMNJBn8CEJwQa60ooAadfsH+1jHL6k8rgc89PIxZcqqC1m8uofvGsg6uXq7DFd
yytUNI3SgUaF6I8YdvRAjpITlXevG3s66p/dFHYhRSoNEVdFJxDCwQAcqCqFQYwo
Hj16fkAydyA2ZYZa2tXxX0f+odQpKwnfStNCyTwXwPtubik2Fj3pFT8riHF1SWYA
kdeXbVwkV1w5iWg6x/frNpBlP3ZRz+fIOJ23cw8nnW5iS96YNj0w94LuxZfPV6W3
gxCWGFbQTByhqSc0HrsITBwaHrs3ujDPhMxqn2SMWwh4Kfeli6YY73bIjY4OliVS
ooYR2tWHzl4f+vZgoL5OqxX3Rxt42JQDIjrb/LjP73BQiT55N47p56u5xpqro4H2
v92Z9sjmRiNww8mFoqKEpAK8MAnxOOriiufzxWNnZ6Q8CyrR/ywWVwBx4e+UARX6
EjMWumJRl7O0lsu/N40dYDzBUQmGZHHh94NtpdNlmQK63ARl4Ou4YYqRTnxLkKqw
jap6/f0/XmcIYi0Vs+xChL1XZVkyAUVO7BfjdXLfBugEUfW2pN5aso6V9/CDKKPP
M5JJEx4CTGPthFZxptyuv9ZA3QY8rIfigAniNcFod3g3lD3Y/zdmXmhLiecwuDZ+
MlB7TdMaAJ+orK1aT4ILPYhLRNORAv4bB6r9OZ5XK7IdynT8lEyVlR8KlZj2KI07
r0St6vhXmGVJMH8+lxOsA40TQn/At2RL/oZSFkURjNTHWdY+jlSxO+K5FebnKpAM
ohBg8T0e+GdlIhsOLmnjDLvf6Y+ADMfkXk7z9sWybZaH5CR8c4AfoNv4yBkyaDQh
U7sTN0xEwapLBvmfte0M/U27b2EMFGAYqetMJaRfwJ9LRflqLuLHVB6ZGw5WNH94
TAGhm0yu32E1QfUb/HD6V/p2LYmqxGngKy95FetUqaTQUNHZxDHZWCprcu2IaXBr
H6/936YMtL0lzGQ+IDomHcv7+khjwV+bUP2qw2YpRSluOVFZrqt2SAndsKJsEdMK
68aOLbKrrW5t8VzIf/cxzGWg45ZAvst4EGupG3zuILxKIvW7r48+mjCktB9ceGv3
fgXvtpphs1WXelZ6eKF2M3YG7PYKQ7hc4E8nD0RVue5I5U0snmG6jZTjeGC4S0ef
+Uiw7jwTERXzGMBFaCYZnZoteje7mYiTLCO+IywS/jwMVHxtgPXShHUZezUc1TyX
NAP/+FJeElHedQ1Oyg6Emt5lReZuxYdpjot7Q+WyWW1BQR6lpRzLaVv2pYPtZvFJ
SxVHgoFtNx7kmil1+XKRP3N3rj9iSSZjCUBmVOmiWTWSYfuH4uCN5Q2vBjI+vhFQ
zQNJL50EdcQkgxBNGlAzN+ccf2KlgaYeEW6h/mV+Nr9IMhyJ2wSsN7INqgcwUbtx
VPCh1tow97adBchOUN61b7c9RXB75CY5TYK32YilpBo9+cjcUdVix3whLhkNVgFB
CYiOb6MAP8wOUXFHdAARkyh8qLanRS9Q0f+x2HxDrTtahz/R/zl/d5bnp2XMJiQ/
/V2+lZx5W5iAKOo+VpX+O4W46peFv4c9LYOBuRCAah8VzuK+LJBhptxBuz8yZs19
6z0ygqK3ofK044D4QkFO1i7BZsUhx39PeCMlzNLeoPX7rlpmtwXBAibHy1NO3lDQ
OxJsT71jC0y8s1bDFjMLqfqweuEIP5wfvJTgVZMkZO2WeI6E/LtfoPbz3LSKwoPu
J4p4Q0CfuW3j5gT/ToezO3rbHQsasJoG42GUeE+wq6PIEM+q3HlTnGafSCWNWep0
VFsdmUNAT/EP+PKmHLUOzIypUvfqPodX8b7hxFcwIikUot0WORYmOyA4Ov+DTDkG
6J3ltC7uM42dV/UiR86eMU6ZQE0s0g0r0hqL04owcps7/8fguTGDxqBgxhTWNaRb
ZQGbRJCEN19r0vkMaFYOg56lzDpLoMdNwr6vRHV7UpADRDcNxzTwaqprGy/FUwXf
b/Aq34+P1lf8KGLtCpC5C6KAQ6pXPHdL5sBWj+CupEMRV25Vz4vaYn454Zk/Ofpd
P37sJeoSxVzYl39kyM5FX/dYB0/TJIUdqKCq/JrURc49V0cq9fgEQ2ww362RTiX1
wT6V1XVTzkXxlvniZuKmMAoDRTndCANDNU+mZtd47PSzbRnFe8pqdq7S/DBDff9X
q+LM+fyDEX7YUPGFaIKK3q+fPbHz+p8JtXoiCBPX5LqmXSeGBoyqYoq/Wgpv8k9M
ifuP5cBJAAV9v5HV5n/tDiINg4DKA6GYgG6AJwSIS99wSHk/5naAEqdTBv7DE3qx
YJlq8pGAHGRh8AbyIYyuiW7qB6IE4StCadVVGDXQwWmR8orh2qfu0z6ImZL+g7dt
SrRZVCmfR9ICtjXyeg03BoOSCV+8Qwx/myRkRJWKbGslvlQbssQ4IYPV+cIa+ytw
UmfFH+qBdqhHthA2CRZeSH/ljMh5ZkV2OnmrpZNmRWzzn3Qu4Nox4WJU54nTX3r4
XMKKiZqK0MKpyQogoagkvS5oIxk9IrKQ2qWBU+IHD2sRSPal+K9iz6JW7yud1+zb
S9kJHUePOjr9jEPaGd7IOH/ah+6Ney1av7GkL0WhzfpXBz/1799YO1fKocW5AEvg
O6pkkI6mB8wui7VwiYfAQmNpbUdBfcAG01CYWOR+2d9Bc7mtsOG7tkk7exfiSTnR
1G4557kWi294mEAu/1pQK+fd0YQ3fnDmKfOzBlmuoiVkpty4BRysUiqkC/S1Iosy
1RecT7whsnKwwRHONLvSJYiSslTH4FECqpXRnwN71ffrRnMbULf/OWlUVhqGWnu2
asmjfZHfheCCnvO+nfmZ9/x2ikL+VxU4hYpI1k4Gwsi78f0Lh3yp0xhsM8MXYzut
z/AX9srYAxtSrYmdAah9PPUVSmeOhFmPsR515lmwb4XFR9RWupYK4x+lo0hyf4Bq
1FTYRjnBYYKPONXvuivT8icybIlLugHyVGmYVJKLDYw1zq3q3z81TiKGKDUV/yoc
WjUDo2/5IGQ4DPtsF1PIiSADYiU1YO7f3bosjfLEx0DBYQ6feHvLqSW+vd91NX1S
HVUzRF9tckM9WPHzWkHYP2H4riBDEFgG8VMMtfFKlz2cSj6W3F4UTBd3iLxOn9vX
ETeiToTWWWRN2MIDhfZ54cCEkIPWGghk1i0TimG/xlt3pEW8fAPhz2huNpxbhO/j
JpbZi/ParbO+gJBRdPS0eGjwtGX7hLgzhBiOKlu5UAE6G5nCuavSsOGyaeR6EWpL
VZW7ztTKtTmlETmIABLZ3pBScykEG8oxbeMzDtQWyvpZZAZ4MrmqJnawtejXeIP0
6t7qLwxP3Ywm4act9hHQYdNBkfPYEwS+u069gmtnep8oJw/ThMpP2dquylgSl5io
e3SJKSaoj9AUxim1+zw6ErPP6uCnJ7VwnNLRUd2riv82bGZPh+ZzD0BcA5S8zQbh
MehLgYk/kqhqrlA2ihUmv9vkTnHMgycZ0VFwPaDr+tZvXwMXde2eck9lObVnmSWF
Knn9TZPIK9BScyNQtqR2wdW28ydahb7crHvX76ZoTGj+df9buIuY92h6VvF57byu
YmGhWqVv5QW2JJqSkfgQVxpThcONtQP7VpKeJF9RqLHReNlqNLoPdkjgpfm+iOCC
eH4lnUln6fr2loLPFvPqqW36ULy5HCB3PJkTVncgCaM7igM2VpSPkryTI5jA001X
Wf7ztRjiOkki42vVDI+rVS1wimZMeoVhFQEGtlRBDc7JnZlHI9yT7zFLPuBgJztI
8tP2dAEigJ6WoCnoHl9WzDJ/DfHq9tL6JAN2Urd0cuhqnA6MKBMz/aE5qbe+E0F3
Q9prQjlrPGJR5mZ+lqmDaenQ1+Z8kprGcQ6IplwibdmYp80frF9Cp+PMNwe5MWst
UcgNhPqo4x7kG45EqPPBny/646zm2iyx2XBOri7gZAmdKDP/wjVhN3LklDA4mRDA
V7hbczJ5dnDT/13snMcH4E0puYA+65p1QMJixoY0wbAUuOemasXX4krRBpdbIlHi
UT4br0icuxuDcbTGQEZkkczN7DAaTrOw5mqCot/tVN4OPQzhq0JhRXIU74BCoqt8
0JhM2myIldMNsLvt5FYhCuh9O6cnXqYdMvx7bZZUGMHnfCynfvblWWhTFl9qIB9u
gYr/hLtjAEcl1Ifg1piocVHoR9v+8frQW00yeyorUXiJnaH0NaNYFgxvy3CHFSlK
JRnYODcymmWI8W9LBb/nBKZH3Xd8Q07nLaLY3r2cWjXd4DmKFZ7u+KR6tKmRPE0P
x9JuOXI6s1IhomiPlnAhtsZJXZeHE7UAKCfymL454if/xYHEvAhW50k1HWrI23XK
ON0YuISf86Q51lXXQRXmzBKjpbHwGtYwyeBHVBNh5RZJL3ZsgSpVE+iyNIhYtAPV
aTBICjcM8ejcmvod5aXTMJ652++Qc+bolLIo1KQhV9NGt35IUsgtcDYwh+pMAdVQ
ajBpQ2zuGU/TItWtqfPcSacAW5603rJsvIWVt3+RO2E/Ba4uk3llkpPVi/V/T1sf
Id1R0cQGfV7jEtF2A2TKjic0bHpN9Icm7qgVbwAY5BsAZx4YUjZ78zzwbA4WRE4H
Jzo3YwIw2c8jg25AjYQyTEpmUgI78/R0IfpVvrYqliXwtu03Do/1t+mqzEJN8qkL
9V+B9o2y/TEzspW76UwLdDREfZchPrDQvZpip6tqmv47xFopgSAq7KmLXbJ6IIzZ
gEeL1KXishXuFuPY9JCHwu94oXD3NbSgkX7WdAL2vFcjmKoGPWBVQjj3brCFqdiL
cXJPrZh0wGk54csdMgHOatdHCdxYQknTpKuOKMbB2ngj0dEup9EGJQpfVY5Vslhx
VDXeV9L/J/wJredeNSOegpLqsAV40sh4SbRx+XYrmXpaA4bVlBsX125BhwdlbEnK
BBCqAgoghGszsXDVSLnNUpka0sLac/E24aUQCbnzaPR5H2MN+7byP5MRJ1pCkpNK
A6NH+yH1tFqZV68D1DXkydIB6lk9joNqi9L27n4tdnRQyGj4oVnp/mX89lRWdvE6
4fA+/XkJXVcLzE8fGudoihSO9rs0UbPcQTrUZT4QZHFn6LefHSWLZ9g7SQPxi36u
mU8c8wY/d7yiQGo/xkwYL3WlJXK4B2fqRlPXYFxDZcUXe4nM2SZJYV+lUXVZEps9
pt5ohaB+YLT5famW2IHnflso3aRiNxVolvlmwmzATWIhR5TLp83GLPWOp33afxig
XjYMt+y8e60+vcW8/0cy/PMX9o9h3jUxyx0bZYjyZzHQ9MiFiuMzQFv1WTdZ/X+l
Ifw5XvNXzpCFxbC0XN5ACfMt2v2Tfc8FMadzGfxalOiZJ+KmknO99XyIGvBSCA3J
MjUYeIoFJvvEVyOSLW0wuasQjUlwKuXadRbjAIEDcpGBKunXGmrRf8+ECgArM0VJ
ZvpJ4ezhPOFyCD+pU1Epjfo5qss6eS3TNvS0t4V1s7hXNQ5jPAbtLEkOfuLeuKUL
jLjolpZjSZMVlNoKKUATFrAlCsF1MDYvhWiTPKIkWefpo9DG5YXWb6NsEK4Ty9ix
D9JOjKv4SquRe+bY6CTshv5z0QoXiz6+FQaMPa9a0bv29U3jp9KkG8o18jjViq03
6BMWFExJswlPj0+IwsjiPi2dh43WLxKhuqnubiMXqQva1ENpUERmIGLsNkHt0WxB
aHTFysIXAiZFWi+hn+s84BI9tyP3qwAb1p+jqhz/4qLiAV3ONlXmw4l0vj9Plai5
c+5GBojOJuCRTwMtp7QGsmzUsQShia+CP0lfvHhf3uTa8ktZtfR+VYxYKFEtcSge
ne+6RIFAAGl1QdtCvJYtJ+Wdb7Affe8Y+yEPhbaNP16sHCzkSTewUTl2sFechT42
ixjRBKFCDTmpSITPl8+9PgUP9Ettjs457ClovBW6m08iKxTL+y0sK0emfc4+Xiym
QtSwdAbdnCpURa7CJdeD/aRStigTfHVicQZ9mwcAMcztK1vnvne4qcikNHWYgA0t
4ZDNXFNRaDxOZYYVuPENkVHWAVTmSM2sOC+Wk3q3Yp0Ey9FjrinYo+tbvDpslw4h
isLHkgr0Z24JwmknWs9K/KuBlQs/uiGQ8eipmLqSAKXi2+0s+bq3HwNulOJ4WMka
TO7k2xe9BOXrVJWTdz81WZiK8EfXWZLjv/NnKg24NgElWZtYE0J5gO3U8gJSWPuO
grPOouxgACNQIbHGEZpBObQSNk4gVcF7n6rL59orxhGXJmP/wtYTGGrQz8Dl6VZ8
lW7u60sYh6KXz3YmRAQYPDc3kvKV23RhdcIf8PRgLDoKwL9zS7VFNh541o2X9t0R
2xuIMm4MjrPtv4dfYLqSvxSmTTr3iR0uT1N8U9DiJ+UbSQMVclHm1DpMa26qAfbu
ay6EXHaft1IolvVTP4oR6puG2ppR8O/O8rN3h15gXmgM435lb/K1xU05DW3QOHsU
otzBtluR6ZuFv+rhYlCI5uuAsVH+v0XDKXMZnCTDzqLq2hOWoeTCEu3QRO0Qeceb
ufZsT8R9XW9BdojLnn2ZkpTjPUampKR+5FPxlh/IDNSaQk2k6hcTPxgZtvq6xN6w
YvlE9mvTGJ+cWGuCWSUAIX3tLgeCKxFZEo0Z+8uIgnQIeT+pOor6a5Vs5PN2eVGh
W5jdnD1zh/yaEonL+lzPD4d3Dz0uPJJcEfSU924b6wB3cPgR5XQD2MeolVYARBKC
ywMVf6PsnfTlyKGmjzE2/sDFAQIUw6pYz4vuPcbaU3KASXyvYcVgq8zl7Jj+Lgnx
WdwMaL1gKgqyJee/zaDqE5vpGvedSQaGb9BxTaMKLkfLEcw3pcUKitjNEdfyc9Wc
B2OKbUBFAvu89iwPGpSwjc42+gSrbNlgZE1VX3dnZiJ7C7dNEe8ffNUqB9Jxlay8
fGFktjTsAWjNSgjyZ1GRgGgbcLp4vD5pphucUxU5YDeVlnE8ifsDu6cp5fPC8tDV
gUMcHLWETnofG6ul+zMdIao0j6DNQxBgrob4coihaqZNNMTL/WJHyE2YtFR683A3
iUwsN5UIdkW0cpijzm+24MBFm4hgvGmNMFBn2XBWmmUC5Q0ntcmwDuPIPBOMRAmD
00dJems70XoWehc6+hrf2dImw0lVZ3xIZKzC8+DnUC30rQN2g4qd8nmRqVt3mWIK
Sc9aBSqlhNSmV8i7gMlFZ0SGloF0Q7735+jy4MWWHu2xwjrVRqAqZ1hI8iYcALZw
0e35xv31x6ddFhb6OLHpwzfkIIgZlP83Zk4q9MXHLz+HKzOUuYSqNqukBEkRYx+W
IP4Hfc8tPelWy1qhhT3DLyB8kcl85znJzVxg9VJdo4iGZJMDvORrBYwxovQcUFf9
KYz13NawiayjHS7XceKnTDCrL/lPeHr0CZwCcfRAI/zdCyVv0sVXUF4XXQyqOS13
FsRIDJjKBJbG03uNUZ2DiL4aAL9vKx/hn/023TaM5EgKvCmWLk2pkxnPY9tyJS/L
CcBwwHU+d5tc7dxd8M8zgPxltCS0f/owElBbPq8zh+bZj7Bgvv6qMsWnz4vrlKNx
SDHmfZriW1XYvPsKVwD5JvcOp9idsGFzYko2BIc6foId/qB/wjE3SEhzMjkT9vB9
sueMg+15HNkVYLRJK85DK3yToUonbvtysQcWdSW0AwZrXdySBG8ybujKVDThArop
+w1BjTWgOe1l3cijy1si8o2J+tasl5dtpt9HKjeecvLnM8wV33xmyJwH66RgrKWe
+jxbN0dXFh2m0uYEx9w0fiRF6JpuvPXvCHK7T6DOPuIHkjIvf3LLBjP/4Jj3WaI6
sOlUC8U5iw8zO/olS52TD1+EkWS8H63gcikHlC75FgR/IAnv0IPr8CSu2uYJQJJO
nfJoIYmX5AXyJEWa0oZmasFAWKLA5jXESEdUIJVonUcg/MWHUQxGulyAX7s9y/yw
toVQu2DQUCE/qdahhNOiTmr7AJOh3MMAcF+9Jnm9Njfl1V37NjEsWmMjlfNYF2fU
lvucNFo3M9Nwu2hrtN0DQxaXB2qZ9LaZwESYX45cM0v8WvCITvxh3RV+5Tw/tsq0
bzJVVrGv1EDMzwOKWjSBw6dobsQ3ur3Jb93kSjhdTwUo8fSwYxF0rVcjbBfH2sPz
r0OLGTlGBe00tW+ufS4J0W7WYEnGD1o5faYajW4na8eXPlIG32LLSq0Uw8BtpMZo
RippNNbwQBudna3bZKdiycK+DLMrhe55vbdr2gUO5p/yMJ0TlZNhuEGmm8k3Ke1N
ZkGZX4738ifWflI5rVbR7pG7mGNLBgTqR7roQ2bfBTxILyoCgf7MrVNqPJlWC3W8
V64GrNq4ISa1A5FsUhoSGbKPVihMeInsuMpgik6v10DyjPyk0/pj/RITW81o+MHv
JYVBiGJ7Y6um4Ano3v7yLw+g5jXZ4cY93MfXx2snTTMtn2CIyoTHidUdMSSoo62K
jMx8KkMrVfv9L70usB/yEFW9UG9lF/jZzjItlXCBpugKsURw4lv0PnHCkXvXTAQu
G2jcLL2QV+oykmVGfbw1nObEyuuhNUyin0p5EtjuYFG3yD5FYmHzODZjuQu4n6/z
crVkly7VU/PseW++8XSu1tl73zuY7MmAhjfn4wBusvh0wWSNtxmaUMit9NvmcZRj
3mnoP/JEPXgGWfpWAow8zZc+KeWvk5G80+UUrLoh1HQ0V4JuG3LznqnyjUA8ZtPt
ZGD3lUZeJRMN+v4fn4+piMh8yeKqRsxooEJBYbzbBQDCBp8d9WMdRRbSee+jFvsF
X7Qg/6UWGVDbZl0+C7jfRVdHFLt1MDCdjv16lVtTZhuigaTc641xdozH2on/kj4I
sPVhzVSLztYBPjxVgeTzyj0g7Sf4pWL/9tjpz99ROla4EKeQGNAhcF2rk9mOETRe
7O27thVhWmycvh3SKFrgAuVuKNvsLp0BZhuideJIlEz6lZy2Qlpajk/IPgrvq6qV
NOd96q/Sc+34IRwDatHaMc5svhoYGekVBPuxBDUhhLVcfI8aPmd8ZNGs146lWiQi
0qLtiAsJ24zvS36nnUAtU0rTsd0mhwfhNILDbWoD++aY03/FYmwocwFBaLFdbb83
d//EAbQRtd9gW0smliqQU3tlodRW36MDqxyW1OO99TkB+qsBqQ38DCBkcMpqoqBF
aoI9MyBt6Kd5vBB3w0fYwXoDI+XU+J/bzBdEKq26/7Zsb05sUMH6PKHB90sx/8+z
kx1WB6TiQXZ0BwHubcQlWjNf8bPIK5Kn9DHwDJb5FZc+Gw4ztdgNDoSVLxLV4Dfi
Iio4aE6zAHIPcJIO3UvE/EotlYtlJmwoPSWugX9eL37Sd6RH5CWdKQIOPz9teLkA
/eZjbNkZGmBF80fyCQ45aK8tphGdiWqroz4n8v0ApxBJKy/BcpgMHVkTTQJdQSUy
DTgyeVk0cWwbk0ln4vsxxqVL+6PktTw5hTl/jN7GDXQ3dAhkv6wmwmAxyk6U7Lb7
xlHWnDLivs0Gey+9pgN2vu2oN/afszJm4GhFu9RzGI5FUvfHHh00yXmhgKhRDu/q
mUXzy12PKn7QCJlvE9LX1cagSBPouoOiRmLUG2Wch9jwL4/AzoO6pyY9AlasRHth
Si3/McH2Ox5t8lD96gQbiIYoXnYpEP52kMBTd+/And4gVg0iQo1YIV0F6/MVSnbv
pe+KysUoDfffO+0MFFO6Q1VbB8ULj4KTKhl1OLdF4lWkdcQjABv9JIvOZmMt6+6O
UmuSzjy3kD2Oexs95aj8qQsO6piqXUlDmW4JcMEkxAZ+txL9HEtTowoB78JwDe3W
3UwH8d14nUXKS9ogiKJW+Nxbz/hgNR2Xc65ILYJ5rqkMx9cvek/Orbt5GU2i2Z2Z
ppAljBqg+c7K5QVqbhSWv21wr34TUiJc4wO1WcdBZdmswhnqQV0vmm1ogPGmfQAi
Zp4wN4nV2ZHQgRO/fTFVZHp7vNWmZOe8hVJzmUC89TlG3ieAZu0zfeemx59aXzqu
qxM51GGn6rcR7WEcWKUd7rcn21M1yaI0x1QA5736w2DHuWmkyvxc+6LEx//hYVKl
XFn+JQTJEhqWsuZfAhGjgmiDHEZAUivQXnCVxCd03/nA0nGUdrlTMWuJmLzx6ZxZ
dQWfFKJwn+yZExJtiiax+YKP7RkuKQJJFo8ss0KSv8eK/+NMKyxAeWcVOf3fxd3i
uVcge81KEno6W21xB6MrB+CHQGPUtLUo0GTzNllFaHRGFP/yTMPxxEkg6E4G6EmT
qE2qcy8Jzs6gktJSxOUFybArHfMyxbzIKFH1uQRN/rQjpyP+liWEIKYcfqQAirNL
5DC5a+hMoVg9n1wR83iFYRlSmgjKc3dDNk50eS6Nr8U7mH9Nwb++LJo1yUPTBeEN
1O9dDAhntstoJDs3tCEmm/wLXQByVq+39/NPqDyC5BaecpJSBqHawoyKcrDu668X
r4iiHaYzqFovgD3swptGrFJhQ3KFcoQKJ4EeCZR3wrEHhWUM6n3uddyXP0ag44Fq
kMDiZokKBwfm6YVIZTIWFgmBx2BoUeIsGmdsTa3fFT8N9TLi09Pxgp1PNRVsgZkp
RxQ9nCXr7XEr1C80CMjC/F26FaeBwEv4m191v9qE7WeI+8aruCEaGQW3jvGhmkqB
eRd2njTFMb0sPPtulFB5KmQOzaPR6Eneer/WJlA6uIRbRLE419GdlsBdEGRwe0ID
WLEDIw42/wvUQfTmkxmC03/thoM5vCopovpu3H9War5e+jQgCvXXhrz9d4tfvh6A
qC4WINwijtyEaz+PXewq64GFqmrHf9VscYnUkOStARF+0N+n8UMe5MF6WMKcF9f0
JMm9QlLxy6jeo+VJYtpIo6e+GEDPnnXvAkuXAddy93YtIGbmBfCpi71/lG8nsQeC
4mYsiq3QPlCUDybvNUau2Md1T5Ni0TEa3nkxdg67iOB++5i+JlCzWN6fsJgkDC1s
KUXIfwwA27H7w/w9qAdp69PPBfWqZfMJUKH4GkCgXrqmYAHBzdFjhxEjPbvWT/WK
xEXO+25Ofop7ShlK/fQMgQ76f0gFC7rU2zqPQOca/vb1AIW4VasO4vwmJOGqeVj/
V9I1blRRNM1wD4hqDRiLl5vvFqFh6W6Vx3dMIc43WCoMRiU7oifOAqGmXjwf1Zru
t8b7GO4j9kbAw8P7qw+iApCVgyJkAK3Wq0xTbenZ+PBtNcsNQKceGV6xDTceewnS
/ASk7G97Sa/E05AYX98ugmyGVR5xhx1zV9nNe8VAJnZcAdBh7sIdNZqSJj+bq/s4
SvgDxhR3phkXgFxRhfhyQ18A8n+SUFMRGydmAbMkOUc+Lw2ptXYobDP38mJHhXip
TU8kYx7ALynNmopX3fU1wO3KT76jUC0VhrZm6wW2rTS/1ETEDgMKa7bYwtMF5ihl
CKAvoP3kLTzWx+QC6EoLCGYw+/XnpOhQmsEfcFhEWMuxXbNrrHX0zwzm5M61/9UY
x+yeQa2BnQpZBJ+h6I+PfRCnpVMw7r/k1+tRJFs+fw65xRT82/biB1ylUTQGFWEM
SMKYrOHmrAdJLHbpf8ctBndBGok8GVDWUMmrbw6glHk+hLp71PzsuWfCwuahUptX
fClru5UpUhQcqQcHX+vBqfC125wRIxwSuIlFlPhSHqFCPnhHe1aea2EY3nWst48e
EYqj+4TpEG29+ceTkkh2zeHh4l2G3/S/4AAgoLt8a828Dz+bEWb61GtyoHvtarIV
qDMl9STM11u1XcaXcSsXEWXr+CjMqqpfdo20YZnpuZJVFaSckcsHPVacphCnlnXX
NvK1KXe9cSPFKO3sSksh+km7qXdxCOLyDjXUcpLgbQN8HjXpJmsadyCVm0ZkmEQF
CZaTBfd8fkIW+/1yGNwRdMTiAsecmWQuuVGenSf6fty/U+tfMd8RKzYvTAkVO+Uu
N/kV+ZKI5acA2Xq+C24BkirTdGIblQwhhdtXW8f2Rixdpj5mHBfZz7Xb1Ze9kEak
D8vr7kB58dQrY1XN4hVBhJexZ1DHnjRU8HLVF3SgPJlRYAL409lWLJpK6holu6Hr
KKCudg9tnVng6pNwIJISZVxVc1Ca9YTaW9XnmhMBIlp576WZU7hZy4YqYTQYD8qv
WI7wmf8tC2V4GikUfIyyambseTiKBrXp9/itlE+kWZ4v2KY4vz0AdaBRsH5Wsmuv
JhkIE9Lb3EnkVIvA0jNE5lGGT46rAtx9yza/Hf4sTg3oy3dIF0ScxqqjlbEWtozA
PoQGVQDsHQPIlnkzmZUP7STbFmnpYd6+Y9HVb+gk6iFZTngKM16uv348tzb07+Up
lc64Pof7x1p9HFdZ1FxTlN/1/qEHYwzbjafGKUQ/LWz9+7E1HIuBM3R70oLAXc3x
SrUioffs2AfK923pdzcjpMqqNP1CnSJ/lw1kr894IZyWjad/+u3+ZxsgIiInOFU0
POOkyQNG/IJwNMwXbTrec/m6VCfyo22qF4ZW0bnCRRq2U5V2cvAHsweBdQpLzIb8
1u3cJinh8r3ZYTVUB8SGQyN+29eF7QYJJbc9x6rG0A6dmV7M+X6v0NBZxxLpigBC
6eZZEOav9tok4iJHi59g1yRmkQ+JmiOrAcTCS0cOPZCtXUMttqooBRYsvTt82OCW
nXkR+P9SvlmFJQ03yaThrfJewzbftYFCM7z9UJIOcaEZfCipY9/qsp0EFd5JhACl
z9sE6oi7Ll6sEQ8WJB6cYlEGKu+C4d11RMKPXfsDXZFGjX/Q4zXA9qoMnIbnJd1g
+hgKdJAd+K+3HFYwFATrANDBVhmc0CfX7fuB1SudXVtsqyE5NVhw+NbTCdL97JFg
q8mnCew8uNZsIh2nZnmYLj+5HdiPy5MdoxiZT9hTHilUG0jQFsGgreV1zvJQs18l
rIMAt0PLtiHsgX3YLNjb8Ws1EAQAKpoZ2zIJuvsdPX277DvJWuLTsXLWaPxjf7Or
OP3D/IEhJjq3giqpLgwA5bcA5cCH75w2rsrr+ZzxkdF0CWB9tkpB4Gvo6Z9KuNHh
807EIYBTYRbhGzEvs92neNB9BY5hOKPSZKOBZ35ecWrFVBFIE+r1rylpXsargTqN
CrR00dTy/MQeo94njPn14nCJ6DPo1qqWuhc7sCBONjWygaZ6OMyqWsotucaUPJgZ
C+0opqAQCv8qW3vNbrF/xnu403RqiJhcHqB5qHHi97UqHaa+czmSPMItcH64lT7/
amrYnUXRRaAoZGSQq3exvbVlq4eLBW2l5ZxSIKB0oJTRXaWJvVxh6WNutGSMM706
oqN+1ZKL9XQ1/q7BrOeGRvtkNXlBwjYY8GdsCNczKgJ1nDx7erRnIXfTsNN1cD9J
ChQ6cVl8iL1OPUN6JKXbALkRcJnpz8bkA8FkxGCGThtRmiZkQh8Om8xJj5uh718h
2KnktsHyOqGkafCDj2NA+xRq0jm3gd8WMfjjrqMb2NQjUyEko6V8Hub9jKFaJNDl
SPvk9vOx+LeqrsXSPzMLGsg4LSFZKezBk+2PpqUB3SJxGPT8EakNMkfZx3lsMthm
w5pAJAXc5OA30onweyhyy+sUS0Usm+atPa54qhzf+sBRRZBku195nLSLgAAjFMtH
fipw8X1USwXzqsHHQQAZdjzphEaTZXu9Havfvlk5P6dc/N4JLO6Np1/jK7nlpfpb
kVKfHufx0P/01hRL83ry7SppVPz0a/+R6en6olsSJI8Y4CodnXhM0BBxOlF5XuOG
vUP7EU03urWWSeQ7iCXrYuowq70WOHzIkwgmWvjBT53kqlLyxAHpITKHpdyrpgNI
ZTZcymzZfTH+tTugvL+MfxSV2JSqFFA/fzCeLMkYc5h9Q3RvVkjZmQAVrwem5Yo7
M76SvifDlObBmwiVdJHYi1b6zILF8xHYc5dcPXmQxyxZ6agq+8SRefuyvg7YYpHs
1yqsrzViQFB05uC4k9vtiwiaO8EtW0jkNIKEQ3wNl6WBjtsKucrzlmia3O9CEbvu
W1lthPFE5cOcMLovVElMT3FzjGeLWGaM2I06zOxITf0mz70wt1li9hXnWWwCpL3S
d9gUtq39ljOZ/Nm75/rDEsQng2kkLrb38hv+XUOKbge8wezv7mAqalrs2LVuGfIu
AaMKjDPbFfbRePgDVjOteWChFg0lv2hPiRUPAoaHZoZmHKmlth+/ck10sqiyZsU2
M0eN7Dm0sQ5rGZcgheOAYPDiyCYcPEiYQEfE6DoVrX1tfAQ8F7HiCZysc6Qx+8JM
RAqrgMCc+rsUKuc21LiNlGJr2c++aMCg6kF4tMupUdkO/TH12wK1gtm7RT/Ko4TY
LWH5hqVys1At23SRBkw49neMFIgcPVHnX5PVwOPRJq0JCraJbWxXUYQAHujvald0
YK4b9FxG7fIu+kix9qKu4TuI9ygMDzAit+kuecStTWZTTdtAB49j9eANs9bGy3m/
9/RTLTA2XyGPhIusyeFYJanCy5ER0QJ7GqNGiW7DcfPue9jNhoJSLvrcTeAthebV
JGu3BBOFba2kyugOuUZayjyjjMoSAuvN4okGBDxuI2Y6A2B+JSgqmDbP3oz0/cps
w+kVBoh6tTRD0REqk5ycYVcWrPxJXGdGkxDEOSTxodqiURnvgvShG4QZpLOOnjY7
RkqSDfFe8IKV4nEtIh0IjTfOUD6DA3apUhESg7esk0oT2XReYErebGFr+tRY891Q
8Lu2YPkEw+BSfA3yPY0bhivRPhSVc1zgu8rIwfp97pxpWJPYDQL+6Jtgo1+rDjIs
0kadoiFlfNBLrH/He2GPEzOHj9En1AnKW0fYVhTZZEbl2RRSrJw0vdSZmSlUjPWG
0gyTrcdlXXRE7Tj5xovNk2OYUp/QtcwYw5pvjxgGWCswdrNFX4NX9AFZKefpBBr1
sexxkmBHpsUiv+AHETYA278+34OOfgXEoB/At2KLS3i+VwpuNOS6K7/3OOYdWVv6
oLI5HsNAgidUsAYjbViDq8ghMHkHxzF32Sua7f3xkxjBYRabBbcGKbx0OHs3YlfI
cMi3XFc5nx1RWVMDaO5fg+d62zcr+V5q96Nqeh+I5cZ2vh66Gj3s+g7OhEhm7H/K
RPEGpQhyqXZRrpfVLXeVJifhzK/Bf4QXMxPZiFjGNXnAEMMw1/vTA6qg1tcCLTAu
ixh1wSs8Omg6ssMWhTCz6eCxoAgFBachfRkSWBWQHIVpxeKgOru1NoogzJAaso83
VRVRwivPlwci0TP8bB6mEaJRGWg8T9R7hiK6KAWJ5SuZCtu1nGWZOtEcHztlwNRj
VOVabNPlzkc034dIneOTd3kdK3xGwBzEXANRj0rFKZa+WBNZjB0COC5SDHYkeyaw
3+GLGQYKVI+kqrs2XwhOHqgPm1+xiwhBlBXPRMKndmBG5PHZhtFePlT3PuarkW2S
tM5F32z0nuT6BVPWXJksH7U4mwth7w7gim/1W70U7wf+FOlceAOUIf+30tWXofjw
kXUl6xGTAUVZbl484Ge/3y7fh9SmAfVjbrpxKEFsT+y+RWpmwsRJDPmscBG29031
TbJGzq1GTCHhCzvFKq+BC3xxWlRYhTnKbRNMopU8EbeCu4E4JR5YHpRULj13D1oE
7419sSATRjv9p0430lCwY0/A1WWdoD8j4uZMKGVyIyu1E2MHUHiCOU7T5M2GUd+K
VRCnFBxqde+dFOcrUz9eaKI55+z6wB+4CPFAhkqYO1Bf9OEs+LGz0I/jVyLhibts
lNPrsano2KqPhcJHl0A3Twa+vp/1NSV62Gb/ICIXdULe0BCgZoXQfCt488GjGeux
nxdd0FmOEEP0fvvASVNRbyq2ZvVLXdCnW6GRejMEOb5yk3FJ56gDfCusmpmdKyn3
Es2t/0fMxgsJ2xEdh7bOfXeIdSu8M+RRW621qMyKrsgMtA81VG+sCRWouwMESlsx
Bh8bVCtReVNv4CoD8RAxtOMElhoqdndEKTx+Cqj2cxpWpPwWHNW98HuThb8gTsoT
PJcfqQOQGRva8hNM3v5+0vJMag0W/N5mztJRLIKRtXKSwMdahWZeOi8wlcNVLtX/
hsSzTZ7qD2seBygnXodiVYtnQHujUP6+54go/VKJVUlRZo1TIBwCKJxTm8v0Xjhz
0qYIs61freMywOvDgsNsn0juc0z5npWJ4QZIy1a9P+4W1tosbtcY38PiOGognT7P
RLxHVLfurT33w6N2H633Zr+R9GsRxKeBF7JVr+m28eYtX7IYyFxyRkdFCrE3LSOZ
nvxdpgWSD2/UGlM0lL6Re0LnUCktCwYICLQwo/RTPdHau/NuPQRtK/RgtvLMmm3+
MQEYmSkjM/XaBVEWkR3U83FyJytDZMiBgYB4vAWQd6i1/c7f5Jac8fdZByjcfiG5
Ey9sQzYaqgbZavB6cI2oSzhF30Nv4aBnfoU3pYvyzz6nZvuS2wOWSfjTpqh8RAow
Z0fHyV1JnNWQRpDcOMnutSNmfzih1d7UQfbhkoNM3R/Si8ERqL5g0/2kh0XVQflA
wQdVwxeRww3XoXZooTQ7fIbg2jV8IAT1avEpPviXdnHUMbC5RcR6zgOqIpVaZR2C
4BxKH8D2sgNF/iWav3C4FREafr5dAFdoulMVHtBDXXpWmUCe66xh9WufcOTRV0VJ
dh41UOu/XIGjrc5M+rGAknPUkTkkFi5lX0BYHObLrkFOiYJyp8/VdRRB0/905Dtb
0bva4hHT63p4el9LbDt7m4QlpIgBcPj/yBRDac4Vg97euNeVqdNZMbCJbGqQYpGA
UL5fJLzLIXKGE0OndyBH5H2isFy7ytsNy1GYjzTQzFocoXX7NKDPRBOK8sCdO9UO
u7RO2a+n+gHE283OkePY4tOSwS4uuLBz0rFrjq5Arj4dyhCpBSsJc9/Sxcrc8XbS
OQ2B2+cCCU+rbcTBiDPY7aDPwDiItmZ4ZwK0KZmWqp8mkTyPJ/s6kdZY0izabA1n
zrlK8kmka0x7jtVJLzDrY7L1csVWfQSLakdgR53xLAJy+VxO5U4oU6Nsip2AZM2g
kASrFTqRRBeVqANxQxQIrV3y7w5FJv0unt+fUAj+kKQbuysagJixZaW0SQhGnf46
UFVpBcSyjYLtYvNKROZKoPyJxslr8q+JF5/sXrf1Kb57UMyDLvUOrz1B5T4vBuHp
IZ5qItyyHa370yDHzIEMkFXAJVp/tnSlUBAGqnUoX/i7HRy0TPDUeCYPaCbJAQBW
SgKTfC01HfZgJPZ0IRb4yOnRhxQ97i5W6/2OuvgQdSGcNZ8fwZp+nY8RYP89BaWo
bKvvEc42qRaQZcD35k2O0wIM5d/IIAl77BDhv3d8i9Yz9j/GdC7QZPfFZbXTumJx
4IKf5KdLdannMBBSxv/FC/W7JboZ/eF66f1JqqkvTRN1/U+ohNEzrIijLMUxeQlt
aKQdgua311vcsDw95kNwSRyGr1MpH0WECa0kQgYan1PYY0X6Zq4ekoOZmSHEA/7k
1/xZCXRu7xMPg1Vs4Qk4vYjGKbnTmh/gEMFSfzftoSAO4qtFlK7fPFZqcH3dNb11
7LAHxJus5Mvg3FpLj41t1VVGV2pPoglEu9NSMRWrl4kZc8ynnOIVnQ2a9XdE5iKJ
tmHf08H4Yani7PaR1r67Fs82U9PITnB5QzglAsncuAOnSE6kaCfruBzLKcAteYDe
oFILEW08ekd/R9tfa/XLk7TUPdSxxkzfPPFOYtHu6J6prFX4wLbKEYm4VGkxiSMm
Sv1pAjCR6PPOx2Vfgs71CzimJWch+rqDR7Wk2VffGWI2xc1Um5xJGkG3XFoFBvcw
LdhkpHdOACFpO2fCvF5Y51EdvoPbC44BhK80QdJvys8q8mG7ANwOLqFwhAYRlcgI
qV4TdzGFuZzXQv7zSulY5gR5zCAXjBl+ABECokFfh/kAW+EF820H4pZYCf4xkcQK
0FDg6aykCXB73hs55BO5RFWuynfkBSg430CLhZvwg1MtRDKs2/2CP7v1zAb4hQ51
W4IkUwFm4fg7t4Y5VXbVtVMveh2Cbdh7a79jdxNiNYICOTDnbsqR4m181ByRu1mM
8ET2cDha8p/P36HzB/hJ2MPkbwiSxfh0EXpF/ECjm+mbl4B227rii2+c3+IZiXIc
p+oixL8NHTV9Ee0S7pRXBD8E9MYyjXLkJKbXLdCAhXgd6RbQdMfsE7DkOZeibADo
bJxNbbuI7HglCanR7rVyc+ORqKm+hqgwYxhrExGQUEzedIyaWlmfyVCeEJcbcb+d
sF1+jv2yKhxjGTVhYbveXw8MxoW9VVFvcvmNGK8K2Q2f/+22gLfsEHsGbeDNkO34
v021Wchzz8TQgmr5W6TLjcVfKPKLfw3PeQpK7yULODr/LM1qSGhKnmiXmYRtu98V
pjUAtiofHbwxX3gUfQ/Ag/ynoqKOlbqNON6gHaxfsO8r10QojbGfLYH/O6z61Nlm
IF6uH/IlIpAW3FAcGDinr9x78cLwxHT0FGZ/Z43vzzZn/wfMW1NrTBqVJkEDVJDn
Tn51I7450h6OCI6dymbVsErFlG4dRoOz4GGbbCp0UrxOZcGZFJIps96lNFmay5HV
kEBeJqvTMPsH9OmN4SmdvJ5e3I1uQJ/Uy73r3ztF7zRrUUKBqcn1t142BE1OLIpN
VeCKiKYiqgeqdQB97CUY+G5l9srEGVtpKitQ1CUHe/+sR4f5Ndsr1uRURHZEJvKr
LiojhfzBAyhzCeoERASRafeoVo4H0ndT3dwPycmOYOQxhOoXE4Ylb3NGcLgbYxOn
ftz8VzWlDiBuX2+O3ojf4tvEoOUOkouOqUNoCILxMTB6zPhwYQQxBTVhMj+uk1S5
yIVm/lnkiVFucXj+HHzG49095guDdByI0RuoJ0T+wpuf8U7AO6aE5neW2z9n1wF4
HpTSAc640+CUqjdza39ilfQSOP4Z9l5jqGgEYRsf8RPBoeHZ+bESz8erNzOkMwrz
+mIP7ELZMud7kNS+UIP3s9YuSpi5EJmm1gLOEmvMwbz8LTBrjMI73vDejEyMSyQM
uqSlvhqSzWMTOuc+b4AZFGzOtNPiIP3A1u5HeoEykrJx1mPnwjjCctYnBQsCN7M2
3kQFjd+nYWg47ahnHfOZ/dAHOGRI+13xFatW75mTXytq1u2hfRns/Ls5rQWtEVPA
uUZkFATB9ZyEcyBbLbljXwzfWM5OiXCSGp5D9TlxwbUDW8h23+RefaY4+vyoVIyo
6SSm1o8rJ+i6xlwVBG6o4Cj6Th7l05Qriysu9CT0waoNkju29UMbgwoXP94O5Flt
URD9Q9NX0JYkyld4Eq+RWreKW9bt0709DWx2PDdHQ9tQcFGfEqbpTI6g2SP/0wno
jURcaIZ9lDDhiLYtjUvlA81jsM4usbpShFUseFp9rvIJwGzWqTV5fs3Qc84iFKsE
MsuFBMqYAK8fYfqSS3oxxfVikV6hDaVnQHxMrIreBwmXR56Na02jYoVakWOb5+fa
rcKClDLYDu/ZD1ZkFUDdcql7smkG06p4uf6V50uukwqKFcoC8IHdWMI5yjRwn+5B
SAJocja92IP7lXprbS4uyPZEpnLLQzuK+4FDcvdqlt4u52fyLyLi92cvx/arKtj9
tLt1vrwTKYYlN6t0ntHqOsZHa3L257IP1hRcwZQ7pYyTm1AOmO9IJk+DY/0727jN
NHRHhY/MiGrWeyDZsurMgi0Kz6lNhKMTJl6Wm59maq89rIJheKlOGpX6FWrtih9K
67km3A1TLVJMNMP47kKQUtK93Q8C2Hp0xYAS9eSz8MkjnHvxG8rEfqSTEipk/MFa
onmpTCkNoE2SJ0Ufd/H0fn2zwfJryKU9TPIFDjNgHdS6w1o1yLA2LBrsWBgpLTWP
Qe/YuyTlQZ1qR/WlR/738Z58beUH4U+TMF4rhIDX0S4nNe96C02M96lCv2HfbAoR
TCLV/a7A7Vz0PHRvMs2aN79QZljwOczlZmGTs2jjMT4hR7PPhiGD9pMQ8nxmAj67
xTzjcQHgIMszRn4U8lu9zH+lDBbaIqA5ZiwkXhQO8GOBB3anzPOJztwNDCV8JnzX
FS0wNDLpWQFalfQaHzaybCJSYx+/QcI+bFV/Qs1cGDdLzVMbCKV9EFmPxuP8cmEi
8+Wehffb0QwiveIjTKgo8GbO2Y5TFJ06UuLL8CZWdiaWXXKYu7kNYWq2rWOqZbEa
zDT/2nr5Fidu6Oov+zV0R+BtvdF+RTBQfBP2VRsGvQfTuUEv4A4s+EHmFFiIvb2v
tA3Dk86jkKLlo/7bM0OSXD9zTa/H2BIIeMY7uc2mdVr6lL60NX+qPWDYMCQKlhFY
Iw6cQPCpe1Utu5x2/z7sY/RVlike9prdLQKaYSgN1XgTn6aFeA8fmn3NT/XB25au
LDIuxlegSGrz8jF4cbBEE6jJwolchMX0mISGcQzx05Av09gULky9cC65eZOheZLc
vQBT/4PWOU3ypU6+p0tMrwwLdqJA7Ngr/tMJGpffVMpkumc5OWV0cX5hmHACeOpY
FjoDO+ASJ/K//KU2kRZNaKMFPkBVx4zL+nxeMrn3XnInwGw6cngnA0ATa6fsHMD8
cEeGFi+ZRrHqs82uk+28aHHaNfUfg8UKbgDEfUFPi/wGgtD0vLs74GyYoFCZDiE+
edY8vuE9zKZ660V4adio+H4rZTsMVzdpvSU7nmHuiXSMjy0yEftgc/El0cHC2Dn+
31zdBke4BgevnHrSF4PhNV/ktRs1u8rRxwsiaODSKKQ2ywKmvEIQ/twqPp30wTej
THgwrXCNJ9APAueWg/BtCiLEzl9eG+Iz6uEKg/vMZCC6g3Ulv0rm7vpSFzJxs9r/
CtQdYYZIU3htl7thGqbPS+XXaCOujtSP9BI1+P6imWz9lluzlQPX52TlgmEG6avl
gMtt1LYBbsSfR2ilYZEqbtyo/ascJ7nV9BwYzzp1mFwNdYIuXq0NUHT9WXeOMG57
jShRRfrSxDEU4QUkfb4W31h0efAr445lY5HvLdT698QeA2KhNMOj9Bn7mKXX0hxM
O0Y/A3XmTHOWUZsINf9fTR/cUMQfrLWPhVKy5RVTON5Y61PkXc9udFrqY/xH8ein
is1Ku0IlnPsnKxai4bIvf5+XVIJ5UibEmsIBRkuigGHsxClQBlJK+O3nTBvEL1hV
RCJ0HnCW/Hu1G0Sa8B5hd0W/HyuvC/w9tVtf6Iit+fbXFMf4y/5ovhxfISdGwdRJ
h06Ed1fLN1UfE5s2aZts0kushXs3wZdbr3sr9riBZfQzKgmVg4sBRcrHX9X3GiWc
LQ9T93QkKMx1ENbeGdLCQ8/cCnAaW8YfGBaexToiJ+yYiZN/3D6Yn/7r22X+kKjG
JC8Z7hNMbQ6Xy+5jg2QtvV7TCq1drnAZ7a4H7Mr7KK3JDDcIM+NxVAXLz73WoJ8i
jGs1EKod1qy74VBBsEabjR7fc+OdkvnvMNYnWXCmAuDeguBjiCQnzNXdBRVDl9Zr
ei3St/Xeek6VI3shb6l1Yc0JAbg6fk6yV1Awhd2fEvXAX8kQEjHzilllFKn6mRek
xKjXIlpld/jB8hU7yhGnoJHnPQPjQIg7DnAXfuPQJ+H9T4b0Mdl/mSLNjvld1PUp
oHIoNZGgGpr8xBj77aORXcOsaOHaRSDMBZHfQXK4vHY8KXRHZi5DBGanXiivUPWX
kBaUqww6IjFuKrT2zGI/4ZvK+cvT+2G+BC79bcWCPWjpiq2HFRmsS9IrcWJ2bCb3
+fJAzgjWjfAi+xjHFgirrDAaL1wmNtro7KHrprS7Gr2+vg5QYc+1Hr43uIDnkPih
sIMB5Fw06YuW5k9HeR3TTxsCc6I92sSV9Sw8r95CwW+vcV3nee8t5jI2afp516Jm
/2q5pWLCWDfo2FFP9tn9gT0WWUfQHuizzp50kEhxUTwc3XPDkBxrMe8/xnRsjRn4
qjJb9VgY/2IdCwy9jNzm9aw+S/OuekGP/YMvXpq/nWeyyQuwq3aswRKXwPQNFqO9
BVSKrTZ1N3BtDsObAYjBlW33+wJz3JGv3dSw9GlECMsAWTOiFY5JK3NfnUoF6CPW
4LcnzySO+NobZxNPI1EBpPkDOesXPql/DYNjB9Y0uFLVII8jOGYVx8FqNaIMoNyQ
SR7V0keTK4a2KcIeO5+XTVKYTR2CMv4nA2u+p2uXKEiinvgA3VOz1HJhHHil2wN6
2JuxpbpCvdwHFcAiLbVf7PgACvx/5FWuxgt3M9SaeUNi1ulUzyursEsTNfSVRsiN
QycV+nd/nExktejfZgffrUqPX/RH6Q0Bo4yuIcsbsslymxgnyGG0RB30q3nwf6Yq
kb7+F688BxkZxG1bhy+QZfjfUg23dnjGui5Zgdz98C6OrcPha4vmJOvCU667IpV3
cjN4uQtyIaXMtBFsd5eTVbhbK1wnl3KCoGVpTfv62VAuC2do+FvYnRAAkS9yPiFZ
2b1c+hf+mPBHHgyybZRLqke74mHNnVq55SyzQ0coeEUF8w6SjkuDzL5uz7tNEJCV
+6ZdZTUsy2Lm9I6WvXgmHn19BjUUSS+xbkk8mqAVmBlGD/3bk6NWCfi241sXFu7v
RRWWS23r2yVBmIdwGrekd17MIs9EmlBrHLC8SSRhENBlDxI76S9qWxu47N3ALCE3
vuskFWqcVMKrVTkKf4CpsHC0ykkP0LKV7loAYaJ/Cxn4agIKOmbPyH3wGZIewJ5o
6tHcwYSs2hx2Vrxjczq5lnFQ16Uk1eP8pL/tkGH8cHui4XepEZKQWmFiyYq9qm4K
uwoPpr+oCKY185N9VDBY7KTkfwXdsUyRBQ7gKzluCR+Kaja+0NotDfCtrPwPALlF
kPkqTL4pLV/uzN1QcLZQzBY6g0Vfw1jA3LuLiLTEH3HMRPHDrBKZKCifVBwUUh6S
BJWGdhRMc4btVX5yqhkahPfQqZ5YyB5IuGNMehrOVSpHPLnnXfmuUoxyg/oOymBQ
ceaB1lJdJVpITG94FfFLcH7sO5gjY6E1eQhro1iOLtquDIRUr4UqYKfIwgmjMPrx
OY6Foz5ZhLnzaDFPi/djarwDEQWbHHx1MbP6jlPDcGHOlIqMOS2vs2WvnTOLQjSG
mPn+DLecx24QfahxtgqTeGhzDFC3Y2vvki/J/ztWf6RYk7r7ZNS2/hgetl7tGBAG
hycYGvbHZxUeDJZ9o6HxgDAA8NBDW4dC7x4PH3ocEi4piEdTKyvSPDXLfyd5Nd4p
XsH6i+Lx0u3GxXqp49zdoLD2+WnWedWtAc4QBD0cldBIMJ9I/aN8SJfDHmzqSrhe
xLmTyjo8I/HnOyEfbiu79MvwmLt4NWBs4u95rf7qWkmlH18TD9aGYJlBXNP8MAmR
wdakOtxFtWj56FCtXm/N4mSwUrCBudYZ3M2pgKH/35C3M5XnxczJ0d+Qe/f5x6fu
nYUpSGcPIpbTlIrA9c45MCD88fKn9av9i0n6adonKrCKBPAdHrmaHjyE1x8yKCrF
ndpp/3fd6ZdVlKrjhoqGe7MLk6rKrf3NFfn94UiIs/HyL9N8hmYd5+A5ezwFJ0xK
43PJbrID6fpPu2BmImt3/Qmkv+1QmvVMfaxeTXH7UId4dUyyDVFycxeZEQGnBq9b
g9bD+674t3aTv+XwlsvEmxAX3hssMLN05sdx943TW+tb/Lup6S/z59oPSNc9wfew
DJrVjFoN8fXkXNnItSKXyYGrH8vfaYtS+IVLEczIqWJwlmKEYxS6yGq9E719Sp3e
An/8tgQajAJ4fV+s9QqmS9rAaItiyESFnCnallef6Bg48CpUQoVJrheYIV+jgH5m
5vDeGkxD5Je/Y0Vrw9vAUZ4KeVXhofwR2xbMK/fsOlCuBW3ccVm/2nIXks/Waaz9
ez066aBebtuy3Li7ScqlDzwA9cn/p5ddjOZb3C92JESNwsGBW2l29UvO3CAKOxbA
TQcTPu8vjj9kZP7kS3LNMB5b6zvSmdJFdmSbMQvDLClwaYVA11QYc8knZLvAz2Fa
50Bn14QeLO8yJHIEoM1VPM0SI6z6ZLzAYrixjWp6VwRCpJBg7hg6N3dFavudafIc
A/3fN9nZoWs2lZctAdIUtoz7yCTL1PruNddpwH6MFUHkwz39Rk6ZD8Rc5iYNasFU
WZTo/HmNSRP8OjcMVMNsWX3t97fzX3b0dUfJ5bP8Pi0wwmJvyaIBy55EK2bAuYOH
1pTvcn2kpgmEnmgMZwz9VR6TMfe2rn3Nq9fPI8gdoW8rM7xdNpDzmZh7MXZ8gw9T
wi5Tq8bFDDXJY/4rDwjlKtXKBVwbrN7W9F+moN2Hfu5JAMSVGLGz374PXOJwdByq
+R5tJrRNHKFjKlf/2grrNu12a3ZbmSfyZw0cmo/ACrnkDivRYifXp4CjZZ7IO+iu
bK1HpP9J9ij41BuRL1iRv/YcFzKbZawnuL2sbcCXppmLnKLIFRFU4I6k+zuHxWNC
hnesw5JVfuu50RZf+xqmadKOQTSYDafbzFM3Bc/NKkjP8vt7GAkcJa2OCkg6CG+6
jRlL0RsmIVfzC99QEIbm34tdY8/Uc+1wpaLWJZpf0+THDh9Tl93orLdw+3545Cqe
u4tEjrNP/1broLSR6VSaxMyHtPselbsRmvtSyWLSu3WcxUoVcOpPovh7e2DOkCU5
mshX8K/BTlp98TXXQeEP8yPbr3V4n8D9W5sLaslhp4DmI8LGjxhTmtAE5pJiQv4H
ymMkPDK1clgyTyGB21jTJUr9+9nXlpgR1THGO36XVVMCevZOY4I7IsWIXS3XXQxj
RR2MRXo+vSg/YhJppqTm7QAG6Tg0wmnpJm94SMYh3ogMCr+asjNiDh502tvOO+Ci
j0iNqlLnbOlMvZQ2nSeBw/7x/ktbau/kWfhI/5qqNvGBm65dVTNX8CNWmHo3aWIO
TVvkMdcrVRkm2aOk+YaPzNi0phYWw6cjDFywTyvobPzyjxgXg8F9gPr2qQBpX+Hk
k3LsvYaCaaxnPCnm3pV9ZI5CKdwwknY2dadjZZW0Wlzx5WGyYd03VfGLfpFBZDJZ
Vx25m5+Y5xEM/S9zULr8vYivn0+cU78lG71gu9SMa87918o8m4QRFbOXWnzXO5CO
NUAlBUeOMJvPOsrn4m8xllPmUOV1n1ODW1BYnqHoprUQN/NjHtLD/zwpel/xtCZj
nBGMGPcyVszdk/L4qx07mtegTzBbTqW1QjKawd++1Nh32ecF7N5ulOC5X+FO5eY3
hSGbGoMVdnubywMXJsgGoeEF3ehod7X2kyuRePJ6GYydQrFQR3sVi2cUzEral/mf
a2P02/Tw7slo9ZHMPwwO4OVf2sjAwLBv7RD7G4XMTks9xrv49251aOgTg+hONV4c
zcWPVnBaTqOAsicaSZ+qmtBDwwU4uZNdNCExu94yNm/mdTOdt747DEgwD9pVZdlD
fOZDXwVXqMHtcye1f5uJrqcqZ6M7H3QD3v18KRddIrHbqs4xZzKWKkzTN0yNBZCA
2Mfx5r03olJtqe8c+molAi2UzE4ekSfOoiQ2ZIsJB42qjUIipk6+JsKPDQDAI/Od
G3tmLvwC1bz4R/odDNAuqCt760ek3GY1w+k8fiixPUcNLzV2p9BYRnHxf9m0kGcw
xnu1pifm+PA61fyutE0SoqY0yGL9vKV6Q22J5dCuLTTyMDG1nakaGFppVuQQ9frg
WvtzvvnltwSlhTOqnTDwt+nI85wVOF4jHAWt4dMGKcM2O28lKcs+UnAtPYAVNBeh
K6XbuVdNMTHo4/82kbOqVDj5PFCciFa/LH42siMtRP+ir1vHQZuqppuS4pDWn2US
yq6P8zqTYM9WuaWCBkBySKzJJrMxEpm/Wf37mVNoyRqccz00a2Rti/BWbHWD2Qrm
xNU7ZxjTcssL+I1ijj2dKtm9Pgq8AdPko+VlFFmEazqvqT4RvzwR7Rq3LdWzQEsq
VzC7xgGt1zwWL2zaO83FBzlILGqG9GZACrJN8FdDx/pdRWaXBLvEDb9A0UtMK6TG
NWNu44mrKtUoK2p4lCW1VkySULn5MFPHJ0m0J2XrPQo1W4ARyRruDWameejpReZK
7nSN9YRe33Ox/9nSDLPBmLrpM+Ky/qG4gyDW5fUQMHRp7XVZcNkX99AXk69oC5zJ
n0mnW+1PdF57QiUXrNndYC1bJErHWwijcUQO8Cd1Cq1v1PWK7L4XOFWZdSHlEO63
Xcs9jF6AWEWTMWx8znEGYrFL4abcXETJnFGR5/EBm4j5blVVHDCqspp0k9yUh4bM
5suhtt2ji26gx8zZJNAIoqXOIpvB1CbgDbShTdzsAjErbUYMlF5mu6qJswJAwXh+
xOceR+xsLDr4OczA4WL5kg+xlEU6x4ArVAyxt744jvEUJh6SAfJKUL05S2h5Gcbj
QzMZVd7tllGCC6FHNeyU5fQ3xkaoQ6S0AE/CZzfjVIpK0CWowJsYzjbYL3AUgxR7
eAD7SqPCOmP8DxkMvU2d2orpSKD0jAFmoauCfH+KAKG72kj2xn21lfYKXI0Hgt9O
a5JnH3NGzi5L/Yxoi36bDwhbRPm7Q3RmNVxgqn5rpQ1C28OfmDWwEORfP/pSfuc+
lJUeXiNCVJ5Z4yQZFf09ZkIkfjb0DX+LElsByLJs/BsFYoUnePqFc7vOJG3p12Me
YXmAmK1MwKDsxKdbAEzxfbakKcvmOH5uHwVspSzJxuygCuD4WzblEbFqsFYdus3+
KEJhBrA8uBjXLRLoh5UIZEme00IzeXw9qwaqlSizc4c3ZZDV37//Sja3rDsi4cb+
/XmXpHUUtscNJEdpL8OL70iuYvN3zOICjwYbbjoVTv8Go3otM7XWCLaNVFPzZLBz
imTGTNheuaob1Yf7Kjf6PzVv/B4rzAzkdUjNfLBMxe7BVAcmye/rPulejzC4Ympu
SCNoab4kgyvAdsFfry5ssR3aVwuvErGXEm2BClOqvFvyPdVKGl1pBj0jfcltR5ZW
xvOc4urg99KluoYYmZtmG3SDS3VfYr85PnLYRPW9XNAhnii3cNZYMEZa72d94SlW
0Y8msLJjvIurSnVLvyGvO4bdH42X3bXiBQW29+B9tqT6mzCjy+Z5nKpsLBlHR/0Q
mWGT49b2Jg1TfoAA33JHtutq8IMeFYKACEGFK1dW0TyTcyNO/FI6oIXR3KWpDKJ+
AcW4GZuvCd7nirYjE+8rJlXFwKd+FOrqCwzh6yxMR6lr4vnKRIDR6OeNZU3bvkSe
jmC5AA0voZRppe5Ks4Esc+/EtLjWItd/Vem1oikQMWSbaesh4vlqEWQ8Ft0LmuHV
DAda4sMi3QoM6wQgQlXJM6OjSczakeoYAuzY3FpMXLThQY07zcvPVthqncAIGvjw
XTScQdVrd6U576Iho0YVcI/N2KpClfYWu/h1UcaPdT98LaIcqC0wKQQUK3eZQAkO
/FzXcmwuhK7W18za7i34DIomZMHxzAekSBCfL11oijWOgl9JmvCVDCqRPy3ioDNr
jzKDhCHZ2rfJr5yN0aNlrUo9QVqwgx/Ts1S8fdYtPbKxlYlSp2iKe3kHKoecHTYD
9TZ4boVzllB+WSRX10+mkhYuS8M8LeBYWsAayKmI+4RJU2KKmCTpTiyXmoYnqxhf
kg9R33mRXrc8sex85G+xpYj9yx1F5oWohav64ChEYhV3CSZYpdfNXDgFImGUpCzO
Dj5m3lTr3GV/uy15W199ILUt2P8yIG7uSwdZnUZiDaTuMyDin2qaQhJQf/ysKv5u
PGUWcbhG7FrLg7XfwocWd+ll4JmUbzJhYMuKVm/ZRo3ONL1Wzm83DpAMQAl/Bo6X
i4KprQfSiLzJLimhA4FTtCuDDfTXcu6VujL55AySxZxTWez463XOVOr+fLHdWx1W
t+qjaYQg7NP3mvGcxinl7G3Mgqh+S6vRbswd8QTgD6wWF8eLdEy+Vuw2zYA32na+
2FOCGzRziHuF+5so2Fkx2IETPreP4vaUT0RKcmB1BCOSHNt0ypOCRvtah+cb2e8R
oj+r6G/q4C3MHR3aBifMCt/6kKlabxigcmXU32iWqlH1Wn6lUHnq3uhxq3LeIADZ
NaDXtqyJ3+pne2Gr7uwfbHtOXRVX3ijF6gqXyrNb6f7osFF4OPOkGDaxpP4pW89s
ACXXaTEgaztnULXf3yLi0+8Cgq8wSpcI/av3x6E6db0wgyTOfd82UTkbSRRolD/w
ycoko7AnLVPqxR6LkxPutHfZ6cRrk4atJwbGyu/FvzTuj6T5beNOt2+ao/z4+WiR
xBjIR0bGh30ZOqUtaWeSTGtes4jYe2uVJ5Lx7S7XqsYC0riAumvIZ9lMWghpHw3Q
8DhoHb+N+1p1H/ry1hae3ET3ylNuMbOkrSmA97rNyxxPcUV4n0KzbVJ8SKcNSIGC
UMBKZCSd8i37KH+zsIf9Uv2udrDfhaFS9WPce+lAT0j7wnA7OrOfYv/TN/RsZSGl
E+Wb2KwVtpp/CewELT7dNhdAlmDITWQvK0Cc44iKXIWW/20MIW7f6XTopWCWJ8Ow
uGmmClonG1rIgzeuofmsn84jXluzpQNdT9M38hR+IajCvXMVXe5ETh4hbD/ZFIRi
HHBXQXb1oMHnKuy42SchSmmNaFs8KH7fpX1FIL2Ls6863DCs2VEB5nn33AeHxwiU
HbvvQJXdPuseaHHRNxjuqyj0mfjCqRJQmCW9P363Md6ITB81c9Z7wSONd5Amf7vO
qXLJrvuYqDIPTY2Ho7m34eRUWto2y0+uTLJP1B4hdWdISL1ge7V6HYlqp+g5u3c4
F7mAysFBOxpNEx12y2wYoYYMU3SRL6IEEMmaLTXKivz5uKr57y6v+SAb1Re+2h0U
Re7g2u9KfJIBgjjydiwMCn3Hj/rU9Kif0cg4sdKHZ0dFS3AnPdj+0cIG91kI3lNf
ask3YhibI5nmXcNFGFjojPxD5yjj+EOk0xHMqvEg7XwFMvnK36DGRcnb8cqmGX9U
8HutBwzh6m/rXhGpnRX5U7wZxWoZf2tZKhp1EngzqW9UJqGZAHRD9mtwd+UZoNod
O2zUxb38w/o+PrfXNSvWXoW9X61h50tQ4gRGYeap1/MydBCT+xVdkwEirV+gMFLa
IaGwOekSu0XkIOyUdgNkyeWu2h9S3UcMoiktRHvSvIzN2vqlloy/LVhLkQ3zqKKY
VZqokSuHQSurrAZnfyQt5Pf+AA7mC6VJ9nO7KUCIH0rate7Ml3HFdlG4qFWJoEJc
mDPOC2ttchMyGU36zpZCbc5M5Oeali3yFFuj6z2eXGOeqteh6xztI2g0gB8ftjoi
i+DhY2EYvLwADakwnvPukUwuURMb1PCuSd0IcLItHJ/f0vSiQ1plhgcDGyVznbtK
ikaC5XtWzKFR+Mp8kOzimBnz7Vh+Lnwmb+LB6DT9x4JxRYnAG+HyL42NdfbC3Y+A
plFJKVUoKHsp7U79lUpwwO1bM5P20ZJf9KGF4eXX1dnV4ovKQq5P6NDR7wzr+F3l
xzEnuUIK4FLzsI2Z5Gdfsyh4gKbAyl/yFzl6pkEOBkhlRDJaBT9IgwqmbNiXHI5z
g26sar/cfLDsw5ouJYbZcy98ja8+S4PHrSRj6P13O6z3WJpnRA4o5opU8z2fXJdE
fKQF0rofSzerWTFDTUHUnQ8ez8YBp8/MKGmDyPgKLq6wuE81QrHfPxKbtQEPTXP/
JkA82gvqQyYXb9pReo3W/Lioc1flMWsfelqih7RUdqLuDjKoe3AZ0wMg2LZJ2FSG
Vd8vs2Oqfb+SXy0gxxqUidt9lEemsF/3qB1LdGVMCeO2ToeFRDULA3LwJn32Kd1W
QV95TF3ZfS+oQ5mbXKs4/R8Yr0HAutqKLZ+3QUrJm8TMwuFyseDdCH6zHygKdOO5
TBJFtUc27rrGzt+rwQAQ/TQYq9tx72bB+kydnjOEOm68st+V3oCYfEAMSHRoAfoW
i+5yu0wyxY761gMy06HYN3wbqgZkDzp7ZQBNEi+SRsBRRzJCInloMcEigIWJbqPn
+CeonuUbr2xke0Q4yKfy7S0EAEtGXYhjkimnfDm8JsJGSO40jvdu6lHTIvv+6x38
0v9EwT7P+Ud5LJvkg5JgvljDjJ04pqksUUMLVLc2r/l7MzV9c6DXddBhgQlUiGra
DS1ZogbyAvWuHufzNzoDB/3ZQr1BeVkPEXqAMGhnLp34U2mK0ggr1LKp0CNJgoE5
QBnh2rJBY+ugsHpmCL/9Ko4lJxLzvZscEhONedtRgIwX16UwZCPJ4B/LsILwYGKj
6y4ZzSURkQfjhkqVPjagXieQXSMmEUrUhKE+IO6XZukyw3iC+W3Pyxra8k9Tm/75
Ccu3xbVCIexIK6YId1aYvpEJAbEAcuyHPh3tHjIXikSAgHJgCUjT9FglbUVttV7o
4CnFwfIv91+TbTTqTvmJj4biM4jQUSoNN0IBIY8bYA1CYMbEFx22e0D37KemI3NU
UgckXjohHlXWZdvd6NWFwyqFMUCn4IpDI+lq2LQOc8+/VAkwZu16ssMXAo2HWr5I
amrjkCESHtJbziyMgDNvB4rLHdOmL0wIOkF1qiFlxHIHkScdvJxRHHgaD7lSzFyp
ILiRMkA9GEmur5qfdKEpiip+eeB/xU4/tlIBYGi7mJJpEIBkWUTgs/5Wg2zmfDUk
uBII3rufx8RNPoOEvuXHUSfwX/T9AXNudkYMyHxl44cMSSPUXbHxezQ4XzDVmiFr
ZqR8ZbimMsVLa8Hu0UR25O4yxjQ9RbQ7dQl0x2VFAryW1OSRauqOwoHIqLea5jf2
HilRU3kSIYiG3jkNf6At2Okn3tbUFJhWc4MNuNy9bllbyG7+3qyOpnh3cSIhHqGE
SrguahzWYdInWPMFDLK60brRCDUK6GPVykQ8JxBEFt2zih7S9P9H7mf5vFUIsUdW
8PJXaw4p1g8KbzpGDrarEDJaw8YERXgTzWnbIad+aB0jy2gzxDGPFRabLGieHPFU
W1QT+ki7K7Ef4WWa4DbVPCQx174SqxYfdBP6kKy+XbW2t9UT54ZOr+9D5XkNlpJm
3fForkaRQYSc+6p0AJo3eQ0/MPYhqHzclb1dJh6jfqHaoH32q3x4ph6iftqsA679
It5Rex1KGfYVMEELzTAJlXBjNvz49gTN5SOXLC7nUOGHcYqJUn3wQP4Dt/BM5sMX
oB5ajIvoY/HPuzXMJ9xYLTKp3omHOS0q7nanHSjAK1zqmNtDJ3Td3S4xjxCgHxkU
AixcuIvhAAiUAiGVvOSKD3BrnUsj0WNscnD5HyEAUMIW/U3M46JOZIVLwAHR/1lB
7ah31iwnIB2kIngMeR6UPS/fvFyv/7nVEI2Z6/+TkW5R/O/X2gT7VGpvegQ80luu
/wp0hIpgudW4PbjZjwRulsOCg5olPPZMHPdeQ76422kGaBGKK5FXfG1/Z3xYqFsV
CgAv2bcEx4vFmKUAB62fUup0QOSwDrlyl4yWcwbq6FLMD5ofRuQR6KQD3ijVnLwm
6yfMpJbWfgnw15RGI0/uuF1oPRkqHFx54nvGOQwJvN1GkD1Wx5wf9e5pckaHuluZ
8qoeKmnPvOpQrejPa6kQpM6SyoXMav+nw2Nm05l2shsPCNhJEbSzaegkee7Ld5Dx
tA96N5M4xV/lLuGMVOGpzwEszBzc8smOg6asPdpzYxFJUf2fF3lqNAQx1MAkPH6I
+ExGVQxPPXtnwo1ZJkCD0E3yedxOMF4MvMncVt0OaNLTADkKSQhfBq2dXJikbwIp
v3OHO9ikYdfnSAT+Pbqhv/OCbZshOx+lsidbNUQpIXCOzw7wFFM8PdVnZqmvoOTw
o84sM00gmC0fL03uRuCp3Ytd0XxWOB2ZryHl+9+qcJvdNbd2xXM0mRZnET/ryPby
AzmWatBFvmD5tAT4WCkEAtxp+q3rnBCLLWXIGqcb3vYjg4wwErmpU/ekov5OE9DY
X72CNW6dz75omyOd5S3LUj0kU+RnghISpxpyMZbE4RjGGeHBlnZADpvBrQ8yzQo6
q8kE/bCcxD6DbM+Lenm/BWe+fBCAtM+zCkaABbqXfvIbBi6iUYm6X3ezht/B+mEz
s34qzOiHuAcHL9N5Ri9dcaTq7aO5Bzk6cjwIWmCzX7cmLnNHEn7KsnK/WiUYLjkY
NHtIfxt1taawr5PVNIDyMfbgK/eKIqCwY5ECO9kEQeS57l4pEJWgyr/blkMoVIbj
S3MFW08mC18sHAgjpq9pVaKKxZOzswXJMPgUNuXoVJEWHKZ8uwINeYjTKVJlxeN0
VB/9TQ96P1GL8rGHYIUiZTRmYpx5TcXxwlI6+qwt4baywaxBf3Qmyq+GENx1UGp2
nt7/Ponr6eZJqXYfD98RgtwNqhX+LFeX6PJz6mHWKt2Q+QbSu8roUlWdEWLjoShZ
8PdyCTQeyipgExxNhsae33i/6JAJj5URsuRpmncQLP0aDjJ9cunTWQjSRw9OHKzS
Hj7B/Le4P/MT5Z28lgIy2Bh5icfLRVbUWxLg2lNU+Tz8rowaQvg2pYC25u5axTes
xvUZubMzCB/x7Johe+jzNKvuUWK6mhqG+oelf7ugRrKqTy72HARu36uXRM/S8Enq
FWq6PqGhCILs4Mlx/Y7vmC5NWP+5V1bKgvOdkcRPhemOKdk9LUma+iRFUXelPx5l
FL6hpDTsxcJGJ0atR5IpDoaF4pvWeJAssIFt5xo8zA84PARG//t4ymGgFNBMUhJo
UJhdx23AOwpEHP8KjJRv/FUmhApuAACITbjy+ZO1q+vWTBa0dktSG6vs+iv7KWDV
MjU4eedy1v1pPl3TpOl9/8sFNTJEybpb1Mz70dfhB4RaPzDszMSZ7PnCcdeYsnRq
w/T6xdHSTleXlo5pcyo9pGJFjcTj7OyzOgTnTD1R4Hi8g6nsxytHGJykpr/RS5Rr
tU8wGCU8aeESM2Sd0J+mF9kg4gTbL4Z6siHLxykcU4TQpuOKWgC4mFKg60nD48CN
daRTzKVdGo6qW6b5F3/zMNifQrTDL8QWo21/gKFgFFrqnXzal9031obgPCbtiu6L
jjUus6phG3nHm0kEN2jT5ZwV2iFDFRigZ/+Rx/+eZlTrl7L+FrWmtQvhoM8+96TF
SXItchz4BuViNe+LyFLaQTXC4gMcpQk1oUjW/vcWO2zIKJ6iBXHpO/ylJOJPglbY
IdrTdWr4lLO6I0Ad9ToE1pADMiDXdCU6fku94SC7SMX+WaaWpLcj/39K7+jE58Hr
uOUgvDTAd4F8ofya89w6SXrILUaNLAa2FgSwY5QKp3JYKRE8hzXqnGsUwvMSkGhd
f3S0c2iiLt8IQeT1L7gCmDxSOwvXkdH3D638ehlPfQMrMiXINCXW9zsp32YAWW6g
7ONI79goRwTIq87u5UKIWGdKyE27RtTq4Nf+sVRuaj9mlfT9yEz88JlSPm3cKtJm
KiXdRHxCCp7QZ7OuEJoPFC5te3Rpu6lCvnX0dSzvm1L/vDoFluPEbUUNZDHUzztr
Y3a60KXThVENBWAmHBNWv9qB9Ka5QNl/WmajJfSXmE6ef/dL7vKlLdGVE/DvlIDB
Wjga0edOXAGUQB8WGOtPFRXXHKPmHVJJ0zsz2tOQVVO9PqaaJdbz9L3GtJNeduzw
rn54E9toacLMfqpgOVNjeIhstNuuKeJ9cb275bUqABECSbMpafNp4eDWLftJb1qk
KFLDRWERA+4Qi8ohk2REnJahm1VY+tP3BxmN/EnKiX3mwHZWksfGerEM/FhGzKGM
/JVD4BV0xa+E8IJI7yEjVfjhP8z4DOYn91MBsCZAww4bZmOLs1J9mG98AhpyhvOr
My/xbbaXcd4TrKVMGZhgAngqRYZRRZzlxWE5uq8N/yaeKbq5VcMc+h2R0KBkoIiq
4J2EGwL2pt+3+HJSrTTA1AtHWeliZ3hHqhFlzFqsEq3XNq+dd9c39H1mnKDl4Q1G
BIpcL0EO7ZE/Uj37xCLx7BXV0YBUjxBNvjz29+M8u4+bjw+t2Ohv9n5Q+YDB5PxE
R/xNTmDPs9hyR76KXXD0QqDPblIS2ytjDfZ5noURHr9IPVNbpYp27pJrRK75jKI0
OJkOemGJ45SZiTFeZXRCeXdHVt2nw35Vet0f8kM2i+8Y4irFEWUdZyUe9KKITdMi
c56BzzMdeNgp1x0EuFAOrXI2ekMCcmIjkq6NkopvGBochI004DJbb6h+S55qViAl
f4e75pqCi4tFaIEoxskDMkFLYzfjHpJY8mw4ka8MvP71sI62WxlXaVrfM8IbiuIf
hnVCNwwmYRucxr+2Wq2wzpYpmLlsYlvSrxCtOg/YItPRMjuDerEBXEVRux8oyxoj
c17FKlSZx65waRdY128pBF2k7ToHyciQYXg7fCis00H1hRABYOGN1K3oHp6+x9P8
3jdr++4peDNQnZDJCP8VzoUJqVqs1fCod5ZufbtSPwG58h6LW//085WRFLps9S/d
QecMeZToM7pfFhPB4brWKLIQB3SLmAJLu3Exwlu2T9gw4u9aIuM8SMtdNdtsRBYW
WM8Oj/pzYsixiRvuGGsUnLm8YKxkTS006c8Yu3Q/KPmgEjCq444O2P/4cUCgefjR
ROKWPwpAG5uZeI4uj4p+wIAAA1seJAk1VhlaXXrWh4ta7T+NSqJHi3ssX+yhx3kL
0aewUeWA5GgjpzKw/b6nrXjCJaVigS5KTH7qd6sH4bWKBSG+KQ5Rjc54sLYHzQuO
S1eAR9i1ehmv/aXBtGrXsvZfvRC9sTO278VAJHCDq0i6Rc9zfbEYsW0QwXxda1pG
aYFkpMMEWnAfP8l7xTuSuGVhV+MdYepp7yyI7xIlWahc9bQf1qOS3etd0eh8yjvW
TBMRDtrxpC8/H2JyW2Rgqd66NZ5itauO57NR9YGhA8PhJ80aaz576KzQyt455JsS
mQFbz8WTiKMCJwjLKGZ/5zkdBJZXUQmT+CM6v9o7ljI+zlj5+FcfoeHHp4y2PMdD
LX7k+eg2Rw/tiebAMng5LC0bEwuvyIPhyTgfr48RssXMCiXlNm0WYEycf3dHLIrE
+LfQaiXwJ0BM26P2/zg0ETrEaKofsPCPZilfq+Sqc4dIuoWNqiyfzt8iiLEfZVDl
iplnCswQHZObwg/xEVQ3LfGJj5Rjv0iEL6YSU22e4ldg1unPTLrRBLWSh2xQztom
Ef0VX3NLqVFFChnVlIDDc3kbB2KjbYpnc7PmEPmF4yZyBkiLyJdWqrMfxOb/9xhQ
sIe4yPm45JZnBhwf1+MrG1BFQqtwK/Wzv6daz1zvebudMxcJgbPBz3zZKG5L17MG
3n2CGSWvRZwPj1vvXNHriIXJoC7hlegAm8eFoQp3O7WDZdIJtT1Y064pAzA7/4+c
uvKTV9duykXvboeLfXvEtxX7M55hiS5zC9yXG70BhfIqOafdH0OsJIVWppfPLwGq
L/lAsHlZUmUBxWPjFdZ+zsawQS/udabNKLXkk3R/ERbxk19/5asiUlCB7sHEsdQB
wJLbR1axI+dXXByAzh5B2qDC3xUVlMK8K2mPkDTEvBu79WF3KiN9CD/6ABTbZo0r
JS8Brj9IUVEOssaLayuqCDpbCsPCi2F98/i6UaAx+I/tw83IcedWMb2737h8CYVL
lWAeR9PQUwHqvKBr9QuKvR8M8HR35xU3Bp1k8RPcfsHX6B73VKcNWhJqcTKWjFjR
+JDeeOI+XyVSQIDhqoEqPBkGc8FygOQcp/Vmb5ivrypZFflsf1wyEUqhs6Ijzi2c
Da10Xsv5ZiMjHOBQQX3bGdM3tAh/v0JqYm4qp0iUctG4uiPDzNRBxYPnvY6UVK5l
eRytL2i9WxHzHqEUTn1gOZeVUwNUHdcD5NM70OcKH0MzyvY/vMf6uLW9d1xCg6qD
RoFdeaO6773WRcuk3zzJtyTGWQLWJVgYj0jx7MUWZv1zRzwMgy07imNxzI6a7pXe
ohcQ6GCMA16/3Td48bCdR6V0PnYDovZolUCvkxCiA642EGW8XdiOGlUHfplr/69B
J1hFdxdkAhZRLvjkfC6FN3r0eJgMWMLpVz82z3kqNQRS/WuayO1y5tyaP3dvTObI
oGmFDNDUav226WPJQCf47YK/dTTj5ScrL7HiPQn0y05X0OsG4xFc9QlaYK2BxLQT
m4CNPEKzrZY/0P+VQA5oHrLG+1QYuixAAfvMhme6fF7Oat2ru+1hsiNJMQtb95Q9
6nfyjG4T1HtoV5pEBa20yUDbXUsCKl2WR2+A0mIgPoBL2hpxsJPHJ8Ym4gtx+OD3
vuNit/SYB7lYnX/f7ubpW+NhE40HBn/5J+k/HXxpHoZIlf6bpKrJR5uvk9wDILim
2FvPr8SWCoxlCeX9uJPm7cngdPcU5UU4XTlZHK5cg5rGAfxWfgXEEBOQXOzZ7rsD
5jjKM6HgaxRhR7jSpAFgxth4ybJ/RNXvbo8oh1USXtF8vRrWX7L6V2xGTCzxMIvC
2mEpgXLoC1AZzrEGkkiUsezisLP1/DvLQZNiEATSN9tDgwrPlFZStautzGeB1U62
D9MzwiAWXhvQn8WlkEnws+IWPE2cTpFM5yWir9DW/hg6xGHtiIv1WWtiGcTexqaB
QoduNt9wQqtcOxrMmXN7Kgs05lyfIfkfzx3dT+piytBw9YdH9jbhWwz2QLO21l5g
JySJ0fhggd39WWZhagm41IahukCub1ykCz8CPZGL19KdWFmto7eHCjNCx9dInq+f
wI4ifc1fp59GCSA9MKoSNzyd/oM+AmQAua4Nu6JFA7K8dNwC5h7OJBVuOJmTwUeF
UO4TmaZ7/fent2IoMkfx3K/pL2Ry+REDcvW499qb4jlY+1EHMAeRVVKJPSQixDIa
PXhF7nPCMJ+jIZWCCsAI52RPpMcZYJDkeTNHJF2UOhA1KO15M5udPsk/giRb+2UV
atcHFV64IxTqjH1sCEWQ5V7LfaVr+g96Z5BI2UwzDdpd/WqcabV52WHz2hFopxKc
kcrhDVNy7wHQZrW+gIYouxilSYpEUVaoNkaXrYINRfBWOmdVo9f4BHLdt/c0Z1q0
PFXJO4cO6RZVYszCev7gLDfcw0Ck4pSI/14ts3q3qgwHwEuYHSK1p+NVjCUF/h0W
+1yOy0K4RY7k7q0X7FjCi80l3rvx4Qtgq22uHCXV22HzVkVcyISnNN+GMp8dlw71
AuUEmRV9fxcHfWaOcfN7WIpH6JZGI9R5vJqzlsf8RNPciSERpX1qQi6RD3lU81Zv
3Q5TU5A6ad/fTQwj1csVTQ5n4UzgbX5CzNNN6gGgmUno7BOMv09rpStAQ4z6MMRk
5q7qt7RceaTh0BOW9XL1MK1EGXvuNpr4loBpsnNBJ0TVUde8TOgX4tUp1oRDNar4
ZUcOZlbYYiKpA4UekXQYe7JGUVYFM+gpzAGXljJdzgVzsYZMmYPxfZV8FasVWh3D
wuCW+NlAG8BYS7kgSUfwJRH085c1Uo3+aQJbmGi2eHyvCQr+ARPE7JSj0cHGbspZ
MLtfNjdrDpH3dmcK1pfz0lvzCIiWMIWEfhShVt8d3RfdVdRKFUVTbD6eZ/6R3EA8
WxR9KUro1j2Dx08hC0aWfD+fCrgTEnPx9zNjs+X8p0vLC0Ifbfxbs6mgkMpH8n2V
Y0G+XVcyB/FQCBkFr0Wpf4ZALqQIwmW4xN8N82YDyu43+ZjjE3y2qLXpv5mDlOwD
ALzcsoPC8MZsWVPcAbiR8cCEhUTgbiBA6uve04zchph+Z5ppQqMu2ay+ku1MAEYk
narBn7lILBdDpGN6luQ/5rlZ1oOHs0scfL0PB6MsSukAp+9tlKYjBte2h51hW4WH
rQxSIChUO9ZJBmGNQEmioPbyTceTa7vY36dJu2R6a4MQrvGGkCZ5QXPmk77Jd/mj
VO7ZnHjaVKX3gD9+OxXlMvkoWO1O0nWnliVjosTRJQvDBmbN+DWKrhDbECMzZBUL
tYj9DZUFzH7PWURkjmlFgVNwgdZjbD0NmrQ6Iejh1WFjzWyp4NJqErFkH1LdT3k4
gnKD6nNnDqxY4XZ5kezQtFnoPrld9TGXDY9F++tYv4NICH07yI2bJ6Ng+NlOYTSO
4/MppNXQINLaIx9JSifhjmr7Nl8IXch6p2ycWlygDi0rXQADX0U2/em04Exn1xZL
UBnFMvF+iqVORFRnqx/k1sC+QKjWjH3vOq8WMTjSII80wyLRvQtDh4uKo/v1RpDG
fMJwXXu0dIWCn8/WI2bCD/iUCJrP6Am+5MAoxe/uwQbxORhcEqFevD+oRu/9CszV
c+d47w9hGimFJx/Y9HZvBD/Bf47pczG6n+O21vylZ+8LGSOgoSPESKVBU7eVyc3v
GllgW1u/dZ3298CPKLWia+kCfzul0e+XFBw488aJazleldtzuoDpCoCv4U3/au2T
PZ8tVYSv/BwCNmHFV6I0QSLCbLqMhU8unE+zAEuIFHUid1xOjxjopcQSgcxmpRoQ
lkzxDo6WgpQopUZY7/1NMHmPcHoxD9ofeH3D/L99FAkTlUdQAu7++kbsBDpx5AmH
oGiXqeSq/C11tEyGe/YQ96uxJcrv+7T8nGapa0/2abfA81osVKsg2Y8RbHk5l1LE
cU67mYXI3aTyfBPG4VwIA7pAlmbEeUVyA6tv+/vL9wAhu/y5bjOHkNDqjCRds4VK
H8dkkovOOoHgPHgk9bjns1glKWgVly7ErpiAzjCO2RGcL0e8iKwf/msTKdB0m5Mj
bDtA4cbYLRUvmCaaTRAK/hko9MnwtVYEyLqiLw+H+Fv6pDKioyVUl28Wp9ssqOYU
TJFtV7NAagMXonPJSmmQTH8w9GlW20fVGRV83Nn8ZTcE4ObDHlDTSZJRtnbQjb+T
SW0s+xguyeKfp3mmIQTCmdzOmAwkuZTHtwcT9ThEMpFvTkk8bNK2d9BjMcIbcVO5
/sG0ig1EqutYZltlOm6V2ggvfG2uSiuSifz8ht6Ew8iLujL43rWCK5pU4zEMHCA3
jsepHsw2ebGpT9S0jecdUHuFv88C5Kuftxv7Y65X78HMfpO3gqRKUBjockT8anu3
JkC4DRFGE8rKV6v5pVHDmqRpaJR/MLil0nQZ1R/uW66xWy17c8uoxqKQ9lJJWbW/
6wHxlakGDYslOklnf0r7b7Qt/IZ6GMyj624/mA6nIZ4ZVQJTgVKGinWXLKNwEmIJ
fzxpJXTwGwIJ9K6XjgQhedinsnQRc3xHFs6vHQ2EcnoMlUeIxra/8xJN8uuR1Yre
wqBMV8C8EgumqTXBK4lB31efXcAEUNzc8re0/hpXFT0lutLFQxm9O80CSX4LVVu9
d+S6RkoYZBxMLmpi+3Tsq6SI4vx1VSvam6Dwau974hY72p3XP/1139/kf7ppB9Hy
IthaaALDjkmNGFoWta9XfLVJwxPgRD5ehb0XF+BLtZa2ASJLIH6uBQ2gYBklO+is
8T3TF36a4uScV8/iSbc+hlr4DAeI13SEOYZFRlpehEv/YpaeZcWwvNILyfZHszFA
Wrj2PmpIO7jUC+m/waz0MUrOU0MCft82Hs3/oRMLMgeBKPXrT4CErivwG47oy9l4
FMwlNJheUEFslUgFK3HyrKS55/D11LtRCwTA1A993UvE4DESED05uml7MdkRB/9/
GfZAH9sXQNUOigMrt9Sl8SzhUJJi0FSOb/voFsIFTvddnmB7g+w6TcYq95gcQoa5
zEPvcHOPyM4g+ZjalRWL2M5YrtMEPiFrOlszTFXmhHanAaFgDWAiuMjyrAsEgss8
X49b6b7MhsRtDawU4zQAkeKRunRbe3HSIjdh+JHhvzOE3l+5/1iTQdnY+1B4GRcD
vQCqF8zP5Y5Ex5Bo+hUwi4zOcNInG+D8hjel3Y8+ZNjCEhOyaw+WSJvWEaPzWlBD
jZqGbh19upbYip9vtB5BN0UfUrBsE5bgzKLZi22HwWrgJ27nW7oHCJwajR8ycQiq
7U8qM7ng2NF9vjZk1wwqvefoVCdIl1oRK3bylRH8eOhlwWZcnMGSU3uPsQlGE+tA
lrjTR6Es5J+CFaSjKnSbkmuLFsNFLIFS/nchxmvchE7NwrvEsVdh1vReVfGH0iLx
psTObugkRnmgYJLmH4zhRXJX3Y5wE5yxQowN7jGLlslTHkkkXcCZDbCWT+WCjI7y
LSHfw8Y0x3AEsYtm90UyqvA5ZMaNAXPYW50bIutNRWzCPbB1LMoxmdBHReGJeQCI
ioz8t1VxdR7yY9FBI+D3OlrCsO8/f2Jmc5+4ez0WyFrqmmhXavjB1QQV6Kfq3GB3
YY/uk73XiuX2yE594God3Uj0Wc2K3sHjJaCsbtUSpENTXhFzPFY6H3C7Qm5ANTvZ
Dsv1mQbQdyqtySXIbIiQE4JmIOVddyP0Vtrg8Pk8GNWegugEu/CfWLaBlS90UwMx
PewrCGOYOOsAMl7Q/DVvIPUbslW/S0L1nsdm2ANReCR3q0+1P1zafbAto3+wSzdB
1G0JsIHp4Ap8tXrEQBgF3sFT88nmqqUnl3taED83D+19b52q3M+S8YQFcEavXwSR
xBvFiIs9KXqvcarmKsHPPg6G/TvSzEZgd408s+d4l5qxdwDLOzx1A2NsCDd4vz2V
3JuHeiLyRhm4ibibeDrE8X4Zv/Oqt1UsokabI0LvazOsD2UdPM9KwGeVWiejHfUl
2zvp4idd/++P8icCNupd4tuy6UH47gkBmfnhZm3iCTAgnDkMjnrJCExLLjvhtXI4
NwnBdNs/+7E/dxE/beo+8LcEfUO3ImEZxal74YVwQvnS2NcDZ67dxMX21DbL7hP2
Wu72EqSDd+BPC80EL9bwfGhiqNAowLyvZPIP3J4QWdqUsCcHygV+oukZYiSb7jBK
f1uDhjUA/roQvpPx0bILPo/ofyfdfIDW96LIdT6UwtbvcP7mLL0yxvdVr1/w0tIh
c6xIHeKI9gWGWiNjMIkVR0R0eARfHk6Wp+8qIXbIBNLh4KxEJjK/QHMP0s0FQh7o
eLsY2L6TPuJQtMtPejXNeHiyV7nqGE47wgHo3+YFlFRsHqe3dyn9FOusFVTPyiSV
c3nZtfACSh0t0R4nE/wR8gJZaEzS4X3M7um3vTqB3JceTxMjm9HaHyVK1VLYN4Nt
YYbb7+YLhTRkhVPleU7//YCQ71TqdiHRLUQBpWth/Oy09AFdVZqtnKQCKoMSGDTo
z4vKOcwOM4oP0TJc9Y+IvM+xOboId4OQNlFTjrwRdxZ8Ff9UpVW8ZtsWwrHE0ELl
omXE6zrb9J9SYh/kH+F9njnDzzZCxso2abUiKQlbM0vjQDVzmGhuliAIKCMI3Moc
vvCj5Tn/W85W2VyKtzLZffrXCy1u+4MLdiD0tParqibUwqMV9vfemcrier3Vs8O4
+xu3N0vTosidQHJM+9ktE8oX/eNixiY6duKoXWEtZs6JZzqqdGpWtl+IQx0Ze3u5
lI2TnUlkKwxpRhFNoFmSr07Jhnxzqx7TSJfaf9k89tOTEKrGZNvexl13bOt36yuW
yQPrXelyZ/qmTb1JOsxMPtkNCtYvDNtia7Ka7RhdxaDB3F6eIkvc21HnUDJT7nPw
+srklKW6dHyQRZ//X/M1rFal0W8s5RnFE2Vz3AD7C8NfRzoJ45pG6EWPOrzqx4pa
fz5weIgODxP8mz/Lfnn7zzCnTip9wqnDHg2Q7xHGEJwCX8eHcdq4yWAjBY4aLUqG
9Ljsof6XBtUuyBerLUaxYUwdsJfYJNSHS6g0XjgeiT2myglYjKUmeD5kwSt1iLfB
yp8Ji9QI0kxRtj9ubiCijk5EZzVgUbIliwOHNBuEIAZdcxtbXhhaJpPiVv0VLhaq
nB/4ga2tDIhEq1WWsleBdLzoofHmoKoHaGv3YlO2DQr7aiZ2iXST4G/rTsYXA/be
gvXpU7fca9sgOi2KnBeeWNmXr4w9ynGYWm+ks2loG2Jm/9bTU9yMNdEDZ5uyWevE
a1G7ec1mVJiWRvfOdze0N6tDZmxUl5tMjuICqeucFTVpRqdcdMka2Q7unuaOQcd0
KWFJ9naLXFy1+1CjuDUp0rw/lT3tJBQOxinoB2p/Eq8v1uEFLWyPSsRM7IijcxxT
Vze/VV1A1NQRLyfoG1KrHtNUKctwy72kzMKrU7Jq96Efi/V2pDmqtS+ozW5dYwII
Myz/jSPawZniGWerb0Ivj7uy+kP28RmCTxpa/iKh/q1nh0kKlmTDjosEq3bIK1wx
kzIkLwYxrRL5cfFRn+Pq4nZF3yXP/q56KPfMsY5OWh4weruaULtqcE1UwypLIhE5
MSHc1xecjsN2yVIP1KB1LbVSPqRWHm53tgD8j85bzNH0U5jtL1sURT1JIME6aWM6
JdR0QlwQqXBa6tCYTRRcyl2qyiHuE/w5grs25pn8EJfKuvQY7EKCZpYSLhYp6vAK
WG/i0WxeAUFZmh4DzsaKTGoNuQDdalymplTLn8xb8R7mf+5d+xDgWwjqJOI/GbV+
G9FI6KKL3EiH6JlvDKYs3ZEyJRPA4xFyEgkBNRmt3wMgFLHltG7dd9nS8aCf8rDv
FtGD9WjGKLEQ3RzvUJpYYyAjOsjuNnXb2WXyivvy0NfFQdajREFMJWjldlStRzTc
bnXcEoKcNsZ5XBLUbvkIB/VU5HkgN4cqRcAhp4tcs7sELImhutuoL6VV5d8+nxjg
fkTZVXoQzgXJ+AtvidDd0fwHpGjBf1pzBS6ixbwUpGYLoMs7ddccfipBg2tC1qGe
B3IlnAj0DGrtVCmKQ0E4o0vlPmxONPMxON8J4aDT7X3PohqCi+gEjl2DBdf6h5JQ
xUag4grYBaAJnyF1Q3BEoKMoZvb8vip8nNZs6bMdO8Xf1+WLwAARL5hw5MxgeDfB
ltRsxrIrBZwdET9wxv6BjvWnrjdP6wJjvfZA/KVPi5occaqtbRZMZGdY3SU6cHVg
5hlK8TiaAPO3H68akpxBSaezm/KSyScJdzPCcbBFCJRZC6+FskCYx9BquMldJXfj
2snqqZ3iuNIjhH5XiEhFiNbrGwzBkWo2uVV1Sds8sQbKwjDdf2P/KZGncqp3IRTF
oXyTmsN2CGr7lOhBagWcjfXJRXsnInmGSFPCrvN+OCJ2un9OTk6EAD5AXaGbcuG1
6dD5pmIENQvKz3M9Mwi/UeLqKk0tJwHsesNQXncMwTVpOvI7LVZMNObIpkW50FlH
vodmanpR8BqxKxbCzHbsyAaXWrV3QZjg70yvedC5fpQqtof3C4gyIKoajlyS3sXk
6GfOZ1YEzK7DBowY1Ew2Mr9A/iMYc7G/b9rNTCEu9Nx2Lp82WqpGA5AF6TMTbnPJ
RX++n917aPO/UaM0gtvRo/vEnc5LIssIkxa2m6nCxzkdl64/UG7z7UYwmZZ3jAOB
bS1smC1TeRFz3ZT0Ablx5X+0MdA15t0WDKGnZP3pPpMr03hsPwpqfb1z0wlON2Hx
/SB5L+xcCXOb7U/o+FVB3soeDmDjLTd/nc/nlVjKSdufIE9J2kfmLPSxcOjjvTYw
Ddow4IShnECrL8t9I/7mAuEi7+gH3ci0IhUbn+doIL5AvrF4XqQqAh3tCGP+Xpxe
WOavcCbhaG0RXKs8L0kNHVTQev1H4+9TIydBhkuVXWtrQnAdIcmtkbL5FQRHZb7Q
UmUTOYzmV/EtWedrqx2M280BWnLJMbm6vhi9o1Fb7mdEc8dEAZb6NiQqAc3XVCSu
vBtgDTrBlpVZ8C1Up46paIBh76IRCuu2VVC2BHT4pTUZHl260BdtDnfofLOYBsNW
nDegZBxH1M+nKPu6Waf5ogtWL5952K0bgwvd6jOGZ0AKuzvQASQoU4/Qoj64wr8C
daxztc9dJoG/d0ydITSnPpLSZjVDbehYMZ5LZ1pnR7E4LHOBmf8A2npD6Osoj1za
wnROsQ30O+qjXts6FvkRZJcIM+SL/t7rnWgaTv+78YG219iYJl4M2DdxsQznV2Bp
87yg9hncSNYE3mb8FS74r3y8tUMwFbzbCsXlVdv5dQr+nGFZTmjPTO10Qcp89IFD
kXxw4wdBvN3xIEmS67FmrSnk2LA5CYvVS8ezEd0lGiENVM3oXurM0Epx2FE6Gce2
UPnsinHZ91bGu4q3iK5lNq+TpckZpih+IQ0+XFujIKGNjJI5H7KcfaAc6zWqnNT5
x7rgJWV9ds8+WgiVzz7w9bu260/cfzbBP4i3MlehcsKJhFqHfDCu8eYrSYKgen5q
DyV27mgRhMLod5HZocb4iBH1HxBlwgU4F2be7Zmhx078FQuY2D1vWSZJvDtvqG35
3zioJICJkcQv7e+SGZDiA3sNGcLB2GASaSoVXFQoNamvWk1Djqs2uhTJ6NPeWZLf
JE2E78rh4akC0fCRWSkmu8UGCD1bCZhMhhYOCfetJ/0ne4m4bzV0fHFTZWKVSQJH
1bJPneQHG5YeLUlrPy+pz/amT/SlQf+MW2nYrrpK5JAdccFSaqD0BMm8TvUqbFAR
TYpKG1G3czm6jWujg95guHBqMOo6e5rKcsOB0rl4yas2KFPtVmn7aAn6Ax4CuBiA
blokAZGv5kwWKFCUuxsCTy59P6Z+y75MeV0CnHpkdymIBK/YgOHz8bqckqXjanhy
TbHg6SHmJmZr8A2aKpe7+qv4QfF8izrt1u5A9nAuwonz4ximMZsu9+C1g5GZ/YK5
uv6Dn10ehJWvDg70vEBAWFyOCf4f6B6F1kCUqgM2vgm4zm6Aw6mGGnplyOg3BsAR
mz1m9J3UkCu6Z673N/Gp51MYZsaJxZP4+IHcHv1pGx5Zvk5CRQMLedYb+yu5RxXk
SQ+rH71GYd10ID7JSbtm5i7s6u7p5zYr4xyjQRYF2g2sxeUUBt0U+1MuCtzx3ky+
ypjuQQiKbGSW81dd453dyknoRO53a5LkXcaR3AM2dDpof8KjFs7RUNpHzxId8l3k
AwhKlukw65zDTmJ6eROx4uC1t98Mn4WMZL7sz9G+RB4BKUDvvpFUkH8TaPOcE5C2
miwXT6s7TFEt2EntKAheTodv5EXyruJY1OY7RudOFAsULiP6lD72UHcB1z0yIP/o
OR5ymNxck13vrgHitfRzVfr+hOXBxO/I2CODSvecM0jdtOHRRYu1KYWZtgvvbifS
d/VKCKzfntf3O7rKObbK/9U0CfwsCOaf/gf51kLwjdkzq43DxiUSAK4Nr+2Ih5q+
DmcgvtNOtQUSRfqV7BYDMwhXTuNxRZrRv3we5nIZYFwvbnbUfi4sfK8CBTXxBNzP
7GTVx9iRw2mHRn3BCYLJ3ufG8igN7Jdfo2F1/ZJdMWE/p4SoMsQxpKVWeSKsxYdz
sxdLCIbwRS7jM+D4HjU1WStDP8LXrdvvMhQUhtGJqLqZvZOXxK2NHg1rUZJoX/ua
usoPdSrJjIuCcQerO9FiBNxoETMYnfvIs3bic+upqwhBNosVtkrbAjs4AfdHeKHZ
08/e41CtUoP5iSEAxfaLKShPTId9crlEyYcVx0fBHfALoDaYgxOYP4Z902uioFQe
3TVxcKELUnFfGRRY/buYBKJVKRFgE3FWydQhsVxMFxMPkP/RpVnSBXNCB4PaQQ4N
ndUjAmK9qI6Z5LnQJVfKCnhXKGkINCCdUT0vIUrDGmRYBwCTC8t6J3hWbGMwLUF+
g93ZTn+SEvz8jHUf4IA181pH65hNUXmZZxYo4Qz9F1VhTlxHMCJqmCVtGljM9F0h
o/tXUpSYu2TxNTv1KvW4hFAg2c0GWb0jmnV6Jr7I3X941sUyxjpwPEfYyyYckK4P
syehKgWLbYH6BBdK6EjPmAw0WqQWyCPoy+PLneci/A5LBjGwJHG0Uq9h74nvTzu4
HOnyVsJcRviWAKq+jm+s5bOHAxLJnUajFf0OqtpoHKFuZX9YtZC6UpZhhiF7VlsB
Wrs42w+Nvwa5okg6GUM8UtmgT278bLUd9ENzd13HpwIln5xfYEn6g2xwib3VQ47b
jaHBOVW+snG0ZdtbjAkiiA1E/v6uUdy4iEevN53Oi1lNy8slEoXZ+McUyULV5lOl
u8MSGTYDwdZsUSaJ62+9AH1H0jr2jUWv3cOWCD1b38I/MsovMtx/dWpAe3sDWeuW
WcqP2aF3Vk3/+pYhdvjjpvAfaIcz6nfg/tDSgsUdwRGNHeEDVMAG0a/s20QvZYy8
kAeo4t/BPccAFA4hxUTWRFFnV6rsUQ7xjzCCXyqeKO8WcT/t48HbxEJYvQkEjcuU
nfT+GyUazj3Y9//y2EUAbVFosvjmBMkq9iZpR3fYLlSL2YxdMejxULb4sX4tEo73
lJwjuemeSLfbbXzydd3A7spFlRMtC/E9BjJXcd0hIHXOC+KaLJTi7ih4dNzwVDpV
j7iFeL/mVyGLVfEx/aKKLRREso2ohpCf0npyB844FtOh56dgkw84Wj5D8CefSHoy
beOC0Ksf5VMz2gMZDH6zAPAV4cFISWHnYDW0S6UMHRzBa5iK0/BWGCUCADnfa1vU
vp/PkuQYe+gWFDf2bYk9uMotu2VViYAF/SpmB064E6uaWo7SI/HaR6/kenxT9oFY
PPwbkqe/PWD7hb7zXz3UJA5lS+gCrhFC+2q+HfBnTXLy3Rdy4HAUpIMVpUvp4jtt
qSRy7aOvtfNHKZayP4ZBC8Ne8756Vq/rbvSZbcSNTc4d/MWfw66QvwNMPEkFCqSx
7J7SKH8yB8y2jKuSJGyJg4VqoBQ7mv239mcZXBZ+db6xoEngxiG4gvnZ3BOKYbMB
t65s0iq4tLNDiEiNi9718l2pPd4VlUsUMEeBJjNc1gVJ4Pd/3DS2COg7WUnSWK+1
Zp1317AyWitutq8zWs0S2nmXBfQqRzgQLGV5BHWXWe/siuad3pixQFHh97IcVQ5z
fdB6WzAy34dx/yqsoEBV6DA5KShRXQvSTZ509Upy1rdoyBP8d0WkXWkHieeJhBkX
A2g1+bDDx2NQbobl5x8PTfUEXPK7M0zJ3ujHU1CxodopJElt0ttkyLMg425tFm0t
lrb3ZmcGCf+uZcdXGsJrLCnHjSu/TAMRhujKsmka4d+9MSNVstmpEdSwYA2JwgMw
cqDZoiswwY76Yjinin0RHcWLCLOdOlgTxjkAIBj32PwkKBZs1osT7uXtnRM0vGVw
TOMDRRNmdgZFlqKTCq0t4W9VfZGUnIjsIvNScLTb4YiubqxHTgn8mE2ZZYk7NJfR
t7elHidbK6VyFRtSGOmP/deiimnkSNeyLPWjvq7SGOUd6oL2fBQNjUGBF7JgPjPb
+wXnBmLEu1pinhv51d+sprJirLVJOI79PgmZR6bu1/XH4LHIpRZtAglxYAbn7P8f
BdF4xot0L8J+xzcT53Su5tnmD4uJpPduDJEbSuSqSfKbeyNF8ysH9voHruBSfA0R
OnC1uhcqdIn53y4ZiNE8IElsBT0WRL8qHJd7XGj51IYK4Ak5wKs5+Til2gcFSNRu
Aj+NmlN668FFAoCxBOddiY0JyBrOg0UZAxnmNie0Tc7wluiMnx6uhm3zvT1CKx+j
M/c1V9A5o6OSUbftEcX5AdierphHOn8SGuZEoIH4m/U9Y86K/UUor7OrTldBLVBs
d5Sau1ov4ynH1Rbx+Mpc934Nqox+g3OHiHNPofZdDQ7hO7ATLIgvTWpwSyz3doUD
7AsTv6WqG2PR/uQ1mYV7zFR3EyseHGa0MZag4FQaBJl3nL1MeK/bBseZvSyndELo
p/QtsKjqILPGlVpGHiBUOkF9cFX2IxA3RgpEYeZdNIA8gXB9Q1gzFkwrD8lILYS1
kJ9ZffMQ3b87OVWBwZtiFyPJML0QG4fikfvmtZuaIhLCHm8m8cIc1ke6xiRXdlrL
NU5ney7duu2SAtSBiZTQ1spT6cbFbZFSOjXu0w2iMppcqQD8m3TuasKmeZyU7m08
kzqY95Ae+ltzBkj9RSQ3GtIqSk9w66X6T2e/+h3CbtNQ+pwhZ5wBj/to+xNfDxRh
q0X3xMnz7jp3fKmw8eijUKi3OjZzxMgAyJxbJLpNCnlw76lW7PphFhtD8touDTfq
rnqBMG7nTwSTGyNiCTCxJ1w2ngik1x78mnEue7KCgFBtQfBiwkYuonh8LZ8macrD
KfrlC1720p6Bra63HRgRWen0MC5TkzCcbMTgwocSiDeEXS+v2NS1g5aUX1psgmNZ
LCfQjTFzl8NQSnBno1EpPbuPCWgtY7PSPByQaH4Eb1hK2742bU/VHZdfUbpjnTvc
BP6UBHS4+GLGqPdI95YxrKMjkdxLdbvDV11PH2Ovmj2xVT0IYVInJDgaSPbGigk/
h0KONgXONkPSMf0bbsP1ULHQhhfqSxbyj3wOBIYQIcVem1/8k4y82PKLgt1xkfN1
RFmp9J+ynAOfLlbXCjg8hUVvoZBqhYGspgi7WZYDaxpu8h5FPUn0BgJRPjQMuP57
A6YV3I8sxnZyxEK0FlQnL/PKlRXYzKXvuR3B4m7psORUW+tqt4TK+sjB9B61Ay4n
03gHNFLccUCkrWLG7Gyd0LKeUBu/GK/EVpFVnjjZpcX+nf3RPdlWBgGGe0KJOc+u
TwWCt/wGRZd5H1SOrUZ6n48QMRxgnDpjlbo0kRjl6dYnNs6EW5RMtifWLgLz63sc
rsfHT9axptb2lU2HIYLL15CE+x6ovw7ueHVt888JCiMpyAccBduojlErqm4iVlOj
O3R/gDaIg8l5MYHfwPc2PWjZblrOXqQsoBjcWwcjsBKtvOPFdufWS3vkyye38Xvx
1BKTRyB9zAP2N5EN7iIbGwcE4456Tfh8zKFBcFcEZ2M7FD99xSauD8WRf3IId+4Q
GlfDacBlr1HxD0PWW61fZQcqJvJKs3w23t0eSMIe9zoIQ/cGFQBsZPFBu6cHwYjf
4OuIW1qvKDi324OZ7FhXHBIxcfMNoCAs7kvL1XFW+kkePF3gburR7hTMJ96JzuPV
xzO6DSQulsUBuyZscmGKjHFU/i8WoHCzNRNsjxcbuPxuIEXpoZa5YQCpiEtqxK5v
c9eyQSoO5CqXwhpVi7cI49wLhGPBlahkuft7+tLsuMfelH43JY8RTTPOMx2ZdI9D
GZmQ0kvrjfzsgPh33w/8tTvDjkMxxJDnF4g7xVQ80tYiXNT7yqLMsh7JhXavWPR1
1S0wmf7e+r8/W8Ue+/s4tl7hiawRqm5tgYZl14Z/AQLFt8PKXIeCP0ER/MP/GrU3
j0a/LO7fOpGhYl6scHXTtMA59tooa/+N79hMtNeNFR9CDmRlExmO1dQMWWHfcMU8
PUKpcEhhezo+cNfOVbMzPeHRGyonkcbVELwOqrU5+FUAFzyTCmtkytwU4DSgqKyg
IMDw9i2UcW/rmU5VLzFExO0PXJ2YNChL3ck61vhPJL3IeuzK8kgJ7ZDT1jpCL3/c
YKKH867yQA73FE0R6RkdfnCwHNYi2bRC93yr1k1Qwdr/mS3GL7xX0jWI4/mNF5JJ
E8MKX0K8T05CRHDicVE/y6McdRRg7eS4DlN+e8jvB5p873InbdQJlDNEgNepG7vh
7IHKf+vFZbSZmjQzqfC/6zDFWEpRMSAPGfOVaaODcPK8YRodtEv+fMu2BIYVSqxd
NAq3ebuaJ6rXo+N/GD6K7dthPbuRNehiqY/lZl4wYunPeAhhRN7Redmzr7qdwq1P
Lqpo9nHMJ2+hKoWna5amm8Wmprdsb7ITmbzQwtVCQfO1KZeQpf5VdP+lxxVFauDS
SpSM5QcjQw55qbVXqAcSbQPUNpt14xHn1fOaGOupgi46IM3J/iJ/PPEx3aF4WBhC
5DW92GkfqbL0nBGeqlDYCRzFWrYXVxLgJfWgOJ+0snKUw4gjFs84MvNRnpEGRnNX
cGP8YR8uWHunOHbQ6S3tAD1Kx3+jEbxLmej0xcHCop/fJtlGZnHrhVme+DqSxpxN
XM00rI0kUUuKKqX+TUcZk7XxuEzH+V5B2JdojWq0BOF5z4H8eFyx03SgnLjAttBx
z/KZhah/TxFmJ9jUK2ly83zXKuMTFRrIOPjZ9+zbIGTzjx7x8xDD6FCJAvSJtME4
8aOtHJ6g3sZ/XdsGelY5X4AoOTs40yapkNYGGOUUJeWNCDhqeFk00yWxJ1FWzgU9
hCsBKrew9V7ihDBbyB86eqLGIv4CIfqLPLD4FkhK3TvJRzuIuV1LcBI1qvdfywg8
VwHNkRkgVJ97BKnSpdRp7Qlsybbf7ng0/ei2EljEMssmadtZ+C9OM8Tzc+RlOCo+
bikFvRAPaQT1BiTFA8qaJjm0pxMxq+ixue9aLWZcLY4POpFTERnTmD/XjP+KQxjd
wLhjWY5JS5djy1uCAJrOpY8JS0itu1eohV3UH8PVRQVu268Foj7x1toJf37m4FyG
979l4WniAKTPgVf1YvGaaIQGR3WzidC7aI5NnYtpu0fnJ3aMX/e6ihHCdy0GfNM0
9E/V9YNnv42C4t/wuhJpEUBeUs23T311+NLISKqH8/vWiPrk7SnhG9kEXelpo/U3
1V8vqxmNqTncCxSJTXKuGejrNXKBv9JS+sqTlmk+wtC4pEPi3t/8f5cBeAx5k3Ji
ZqBj7NTXN88frJ6KaDWLvGATkJ86D/pcOwxc9vSNZAVQ0ttCj5dY78/K0YvnuCqC
qY7ZRyculrDqYTz9Sby+bDMjL1M/mgyMGPVjyYOKlZX2+hEbsoLDUFohdDHdGwNo
U5rdoKGo9Rjhk63uQTcuW7WJbsQu9f/abTwPgxMF4u9vei7Bq1867f7MHsnluWri
dx2Sxx4MQSnlI7EOmP5+eoCoNIF8CgBBjp2ctT3Bhg/bcArqgIqO/xH2TeoIiIBP
W0UnLdk+sP1eUyj+itl++cNDNi8WXx8roQnrsGbB9s/wVi6QQ7ohj/zv7QLoAx6z
oNIT+wIH1miojMnw0t4f4D2mo+0dHYxsb+S26FpaewACLznRQuhlqSUUHyBs6Ho8
ibZzYAqBAXuDPYrnk+x4o5vC4TYnCv9pT2SR9rXI8TgGA7DNyJqW4/TQS4CY4N55
N0Rb6qqj/rwUwvyqxMujhLupyGuGEiEPix+BbEGbhh8i58mn1BVwAMiPu4pezCMh
1Pe4G5d7V+/OuL059oJc+Zln8/P6OFwfqg9YBmxT1P+8gbPnNxJtgQKeXbjz5dXT
zN+1h415yDp6Msl6fRk/PVb1SwRjsM21kCSsOl0o0tPimJvBCov83wzpOItLa+vT
tr80iyp9Zi5cv6KBytcopfgjxkYf7LDy24fb9sljNrWSqyE738a++RIlu4cG6u2G
7c1wjT0nwl9JV74pb4Np9cXJU+AvS7aGotgccrog8HICasi4WmqSYSNLphWq/4nr
aI0F6+1HqHyXzXeqj9VqSUkXjM0LwL4vbPRbP+HRoMOm1UOYoWj0heBnxmCICbBb
Q3L25Hf3VmvZrIne19Rz8RWj5Lg0QiIWLg1gcVUFUtw0FaN4LmtJs0n/8SEd7gkp
iu8jieJTKANU70R3R9UJy9NkNcNtbnANUbzJP9/pMQNAGVoNuYoKxS32da+gpdVl
rK0L43STR7N8ITU7DBzm9aLhy9afBcHj+Rtc1yGd+9a9sYL3lmJAAIAAzDhVd1NW
J5Zl7PpzVb2a/GxEHVy1aMDyNSKNaGg4JbcgSLZciWGxjnGxUWtQN8q3heaEQtOF
d51p1vbWHbQ5vFFf/iNesdbM8YaBE3/Ig+ntOV68NEqlfySM6M5jPH9NpE026lod
oKkNtMFHHqM2W3qKPVcnUINOUXK24ywNlymFRGTElmrfkb6fRGsoKHAagFAN05+M
1iLTjAncs4wOQXpDyVM/w8JesWH7X/e4mNdg3Y2B27rNM06GVopBgJY42LvFQ+L0
ABV4z76EDZygr4rpCwQ94z7KvvCfgpbN8mBhXYcgZ1TKdHbqMtlsuTGrm56saMcH
i7lGrZpPk36/zKZ5qGzWAQNt6j/7Ctprk3KDWFwtK6s9msjyADh3zBpqe8MLvFvu
3sI3oll3il5QWd8sEhL25G/bsIpbSualFEtddX9UlrV1EJpNr6GN62RMRcjQ3Ckx
zeO9tAo8DjG9G+3jPHKpZ5gSDuFjb0tUxi1G/0WONRzhgzRxW/zRTbE6DhxWbcac
b+EoIbz3PNEgtCMG/WARTve8zPg5TL3fgTgS3dN/oyA3nPK37cy3yBr1A1equ3O0
+Bv0GqVwpNyXXsyb6f/VgDQkPvt+cn/VRy177QiU5QPASTTeu/QlHCUrkDY9a2dE
lToGnuk4w5xle47TwHXNWTuts/0O63R4WAiUKYCCYH6XjqowVcUephZiqfq6TqR+
PivzyxuKSwOaD0xPY5KLTgmP20F//ODT+jPnEXmxs5JGBgsF8rDS/qXdUIzDBCju
ERMBQbtAkuKgMBxQUuKmcqvdqeAC6sAdCNGWBe07kFXyqpVNtrDuYFyZXaL4PduR
JygBE1mqmcTqiOxJOB58FaQdoD7yyjTVi9kW3jrFK84GrHTxEwDleRcTYTaDEfTj
zc9rxizVVu1PcLbjx1G2zlnlL8ZrK/t0MIhpZbznS51Wk3pa1KF52bMP/CgBagc7
tW3/7U3SjRe7UF9MPfIzlXmwQLxTD6BC6FV4feZvPAN14JyC99JTCz9VrVBMaPwD
Nf24DJvM/zBJI3nCr5HXQqJ0JAfROYIMqs0AlHY5x6L22Da3Fvw9Zee8PU3niEI2
yeWHyoMkyCATuu3MvGGZrrX7mBeuWK/yAPQmZNP241vhwpUB0lIpQOpoYiVmn05A
mlktL4eF07wYPyHeV1RBZ/DytoOZISc2O1tHV1p1obQAeKtZBOEuYh3+ZSELrVyh
l6+Q7cONRZoeDCzPuPXNWPE5INoVGTA/doI/OPdrMl1+tieu2ysZAp7FDu+izIUL
GiwqLaplXr2r80jefsfZVu7E22cPZ8n4C9lbNzDGZdD02KVvm5MSICvKFtTJCwwu
B3ri77K/A1nivfdZIkxXC9LzBnmOhlVg/e4hFo78wiy7oKSx8XWJUbQpqsQcTbi+
abL1tFMwgdBiSc4DpfdcERuvoMp8st+j/S5E0CqcgQ1ENXBzJy4dZecW3GR8HF43
Ho+8ZUhkMpbHrk3m1LC2vOAhRBx0gGesMvUiFJiZdqy1WMbH61IUuXFZk30UFqNt
aVX922iZkUz9NQE+TjQzLwLzuYgQyxeba8tZ7qKUY5cHI5YUdf/twrZFiuC84Ozy
/UrOKO8wzXJJ/K2WWKmofPjT0/6HsU+9FU8KjQKsU4vmJjxz6Yn0Xrs+ZSS3rEn7
TYe1GWxdTGNO+ZGrQThAJ6Ylph0iNu423aExC8iVjgGFDkpKNHwP2E84Q6IVgGOU
A6KOw3vqmuwkafX3j7GRQAC7v0GfQZ7W+VuCkWItyvQ6ROdmMnf7oxxmRFBXHu/U
ulpKG4sbhc4Vy4flSL93iq3g9CyEtFv4wCd7TzwaiIagYRXK9y4iQCDG/mLWyBR3
yYXr/eRKR/uPqrGL4uN9Ba89/Z5pMV1HmxQl3GxfIW+VtkeMu53XhZS6h+NDIBoC
t4A7YKzf+y1mib7JUyCjW2uERFGIB4kwWAqwwXFb53hO8SkagixWOPEKo/OseRum
dZ78xAk+4ziZx2O7+Lyjm7Hso4dlobM4XEaugqCaUjHPQgOQM4oQ6G5h2MWBtM+4
o6QlbZ003TyIS1brEtm4VR1MDpWDiMSvZ+ZodjsbD8J3EkNh8uUJaoASiyd8zw2H
j4nhDuwGhN7k2VRYVrgxdjDUXL2sE1fwuWtKoX3vQV6af62Xokl3tKNdSz6lmh5c
O1LzfUKzQj6IWRczc7lQUpJch2PXA2w8MIMfd+G97Y+m6pdBkvdF+HCL7s6iFBJX
o+EHwWsX7IEpd+hzcLoQCdGKXY5kNWTh6tDqPJDxDiM66mVaLLiJ2truW/UQ4w3i
Q+psTLZ4GMfwoiMcf5WAWI3JlQM4T+YWKS8Yp55Mpn+5E5E87Dv/+vlcTcwXxP9C
aRAvJfVzSfi/PRpbmMQnbZpQHxlStxmAHCdFa+KE+Xgxogj76UsgasT403ZENBsZ
pWyz8O82WfAHaYoDhI2/rktqXx0kZtC1G0OkBsxqXsDcXVk7oYAlOtRv7OFkzRgw
BkLG/e+pbmXX24JthSjFbYg1tsVm8Sw0Uw+XIYl93PctDMOle66IUE7HA8FmEoEO
6RaIxqvBf1MplSufmpulgmy3QiyGYUB0mRxqiahyx3hS4fkudBb4TRpLxuYDoZf3
vTj22myy4nzoihUWgItOibS8UUKmZPxYtL8EGiQ+KMo8JFkE0KlJQkL1iTuUlbei
TO/VTFZK3RjKLd+bh0ImwkIIiC1hU9EQYmEwny0nvmxZawYLdqfCWvhqb7xuQrrU
/FJ/w0CtNpyGVnYJVqmB07w2kU9p1NpAmnG/ZPjLjBinUeLN9lVptmSC0/f0L/cg
+3X9KGVa8TnvDGMk54yH2JOVbMA7hVxMykdAL65WV0LNDNWMjQSWOoCyWrK4XSg6
gdsH6+Wzkf37a7h2zdvMKveohVF6EW0U2YFcWoiH6lF6Y2J47rUMN7UQFCQixN+2
wx3VQ76yg4EYOTHIjGp6QAZuWn3/vamnF7LqBm2ix/5L644HTlL1F0BZx4Fxb/JE
AEG7pUCSmpTf9EegbQjTfXQsZHdQc56jlFKEwe+JF0tFrvDbQMSKiqciGiVz9woj
m/Eiosu76kDejs8eV8uaic/2Lt64RI7escGZ/4h7aF7UmqrvPA6U8izAAqPE1sRC
BoQxYZcrZ59BIlpcYLSlLJc5XAZJteaTJqPPmVCylIDcEnrLe4P616GBMsay+a7I
16Ql+RlmuH1RjYReumpLiz2KhGK+jEO+3URVWhp2VpzNeScLOkZCqbkEJ15OTDHP
a5AuoaJo0CjS5kiXYkVfWkf41wBVUC2FXf2IiqBxCCr8nK+R2NHHXXU3RYN0NNbr
vEAyE+JcoqTE8lEEYOVvQpRoAM9XVX6OFmm2FZPvbRr/QX122svSNXm+6biExlwi
5Bfy+FY7gcsmgYllYzrzUaysEJQu9d+fOgk1GgXjZ5RN9IA9oFtLSV6j9NO8oZ3F
ZbWiF9gRh0w+vBLXXBxgk9o4QXBemjG52mr0tOSH7ROK6hhPw+IC7J3TWewLNXDf
sF74aO2fF5bkP8SudnF19F4i54R9jXYnM1RogKWiuMngIt1y5v4Ay3UBO5Jl0CmM
lTOEDhEQkRR/O1ZYtbzu9gKRF7mDqALelCDtIooF2q0SqqkJXAlkrt+rlKyS3g9u
R+xlCWmb7DhYdXuB6mXXoMiB9P+DdIvdaaj+FlunWhwBW2DPvOUkhyuidwX9ADuD
rxSvLKpH7jkzwbp1cqWJxbzRwCDLUvNlei0UEsLLXdRicDDGE/XshFbEuv2hTke2
2VfPUHqQudynDR0a3SgNqoXHjt0EpE82jtdZeZgtH4ZQBiSQudDeHS+3Xde4OStj
tx3wuZ7Dg+14XjR3fiJrl/xEiyruuO9Iq6Ki9U7bO21zMR8q3caGUw7XjKmUxRo7
ENNVUuWj8QtH44eijBXr+xP9fZgVDgqRPcFg2iYVwChXQY8tWecC1YAn1xe7uxiN
P/AgprLW0WpLvM+1zw9Io06DSm7gb9em4TFsSEnezNQPckQKBClkEQpDJqovxl0/
+pqfObPIA84NQtxjqkzuPfCQJfyB1SF6d/FQqpMjuL0nuOCQ89rpVXSOTnYW4e5v
5adWRuy/qrVWx4HMxJAWmw1lqP3cGWLQkImSCO8SNik9dWEa1XQcwoWWcYhwx1ku
2fUEOMr764YjoDfLf5mrHgYvJ0qLyQgiSBf9MXqzIxx2BgRBJJz4D+ggSt2+iJnP
kQ41EynJ0FRy1RP8P0lxUWa1m6Kh0Ngpi38eXrld+8EV8tiMqhrIFhUaCR5djQ9a
qyo2g/Zu3r7WU7tpztux7K05OsbgVhPjxT5lrN4ms54YrM13lA6KHaPOpP5qUILN
BAWzmhhd3XsUnegmUH1NL9s3ZwOWX/wTYFz/fVdKUsKWCkSDUrv9lTgbauVL+NwP
CeRTRM3zEiHSciUsymNw6Xcfkd7ndzlkm/mA7l4kH3SZXr3qVzizBOOfsw/XIT6n
qcdxXbsTlePUSO/mO5i77sOKq4gZATmubNePbtnogFQsigldRkV5M9jW0NGs1eoK
+ZJV8lE0RnfZ+5UM1GPyvkuNaphV96MVqo8SMiW4FwWyVPHeSu/Tn/4Sgc/Rce09
V2IrxBnm0w7CJSXVq6c81EgskhZORCPKmtPw9hQyi2y/HJHY6ZxSpbFv0vfTDcOD
wkmL7bdyFYIRql2LXaeg7fZBA/BefDX6VSnjTdGRFnTqj1cKWIN6Z3Pwrjbd0dnf
8Rp50x9Zc/55tWY2oPuUiYSxwymIwvnJT4zXazkfZUnUDIX3Oe//KFj09mfF7hPZ
R3Px1fvLc7pjNwW5yOTyUNJnHJZ5KWY9O2OfuHT1JeVWSjOHpsjisPYRWe0jbvo8
Cc06aV1Yah6pIsmhuHXB2mhapsgDQIEm6/UTMcLRV9Ux5DMcjRKZnUhNAhDmFG5/
hsLxp5OOogVZ7I9DnLZsH5dGPO/mPQLOWSQCxhYP/lw5sbjHotJLZNBh7eWX6pEG
xlva7QNmJ97JvgtagoheFPXI5BC3Iez5Ks9NCozGiwpQJX8tl3CQFYFgNnTQhL7w
tNA8FeMnqzLDRLLZGGcO97neQuYEtFFnybt7YAif6u7B/NVMdmj9veHsP2qGBghJ
F4pcnvDKJR+FJkkvNaYyAQakwk2xtijS7oCv/hcHnrl5ta7xjsNNK8WGLbaLvQTa
jtlbL6SaS/0y+y8RpBHT8FTidlzECFVw/icAfJ3YuxGWBgrIwns13mMhtL74pDgD
AXD9XAAJxuP/qq9jWUasbiE1MwDLCUljYQkYarl3oOzwsrqSZ2q+AxzggeU5C/c/
BQHrIXh5WzSGMntp9VoYT7gLUYyTwx0JLr0L7qxaZiPwgMLwoPZ+uRk+k94+S9cV
MzQv/CAnq2kz8tV0KIC/PH1ldhDXhAJwvj7+KyEzD6Ap0xkdXHSsmvnDDHnbSr4F
krC8PVvvqdoAflvQDtTQRGmR3p3poP+BL7QQlCxX22ghdn9DQoygzLPWqd3RPOfm
WuTcc2B06FBuO6pMQOS0gZeEhX0b2K0diY3OwLe9nD5sqEHmxnFPx8J0BVUhpGTc
Q6fjaalgcFh1T12Jgm2tGuVG8aXsZNhFE44Qxy0OjR/kZ0TVV+S1OUBxXs7R4Eqe
iRg0PmXDzF4bABNKJuunB9Bd7yxNoIXMpltt+ddoyK5Amk8g5HSGy4qebj66F+mU
rpXieixlrEaf5Sp8ODcpB9tGFPKC3khMW39F182ESWW9DQtgjEVuAt3Zs/S+MUxW
UjL4IqjiYlx8JjS0ggeCoBZ/u7VbG43H2anyCsKgI5hnAZIh+cDeTkPVc/c7Rl1r
fmUlMEcoBbYDikE9ItBM2l+swXfuYXr+4eCH1be+3YHK2kGHov9Av/6NDOeceJbT
7Kj/o31Mg37dap6saYEsCfX05LmDcGrs+YEAifZ9EK86GHE4joSe87WOFFyxfpfJ
f9ZrW3g724dLEEvP9ultBBrNlwnqKcfn8KCVrSKo3F470D52XP2v07RxWNG94jQS
6hv5OhyMCorssa0HeJBtrTy2UwL4N8KMFG4t1rpg+EOG3esKIYMH+RiCEaMvzVxz
r5cLmDzW3xVF4Vu9jPZzmA1O/5S549TuIEB6pkpsUxXulJlsx5kw6bK8hueN7tuZ
ny0rOjqr18U2yG/KpgqKzdA7QjYZjtnTDG45tv2OZwsC3u66z+44T+GzI0CYOAO3
9CzNivrkWcDuLgCdRH4IOk6qijMKmm0yFXex4aVtDRiCB+k0lOv12XpGLoyhTZMQ
2N6FhbxNqWsWD35Q/ySgAjr//D22Fc05+ru8hFCJ81uyCBPvbeqXGUrZ39XTYxz0
fxH2765F5snQmB+xj6a+KwGVdOJdpJDX5ttF5V0bVToheDHRv19bzPh84Z/b43S6
gLuSV3AdySH57Q/sk7sbxZCfbAgFqXDFQhgXHkBVnskBGF/DhxhjcBw8ExSP9UcT
OirmV7aLwZy8LJbV45gBQLDlTjiviYeISLZ0dOuthT3hDnkjt6bVCjFesi1KWpiG
t0Ps8nLGNLZ0aI16lWyX1sfgfigsT3HDDR9FBCykV7wcTSy6C3bNYUSiIAkbFlMH
zPnkcPgcVOuO7uRzbUoGd6cubCvHHdPMpza6na3mpAnyQKsDWwK/swbLNYgJDI7B
QHm1gY/sbjxh7Ddvckhoo8GDoq0emXDL+otm5lh1idzIypZXMbRY0iq0eDZ+y63N
VnG+KOI8gVHajmKkMO37dngMUYOSDOfowBgOkwuZisf9wEQlsFAaBvzViY726lNu
mqRLVV0mify+MauxsJxiPLuomenicoz+zyrZQ/90ikWrzgWD1jTgKntyckFOLzKN
o6B5r08XRUvzSLgQDFBjCk0037wc0mMvUbbRv4a2iKCjkx4lKYFuH5r8dmAvMG2S
vpC3Gep+FKWFV23adHtW2sVOb0rqBC1E4xl9Y9ZBhU/5uGHNJT5neWdyW93aKN02
YywrB4JshqBHO1Cx1+Y58YldTKXBxTc80dBKkrcMbtqLqoYNWt7yvS7BPn4kJuku
cwxlp9Zh3aoWALgcZ+7UMO35IpmNHApvMXjavBkUiZyJo/BDF4y4huRl4x5nL1RT
DWkz4ALjVcwTVYRRpweP8kYgEGh/+NQIqTYQG7eM36lj94pwJsdCf9PpzpQebRmQ
kUOIor3h8pdxc8QQgNinUxJTuRf74pCcgjGGVzFMM0yErC/yXqAID9E706/Eq7Gh
5lZ1mCSYL2T2sBNJOvOaXAMYDnFSOG3qNLNJhcg0UyHR2DgNFQnqAATzj1xhXYCS
jgiCKXVLRONF1pcdXqlBJyrgt2Qqq/yzqS5rxhFiu2nCo/foeYovvc/tecTe3Qah
XOpUnm0AQst4hxhLvL+eKvNDWWMsl2evMeD5O+pi1ILKbKYt1bmSpcD+DttFlAWM
zM3y+0iDHHShFYlApzZ2Gno7icKOKeTYH4fBFSup+49oNk7t8Z8KLFRsQ9Jza+3j
vILZEIUlkHX+iEFIB6Mij1gbAybdJU7SlEwzhhgXhK6pzrB2NDZEjVIEjCDGYaiK
O4eeq1Cya0eO/b6ahGofh5Ej2NfzJGXYUqp6RZLJuYL5e5aGslbj0xb5Ps3ynUFF
MEwey/XOMRk4L2zXvY5bloVp/I7/XJzlb36HuICk5NIJlC9sFVcBtb1qM8yVx+aF
LltoXnDqXxqYZ08+SxHnrozAyJvz1WwfeX35vrAUngi0x5iqbTuzReMKxYRHLpso
FIfTIRcALwx1o/cuYcuzIpGGivgkxWwoka8Ij9SGuGjTQu/OxVCzpEFLDci9vMmP
CC7MihY1NfH8p0SftujofIoxrYbOuZvJDWRFq5l7k7BCR9cjDpInNO6re/by8klz
xkZljKDsUmNlZa4fWIjyapy/m7BZ4R6LP7xNO7s6VjtVt/NPuU/HmfKJMH9JH42/
SxECxlWDnhzfdL8g5RGwdKEPu47MBCPr6w/bnRw2dESCY+HcUE/KnJmYThF8MQL0
529OMKigv7ScRUJma/eDYJLDayQ1XutK5RgIOqGGxmLLyY3zez17iY7wBKW6/RT2
h++BIOhIptXcDl2+1t22VHQoOgGDo7gYhA9/5JEX7PAeuwS02J+kPuICE4g7dBZy
XHO2fBcfd0Kgwcsy3ZEE1x/uOViZJx1v6+/Nfk1+NghFfA8blBN7QgdaYT+ppiO0
BQ7fP+FJAJr97jTx3raISHPSX8QPu3BNrl2XnFpI0Pd8h8/KQBsnTunBKEMQjTPy
+rS91YgCWLLzjEXd6vITCspeFxuUC0NgCJ9y96LS8yi8h2A/QHefCSRd2Ree/ZDt
LLp5w3PlNah7hSQ9O60DHAb4Xw0D4ZjsshFiy9K/itMTIc61qbY+YX+p8aF0t5EX
1vNXhwLlj/NTTFlDy30x43NNEr9JDxsd6GGCbr+2I7GJh4uBBORJG/ntcbmxnlnQ
Z3msFYHKDItHeTP44hoKTWcUMrNRAiZKzKhNgIxESCqLtH7YbYK/VEEEAA0l0/PE
vvm7X5Z3kGGcAapH3t1m0FLoDK8AVJ5sBQA5DIsdS1oXSUF628+yAwdhxtcypNKJ
2UDyCuS01Bf5KLANdp+BtDzSSmcLbhVzq7Ix7jZT8lxJN+gC/cfWpJYvdMCyAm8v
H1sIJSFo65Mi7t36OgxKI0yc2cfJxGFuVOhnImA43iGIsYl1aJFTYQZCYcK4+7eG
JnE6az4zVpC2p+wAN6jSlL4bh5KSku+j4GTciMpPv420/wjnvo6qqui9xhWmhVkq
HexYGz3MLBaKLdEAK7hc6zyuOvADTErvdFlUsYDs2MpQej7PsPQkZ9CrX4NQ8FTP
33cXlkORG5yBqXZiyBUtB3rSfPT9I6ByRdTixhj68h+8Rfd84pICU4/yPkd608J6
UtEGHy8XZDEIUdFC9YLKznV2n8VTL77OX3bwDTDIVAy+hnEpx8+0zOkhcZTVAufX
FLZf38lMg+3zXWfmuoVeVOTgqUoMAzDVDk345mQg7JROaU8vrvB3rsH1xHdoKqYg
pC55o0yRwLcttNk1Qh/eFPJP69QQWcaXAh8oJGfUmpk6X2Pj77JD7L6pBbv7pDjS
PQ2ssS/UkxFnCcyej5bNEBehiwR189IjTgUKRq10JsYUvWwuTHR/4pMJf/v+hzil
ESoplbRLITiheW0hru4DdSdNwbna61LMZy8BAzZ5cn5EWndjDIbccor8gBVxv5ZN
UEP/WcRsGEySiu7lvplbCAtxxi2I7StwJhrhkRESv5kuhnADwcUEOL07FuOz2KqB
JRkV+SGnYw1vWcLrBMMwjoisTd2+glOAei8f6vZdsQZD/0h5VuVsFEvjwmaekQbL
k36f24rpd5MRhDBPv06qk6drI9TcdbmtWs6xuL1RHmh02VKSrlAZVLVpmuxvO7ZZ
LM5YBFCI8VdUc7rPKkOsFt1g3LT91nDYtvVV+Z6J6nFx3BkzG9Cs121vOtH1gtS7
UmR14w4ihb4YkiL/vQNIT+M7SmpoMrbWnCcDnaToVfMQJR6dWrwWFAmEL6Oi7qM/
58KSDYGYNxWLGRCpWDZUOoCht/dz/7tNvzrvImxFSrlu35tYjJoF8/exF09TGqND
ld4lHadR9hdLXE7AP+MhlpPbx4datNZeZ4k6jI75rAbfMRqTR5zkH5AOgbhZkkeI
cQ2Vp7ls+ntYz5Uz76/tI8HPvbJPstpmuhMn2TcKtMPMTCM0D0mqsqh94xNpS3l1
qfKrEDZUdj1Z/LrioBql5LAHjrTSOOG0iYeuS3tb+DemMKvaRUtsF1jB3OJJ8X0c
pWUejgT0v2IdMpJeOguDsfYx6NEB5rr1hp3DZUhG6YQgg+2ZGUBEib/OiGXucyvg
7mt89nGzVML4yKOL3ViYWU1USGf2JmF/FUOWpgdcSiTW+kwwQ1y7p0IQl4ksBWvH
gbGi2qvsJ5n/6VAiSXSHa/nR1zrcIwrY0BXYyH0x/ui91PR5dITbk6oudKEPNV8T
D8qU1c1YjN0EPDVf2ndfLaHr6JUC4pwDpGpAxX73BDZJkavKPUicj9bIHxP0DcFZ
mDl1vHCvFvvVPO+KdFooEQGkdCUN/9OBshllCNOcWJWEyuyzQI6gb6fOg7jaag+O
2uJTqkL5tDK6FLTFmrq/OjB0jtf9wwD/LwoYJJjHtZyCo1+D6pvlTwwfqADV3ai2
lCNoxHSXUYS5KUF4EBMBOsl51YLAc37qdePHyMEKT2F+MCHBFj6ulUWY0z4eGj4e
dGuPY9mQOLGwNhyl3vAw6Hw/KpmpKl+JVCAO8FCmwoemeUjLbgGVsMR8/evOAkY5
gyzKdRNow8mgRmBeW/pG+Y9R/WAunOx+WvVvCa/uxFE2zHMqudsE9vnLI2BNsrLl
TU+nyK0WeJxpVZKonID+hKH5IczacpMFt+dHLxbEquvjiNrud2uO/qRUYNzn2uzT
aUqgCglD3uYvuO86Sxx/gvDz0LqaXm7kI6GeIqgH5m3r3I2IJi1Qz2fXkVPRtoIs
aquRaMUHG20Rjie6XSK8Qnkoa3Zp2yaOp6jp82b+8j8xHoRdAgbkbBGSVimCZQqY
PqHM18qPPFb/mBEKmmqhyDCeX6Zp9nlYiWEmNX2+Yj7ohCMN86Ga3m0j/B9UtIBP
vVUVrs4xK+3LndvH35fuNJCikRqS+5kzqqGaVcMk93wmHTWl3JpCq/qi4rGYrkdn
59n6EBp8oI9iLuJ1YT5r9WyZ9on99RWYtOWW+mm2J3/1gLdBWAaAU+AJqH2+6Mkx
Vg5xUCjpaAEO19f6H8/Z617hpldrvcG8gvNIelZh5f/17m4MSdR2jZv+Vkhb0C41
iM1ZmyE8cPUMBSbJtFsdq8h/nyXJ7DJwjp2N9rDALT05Y9KCnlWjtQn6ckSYB8cr
rNhlxhLDbANQCWVxsh4yLMN+KjItg3+TweQEQfFEboCzD9gF+EKqVStDCZ4Fdy/w
Cn3VFuHBT4yxoOrs2X3KphKc0ZzHWMdKt8rsSShEtaI2EKqnozelm6yO4YMsZMHM
YlFAuEmFmPZbVrufC59c0gSCUJNZ3S0qo1y0uNxu7A070WTmd36m/bao3y3ZS1SV
GgFMnevp2OxcdVUPs+DBwiVzo85JwDhBPR/ZH5c+OmjSN7JaMolOOTspIL5TrZFl
K0y/txTf+mPJOVPLuP5602kx3KEk6vMPXzhbJY9otrJZGY6ooN5Vq58l/Unmgj9J
Y3J6pQ2WjTgosG/c0JK8Z/YVvPS59Ob19F1apVsQ45ge2bllvTWeSnsPkDymMenw
4dEDywdqyGeyTfJRY/nNhxq8+zAba/jdI6Wvkag2CqMIlrMllN+uZ5arFFkTiX6J
bk4utHiziZW8l5zfgoMuyNwKau7wvXpbSaV9qrq9+zivPD70JFrO5QAaYMhmwnk4
17NC9DRX5Tw0FL/QOZZaU6mDPznNX1Fz7V5xeGe2/Gns9MwBPQNzsJYRyc995SrZ
FgqnOXmAzA2FWqwkzMA7QPHsUCPwBJ2jOd3z6SKyU9MAW7AiIKwtSqv5gZHHpwYQ
aZiFFYtfqEBR2Ss8NWeJyFBFUbFK4I+bbZtKAavAuokhXdxXeoqT5BYxRoOiKCsp
mYvTrHQICg30fDwrQ7WPkWVRNR93lcW8IGyW0iPde8GpEgX9DU2SjM7LMeJYGGRW
RKYBWPe/gpMR/ld/HtY1aCFK5TlhT4YmFjjJdFUGEYA1jAQKmnoufGEuBDXLyX/H
5ksJ8VxNi/PiNPuAM/VnmLDlTMxvoqVqrFpg9v/OXl5618kuvu99sisjMS2vXgwk
eCJFcMEIb2dBbrS8EOuJZW1nzQJ3FRZKQ2lb4oFxx3oIs+4Hq2hulAxL8MiPlmgE
RiWZuUOtK2Gz90szxTJVMSWb0el3+iBZgqeAvNjSF5kDJMN19SabCIHMV4EXV2la
BCnGmk/UpRqkBWM+OXGCaA4gXmwsx8K5JNZbCfTXPCYQQ/cbQuJFX0YLGSNznG3y
UwKHx3bzGgdXFuSuhmNKg8zossgSk+GJ/YeVnI0xAbZKD3tXFCFf3LfSCXrSytcr
F5OVbzJKN8toAdCb+rO8rNsa8VFNq1r54z8FZ7maSDt9Fn85dIX+p56Goh6beetx
BsKLl+BIoCMDUvdc2/O8BDT45kwtN+V0qNrfrNQv7/Tm/vCIaHyjKWQAy2PNoIkZ
K6N9MlvuXaxYq38E784JMSXRQE5otE4m31dNXJhpZEfe9Qpt+BtHOo2nu+IFnmyn
z6DiREQLrzv6SRrHYwBw8cEdpI0Wp+1QWaIROBRkWvb94yInXqBWfu5Wy6XvZnPM
YH3SF9gphzNax1ADkd7iDeaVXD4pt0D1L8sBeuWBsIm1iTg9PSoFV+zBJjcIybWp
Pt++KVEoh5kCso2iqUwTWx7gXuUAIS3Msz43rXxL3zoDCzjXncLqefG9COeT25wb
zqKz0jA1Tzzk1KkuGDv+Tso/W+q0DoBfe6uA960uoNpW7vEeLtv8Bg+73qAET5u4
bFeoLGMvD0BB1EJvYCGF9eR17yBD6j8utWk6zfebRs/lyJ2ltSzSaLD1gO21jB/h
BcNbTtAljJ4npAg5u1Y9QXaN7Pe8FtoEoVkzrQI2k2JSSByJdJSNvL0YYUTn50gP
SXYBS+IidnmQCMVZcZbqies6JdJy2s9Z+wtEdCcNEJbL7hT26B2XmC/yBtLRqg1F
jygY4IM7Hd1Yeax+aEEU08GXweBYf2joYnqe7kYQOttRdHT9D0NtRwOnqzP1Ang3
/ZFw1vVNliKl7cffXhcF5EcW0KbsNvmalhoGhx361PgV3HmP/OSn/0GV9XXOeQIZ
7BE7FBAzARHXZ4LdLLlSg4eC3UnU+YEcRwSAIJTFsOf/SpNggNaFsydBxM/FEAtu
wsM3RzNf3/wRxXE4i1oDKpN0WiaknK6JcqCCkCGcNHdG3ml2ZxXLKJRJW8pElLf8
DrpJVfAVEH/GKESFIK4gMxR7HxRNpkCA1nl+VnrW1Wis45LxcXBu7cecam6quq2a
WQay/VtrnU92eHxwVKK7exvL1dzqttoFXTvP/RfRnBuAOpLYMmDcJUwxvdDfKSRm
kiHFNd8unfgPre1labG8PoIqlOgWtSOO++n+uBMc3ARyxv2sHB5b9QdMgqV6+shH
OM6ULQ8U34mIYYi0LuYBCGT9CckD5IEeXjGNikOoPHz8xEh0KLEXbm9wi/lLFQgl
UaRvkrsx4b+0SyxcoZJSFqTngGmZvgaV3rNgFufg2BSCkqt+6mrdYccj6+Y29JCd
vUwkaTgJUC25UqYqm6zZfKjbdvt+Ar3/ZvGhaZb77lT/Lif1MdvBLJTQ0kH7uUG9
UDZWs+Iri03WDvcmVGnN0oriB6xvfwbtumSvzh08EssiYuZA/OjCold55aqja9ra
vvMyHiK6vIfTG5JU10JP0kVLIgz5EH8+WjZduedAcWpY8KtV68+0OKPh5n3F3qjW
kPA2rG5gUy3vJuF2fJ53dChzjhwO3NJlpoNfw4Oxjywu2+uPZ9B1E+TPEzizwX12
0+iAsOL/7zHkVQ8KU2zIrjbeBlS1xHvowXb2YflMlLTa6Mfq91/0PeDMPTJ+RTw6
GxCHkpfl4M7FEguAZN0yHLZQHEbASUfRB2WHHStOY59LFphGeOE3x9SgNezTh2dR
9GIoYnpaThsTwpwSxQD12Fz9u0PmmZ5UPf62lvDtSn4g5inqiEtbxm2FchyFKMZI
3VdEorH9wLzB1/XRZoryTwIK0bcyGBYGlC0diWrGHZCffofZYJcZzUWs7nl3z9ju
fTJ3nlzY/7Q7GGFc0n2hvFylr/9vjeuOKgdN6NVjoZkqPbYwet7Fx3/3LBSUKQbJ
D3avC6ARYYvInqiqiUly0GdRkyMtJRhXdOQgcmx/VM00YFl0Y5wQdqkhwurE/+LL
ztUzIaOduil30juHUiZ7mdbiQGDi5EFFNB1IkOEiLAT+Iopr47MhjEquaC7brFqr
ymM0HsJrnYL3b2eNXvwJHvwalFxiY4YDCDnzS1vzqoGOUN8SuIwabb1fJPFm4OfC
CMtYOOO19MEQrYryndcImYn8MvJLqqhXXFXDcG2+H7587HXcdbtN4myqD3LVn0U4
e9UIDRCAd//FbiEoXFFtFrvX8rla3nkyYFRhJZz8mdQ/MeEfeqKWWlYAXIbyZeH9
2m3+0GSuJyGYvG9KRxYbm6nUnWihQ68+GDRLwjkhxnswubEajOTvxNTpeenzbuk9
6X7pAeqX65b6DymgM7lnWyXzIc1R3HCVekzA/L+rmn3DsiXL5gVTx/QGMFSxUSSC
LzujXp2hN8FOkCS438Fj5ZhcZWNCN7TyKw7FnaMD8Vcfd0p5hkYyymHTlLti0KSO
NrcK+La49o7nGrLJXliG9YEb8fjKl4uzJjQ906yrCbtG6YxUcYDq0UyZu3tnRLoM
P47Sga/chSGsHMx6uHgGf/LxQSxjxIwXIaRQvkfFQ4oiqrAV8f8v1G22oe+lXNqn
IjUiiWiQYPmoXMmRmu6jRxgM2yMpd90VXUj1PV5sh7gpYuUhbvayet06z2tyLbAT
jQi88Rf+Cwox41tg3eI6NjKkZTYJG0JOQxhDL24CjlgpB6tsR/bpP7BfzuzH6kaI
4o2cTmuxYT2xCPq8tvK1i8FTkne24UvafjDlNdMF8T8J1lNX7moBM8AS886EEZyn
HwOHLe7nT3doixlE3gbaD4aAO96uUcj3XfcxXN0RNBxScDgrWPU8QXCHLDPLZUlR
1M5RhTnSKKs4M5jjZYFAkOm6ezd4xvWOBkoFP24bTI+Qve7g8VqodWUOTJQ5GoPf
Fk9hJtw3hDg4N50DWVs0a0Q7lm/bDeE/9OqPsrCvq3xDS7G5GCdOluY1m+9/fD+e
v/TjX43MVH2W9ZpU3a1GQz0qwR0tpNuAJjruN049WgMvYUxS8xy0oh/ZGNqIqzbF
nirlF9lssmi1CZ2V7DUIKN4RTrtqubvQr5kH+i7HKfS+cSly0I2CmewhEXtrPh6B
Ym6j3HavW4CrE3w7sRvLmQb/+n356Ab6mK6PVr0PdxogoIjJ7NfHYUEFP7iL7GRy
rE5vq9J4ovS9iqinuxEO/RMp5G8R4XqPdLsgqpJz3PKWxy44mkqUtznG7pz1wAL6
oYKXiVonqlpzxdUuo6Zlo/pU7HMvxwuFuDVseHII5x9Rowm8mq1fx1UcmACF9WOB
Vr97kvTrT9CQn6Idw85PcAqUMCdtIel78IkO2Zb82suwwIaporaFGa1mgKk84dlY
ifDAcvyJGaEzvbJyyAdHsikAoIaJHjLLpx6saJSpu3re/FY1c/SOIPKDyYdCs/0U
m9P5tmChZMYpubuQ68kkY0twyRqMWYkCWU9kpxyBjzUUjIc+GFcW3/PpexISy1AM
DBuGHMRQzSaRFspXeL8/6aXRjWJASVmup3inMOU2XBzyEd4mkLCZAB1q15ZLb3G/
Y8/XG6NK8RJsCdD+0pLbHrzF9nw4HHgYk5BpqSsYIp/gDVjGyfadZg49TUpBilgN
uN7Y0p8LsmY6Lw5wY44YsMNkVlZC4fIEjaI8snPsRxFaM/VBJD1Yw4/zclZSS9Pb
ayLYn7V39lB7EKwSo0KpzjfeHSiQZo0T8gQkb++P2P2tbXkJytOTCkkK8cyKGZ3P
OZ9Vdsrkm0IGI/XAUfizo7N/CAnTZoxlEY94hqKUI9RuihGHVImKgjPu4TXFgKPR
9JGqhL8HLuLi5OlMeJIYfPBA1ELVyjxXDFhhieDPVtYdGshFTROy0jl+CNaLkkW6
xN3o8ODyhnQm7bEMtHc0xv36Dcq0uMWleMw8N6oGHl9MDEfzOGs5/aJskkW1xe1D
hDn4v8HxY6u+aw2n5XGac5nn5p7j/Oc8ED1UPQw4Xn7I6hLqmTFxMcPRpInW06s8
QzjZ8kNYj5SOqm6A2/CnGuSOG1oAAh/Z8XSiNUss520BWLyufD5QbjH1zaaz2bxV
8iJJdbKEFVroTEH9x78ANxeBYWAvIrWgWUoSMX1uPsm0AvAukgjBaMqhJhegsYFq
wGc03HvCeGa5BpRnoCKOA5/s8DB3ZrUTY9wpzS25coh6xLQ3/xfMFnYgPGYocQep
wFl2ORXoPANCtD9gEvkXcf7sviuhB4MLq+GkLQCfoVYHDmCYW5Df2wk0q9XBvpCp
8WJ4QOcng1hIEOvWb1RJYRvpJIHYyyHHt71oD+n1QAlGgYF3TM3RIX8gJHVk9YJc
7uEOApqDl0qYUNRbNiZt0eYpX28D/LYP2W6TNEtXO1pEs0M0byR3YGmg+DSxX+6/
YBOxtoqJ/VDp3zVjJMtZH0OwVt7OReJ+vkrVgCA2NwXqv+UUIcT8T985C1muuNpQ
GTYjhwA33qWcsjbSc7JjP6wqEvlbNTU2JMhp9BJ8fNBuOWgYrjPFb67Ait2jUYuN
/FfyvX59OasE6voyLXJ3+Rc9mQ7JBOJzsN6Gz5yE5E1mqJV8CoADVz1YCdWEMGgq
EG/COnaIkDITIzni/eEknI/VovoXJak54SgLoixGfceMGjD0tfaoEmfonNI+sTKs
WQ16R1w4DhDWc5aU0gz/k23LnOI4kt66DSgvibmqvIZSAxOhn80em3XH0KxrUtMc
8pyHP1vGNtm0hC0r0Z6Y8KDao8WCx1Y2xzW4UrHtLWVkl38qPWKVxEeeiCHKYDK6
bWX7DS7WwZhEsQyQiZ9mdJ0m4DCPjGwbVRfjyL13oJHW2P3+oGI3k7ENzVPazS+k
qCIUzItwDWoN+rMnv0FSp7NGlDO8F/3fHDtI4a/Y4+6UGv0B/c0yATHk0fUZImK6
qpvavK2E+GCN5JP9RdNwK4pTPXo24s5k9qx7rVNosKJBEs8lAr6s0l5cS6skV6ng
q/TwOV/B25C9yLAQXtk8ExHrZza9qZQ268tfU9qcOWXE1IBHnGAeA6TKAqcFRdIS
C7erGFnTFf9yi5IY/RB/mTh0ytTSPWWrOURwgEKPoN7c/zne7+rAuIRx1Sf7O9tx
YocoP3sep2WpaAwTLGy7E3Z4E0E3dGxt+msdfEjLNg8+axtywv9bICUozumDuAz7
6kNzPo6ofcFpgtu0wD0KmQ7qcOEItjPQWF5J1vXCXuQpE7mSEirwDy+wZQZAa6A/
aAnCvf12zkQovJaL4QENjzXufXpJS1aBoD44ON22Ti8OxFuUjT0io5IARIT4B0Jl
xYob+rL7osCOnNK3P4Hld8GfbYFq+8iBhZ1DNiWeVPCExsryaDNl6MlCYyiRXRGA
dBPlXG7NkizIELCIW/BwlcAYVSffGqSUa3Y0M2xOv/jd3i6C1LxYNLCL1z+/Pdop
jBu7tqEw+WIqjM+eYv3H3ihbDEs+s1o89LLOtm7z/d74NTEtL+S1QpSSPaqakBmM
NqNvyYBUQMRBnsM9cyn1J/W6yUrFLtdOEM5uudQwmFVgdwkMSVMzJbuhxB2Otsc7
prpEb43GXpDC6Uy6Va1a1bB2HzEKJLFzgoSFjkxL23bN93LovnFCi03OQEjpBwND
ujysVD7fp6o6rxDpEebxN2mdeYdnLE/Hz3Wazm20HY7E3O8V/SSRnVDNCm5K7VJy
5Ghqw7eI1GXrcy2MpyHiezRcjFhscIcs1kS50gBVH16sy34Y6ReybGwKJmVe+uDb
U7FUp26s6LHSA0d3wzP8j5OoYFMDqDEbLWwGVyVSB4Fw3fGsPeGpfUfD2fjYZSdA
sHg/2smnuGwu+kP7s5M0fhGc9zJP5rIJyvLBDhUetvfT/I0vHKQ7k07N5JHZK/Cn
XIOFCtB8fQPKjzszl6ZfJX/w0Wdy3HyddRU17+1byPc+fhIywcxOZ9g6USJznUBO
PSE9CMevXGxFooBdPilwaYW+RgPqEkwIfgFTxYOtCy1TF75ysE3t3n6lkKXZBWRW
aAnshpD+LCzM5v1Xy3fRsiW7oi3dqDO9beZENGnlsavl9F0x503dM7eMHaWDOl0n
14hWMulxLJI5biFfjCKpQeKCUmG4yUtO6sHXOwjnXMVhIQEQbnlsFHVHHGlk4/Na
XB9uCc6l6mJ+xJFJjexTOCDYaVLdHkuuQeLbBxIS/Cja9V+pinx73xT32By9fhsv
QraA243BEb87d2EG6XE/5FuGixDthNVQG7IZdnQWC850vtef4HcWXoKnpthBi29e
q8GeC80ch4zZr4OdAt8HYyf2+Nv8GFbPgHPwC/UIoHYw3Hj80iSLoJh/HMviKlJn
Mnp5eu7m5PmQHCP5ReQEXsGaMQjeJzG4/JASoLeboHIkhlWUmWR23LM8q4hdDuLN
urC/ZHzJ0qxokHfFkgLRrHRSKRIsLFnUpq9rtNdvLZwQ1akZTRuIHYkqXjMTEdPK
FQTF3BhMYIMQuuU1AqCb34VZ8sDSZ55hDJ22cOCna8iBrX3z2puU+w/yg00S4Ptp
R7iDMMitt9oXjHXxNb/uFVnmNnwZdA7j+cNUKM0Wzj682HIOHiw3vRgwfFnEpfE1
TTQB/XgF9zMj0o+QGOYte7JAhrnZbnm8dKm+nuTXLJd/me1y2pDTubSQ0uibvaIp
5DVRuhucWCuKnRSbyENlJ+Y7eYJ9SBGF4qUZL3pzL4LXaWe3RSA/+iCsyk1xr38j
0ieD/2QEXIQGjvV4yD+H8kr8d5e9eqV0JBAOrykpJ9ODsAGWoTM5cyVm1K1Wllk1
DEU/4BOeuThvZSeaM6/KT/CtS2tG7/yzeXXpRUCzoAbdXFOH+enchGrM16q74qDk
xQDoEgslSDoJ5gmkAGEprFP/vhva4iTXYuVoqiIUSQeZ9HHZ46wyOXrUdZ/6CY8R
Fh4hkzxGrhetcqZsmxNNCdbQQImTfUAhPK9b+1u+ueVgiNPI8Q1NIzAbNhGIsT++
XXfYU5SgyQMzEZpZfVL8MNx7i4ZwcKc9u3JX3Db63ke4reSysnK2o7pisgS67Yta
z9FtY+T0MJDmvqZ4YOI/NXOtytBZmN1nMliwOctUAS1a4s9SiMsedbDTuBbDEm6x
1lx5b0kfKU87ToHnEu9idvEmumIhyot9b3H5IMaN2wAT8J5Uuk5Z94FNuM6+Qhtn
3f2fQvPNB1h/GQreZKAGk9Aho5/EOD8ie2MIve9iveEMmHVpwnqKnkQOoio1+at3
BHYQtp2+0+mmi7s1onXX0DghDC3eqauC3vvhyiGBSpwhJqMUFW8IaBK4kKglbgBQ
aBW+FdRoThNguAJaGCklwKpTujPbWSaumKj1h1opgPUzVCc9SuuwhTqfLZhprC5N
3mjGJZ75OpLAfnQVn40kTB8gGY+rwA0XixxXeKe5LWLp31zUsvc8IvrXuZkBZS37
lNaAkVZbWvu0ktkiGy+huWxtlykXlrcc6l7bqU9Lgo3Aul+G4MyshGGENvWTovFQ
lFNFT/0b9809DK8sTWbDCeG+8k00pqjDP8ySuZ2djy5WW5BMMKWwgxnLluidEdnV
Y7FdJFum9x8Uyd7HegSpeiudkD/QkrlTMPfGC7u12EJcN3FnRN/M+CVLnwO7XQZB
CmPlww/FTVvZk4OvB3V6wBly1ReKvvNU6P3NQEcijdlhTehTekXTH8hnIi+btx3R
oJZQNIVMQH0Ytxgm5zbAZsgPikU6QzqrHOnZBLyCVLUc1ksaFdTpvjblchfX/Mp0
v82Tm3q2VRDYtYFYyzDjvInmZpH3dtHKZPu9w/+CXe1LuCRVHNCPI5iNTs9znIKj
g36GJ0g4siV3sU7TcAririGmG2qFfdU7HCfc1Tg1rF/BqNnkgdwhgFhc2M0RoFZr
bYif2EDSoAaWjFlDrmnumfUW6AcDOr/dl0S2vuMUyTE6QRHNhvmlsCYUSutTgDBU
0KKwcvuYbZ2Cr/2do6U5D/86tsdI5KYU48TXbhoNXeLDVTVjdw/On0VfOBNgSdg7
PhGDx1bmrGMigMk3T4Fiz4I0JHNhocYkugVAeqlm8TyMvtBCG6X8TQX3ANpWlFdT
YBU8EOT6eM4J0cVske0Dp3TzztXMC0ET1Fp7F74UCUm1gLnJ8eUeo09pJj+xnnL3
/WKk6SBlUna21Dev/T4+qNlAFk/0AZ2eB1usnI2hkV7I3MOc4xFPWXOdo8jpj/29
vT4SRmhxo5a1We+e08VX+benHiTsAIYr7dRvMtBdiPPafNQJh7BWMKdNAbPcEn/i
2O7Ko15BsKTnKaQau2RFnFJYJHaAl49d+YSqCru1wVNOZWeU4IVZUlCVUy3v9+Hw
MXatIy5SRRAQ5Bq4IMTbubpcfNHTFUw798NAcnoKRv1GU0w3EB7pnV154BavoEg4
ufB8vMzTFq2ukwR0hmTPKAAwQsRy1sQ5k15075LGb7LXU345tt2Zn+DaMsbao+WG
pcBB7ptPOVmgw5lELn34Ikqq5srHwAteNlrspHtFGqZnGGu9mBk1GBU5WnOAm1dr
AkKm89l5FflzhyeoWgx17ODb+8RLJArz4qTLrzT535ozpRUbFF5s6nMVALiQaxT7
kSqOWQ66YxQmVPV58endORNVu9G3lJyXV7yRQIPg3vAqqJIY7x8gu+QLQSWFQ4Sb
E738Gx6KX8D+Duc+oGubHk+VXGvdzChnA6s9R4jsKGL1emjZzRDLUZtnysFGmp29
SQqS9d1zBKFF8xnAf6T7AVif1unPCfsvAg/sN3dwJQO6EjafoLoGzbsVMKyucP+I
0xiRMbx2PLY8+8MV3NX0Jdm0dhkY2VttfF2pb1f2nue8UPg4XkgWZH40hgMgcj4M
gk59gnj+OOyunM37YOdx2ZgujdgCjwZb5AqzFoohtWuxEGSFuwT+V+7TwAb+KmHo
LqcIqDF4vn4JAERCFk8tEVt2zUnm+sN0OR7WDtJ11+yvTZkJSu4fgUnKp086Ee1E
BDmW3qePx5Qd5jGcB0Dxsbtaln/4IzYCzOedgTUSs0+4UByuYUgxskJLch8AVsdB
VRxiwPN6RFzLjk8tYRQFHwYaqc3hfR0oXsMflV/LAdQliYrDv8uVKKXgOOOAzEtY
3lcH0e3seDxH593pBsr3x3lgOiNubDdy7uBYfSZT0ZjzX1wsGWS+hTUb7GRcgCMg
tHW3y9cUHN6AOMCkcjmWS0DojzLQ14KLUAJA3Y4Wqet2uD42q72WPMuSBfSbOU64
qCtM57+bZ3L8Hli+V78etL8cxGdVL4E0rZ9DE0uMT1fLmpznWVa6XfhQ4JnWwz3U
cWLMdOSy5I4XPPmehZMCyB1idNWk7mx1r4u7sSmO1XSevjl8x9EQcmlAVMLwrAE/
Y6lpfMM9npsgBfLW4wZ8V11pF/oESOx2APJL0Ch2IWxqpFnyDp5dBw+FMTUjveFL
isKHWOXvcfT+T8DYgV9r0RQ8BGVKhbi4RSzLbuna0lxyWv9HS1NWKg3QiGdNDtlR
g0hUwhuVXJEs+wM/5zyTe5uFoYZPa+ydXP1Nyo+1SGGD4+QrI0MnnVEGn7ZcqPLN
ftlemFiTlvcQIcZKQzGz96WVfQuJ/+/NySReSsyfNpigc4RN0pn31icPNLJ2UvIJ
YfM2XRJum3YPMpeq9CIqNzM2dh855y01woT1V071fLjXPBL0ayaFYohJJrlh/oGo
PJv/KVgBZ1TaV1Ov/rAg5UxGXqs5pqlQ+r+O+Ph5eXrfNyFl32cU4Mxfx13LkCkI
fy4rMbWddNJ9kPfQjdIz9T/CvtKlYZfL8H5kDm6Z1IHN0SEsTgt2t6N1OKWF/B7N
VaU0SrZckIcl6th6DKNh4sKNWb6MerMx0CmRWsR063EvjnbYAAPpgk5L28EGoLdx
IcgpBk3JKhpQAnZD4zsQ6PXlsRooSKv+eF3RiQ1o70AILmhzsaRK6wszrF4MbM9Q
y7cKdYpkVbbozlqzdYfRW+s8+ytOtcuiyufRZkZyiT2dv5UlT7XL3EQnywUhWScZ
6e3bqkt0cAsdIpzDdFjzVxJglalh8s6/FAsUN7X3lGDeG9GxSIQ2tODbjIjDv3yt
TRdCYq+sj+fl0bcavm/mEMbcAURw4J9NDRS/c8m7ihljILFOS92H67vKhhv19B+4
6gOqFE+dApSQo1fADQ53NwkiXooH6M60zY6HP0yZrxnKckt0pzQ9x0rMx6QR/9uZ
sCm3AXROu2E5BPbx93DTVJX+H8t9PwVc4bcWsC5H+6cEiCjQE7qSL8drBQXWVPvc
5YGpX6AtfDarbhYBkqiILQ1z92F6xj4OuTOYHljloCQlKu1KUEuhA0FT1FGiYwkL
FX9+Vxdetyo24KWaiPVaGp0B0vFI65bGZjetg9EYh6za6m3pmKvm53C93WjdtOha
rrnOtTYo/+X5nkwCCnSRwX2DlfHlBQDUZhCT2GnXn8ok200bdL1SiphNjuWKJDys
6Ti+tVm+ht/yDIjTH4+iMovLIIzeJykca5K1pdl/d9E1p8XNIFSKNcFodXjLF5Mu
OD4T7Ke+u4t66eRSEl8zfn5PmYkIYF7LLl2xfeM3DZNNQkOcMAbltFLOsv2fjGSA
qhm4LAB3/w2cP03xGgaRSR3PR3dDiKrVR0LIcP4U+5lNYMkoGNGYADup4OtlGhKa
my2SxFvIQSYeLln7R1xiRmYExLkpYKFSIJRj7c1jFFZmc30ClOJokNJSfXZSCzbZ
q/Z4ujs/tqcHSDy0jkwbMIqFTwWzE+xRfBX/WrwbL0tfZJvTQb8kXrS8Gbd4Ub4N
hxl6eAhMRHS/PPg7oqzSiFOclik/31b5axWf3y04ELQFRxpVrirocmSmWo0bzjg8
FkUWWagACWF01+UDszcxlYSRJsGq0EJlwqcMVLDiyOSof7iA6DqegSg0agtEpcdp
7m/BgEMgU1Oew8c7ssluwIWSsK0GpnFdE6Dtow8nBkx51Max1JNDDIcANw1ZlYlD
QaClSp/s5ZI2M7pm5tbH+jAmvn4dEE4osgh950JAPxMpqEtm3LRnA7XDExEfg1Qa
hRbFP7XTVeFzDNYqioHldxB0Dawh1rQb2ysJ8MtX5iusimYah9xXmg/eu9BhE2Id
auiLf2c+XMWBqVll9fU9zMRpj53Rd6D8J2JM+zqYOh5pq+qEvvVfk/XT8lZNwePb
IKw2vcScqytE0d9sdWDkcpnns8+S4liWVydwbZK3RLqrB2iWj/QsQPuITSgGMvxN
0SixCOwxPwKy9xsJOgmFHho15WI7a+QG5sRJMzMkp6UsQNSanCCP4FcY+2ryZa/K
RXEIDDHdtVHYQ+pa+7gErqnKoUOaxMVBcT7m10BjEWP20KICOVa7jcjau1F8pNDZ
8EUk92BolSNn5Y1bYgbgIYCQH2Agkci433HXw2DT9AA+ANBewiViTvunJd8gXS63
DXYp/dzzF5BFo+OfvT2IK9h8tF3n4j2/9K9DS6H1WbfEOABoQYjNarxeA+fTXTMp
XLGcojLREoKZx57az9WArRwuY00KFgzeU1Jr+9qMe+o3EbglvW5ZewgYRzbGqV8Y
w5AOtf+0C6ZK/j8gVxmKiAo5u8q8MBj1MSf71Rh3Q7IvM5wKGlZ/4n5ZjfAo2b8A
xgGvI8R36QaP5878cyMyzk9KNZ81iF8PQFR3YJOZgt7ZJmWRz7WkMF0b3crD0FlA
q95yXnp0IUftxRGER67P2ELwgj4IXBCSsNtSwLV07OaMPHU6IzbpmZmF0kaLeVpw
KI+nfr+NL/w4WU5JcUuDGPWqCfPmBP+2r0CRakwDkdQfqCbDNo2oL8HUH0FqnOal
TSfJvgipFZ5WGcfDD7/g+Ilw+ZDWtjILE1+xSQ3H1AzpRUGaJWbAoc7z5NS7cmJl
k2psx1rGU0pqjJlPmzT1Vcu+EUmVRwoUpcZUg1joJNluG3KgC7b+6EZBjm/clj/t
eS+lNbDhfqT21xIz90VvzIWSZAxcQgD6kpwoU3lyPkhtseMlR1XTOL50hXXCApwJ
R56mV934FL+PmP47bvcJoRGWbkiSS9dSEsuXdlZmAO1IaRqPJFzqy7rS4SXosZ6W
8YK8T31/um5gvHiU1DsJbMuIkLD0r4BinuZ0oiOGyAGojnvKUchepNDEu9GiwIq3
FFYWkLTER63074NExxHwY2Rcj0WAfN92xclk/LlIGd71qabCiC9Misx1BGGTZJ2z
GTKFmJ9638dyNAxIBqGBX0BpTCc5O3ptxYxU87SBUNEBVWyFfAtkp+tduSY2oB1o
CwShL/6zfI4BPqH/f2tH4qEhr9WPZD17Jy0gJNkhaJt1IYHaL+DdMgfaDq9HpmOd
UnQPV24/mcV2Oyjexhx1Bo5gLkHOc8MWQkXoqL9+we9JMlzcv+hFIYwVY+t2E4n6
VG55uW9DJ84tkQBUadcSuO3x312NX6bYaG2w1M+++JZdGfNYOd9jM0KcCndcrH56
FrGq2Fygobq4/qKwKDcw/fiSIGAO806HFShxUKE1uk1bTqveR6b0p90Cwa0La4CQ
ozkTaaHEz+jPqmssbCRwhsqcKBKTxokCEE2TjJVJUrvDdud++7oVoDRkI900fI7e
64WKL0lTN2iwVh/A0hUwIn1e//vYxY8znSG5HqsViIUpklLxiEDyOBk0XYBvZZDS
Fxsd6FP3HIj83rLNzYhVdZ603NiTt6UaHq2m4XAOGrinfqhNCnYFfGXcdtnD53Ug
TrAsKsAEd3otH0PJDJ9CI4eRLdSjNNchl2IHqm58B24j92gb17dc8C7jeCs/VP5D
DABlwaKo27L9xadEUIo+6ZvasR7ILBNih56tVyUN/CmflX16CFlQqo0dDtPIRBgg
wWRrHmEAiycs+Ih4WCfzFUCLSLlKYdh1gTDDL8MzEhevJtgbQL6Hk/SsEIt6ma/S
xKXVjAGsqTappLxqnBQr535s7lz8i25Xwz9k/JevH8nqj4HNaerDVqdUJdh+ndZV
MwZKdQWBWGY+dkxdKrjO0nsauK/MotgFot4ObtSuwBOF/w3yes9S5Mb6MyMBH4+t
qS2REkB6sJCXlz0cypT6JoXmnEwwN1dpi5vI6V3T3Nw59a2O3gGUvdl1Q4hlKvTl
8Ai2gP01rBiTi/MibmCN0ZoOQysIyUcv/7kiHRO890t0SDhqy0qclgSVU08xWjgK
hS7Ap7oNykL2SEtWf/qIaW8N3Cl0GKmrPCT2Vf8JH5vmdgF2WYKNJjO3tBUYOEMQ
+rmpcEQW3Ld3SM3KelR+V6e4/YSANT4TByOXlYJQsJ/kGtoepS6AlLXt0vAIe3pU
WXVXNbPPVo7KR6ZZiD3Yo8+n3aW79EtOHneB14GG62A+qTbNNmFdVaBYoROq6hPU
FML6wK6MeAmIN+LqNuJ9Vhr2jpcHMeKnrVc2kHKLr1xzAFz3xUPxvSro2SaBzZzT
BTpRM63McVQPcTCM2970dOnmJFeizhAVL+piF6jbLVMv6sOg/7fKgJLM10o1hgao
ugg4nG6MUSt7F3/dzVC5AxKflldkf8ItRSuFFd2y9XCYqLOTQ4Hlz/Y+o/ngTemx
PyZ3Z+QxQEpr0gf1dwQg7Cap4AF4lvVUjxS9x6FtAOkBTYvgpgolHiVr7UG6aMf8
tV4BBEkZSZhAUOqvOMQyttkH0CxclHqjyiebBEnYeVGcVSRbXELTZbHvWPbfRJVE
ZAsoqhF5RGf37r5rH04mVFcp9v4mGNmKFZA5SqyTihctQQXA1IaMbXEDlniRqMvU
oxjnTiw6WTdu1Qh8SlnjphUzEnMyNLZWccf3XOfIVmn87MHryk8+oQJ/1d8CQWLc
/BCjYFo1bIq4tCbvEuY3ZvJxXO4NgJRwgk8BIUIuVY7HasTGW2YqIhgNS4HWuGhE
H+dwGq8AXxtoKhHyxJMtr/pg+zn+yWkgErbtMca/C6SPvwv4TbFY5mdGDrpZMzvg
Uh0w6Yj0Go+6FbTC1fIjN1A4b8aoVcwcQIGmvkGaT2KAqSfHMqKWRQuX1R2Pe/w8
pcqrzuB7iSsnCy3OUu4mv6ogI4JWkkkEWSL5524yjdbmCHON59yccYdSU+2C3U5n
2/z+3p6VR0Fwm4XzaQo1U9N5Npy4xASeEDPbb37hCA/xe/CUv9gR9D3/1Qwu4KZN
nDedJiKZKsgRhymz/YUKbAUKGFcoLOAbgEGcrDEqjhw7eouRiE8h+5Z+0u0EAOyN
kuoHLxfIfsgYenUTVUKTXGitI5bdv32KcP0qKX+NZY02pGnmDVtQkOUOCmlPguIh
qW3UeiHqkG7dL5RyloizjwR6BkXnDkT4a/E9qOOy3YXPNxTkzLeFnlK6RMtrFko8
0aBsGPBQvLNrVGR2mft7hEIMCGB6MySOlMqumlfUxEW59c5lQCDbqAsq+pto2Wpd
wUAUk3iR4Ufv3iml03GCrW28oj8lx4p4y3NRHYp0TVnYT0qSIa7Mu+x9tGwbIBlB
U9sQ7HlFnZcU5Rr3fiJAoCdwM9zDGCUUu55QtzoM8oAQQc3rJZS4ZfyV1awp15ko
kRJbxwU9ceVIMaO6Pn10blrsAXScRAjDzG+HWyIcKbBeFMI1uZLb1V7EJVnFV6hS
xkFpgPSkAwyKJx8Hn//LD2YvIT4WzFQ6tO6SocS/DwRtZSHXeVsmZ3cVncJFZmqO
MCanA2x59b9In3Ldz6qT+XKHx15WcQ/7bMZtHGSsZJhZsNKtrq/BXykTd+p1/mGL
Vyz9cBW2a85Q5lb/4SAhV1rtKASNdLRULvmFhDHIZfNyTNAk29epdqNl0tkkd5HR
SeboKumQbpE2sB7sfrrAXjHyf1+AZIBWWSKCn6InEAyhb6ueyd5qBNgayfJZenPV
ksGEALQUIR7jTxAHpGNFc8/i7guBvMidzklt2wH/ElbkcTim+qfXZPMzNlWJ67kN
zyMVOObDTbJ6srJSKAGbADAyGMA2yoQTORrd6f6wT3KD/nYdphdMpu7ggQ4yrl47
JaBjFwovP8V65EVcI/j1VHeCCKX1nW2Gcq76mh8ZQTVptoCONfiNMjd3aQien8nz
Nn9VHItaXeCUroZxhy58ZEgcfY144hMzS8aQCK15Sc3KmJ3Ic/sU+KMYDsEopDsq
54AGEXIX2rrn547u05sv6dywc/BJqIJBd5/VSjf79P8bSwM0VJfwbhx2sIRFFLH0
3PWO9xKXWtve+SkfANTJyBI7W5LRB+JOjtL/SdD1vBSxFt/2LaiwvTqfW+n5IG/B
DlaQT+iciIgUZQpAuPe9UD/GcXJXkjYQAlDLRflcFBKpgOW1DbJzdNvnImsoXpjO
zshezvuuEOj277JZy6IBbA9vVaIVOVCh977WIT03qRn68MMHQSWKzL1HR5d43gXc
JDhJ+SeI5v8EJuv+1rW8CbgyANTwxMs6jfbbFSjNBpvaNcvQjGs6KzkwO3+HejHz
9dLtWtB2Yw1IW2eHyFyDoMhkaSEBdMuKNRC59YcuZU/RgBjWTTd/gfNafpfspaSV
vCUN0zYYaq6ziXG4OxGjcou3/RGmEDMRLiPCzgaWB+H0zg9W9Nox5HrfF77kpNJn
e+Zmd+qwhrDCsLfluIGepmGfDm2FFum9HgfAa/YtYsW/eYn6f6UBDMuSRQcBDDiF
XMqrpnPhSWVnRBq+4MIhFELAvn8PhuNUFGzw9y4DQpY9XMyDahIpA6c/UCqrE8xU
6aAWLlnC2X/su6MXZplRHMIjCLLVZs6m4BEzznFc/hvPdsduacMemyTglJbV65EN
V6knPviTfryWeFI/4/U4u7FeRGVk624DTzHSkDhJFbH4/jg9isrTvfNj++84WV9m
oO+n/V4KDOQue2/OE2LuaJbkc2fD10EZJwRpDmmma0cVcAVphrx2kStsZsK5DVAw
etliqOvBFgnOeIAgaINDpaGyMaaaoXmoeE0ttyqXsHC9/QUqwFLWcynZsgisuvVV
H+txow3dYWhV5xNjH2PA14F8eppyQV9WPvS58ziCO6M3gaqis+mqK9LVKRjQPP65
0zV4Nhm/T07u2xrz6lb0/QnJuZpgkoq6lTxaxZnULbAYMIHdIR11dZGBrARafnsh
P2sA/PDhcaMgjhWXj38yAdekZoXM9Rw28HbgOBT9G0hqxAnN42wC4G8CBNHwj7bi
2L1JhwOwjvAbYb7arfqGZszz6o58C7JkBQTp1kkGURjHxKSyVbqCG2R2lHS5QNRe
Pg2/trBJ9ZUplIKsIixWgiutDyQ9VK/r5Vj8B6MGfcEq4gbVctdEOmBM9VN7aGS/
9Dyc/v0Y9wWTmoJZNRKJ9J66AGPt2KTrcXCCZffukZes0cOUWzhMJNRol/ceXZn1
TTuQdwF9QsyxWTGVGhOQFcHElJCK+dXMiYszcW0qx7tj5v7pZ3eXB+5Q5S1aY2tW
rhbID4J47MZXhdnkWawefPbCb90Cgx6bpEKQNLJJLxwDq3OzdawGF1K5UOCZfSPB
GolOkCU9x8lZ23/1tzV1eYb0yqIlUNaKh2NKkMiOZX0IcMhsgQWPsDjqtGN2PpJl
Z+zvvSDC+ZfzSzCDVHP/sxoo13JshPgq7olq7ynTccoKmRPsi+Ix2R+tk9QsYVne
y+oVUZLgmsw41J/l3ueQGiB6DuB19djwRinqkXDr6HS533tPDEl1gbxlo3Xfph06
h1BDPFiTGav6XURhyED1It8KzoH7MIdbRtWiilV9qFgCuckidfyos9vWnGmH4DV/
RQbCN75HhfxAWa6qbeKN1Uo7FXYYtzuAExQYJnk8+gK75snkb80U+OE5770xRjUZ
6bve6HEuEsxZ49kgh/UqQ0SPYslVEIauQa4M64FtD5+MkM5UatL87PgHrSs2srGh
zYAL79fnhetg8/eOOot/TuePAMzqfWO5S+vuLQoHNq9ja2MeGW6PmQ0laigmBgq8
kwx5amWL2CeP4/3ujauYZEbZsbT3ou53mfxrQPVD3mCvY5dyYyUX1X/dKo1psoqQ
Fd/jft1GbMVLSglBdGJA8fyLX25lfL9MnnQXvJMcUBTiosOHPF2HWIoheKgwaM3f
m9VfC5x/p/yS4u4R3Ekyl3ON8Ykr+cgGm1/4ubkEUmCBpJRP/VDxYdgUbwUFtbFa
8XzQ9e4woF9G3YI7FVofwE6DUZnOkrcjgAlXJSzneosQ0WSfK1oiISDppjIQmcZK
u0c9Tm2JeN8tbu0Bp0gjOpHbS0X0Ngr3kvUKqNE1vqyI4h/gtTZ0Sw/b3p+8ejDH
OxfbGv/oWrqqDBRggYC3/9DxN/nu2lXwkm63lBrXNhDQnlFhCc3QqrLtKMk8HPFX
R7nF/0R1BiaJvporro2aFMSUD5KwFVJwSyqn8iAhSwT3NolvU7mQWPljXCorbhaQ
XKagBFdJQeh5bAzXOA7KZz9OraLg0dfAGCJmbWtMuo3dYFcmgPX1lq+AW5yXeKRw
eOJjisnYsez31crrXLNJ+PR5aQMRdRk3qL+oGBTbUWFMAig3aYKa4/c063dAQPYV
Hrz2zEWNTmmILBMp02+38OH4HOELub1Nw9E+TRYBj3RKxNjY/N6pXuXoX7fBlUbb
0RQSsoYhf+pcIcAiEpfU0X6CK83UoXODHEB4XSkGiVryhXZLo18D3/wysyM3aSyp
hqhI0VHcP+qm8mQzuUKLx+HGNpJFbcYD9vRJIEnPJ1REyeJoBjpaw+2/u3ciWSkD
p1EqP7peAjCGgVLg69zeL/rctCVAkY6pOJLi/SWBhx1hSnyuIU2C02/lQ5yic82A
9qwvrkyPkfAI3ypWgdpjI5SqE3bVikb1M7wUnezdvxT/aqB6+WALauBY56m1BPdW
2joLpNVv6BZ7bs6zVC7vWUt88aKtlMc4OEz6DLDWWF+N7MfTSQf6QuH5HabgK4lY
KUXmnfRG9jf26CCTn5+ZYgQ58WSa1ZDLAGC4pu3NadNGFYhYSN4WdszQMZZVfq5c
1Tn6DMamxM6iPvnqeO3cV6rCU5DeOkDHV0m99IsUUWDU/UzD29nOb7/7dS/hYfH/
8lQuu1zYAsdN4iFGao1xeCyJINj3DxkuYW6N8dgs4G3DShwagje9+8XI04lGrr24
0yCPn/kX1uRDyD2bbypI0UWRxGBNnObgv21AJL6q/fbr/+6UAUKorxAVbIK1Zlbl
nnCFnh+vmYBwKnMV3slP8/qHNg+FoDpJusx+DRDkTEUlLDVzbEJSBBgCk5166zfj
8w6DA7HcoQ7ftqZVathmt1zMN3jD/NUB3ojuT1Vy5I0LwK30pyMDcAq0eD2Yu8n9
5bxViwxKNmGXbXuwrO75HwPrNu1hr8F8J699YWeu/vFAdfWO0/M9/kUAdr7pWwKs
GiYsdtEgIgxvnlneSSMgE/au0eKOG2+3/Ox2IQI4JdFq82EyfZQjSAieAT3gc9ss
Arjm6DpmIankdkVOuYxhYdVNgFosUMGhw258kA/fvtgkuDKrr90GiskCQ675YF3A
wBU1RUCB5Boi0FjuyrsF4fn+dBLZdnOQr6ZXIa04jd8G6Fo59jF6F7ba6gUv3Coc
KaiCfo3+1JGe6dgmVxR6iEfmuo27CGR3Erh6fGFemzJOdcQLJLzuQfJd6fH6prhr
0oYvF2q9LSBfFFcQ1D/H3x3Fxqr/G8SWTrqYd4reYk3i6Vu7mIK1dBqcEKFeaiBC
NPpxEbI0WbnKFERgaR9sH5dOQrOORH7Lvr8enDBEh08vxiDrWlogl8TKd2j468ZF
V2IF1XLeC+SdF0WBsebD9Q/JSghn56AtFPr2RlYGX+DPAoyPiH6Mb8GKwb/g0J7T
0ogzhPzc+/5eTfIXDx3+K8tz56pflJFl7ct/xdnfLp+X6TYiFhQKjMG7fLszlP8J
9xd6AqXIXpu51WzN3yKwO6COroZEjSSFqIS5S3DamIR+8hBV2dnd8z8CmQ+r+bsG
P6RcuD+8ox1Tc3t4Bx+VELrf5G8E0IBzaMvYVXirJRQquAinnzJgkcCgiU6yejkF
3R6H7SpjlZRB3GfPiBkdDRpHGqcsp8SIepxb0kjV0wm/wWjp624aqRnIRXu0YiEp
tLFAURNaQKCIGp0m8mO+AzOBUI9/4KbkNV0eVSVVzskV/xg5An3QVUX/acZxc0H2
QP5Ih7DdFXNIafnxdvAQM2fHu1CRi9096vX1XMAEUCBmZbjXMJu4KGm1lOtHQNX7
Ozw+1K0X0syQhM8nZYXz68KQoQno3Ny8eHkUxXBbD4DwjK87bpmPxctWOrGcYpib
N+QJgtfcMxTHj7TqUdJBn9DjuYuHHotx35hxr+5Q4dsIUm8yYfT1bxsO+hj6y+dR
5EnTrFjg0ooJoBTgzCOfkXFQZMKRYQ1uqumoO512gU2/zZmU09KjB5obMiodwz2O
nixmKoxKi62op74VAYhtmWQOjpcV7RLQU3gnwVDSii2pKBnU4VU7eA3LPZT6olAN
cT6BvKfBxLM6XHKwMeXLsQ/08hPz+1FnAfDSNTnq/T4nJDxdMdmsORPXUY78MFol
gJZnQyyg5p/LWWh1s9nWWtI3fBx5igN4kSgyFRu3d8EZTE85IDfuSrlK4s6JnYfw
S9uOuneZyESHjcxHhB5ZWwZcjOowo2SmfEBYPI1PNfI455dAf0z7s5iHxNPxQoBH
bv/W3sLqs1w2cW3UAjnAhBN4y8HVUtjR3OAiB+79x9QXXB1ZpS0gkPsg5LWj9vJA
uU53sDtcWSyOsu3qYKjROXB3BK43Ht7NnRgisZOMpy3xJKH2kzUPTJFa4A9e1Q8J
kNDmRkCd2DyP8w3/teDxvQc5gOhk39k3maUjJUCRF9JIW3ZRRUIZAWN4YMGStvSb
oGKX+9xuc2FZknjkY0vI9DVvwUt3TKF5bvRqtxnVbufRXZ7iko/fP/xEY4ms6cUu
6eEdVuAXztEB5KrXttO0SY0pzdVckgHotpsoOMxbY2vgddJNo6SkBKAxdGotADyS
BAENaYxlj6qIzIQskj6wMOi7PCJrsWvQxIjMAaSzmD6uaenCyH6w1B1s83ASkXRZ
/Jeml9lSRAdENsDlf+h8FM6HKMbMA8gnk1KAEvKXMGkaAiCIwpaeyEBPjc3AZc0L
7hVQw5w62Utr4MVJcJkoNn0FpzLjdrhTgirLf/x5QA2ir8u5erjzY0M7+3iyQunj
e2CUJrTrluttpg4JX7S31gYBLnHhILj9A06TmhRbLIKT8Sxr/LwJ6wt4BgLS8CFW
T0bqJ8HnoUj6P4LRSe4TDeFSF11FN9jIHg5fCdYf7G/OPqIYht5pd4KzIJnr0fYI
9+5QPXtpxkV9VlsbWu374PbnsTrSkCDubnGeexh0dFr/OSRfMOHb7NUg4c0WIj2N
v1GttIDqoDJYariWSx0MXcMlEE18a/TBWzSjsdA+QoKBX97B9msvoj7E/60i+PYa
9dg21d1zQhTgADEBJohCZaGUMvR+lB7kyajFlI/JtydJ9v0iGX3NOukXIkbqMaAZ
TF5La7E5NVbKjXc4IpzOcybl/oxxLsnbCMVyARf6Dvb8I6Q3Wt1L+tYvjPaQFyp+
Vsk2xx50FueGy94YvpLgMnEcyIoytCgnFSrO2aAnQ9Qj2SDJTaaSh6Dv2ADPxozX
/4qCAb4cc+3wV7/RiMPz/EXxi+3x+XRxAj6msLoSUejhhKb+6JEAFHJ5YgzVD35N
C0lCMoNDNkTWYi0MQ+EP9EqJ+rZ94MvjbcJijqBnz0y61BhWU/fb+X0+bsoflEI4
Lc+Wh+cDfULeU5t2SnTYndEyc9bp0309/Xj9yZlkM+Ko4Kzzf9opIe9KO05d/J+X
wgCl543n4dPN+qljQ5J1/grDLtRdB9RHaUOy7oLyWtcHoHwDMFHWkx8c7DDRUk3C
nYQ+MBOFQ9himtKGVi9ym/o8cuh8Em5BX99DERuYgYx7ofYHk9R2QGOYUep8VBFi
ubDDQi/SbSzgMoOGG2lJigfvhSrlvcY6QLf+BkOY0gsKI2q7765YMokUv95jPPj8
PnEFy986UwUklYIrUecyp39/NNpnCHIFrOlaAc27wH4fSlganpI2hMeEdBU++BSy
jysG8E78QX9D6DedQX0Prb+cdvy7AlEsBCyzfz0Hgga7bFCDYKO6AwhBIhGkWO7W
llJhPTLZl4N/dPpouWCKb9/YXaSh6H7O2QCoViBev40CeO7YoUNW+XgLjDAET0/B
qWd6FPjauEIv5f6dL9fTKK/3ZPgFtrUADLRQ9v77tgSjYZlKTuHAjtbAyG0bLUkk
d3lvH+qFxUYVK0Nsqqe51aVr13BxzsITnOYjjMFCzadhJ19hSJI5wnRrfVdPWJOm
esozhpXrs5oCQEshWjUb6wgnT5y2Dg/1YxhJKyg3Z7PFJyKOoEaVhtOApRqER/lS
sScIqLY1YW5DozS7/TImuG4fjkUPShduHhhBLsgkxu7YCA+y5xLdQcjYb8/BESpl
qK00vJ3Gw1VAZpdZ8ko0f0x/7cEtXbE+Y9dTDNmSgeVrgO+NZN+xKgzExHHvs6PX
82AdxJ4YVg4azr4f4Q6OkM884hRt3cOGvUEdkZFGUKY/hGxO2LDfyT3oq3QDXxA7
MhXV2glDWx3NMGpDChfXspN9sqD13KuDgW//lZNPdYyaF0ayK1ORFS407K/uv4c2
c/yytJ2WKPAZxDwumLZ2DXEhASpUuqwATw9uZEBZeP5FAHEfTLuYaSlK8v99BXN0
0R2uyMQbkrzt4lgemEo4LO1xap883YwFQKG7b79PZe/Sov0tyK7PqcCt/DaAvJi1
T69MG7NbA2sKTmwvvYbIF866UQB/zVigsGzetVRJvh53AOwUP2WoDOvFTkSD7F/S
TDSTWmbeDVT5R/UhTt56j2/8jpGn2dQ/XWNSFLARoPZR0wJkIxBnj0hBiuGKoCaZ
0qYDWqQnOMu76kjI5kB3hW9HBXoP+gtEb8LCsBUoj4HuQnW18QLzg1MqdTqiCHxn
0Hi2vSpSnrXAXovLTLMLO6n+OuFXGAy55rcjLjHEV3itOGjrlgoj2IDBT0smxiJp
+eOx8Rq9cUw4SrEReHRifiRPCE06Ykcvd2pKz70GlxzG4oXaqraddycc8rx2MeuF
UVNITkrih7Gu9klx/GPbwOv3cIHN0nFoxrYF6UtQUmyMDIFuge3nJXl0WBBYwt19
9gbqaDWNLOYTsqRGJeWPyU7umaewCaxqZCiOfQ1AU9Ownwr096WPTeRVyVRl4QPC
Ckog+dHml/8Z9Agz7P7er7gJ/pl3US3ry+zs0Jq3hsjDYWL1IzlRJZfCKbaCCA2V
NTR1cu6x7332bTgjyXi9rPoaabtytvCF3xKRo6SL/WGfT9ihrACi+MPk5pcW0gfI
0+//EsARmg795IrkSoxzHfoS0kLkW2BJSpaTW4UZiTDdUF1qEU/Q7vgcMEoet2Fx
PO/fIDKgCIADZ85+854I2qeJyuxvC+CMtHeYkTKvArIk/vf4sKGXQCjzvg0axJL5
waYbGFh0Ol9I0nKb35XZUQv64ItP+JXBAaLvXHRvjXm716tlpDUQ+qjR5kj8MdVn
BKJOWiGAyzLgVxawIzjekzNw21SAy2fCJ8aYoDIJe0Rxg0Tule9yvdU1UUdWm/vb
oB+DLPPuLn9CTsH6Ak4DmFdyqa0rcs9RduqsO1OiwSZJuT3oesLaCbxFc1y1AiZJ
bkp8ZNxBj56gapTWkmdzAizwoq1mvf5ZP5fUtIp/DfUBB33khu+hnBA3vPk6yQUN
5T1xE61N+rRt2EF4Hcu9NGj+LPf2H4T8SkMoRvQWTSjsJDpBUih3/vU52jKcQQTm
A0miqoiAM7IM+wFVEAQy/F45DDkfe+sdLyk8fGdrn/16mdJw1oepgIm0dWQNv/nz
7+AveWlTCR9KtWQNHWi4ub6vkyNEsXVzYoZ7CbXFP8OogHPxWxnLZVEaksJAEUCW
ws67YiGZHVK4SjLRJgElf7XWLffiGPtEjLIiHz3dWCih4kzz4aKxM4oc4jiZAuy6
+FRGGxWwR+CiXKFaCh1gzEkckMKGEMNjJiG95vBWu4hBIkzVIRAInB3YJvzGe883
m+6Md3q6miUXpPyCInHnPfPTxQYqu5T3xYiuShf2TMoEp60ArqeaPkOb1Ln7pBAn
R4iRakiVPuXNOYf4zbG51xZEQ+x5k+7pDchg4ogAEz4HVw02bJfn7k2AVFgvXhLZ
eIcxqXqOomUQR+av9VesL/yHJab06t3TrteKLEJtaO3loERFdY8ikT1ofsQWqtUt
h5nbrTqoh1hA0ihUacneTz9oHNtdERXPjoTI/ZPsHewBlR5QjzisEXH7wyJfmelG
IQ1sp5osjJkPjNdX3IO+gIBev6IS7TiEOitARwvNPONXT6kuNN47NSYa6DgYuHrV
QrTKcvNNNW2knHVYJDmkXCC71N0Z+7x3XuMjpdZk5dbSJavTASNIMhdyQ7JPUtQ7
k18/55M9UVH03vGF06ssYr0b7V5AwUcrtbH327hkHHi2PBpiPgPOQ4i9D3v3vR5v
iQQi3IX96rPxeYqXl9xaI2DRHmpj6K3+Hk/eMfHwVDKnXKY2LULofohNJBob/E8t
kGR/HMPt6qBgYoZzCBbFMRVfH9Aa8IoQv0b/ivtU0ucg9pV1pMkqKYoC6I+11ydp
WHvzM6VNnDP8GJ9qZRaddVGp4a85x4V2gNpLkPRahaOcnlb7lGN2TRSngxiB4G9S
BXI2rezpeyTAW3nVjzQcvCM+03eovKjoKi2HJpVEvmRrH/m7zUlA/KNwfO53/wy9
+vcguWvyaP1zslV0oD1r9uwhbd5NUHJIniuzgna1sOjJIPOL0/zG/8GAEXAFCNFi
9yl2bdH1zhkw12BPphfoPRdR/ReuUaMhnewyoyjOX26all7ELt97ei8ysFsAOm1l
2PdpCfBORKUbdM3usfirLbjxoHQ/ap1IchCVGyQS/3cxoGjRbSXEcIyvLOenEwj3
2CXJ2zD7/25QOhsjlWebkZ7shb0Kw64R8Mm6yRhZpg2LoKnlaiR8z0z7YhkXTQR/
bZOFnnBXMJggZkN8PlmJi0EiyiAR/XTxPoesq3ETcuoya47KCYfd4X+CVcPwnX75
RhEaoFwhc+aaL4/PIFcWKFbisjTMIlV3FjecQm/tN07Yzd9W4peQuS4ZhBqMX7S5
IqWeJ/3+50wFDS7OcVCW2IYc5z3DNB/VyNay9xPzHFQtoUVEpEdXWn+XFQw9dFnR
33TntaEWxGvJRfjD2u5hrdYiQxqG8QA86UG4hwKJVWPP72f6CtUdxvNkXo5d/gfm
k9I1ypJfc7aD/U7s9HK36aNppQaBOb3KeEQnX97Wb6Em/SI7vXfCUFGKqcItr5ap
KONzI4+SASxtXC/Q2dbsFDwhKv3ti0GsAJimb8xbF2zwbxVJ+tl6y9+gktXCsDRS
8PHhQ5QOaB5oLzpfxneBHI7E1+LXEZGcQ4fAID/J60/cDFFN8w96TIxqQUoxMbdE
Bh+8Sp2embi/r2hvetye3Nhi/b4a3FG/z8/YtYZAkiouCqqAGjussv9NRY9prcW0
nsoauYZMtx+TPQpVZqJfVWe0v1UFmRuonL6QLmhLgI4JjrEckusadAhZofWm7pUf
FkcCgBByTXEHIwWXAw5xubZFcAzMGEz6NnbgEow9VN3o3bXPX+cz7pX32NF/srNY
WUZbKbPAJ6gYCD/5ljQ8fRVF3op0nCs1k0o3vWuuSw3hko3sOmR7x4lzPrGXChdy
thbUGLlauZ33WSr1U536DhhWLh6NVAUJngAtuPqylPB5cp3vW1TwA8WOMrb+txMt
u9YZKRc7mZgS2tOtQP54Ylk0ydR8tZIF0VBbp4ENror+DowpSVjk4DOAZCSrFD5c
Iqvl08os54Y0y9SNaxjyxLWWucCZQCr0s4EgMZT0XYSIWBKkJezxU0CJSh8QHX/Q
AZs1fjFPBMNGsE2GySqmoNzl7QyU0q/1hOsozkr+R9FKw+I+aJEAczNmDwkavCd2
estScPxT4/1vp8F2DjNQViiu/vukCzuLn6G9qJLZ+KukbaEBv4QYXOWYA5ixfDBR
LCAm93dqf/lzcdNguzOI+LJWv/IEBSjg1QxtWMpOCwwwvUZzw/NACvTTC1tX07VA
GWvWBaShflyBEvAOl9cADhP0DCgoDDJo9Qhr4z8ee72y8d1vM2AxE3dbLgavWYfA
ALuL5RQW6D6MYQROLUP7FeZK//fzXHtPe1g5E5cZfaI1K0FpXp843hXLm2BmJ9BJ
E1VDwqIYD0qJ1SEqku4ZJZ50XfENUMtFv12GjYQ9dMnJI/HVOS6nFQitoZxTkvBD
rknnrBknO0k7JUKtnvDUqszGxDKJtFC1Aleo1iEiru+12loinNCFYhJWHK4bqtzn
4QTDSiRYOMvA014gLyYJlPtjGJd/6d+Lx9uEiLPGLV5aj8rh6EAdrzoi67jeOCx8
PYquUKnaPQuJ6vtyIuZF/Ela4BdedaHiJ68WO6pD4DVkQ2WXuyIjr5XGJ9w4naOJ
AYkHWc7x/RKYWh9mFVBg4u/HE4rOBAqQ+RHk1kTgtn5thKO8bBN/EEROTN7GmOAj
2D0dGGNI+BmtG473P7qRREzpAXXbyhnnuuMHZLode4qtu1NDXDd0tC/in4VmOFuN
dOVLhLoyLkC0En/8Uh36EFNZJfSLYoebD9aoK+oApzGQlBP8DrxmGOsJdhpN7Y+k
NNZwluYld9VZ1JfdKgojAnS2LRhfXZ99Q41YRrxiLbzzRDXdAAWA3Ue5k+GtmvBY
5+Bl7WLVnZ0/DZiEMm0ZC7HinaD2F4NfTj9YkMMBRNJ786Yaq09u+urxDIMfCQ7i
ytZNuLleaJjxVvWgYTeexcw2Tl8rv4zqB8WBCzene+ZLdezVjGb1g5clSFndacGl
7IQ/n4t4yAY0Ohc7dsMWG9vuK3C7WLXYSBpMRBfnJfnexuXmTzYGUc7ZrXkQCLb9
09SG5yT6+Kdu7E04+XPN3lM4Niq47c5TqbOL9S6QXXKnKlN3tRbAztQLYKRagDO+
EXR48AWEqFtt6jhoGUM7tPggpM3T+K3wmHkkCJdKvTG+nNLiDfQw20L8geQr+XsL
sfNzSLp4NLxGsrJpPHdaqFXVQUjjue4rIDSInPSQbHPlHkFK2efW2mS/gCnmjbW5
KyzR7D9Ecm5Xf0obVKxstLxcK+FSZjw1goA6NVMbRnyYbnMqFwE8PGUZF7FY9hJm
07Vf/itQI+1E/q6NiliVgnyiojC6IocbHE0WETZQAweanpxoCIZlwTYs+68AL1el
EyTdhBAXjvKEOFGW048gaCWfaGEkvqiAneh6beT9B7v/nWpnI6ruiDGtNfCY/7H7
sgx6bzx941u9w4a20RYsF8tvhFVH8uZATe02MsdYWWfa7Uitq7o8brwhyVOPL5bx
DNxdTf1Q53YMaDJzxqdoBvSX36lenuUpRbmYew/zVR2eT2/mEh9Msd+0ugLurk8q
waIbSwUXG/8D6HN27NCQdwWk1yG7LhSsO+odykpSfmzCv0+V7YT7oWJ8NV9X4KDJ
0JqztB4JmVh+LlqQV5U6bfrSXe3nrSMnOL84p9lHZeyJsvAOJkXE5eIyb91BSq8E
TTUztO7B8daWDP/9XKI7ETj9Et/WM9DmE+yWrssZaPJMP1FqoWyXoLe6XnBylOsU
fAK5NwyQtn78XzlbVr3oDCa5EL3KrqBmgNfgJhlIF2qZ7+eFWAfkILLSHP6Rfjy2
AcNxkYUUe5rp8VjM5A5G3ZRj7jJQRbHz9uj5KhynmVGADV1LRND6zlJ2su0Xn6gq
+I0tQqrqQMbj13nbBtdOhprxjqXGUwMbs0WdLBk3OBfo28evGk6gazXvBytYWR2W
gm8O3bVAWUFw1H5se3GvKNDV00QQ4NS67QQseNic3a96nuAeXnpUow1izd0prHOH
k8tE5PEXh5JmrGUhsbMiMdR4T5GxFScLVPXrkVbxZ1hgvbSB0fqCYV7rGS/7eGat
k1ztqIC9Vb3keHb5Zr42P2cmIUwFWk5Vft3qphDs0gx7iKM94ZG/YF1tSWepngpp
gOGnA7D1EWnvXWstiYiW0/Kl8cALft7xUkpCP0wM1c+1XTppxB/FiyD8DlCd8Z1a
YNUB/Fy/qqN3nZ1guz3FCEC729cuNvKuc8k+R/C+60OT3t/3WNxMaqamBeSmDoOP
fhfxjWVTBNbp+JKyBvsiJMp7GSXao85hOpuBaLltxlg/HMws8rSnNfIagGhD3bDK
udCRKrIZ3IGADgq9SJvZyEX86XVsg5npiseFtuOYcvJdvfjC+PzCkwkfzclnGjLt
gFQNdoxYig3y4wb6Hn4Siz8qVZM7hO055LJ9lvKxylAJ03mL7N3ObJVIwpj6SDvw
PY8iBxAToo5Z9fOPKhUZ8/UY/cOlcnKXo7UCQz1BmKLqlktZ2AzFeL7BfaBSd4jB
CickC1c8oJS8WfMuiieHP+JScmur3ET8DbtjpBXsV7xSWmrI+4nPUg+q5ArUrJ6Z
HE3IxeNhM43KaKEQo1c2fhZPfNCwgKgy99CyU/ADiCOBvbcFpSBOakneIN6SJts3
BcqURPZMuC8Ag2nenIWzAw0Us30+8TdeOUalIeqK7pCK4R5bnKPlzt4Han5iuhm8
aRP4mn4K9Ozph6H1GZHfcS6WNUrf1Z2JliqV42xsVBHxJ1iChCcohYIFMA7Ff/e4
jz3zy876W95NrZkywcwDEcdBSupR+v8Kr3qIFW3joAC0osUZzoqfcPkO5JIFRHXO
n4bNuWjA2B1qeEWeu+GtRjZkCgBj2xhSutunNtVbT16+eWoB7l7tTQLIXXZMX1sQ
wzwMMhZJtZUO7kZ+uhlyFmXox/1L/VdxkeK26pJDjzsbARnIciZK5uBPYBP0ORvo
IYphCkawPxpo/o8GVH8qox8tq5GkriVG26dfWrBFL866umhIeUncE7ysyish06Yr
GmJ3y0uY0Jpotw4zA+lHL8zvOTPSTjsAQEwWTiVB75ST3EIXzil7EYpTOb4C2PJL
UzVO8koImKkaVBkKO64xyWq5zKYRQTr85rrURdTaBd1mfOzZVnQizL3p1+ddb305
liYiXG8ripi+05v6csANiyKI2wfEC8xJH+Nm11qlU3Xu6ssWP6qg2Idsxdj630me
+grDCBc7yYlJgjQ/L0pIATWBgtVYe+ZOG7BFryKhU68xtrdjlPfXhvdl8fmTn4bt
1Orl0IP1AMUeMSzTfx6DR/b1XDSjvIqpMSF8iiiQkWh+L/8LRWojYiQcYTKayN6S
LloliDH9cet8qIAp3qPId51LV9GhqYgWjPNb+e+8Hfwmik7TS9qkgMhPgA/RUKts
xkknOBY8CDzu7vUTmLhgIP3cc2C2oND1FR0dd/dKJOoQ/ozln6mqo8wMzo9BgioV
zXxPYkKOE4y+ef+nFENYzvumQMGXzxLN5kMMTLCrMKbmo/bsipkenwXa7lHEd52i
BcHc3eOq3VCnYnycW/o0XECUpVW2Wb3OPcpFjcdvx0lDshIPawGOdY8LdH+EcOdS
KhqarU7m+jE2n8vPhV9wibkb2a4X446TUYC/kr6yfzKufC6tLf9KspKuUvucCxox
P+oiVyfguXtyUabHZqejSI62nBiH8drrLfp6WoFfn1P9iqc+qUQ8yLhqk8/h0sk/
iAvFolzLboIZVXOqGetWf1C94uPDTRYPxv5E5aviJrLdMb7WClEP1N06c6K3G1MO
3f1l0mB/4aKhh4S77VaGirxg69fipmR52KYidFxxgqbQTSWg6MuGcEj9U8koXQqg
pDHLWj8hupo6GxPF4EO9iKx62Dq85mZGV5QUzYfd13m0HC0ZvGuXZzurrX4tarZB
+bCOLnaWCHTFWfjTQZpMVMXlIvXSoufGg1eWvA2xWrcuE0LZRxiSno4smTQeGfIP
2i6BZ5E63BfdtdCV12f/3NPKORfJOo7rFGsuIjCl/O18l0yp6IV+CHX0xuMEj324
MEJsBDEYnJ8Hv3v/w7OJTjtgcY3zdmhaucRNJ4UoHYJHUuTqSopHgU4wNBztjVh+
OtTiY8ubiburY3t7SA+H5nRkhz3qKkaUuxObIu3hI1BO9ph0o87HP7Jw2gFj34qN
XeJdAWfg9NQClVjr+WvdKbOkmj9zxhh83tZmfd4pJ2Ld9D/cqpSVu9CCQSqE+6T1
2oMn2QFPWfKzspI6OCU0uvJG/nynV5X3W1LfYObkc2yHAzcffzwPlWOUyw5GNOGt
kOcSoluN23/xiLIi/yVAkLmYa/WQ1eXw4cMKA8HTU5UJ7e+ul0d4lQqG37TRdJqL
rEv8WwYUF2D1WuU2Ivoxu5xMagpk4Faoziqyj6/KKb6nD5+g6mONuLlcx+nblT9X
GQbKMeFuoeLFD9jZY9dkhBWoLDsSVx4vHWPGon0icegd1KvsaywEV6z750NYKgc4
tRu6pt3XecggXpCZmn7NYMhyDH3DMLXQaxdA27DWZzpamBQomlcFraOzVMQQkJXq
u+bO4K0VokjZcnVl+873NKkDbPknIzeKV48AakF7U9B/eR+RkdcnUMj9Tf2HLqim
eH37AJrc2QLAKXsnMTjWsrmOITnDy+GBv8q3yoT3T+JJ7ZJCK/rbgwdNgqQvAJwz
bwcf3E/OXtCu9duywHKnjplqYtWN12U7Ph/wPqgTAlxBGRxo7FZu10nW0uPpEgdJ
cSfXI8g5Ii2rm2O6dkPZsOi5r9sftAcra5LsX94v/bi5n0yGlUvhPW7IgbpjgN3r
TPgkbWE28KbW1SCImLXBxpHON0VuN5B0IUYVvu+rBiQ3dF6ejMQEak3/yY8267FJ
Pvo+FlvdokT+LQWU8nSeIEENzFWei791If4UEOGng4o7VgQqHwTirZYHo0FUPFrQ
3mSWRDZMtrVdv7X1rgJYHRuC5MrgMsRcG/7kwwf5KW87DOuVLsTnKEdGPVooqf3z
AaZY0bPAzdxUrvlLz4mDVWLPUryRhv43Z4A3+pSxc7YbFyeHF/wkI1MZBp/tpOFh
/fE7G71nO3WAmsfJ3IXdVSltZm2CfMvsZOnOjl+9a6QtK4XCGu5aVpx+ezzdM7xK
IB1UqcHvCWSFiv7qxMVJsY6F8mc3cuC23dLdn+c3KjV5dPN7UI2aLaNEOQijrQ+c
9rHgApUODLRQO6yl5L/pmxgufnrWlJeixVHobIFKOZ29S9uS2tApC3S2M691mGhI
ClW6T4TOTUnIt5FglbBu5AA2zNhEvCoKAf8mfDITRU5VReFu483vXIVAD+f+xnDV
NUufsj9v7JbBn85mdAO51niBNMRcLiBaMWl9tpTmPDEqr+C0VluYsivdQA6kkTqn
qFOUmIs+7pkWu1ym8ecfNgpUqa38VWfDQZH7/vnlCNFRmYK0PmUK7PDugJ4K5SCm
q5sTDYS3ofsowUXpXTIIAMTDBDfP8D4UNydcfyAxHhuF1It5iNt441W1+i0de9l+
VZ3Gm/GeuUUvWtG68Ev0vO5ZA8XIYYhdeytBhfth3w0ytUg/XmU8DtygmVv2yql9
AV0TxMNQfSOQ1O+kKDjtkg87iLLCl9n7b6BW2gBoS8rbM4VXv8SQg1o6A5RPNfho
h4OMCZ4NSxwuhI9D8zdCs9TsXyMrlCd/46pnYSRCT6M+TXOhx2qrv8pWkZbItw1a
be8Z529+qE5az5xlW8yz8UCB60JOlpOIirAv/MlLqzXufD3aQTEL4QUtAoBoKyDZ
Sh0adQJiyz3Cteg/fZhy/jcgqXCTlLlnVvpLpRC8gJVvDAp+/g74S/3mZz4+vTuo
E95q1ooHLlyey5DZPOqxiLvbMZhVApXJu0aalvJqo16r459U95Pu5/75iBz2guZ4
tNnITfihcxJA+4/CX0tsOfG1JJGFrwhrLopaOtOYMFsZGHkaD0npeQjXgZYv1Fr8
FCM78IGWgMEmUVejsPeO/QoKT4/ChX1lA4aQiuQ8zMlvsKpKKbZqijlmeQXxRQ74
veQQYOGilffzo4qu8Am57WcA0edBeuZC2lfkUrCbab7bx+ExMmW8nIDPJGnAwzAd
qcEM+CMJ4bylchfhO95rvJhYICXibRBsr1EhyktfxsWTR5QVvkwDAe+hiSnnCCdP
njkgVSZSXPcWGiW19soad9KgXqvzd6+7dYddGJ93fFAdOjRivf06QKYmwV9NhzFq
EV0CCgwWfODElJRNx0d8bAytRE6U2Bb9i4WVUOhdRsjX3dZl3tHwY0ZCiUK9nu1l
ucFrCMu/J6nPdZj/z8rRFdX4mGu63uJyNtHOsTOR115nKAah7T/f7OLO5AIuBZ/s
yjTTuQAvZtZ+pM5531aosDvAd2AtpT0oo2VFYph6lcf8Fh7MLCPC8EW9tw3ygupB
dMRl/fPW4E+mog2KVyyGA3IQ0HWTFBo89bJaGdpTZ2fyTwCpmhFYF0h76EmJ3knX
gSkC78c2s1YruyZxa8RBmY/0/BwezSB3r5JUVHilmsG9FOq7woO7mbTYhvIYVd7j
mLiOzwxNxyf0XQk0+MygQ0c1ygpF22lW6SSBOWYDfttGVPTQsvjnEuyk7FjgPIS9
5BR2ooT7VVMSUJ0xQQdei+xDCnohgpE7QhAZ6sKt+howtQewe/wEz2gtY3QYkDuA
mloo1L30lrlUW97SsEd/1wA7SJkB3uwS13D6kQw9RheY2HqY1RNr6EviLkbirKnP
LgoWI2vvQ/OsRkPANaohhQy3VJH+11zs8H5btZFncrlpYd9HLvs2fgtqAJ0eAf/+
pIoBJI6JFzvEVtC6l/9OCo57x5HFRUKmBptlsO4CS6cTyLj7zk0BmW8RgO+i3nmQ
xPn+ZB2sTHTTL3DqAzNvlRYBGTBy5p0C3d/Y7DPdlLZR+ZPU3UAPwmDe9NMb4K/9
Cvj1bcqpltJ1J15N0e5THw6JCYCEajf636v4NbLToW8u//byHVjKVkWJXtBIghOa
N8wEcFtaq/kRqwPh5ngXlJhQNFgpFEXzhX6/VYFnVNeqQJTuPATytIul808mMh9c
a5y3ygVTGFfsJ5AUW/o3rAMzerTtbaOQN6xmKvg/DA9WnW4C4JiXim+d3HKVIYCU
p/gNi8rr4esMkWDDfyBCcO6Nnod17n4bacesUVCgi1OMYS5wo7/MC1Iv9/Mx3GZz
VRweyE+B4C0DjSaUk5qxHoLWngCfDhAa58YUsSgUzw/0gsK4rO0mx4xIX0bNsxvO
uQKZsmX08WAZQKGu/1gOFKBFjgFpn7npZWtv3VUxWFPWjgh8gXjcRTiyLoKtRyU/
iPRjTIkfx5llV29F4bJTQCa23y50JnKXFXl8lZifF0TYDm1ZO5PVXn/mVjx4ou+H
BnSoN/IySjAexxS52RwioM4Ieu4hyYZYClSyklE9qVpiaxcrpIcCRy7vM3FrCN7j
61YdpWaxG2ctesaaegf32d6wSutOZPFlxPwYCQwnd534+pFrAEQ0eF5WPgpDfg5f
Q2WDfpNP4vo1Y06Ql+m90pKHM1wsv5gWCspHKwIoJeEju8+EVRaRXgnyogBtRecO
yH+5/VVUTzGBGSCHtdUn584zIMzYVUJ1DY2R2O6u1bd7Pf3LfsBDxSKFKH+aWUFc
o1NTRUjDx/OadBkGBw5p03/3ZebSwhSFIVt+bR1BkpLCqUp8xoY0R+tvraHLpf6X
eUI/8WJe+jKoiDqYsLYcJyrJz11/OhVtzn/kt4iHD23btVDfEDRkiT8Mx95IKE0v
4b/GWE5pRzVj6WmK5ZSSfWoE1JsWaEO145ynPt/syU23XdEdvPn8tH47E6EMO+A3
81WGqoe/KD+Hsw2ekl9YghHKD/lhHQl4Nf6PZSWdzrMXB6gxhCE54BlNIZaiVFY9
dto+khD+VpG4f+siDZKl2RSFLCogO8Yszfzsff+YVsrWsjSLLdxvImBF9y91qTvG
JsLQey78BQZa8ttXUEjuGyhaHCHb6GA18o7vS8q38WM3pA3LTrmZpy8q+2iwr6RR
py9UadMCaMa9rrH3atWaBeqZpCWjz1ds5PdjrxlMqEfqBi42ltWLs/ghcTh2U1OS
EZ7CCKrQygDD5pEA9ala2QMWVnzB5iUIwjZbyUnLGWdt5AViDkgU339DW8oQkH5c
fqW+lXuVJhm2UwwhP1htgg1zPaA4jwfSsmPSJCR4viDoBYWDO9QqJPUk3rHxoxF6
huEW62Ca6CF9AXCCRCH1qwLAL+9iEtISyuRqmpVstdVCNVuZHmEXl3HE6l0hSV8c
K/ttv5maluDAsy0yZhP/BEAYv/PZNC4CNIyo9CYQ2RWOBvvtQcr7VZK2p0xLq9RM
DYKV93p3BKALhSFcYxM2YGhtMj18y/fcihvE5VMjNRWH/XLwS/z7XEyJx6ioJWK3
GC/3cMbF/Ytz7AJZUzA5BReXhhSzaitv7sIt2Wgk5dXJ+f8TM14RDWM9iRssrHvV
lNhBdVUYhkbgtvsgIwEwl3rngdYJspsUbr14vDcehloMMjLyqmZAHM27fZhYKBwT
6SqNTlhH4KTz92FNCmGXqqIIgWQwUVDEKNnbrQN7m6O/BVnhpsB7yrJhsQiQHU77
ofCIwRDgjGhCKkN1H+NdJ+Mo1jXWGMcn+jJJe7iSMxmgf3KgnVYI/x2RxjlKQe2v
VLYxSVVmcTSQiz2kNAZ400vC0aBbEEmqXQxoFcahfCw7DzN/jBm+/9nY4BCaUKfE
cVX45OfdDW+IWEXZV5bxr7qgnjtiTshT5cQoRuS/e8YhQVQu0D9kZO977uO5aY7e
C76uGjwZO3ORp8PRZBbTipD5Vdr5w1SRW/2vt0UUx9yvjhgK26QN67aBukmn/rO4
tWdfRKVducxvfYyKt/LKQcgj6y7SdDIimbGSq5pdXE52B782oAC6cwEZgSwLWarK
NERHGLbzFMZdIxy389lD1v0tm+AbyyuJz2lDpIIPiiXGg2wJXsHyER1HZSKvHJs4
ACWiXAvVwUwnielcd9Nv4PFFmMnOpCV7RIh0wwDFNV1vsdL9FiEEmKHaq0ht/0Oo
45spGM3IBJXgHOKpaRA0G5OHFAyx68e7XngM9Zx5nYukFoGMhe3BKlwdFYgTfsAt
Mq82LibkvieAlL8gfo+sIUBLNKU32D3tc4HZPjTPDRJmudALymvJMmD8O3+UhL7G
Ta5ZL42V16ylSB/j/M1VJX0GSkuZKSeTPc7eaR3F+WwZGrdfQW1xybwU3FpRoz0U
19PLU+HoqnAkYZ6Xeb4WhDJglmjrjtQztDLgJiccjVj6Jp6vdGmCX4lGB+jKrq8G
Zy4ymaUyd1oGtdriG5Bzhk1pyH88EgLZe37y1pUEr8q1D1VLAyOsCvqxX8ythx+a
imFmvSvvuTnCSU/nb6JSDH8KrwFyOW7InvHRu3tZeSKWyyxW2Y0Ffibs9JLdpTP1
hXQzHFkzyoj5h1jKNMLCvEnQU57DILBqKeddsITBhsDPEzF+/KD6rCqurQ6JV4We
wkWv8L2wPj0F6v2kpwkaH3Qi6DISUhnA2bPQUIqQwe866BOPvck+xwlflHhi6sJ2
BAL6VgQuhLiEkBK7jL+oeQg2wN+nGsuPjWROwxAwrrE0Jfmny5E6b2efkeB3qwUZ
VxFTDfhlz/dFpC0Kh8Nqc1h1ywEFRPKgprsUrEInv1ZRRXCB7RtPT3v2OqOAx/0F
GdBk8GOJvWTJEMaIN4wuG1gfM1iXJq4/8ttPV5WDNwXqJG9/V9EEgi21SjuD/kq4
FRuNZzvjSi6FCAoPH4eT7LGZHTnxwTwKNHQPndYDRqUOGcaYSPS3MiIBGSQb5QXN
rDU5H8dJpQzSy59A1QK7JIy3t+8zCEapgxGz3eDfIw6UGGiYDrD9UWEjhqOovDVi
VR3S7zJjViKjXCssbp9BlZ/DoJGjslc0ZPx14T3EeuwxU64o5J8/6gHCk3ncC/8M
RKMmn657za14mxY+jkvFnp99SWjL9i3btjJgV9XfSvScJNLgLWuY65ZmP8aCWBRR
qAyLat8M39RF9ibIBNwFOrO6in96Q8yF4f08mlU3YA0sJYDWbuslALw+iHlRjZ69
XyVV931LRm6FFwWTjAW2xjlxTMNi8YARCKtzjZMsmcQ1H3IvUEZwXBjtzfVbpoN1
S5tI7+sywSOJubRIqavlgTzrFIQdFC3YysXWJ6NCXEuBfxKeD4AukWykV1iNQwh+
rVdtGMRqcVjeGPMYVaTmKgrwlAKGiF+WyIC00YQe/sn0fWf/X4hGcCUvFwyOjF4m
a/oYycxXRfkc973Wg6Dc9DTRdJ5gsIpkir5WArnNY8NzL55wBjIH4M1qUJre8oQZ
yDm93nPDVU7HFmosvLgeknDDN2DXDeerImdLJe5nDYAJKTpHYcMUSfGYYuaYfalW
nevaypAM+fTEOZ2sDGaGrtF1TEAwfOIXlX7uHHZQxR3JA3GFgodfNJEHtl++ZtKj
k50aNT2CJvEuaauK4aNc1Ai/MDNJF1ijc0iLC0L95dq6tROoeTZzk+vaAyfi3yja
lxq3RtL4lhEtidqRXVtbEEInShHSMOgqb39Jkhwgkl8zg+sKizdSavPSL4nKSKWJ
mlJL2WkNdI/CKRTZ0I+cSztDPrqYvxEU72uHgDBE8qNb3y7QqoQQwXcxezcDP0ww
kzDxYceSgxQZ0+9squ+coZl9Ih4sna7K9nqowgEQh40R2j0uSA5wDkl3q3MWdmlD
qJbcS+igQlX/pLzIs8YVVXlg7nQmk5vLCDAkJM0XM+AG3xFhpCpvIlnqvQ3JWFL2
DTzwMohD3oLGmEAxhjOrDr7TSBBJGWQCDRuRWfX10d8DNbXCO5kMn3y3xrW1Pw+7
nFuoB25T1/bPxRYUMHtTL1R6usUCChiW0pXOtlT8mNnFh7QjqhlsZPUwt73zjsBJ
FhpGm3vtdjmPTcveiQWNmlV+fjW9+rdXHL4qIQPvotSKjTpoctRr+eFeslcEsbbH
RsRM7qSs6Pza+x1+8q1/QJ4OnQYDp66dgw51iSVEI1kb5QiDeTninwwDfetWta52
wjYVkiVgrws91/w2e/nc9bv5tI/NQ8+MwswgOfBfTmzkjXq14NHg9f9ykZCmTZCm
lmUqx3ONghVCfM2wkrqc91V4SKPKprP3Fvxe7Nt1DHxE//wuBcOjo2lHGgK5PuTX
U5BZBuxcuwzcdGr9FP/ip1wclTL4wa55Vzb+gpM3Q+fW5nwRprWvTb3yGHJ1U3OC
mO0zdN87ilSB0yowbQpsst1vcYkNyIvYceS+VnAzGNbVNhz1wOIZAqOPEYYsClCY
WuOQ093fmyp9aR0/lUfRlql4lY4Iv+7EFUIPXJM4WYY0tJmOKuPgKdngL8sfh93g
dJlzOMmhDh6YOvTjwUJkMEmRnafDcLTie6wtC7i3Np+duF7kN3TnREEZ0sCFTA60
f40S54i0cXOL6MWPMmNB0thVBJKNlpzGN7Vv7TkcXiDBnrERN3nI59bGnlZtfHuw
K/eX87QYNxV8EUdBzXce92+QyldErwJVRrnUUZgJ/dBHkel2Wrflw8gRDp4lNw7B
rMydMhlYQvxJ4PFut33J2eWPnwb6RsYSdEiEwyi2saR8nnTy54sUe8HmzMtcg3BD
unJhM07G+ZBqPBCuUeKeFYcoZkuOyzqEfuwhVA1m3tJN5ba/mAbF/7D+QxuCL5TB
12h5yyxywDGsz5I0EfVGsRXtHBdtS/HMWo5lJu850FmWrb+s/cbkcvIkiiIDSYaX
TbdHnW1FTJZGDTQQN23gWGuk4Z0RkO7TWC3dibbXJNziZGN2SeY2cUAzGkMb6z29
3Fb16M6vPjcAtAEsbdlmb9FzEbMtYZX0Be2Z8PG2nQze9kigISHM1ouqHWeUWvQY
xV21DvQnHKHJmQUALuKKtgo/s24308BeCu6o0nAbKODrNbcnJQ2hgP2NMwnC3UhG
3hViZP+DMIrFzq9ksOEotQp7+hkzhMzIqD8L7wGlDOJiMeiwolgIpgMukQB+sNuw
ootCl8maJOiXs/wJI+k85DqxzODmvGbMUEtkzPHP+M6il2Vqlisrx1fLSTUg1JFG
VUheNrVFiJEmi+vpailcXG3unyY08dVQlao1cujYkia9Ljy5BqZoIBH4Nq+5GADS
xmw/afJ3hWw7oTuNowPWe639qPJb9UtF7JvCuL/dBJ2J0DkgiT9CPH/gYOs6keeu
QO9kEymwc+EDzBW8cmSMnGqlgxUH7Zke/Cp4AsJ2lGCEC4WDJFjPnr95h749z0T3
zXVCxupTx4ZCRtEL9XX4y7ZGoZznDM0MM5GL1Ms/VkMR9o+ByHrELZvL/6/0NgMy
ETh4mbO3Tr5nsAhS04bBJRzmckKgkCtjbzuggUB2uV7EPGu5ceKSDbHlztnLj66c
R7ptR2P+b5GgCmGSyzQQYXFG7qRzsvV4SVyFOBnKVDpGIOgQgkU7xtDBl9/9EBzX
GPVSzHkhlRQ99f2WT0YbBnwNgctHQkuzW4tlB/IbeaSnIKKo2V8Roo9oy3cXoM8w
fDGyIQryXuombUWE6slPlLf6Raa7peLq6QQzfESPleVYGxps1N4cZdzAhLV+YgDi
I2MB0w84Gy8Bxi5BZGa44droISnK+/gZXeGKUN/g+fMTfaqddkXgXRrbj9Sc5e36
d3mmAC4r8Gyey7uy7y96L+wbSm8ZZW6ikts9TsBGTwKX+l/IObdyhXcmLiVT8uHT
v0nMuz/3E59YoydXK4Ctcy2QBgDv1sCahi5G4b+9kZMCflKWKjC6VoddWKy7TNG2
mJytcPA7X3lFon45ooBPUDM46+79u+FW7YmLiN8gpOg9SZG42IAO815AnPpnzMyy
rdNi1mW29ayeBxcx69kfdkvnFNnf6ejCWzxIfnSU6RFU5HRPHlpZLb7QL3ZUXOqf
H8FzhjXh1USanx5VGZMN6nx9ZvWIoV26p3Tnzcw2FZNft3J18OuZ+pAvVLm0KJP9
fwS5sNGOYhJhRPjK/gYjm+pkQ/uamQNZDWOpZixY57wjgWm3k5WMUwPucCXJYhao
LHPf0skJbhPe8TcIb9xe9nrLLlPO8fW+NAijNWFoVu8kYokVOoDUltKc5PALtfTu
yDofvD7mkVqWLjwSYdSwpPSTqI4TbtLccG2fb1z3SLZptSGnC8iRzzPavHLKKDBP
u4CoAz3fXR1zE32hnHKAwJ6m89joNjFkxFP1Ac5HFfnQVB9Dqrexc0MagR3ZAWbe
5hpJ83suaMELoLAtL0zK1Sni6WW71tUJYbJ2zG7HzBqQY1+Uqo+be+OfKA++tv55
RLCUyE0+72S0a0hoQRsMrRsWy/phzTC1HJbPN4HPGeCDAeBl0U9cbzHCzoWdMiLn
B6saf7s0Z7iKwOFvJx2mvvwFetb5oRGIwL1PlnWaKV4YRsbrk1cjJ2zPgay/J9/U
rOFPlF1hOQBPoXFjtSfDQFT1FBztZyKWaoYhsMntJQ8T4ObYtnBRB3teRIPFqVW9
6RcKFm1sSEdM/ucMRcH1oTFWB+jNl8GzBbrHcgyOw88S6C/iQtf5AkKYGysEF3Hh
ymJxSJHiAPPWWrgQx5oMQctp/Nx8rap3hKhgdI/PaR6CoEqqGx+xWh3Jeg0jeXxa
O8bG7lKboVy68pdZopyOsXsukpb/75lZmXkNLN43yrVgb1Wra8QvWj9waZrqWwl0
dDpZH8QVFVA8BQE2lOwypjHHBsZvVz09DOmEvfdlkjScxifVEQVnCwaLSVaUIw2H
o+hBRI3+2iMjw8Wry8R8r8WEGOtZGgwcY6PcewP5Q8D3zGOnvnt2j/PMxmNugA2h
HMV5mJJm1zyTlyMmf0fImsMRs8BKV7OiZcKNazVZJjA8lx/5kj/FydS/nHVdObiy
+5V1/qERGNXvyjX+ZQe9s1bGQ6V5VjDOsXjUE2DyCp/CNXF0WMw0UQ/akyvEPxuw
iX4HsUUF40tXTYriR/Ds8L30kiZRgmd8+3EwuwDZ1nFJs6AKubx15iDVBpZ28a9M
V1fdq28WnhEzrcMAqu83BVsACXcPz9PX3EUFtPdTDtqb3ISibjC/BJPiPvTdAemY
f6aQmjcH/tN3is+JAhICBHS3jkdhi3tFIGsvE+RnE7fNAtJzo/TFRRY8P1LIthMi
rlvZ9x9PkuX4HD/mE1SmLIx8B4fdn2LmB7cWRhMiu8G1Cc+DHxUpJkAj0HTWtOPZ
cTm93zAyEFAHz8+HtHtsnGDD/utbdG1nA+4wETizayKfSSCG2b47mXhdp7Sc0nF4
CGd1s8lXx91IqGIDfLYwKc1JZ7t6KGTgI57WLw5z1fysFjQ215bG6vIYjnNiuOQg
L+m0XajDJ4+GCqZdUE27cHt7RcSkMEjJmTZnoF8j0BRBtnmycLV+GRg0YVpxPbuG
7Y7hWCOVWfl0WYokA9Si/0XXSKWE22akffXUsfMRHljZ69B6wwGgghk8jtNc9hoG
qvc2iDJgj5PEagwSLrijexfX1TxrXqOVsQPyqG5fhQc+9UI86hQUk33nOisNeM3t
cthZjUcD2xon2/tssFLGP4O56sbXw2A7FRk3BiCpCzuHk0VEFtpx2zLgNosDtrJS
RiFJ8sa7+5U3X3Js+ZYqudee2Y7hi+qrbF6HM3VzGL0OzvhVL92lM4PqyMkDo7tY
JXplQSmo8l+HI7mw4THuQHySfIb1rohCUiE9kw0Wb/VeVEcb6eCCkZupn+w8ZYcE
purLQg0lNfbQoOtxWDvI6GmSiakUQ5NrsZBYAk9J8Trcgbc5GTV/dEI4L5UTyTb9
KNHVNB+3pFMe5ho+JqFdF7eRfCCq6N1MW4RsplLO9zeaUuNLsMc2bw7awE3SKhQE
4JmCVPWX4F0L9+CBEMRRk4W2fgs43BEb+hLWm6oEsUFhIbsZwg6hNW2+IlZ12aJe
GfPeE1N0XVt1NiuxoC2sAOyxUE5KOqlMFbRfIkVRL4PGHzYXbe6qoMYm7T+E0qYk
uLh0wgESxBNHJswBxHCjvuwifuvD+50VQ07kuux9d+jPvpVh0q2RLnzoRfxqXBOg
fEocuGGicX4UxtjxiaTE143mYH/DpCkdTwuzaMmUDc1mzcxnN121tBrTbA8SDiMw
cEK05hqCsJIn6VGF9s4elX2yQ6wapxKeO8rPpcmRdEBaQpls1clcpX++R/jpsHAg
+18Cw/9PZxkIr7/f4bOMUmhSYrCHepwMSs6cVYkDU78OfdxrC9v2XVCYE6ruRfOz
VApmKh5QclE7irwkWQVkrdU7jo16UaK5PQ4U9Fdq5XBJelllEgObi8XB0QicHGXh
J1xCVndLN9/iAdUUF9KM7mqx5ZnCSvCZ39lNBJelXaS290wuxkAaI8mR8JKRfgnT
zM4+ooUEXQ1Lu7kLFsqeYBqaVrr7vcpjzhBANblSpBUSTMlRnhEW+Y4ole1beJzp
Bwi2N/lLLjJs1owEvz1Gx6nnbCeif5Mc1t8CI66G7MMuoOl4Z1/2Xxw0s7p9fLDJ
fh/DXdLvXiMWawLSG0NxMpx+/zbztLAaReqRZwfoOHQv4Xq9n5ZCwscNpbgfMOFJ
M7JhVdpTCTOuo6vjSfL8qCmi+ANRfb/hnvJrHvsrYLc88ypPoj/EkZELiAyw0aQP
ZV0Br58phDApbmhycRXFMbGlKZhtmWg+Gm/sQGnicVEAbpaMexFWJUHGNhQjZnfY
TlC6B8Of0xEnO04jDrmQFVqbCHW3I8U+l2NoWCDFniI/R8uGe4fdBYVBby42hPBP
hnrtLtXO3yNr+7slmVkoyr4P3QvSdg8guIR40eU0ubfsLOZZwAQJg/oMmD4G4OuX
QfVN14/9MtmnUsEGrCzME28xfO5RMOs9nIhEAtb3nIabsUtR2hmgiH1uT+e3Xe5Q
VjOCR6Nn8Q8/bWPVF4FBWfBqYKa9pBGZsdITNTbgIt7vQrV7GstN6MGeWJ+tnyn8
ddnmv32tdWay1OJBj16dVZjhPnqLeiDMULM/jxXzDtWq0E7b1VSWDHyu3jNHN8mS
GT4TMjrWpNcuXpTEY5WkwLQ9zsdtnmF7IWbhae1LQNy6b8ElSL30AbxOg8hPEHn8
/Kk1ARKV8vz92hekuzH6gk/w1mt7pBHJhqBQKUlln2JAI0rjsBqAVFD2nqr7KtAE
Jr21JTFWzruOlgpPHjJ7MGyh/m2U29cnm+m1/iFPS4fwblaRtJiLQAPCN4mudnVk
KmHA7TJ3AIkVhneg0zWvvkFLdOvjYOkq/J+A4irSx+w/JyMSVhgQ+KkgRP5T/jSF
Er4IuOgymAwx4gbiKxkdqZgdFmyO/nife3FfGgBFuCM8EsJmm/x7LgAUkDDxtAMr
3BrTvGNRJ/pFLte99VZHdn7048mZpTw82ZyDCuCQHuL+Hw+9w11elDGD73ErMsXG
qX3nv8sOKvj6x30bQGIfbN/sSI7QAIXL9q4k3G463V8kNEAmx0TfiQQRvgPkbn3G
qZOvaRcNSn9xd3KZudT8ropvhA8CU4OQJ6mVImidZeJB1gaDv9DGwFyjoua7+Vup
PYEY2L4pBBDDZD31HJp/o75BwCWNO+XV9AjBMQ+rLp3j/bOsLbPY2+nhjvziYL1V
6gJoMb54UDYKKRQZbtHAGO/E4z6vKQkx3fKM+dXqtW5c4Pv19CVk4LRVOELp8D5b
U5MdXJKsHhCFKbW1BZJE8LRMfBTRd7Fp/ninHj1sho+YXE0IKDBB8OH3d0kV6y9s
oXb2v6s3Ic+RyG7sLA8Qcd6ZpiHKnLceyS8Q1KgxkVBGiVgkYXxoKnCTUd242emB
YekbcRcLfYjCcKhtQrKwxTCsxibXmLmXQDr2Hp7Lp0tFAgvaVTG5olSNVuYQOsX2
4NP4bTloXFM3UI/9f4szZtWMt7nssxHM4faKeVYunFTy332YJ8KonPsTC/1dOBL9
8d+nejRx8tjMPicAqinkNp+QmbWNmbMif7bjSd0mdvCOLho8Sthflo5vaq9+ZEd3
HY6r0tECJBaYmSJgfTJGv1/ArhJ26wibej48a4SBcCyl9/rRLFFFkr5REDlTU7aM
CtwLUlcOegzBym4nM+JkXlMD4lmg7DoU293yzPYoqwKWue5nb1X0nqmQbhiJnEcx
aCaO8Wqi+k+YvL4b+GaXAorTKGsCUfvQokQesiRDKlbsI9v73sY89rbCmf25m2MN
KZrgS5mkVHYekpEs6aDjVxE/28MIVKsNWKJRBFTZtGuAzn5ys7IC+BukniGWSs1C
0tzuRBdWgTm5ouxF2Z2ol5tNn4jAHMxbExPaCts0a6T4CaPhusPtjA/037FvBUHj
VBziodkwRxB2G48l8uYuYhnXivvZEfVNyWFBUw/RRwIfeHBOob3zA1LfPRTr8sY/
iHUSw8dt9aOBK6JeJ2Wex+BjDK/e3kgtSK+LZaE1/L4jw6nlj3LUYgXNnTrXT8F5
GlFF1Duxvvt7Mg8pcos7PYRl2drB4aAZ3v9HEseD0czmmwdcIs6131RYRvpTJ2U1
SqXkrMfjSpHmHLLa09DubdzE/9aFt7v+elLtuPjErzL0qz9XKKWziMtLB0/QlHw+
VfHwuZp5dYSCRrb2bd8dMRwq9g/pukhpAM2gTnmkRjw8VdcvZUs3w5GHUNNX94Rx
G2qNSY3Y5dFno7UuCIijHhZ+OMAUFjFAKpTVbC4GrRmlYcokmFVs9OdyCOKr4zlF
qpNVa0qeGdmgFQW3/mILB5rvI1C1ECS53ATAWuwkfH4PbKd61K4f1r53H2QotdHP
Zskr10UNG/vJ1HRkopL1LOtF6D3K4UCj3vii9tT6TbcAr7p0yeMiPj9UxuPT28Rq
osB5+eaKPalPMZ+tedGBrKttcTYHzLdpoNyaleHBVqSk4ve0PEsny80cwGDLjSxG
P/vUQyBGLcqmJaGUzqyvu7eWW/RDcoSkN5/xOXuOCKBh2hGzJwL2cYUIdYP6sINk
uf/FAT71Q6ECCa2RPhktfi/7x+RCzVIgRwukpOhGA0tmG4JUp4IEpzTFZ06Fro5J
Ys0aWDPBdRg9fL6RqwO+PSPVURFlz2dpJZiiGHdjuHXGlYb8axRmNYYuIAKpPHJ1
Hg6zHSggvbldDb5b762oIRKmHhU3wHclUCvcn0f/wO11SUOZJ/REMniWKwTbYZnz
lClox9+NWsaYuj3Lf7NZPIrcwz2o6UdlWPGMgGM5LqoxG2WTo9QsaszcJbvUznfQ
YW6F2rPEENwAQRzrvXRMkeB5mJSLaqsTPZ6ZzZP/RanFw77aUfBYPgAjKuqeYJ00
Y4pZRvieTujO3x6I/MqhQkvGOGy0kriZSoQk9PJQXagGaYoi8PEeLFSaIL09TnH5
2DJ/MoIarPxZ9NPhMx5ZA6Ox2zhhBYMf/6jzB4heiY9WLn6LfWybfOO14XOIJqAo
yd3/dwF+njjhOPbZkmFMyluEeRDeVPzoekqZUUeSDFav5r6LTFSHzIXsyATicKjb
tvtLj1OHhxxC0q4vqdo902zjIr5DaGQzrUUiAreru/sbpZ/246Inc0ufh4iPUK0x
e9uyCnYv9f6m//QHVqfelTQEONYbvmwRJz6TiyjB4EVJF8yyrwyoHiH2MRzOJpnk
wRUJksTywl+QKncJLlZQwZUL/M4m44+qG4AxQ8iU0+/j6HYKzRqzbN6CqNU5Vw3Y
2Zdh2sJgHWN/wH1h+7VysqidcziQv0erPlZz1MHjX4e/8TGCB1iiUbDOfAFw2h7s
qnHRtmJQZ5AlZAaOtHGOssF3fJ+KfublbPDKY7j7Ehpmrr/S2nb6sCKSlinTWqYf
ep185DHyOwoXrKHtJ7U8iSd52SjlkpW3UofxGQ1Uik6LrhULwiH3KqJLHOLSDdBq
iCcTpEspu7JCD/uZm2fGLj6rg8p2CVFlIVF+WSd5mQL3Jwxh5sDjGaABmq7tncxo
Il/rTgRCMmj0uD76FiwT6jNwrff12S05kzhj+fIKkvolJxgHZvK2s7zg/BITsmUc
ZPqXejcI0eQRmw2nuiRblAk9oSMRs1a72DLMR2mY0tFfdWVcar05WcB3i2ZB6BAS
+zBdEpG45Ip2wvDjANhRJUvo6VD7dukPYRuue1iQLCwvmI5BVICDFoLFA8JPhjxr
4DwLxZMiEMREIq8ihnK8zOeI1O0Um111npr+WLBvEdpzu88nU9Yxj8H3IbguP/yz
+vs53PGQSdUrpKpyzYSfM4HuVIeUjqW9Akip0ojkPD3RDRb9eyviGPemNl4D7kx1
p0YjjbpbLDlkj8Z3VfM9fmQRwh3oj2SJPCI2tL++GpLgOPSGZhO/tYc1zzuKg135
ykTfiJIi1OK+yqH5CkBu28LeseA9BVmzyUtioOU852MKNGhzBAFKDTqrNNJpJTJN
GqnAFmhP9tk1ptTWrCmO90g8KsZj9NQE3c2f3Ww8p9l4M7mEh+d1YvUx6yGzD2iN
0QNSeUgjomvGBL2VdL1a819S6ZADuEFNV+u8T0R291dEszE6bbF0dpnGvkG0YSBj
wnVIdQ4XwBUVq08k0vFdlwLTmHiXPBI/qIYYhB3/UFBrS7B5QW8lvx6zDGx8hX+a
9jUTo9fIR1f8tAaPMyzDXFfWM+4ioZvfLAtzWA1ObDxm3kxATjxVNQIE7OMB9D6O
PaFdyJ/lsKcDLfcO43lIG4H6nRJl7D68zFMTGliCBscPXavCXAcn3uiU/YHJNjG2
MLCnegitzPGReGZCQk/v+WXEzb/yjUkN2v9TW5wZJStW95hpe7JGIrGgsIMjzIvY
s/RRoq78/+CZqm2WAs4FbSfZcjlzBUS7X++qkiRNul7rUmLwoAqZBVAoDJAmmuON
gqGO51lbBbkmukhz75JrZdVhojNIuGFUa+8m5W85jmiCMNd/bwts2ws7xy0c0Ydo
iLCvsEyU8/B3TKky4u6iSkX5uCWtXJ6LEJbw183Yr53xoWt5ND4L+uLZUsOf5RNb
zrV/cT1KkPF5rEoclTX+WshA+eBHUjC7k4oi/1/RXstT/dayA5QzBaYkKLqkmAn4
gO8aYbYPmPE4xz+lwMDfp9KSbLwGbKaFeWmkusMqJZqBJj6a+Eb1OO0ZNz4OGlfF
DdVlrPp4SS4/HBMRTNgF+I4IM2wTjuYJXQFntEnfffIjp7uTkKPstmUaajt7fPhn
PgpyH/3Dmxau+HiWJJkKZJMm1eWanimFbfwGZ34/cLeeLPHV9w3LPumifNDErH49
cOarsuNJT+DrIKg8+CvDRNsHRLEFTaOEwICzNb6l3XshvjwvujyKGMSaPqnhloif
z9TJZZSKjj2rgbFnJfQTLw0KqazceGD46OxIw5A2TzyXk5+cPiqzG/UGkErKX+nB
iNj9//vPyaz1w41y503wKSBY2ZLhEbTz+CHFabX2PT8bUlFDLLTfg8rsrPkB1bzm
rP+J1E6s6c5o3UMzxVyx7o/H/+44skSiskHOQEEKlURJlJTRFwCY39X/6twSanUK
nejyLaLaMg2htON0iUVuMfJ6Z7IrNx3I8WJtHWYFieh9c0DwGVRaxTF00D67TkVg
Z/dJhpW26jD7PKFkLGDkPVQ1eFIUMpiaaqXpyQJVfpD98Xcz3cNA4OkKe5T+7AgT
DHM30Oqig+9XWl+pNiXWrItdAKhtg6La7xTkvzcX5MLALzHAoz9e7+Ay42K3cRGp
fLoouAcbA6KmHTDvU6dYn+fuLaI4JN2UyG4xLyjmHgHfZosEeQieIwGyMj5h/j1V
lrHizSLWH5MCqFM5VWXKcjwJUHRSZbXoh5tKEsU9tScZfwlNa+iCTKP34OZFA9Im
anRUHvQ7TNLr2z0mvsjb/2nu7SDrHJKSLKW0mtdewSilw0TxUKjicJhU6Eob3W+B
fslVzF0KzrvrjQN1+PsHoZ2OQky7M7O2qd5MTikuyQS1UGdN8MavIc+L96KdcNVr
n3VCMuoJ00lP70DyMqB0ZmnOiZe24cqU0nii/KUd0A2pH6h/732etcJp9ehXo5Lo
Tfb3BNNLoL6pRshZzpg4ioHc3ur0o2KIm4JPPZaJMI+qRrHl6C81KRRKLXXksJQq
zEDBPVWZKOnDe+CWx6r5T2nLxemfJTgTrgmAmBsQjVNs9jN9hI/sijXICnGGA5JW
KXaHncV3HsL6iP1IIgJu46Bz4Td3eF+llotXxV5wp9Oa208Fl/57BXFsxbYRCI6P
E7meVjsQLR6LXc5lLcOi3ugkVPwH3ocMJm4NpfEZ31iAr2NbVMgUkNKcki6zeVAO
ewiqOShTAzIjkn3rnKHjjq/gb/yO70V/F8HzqNrHGBNCts+kXYIN9EclSKY5Fdv9
NbMjiNxfsrB/XtYCG0FWcZGSs2GyUTJpJ1V04dIw8TIEO8lUqN21I4VRmJvdptCK
ySr34go9RSzlOO7HGqAp9or9Wvr/mV/ow6rSG92EEL/zHvT36EWgLnmr36SWavnm
bHQO6jiWfQi6M/3Jp12Y8MPOBF/64AA+AxQu8zJoFrhe9EBv3Q//doeUmf6Rz3Ft
OAckYhNPL3PVnPlziB+KU94UX4iVvZNb7Dd+j5g2NKxWu1moBIToE/FmNarcE5xq
ERMO1xf8h0VvgbqYfLSSYfCbKd+PGmsL9dMebmnf4eAtAKU0zhFLBvVgW37vAquK
788KmM5yCPRb/I/3o6SGX1R4Ntc8LXNZYu3cBKjL/Nes6h7PMgvb5hvyx8m9CA1A
evuGKDHzRN11fUkomGzLdPK2XQReS/rWHsBr3PfexoK8/3UzlN1trFMU/6pwOjiw
1bKr9PJNn/TGbHeRcjhYbPD6EVVKFx5OE1mmt/8efdTESlq7f4E/bKWnUyqPk6pn
LLC2/AqjXX5p1G8wqcLA2StkVLZjM63sp9O1Jox/oCqO62XFSp8XkMg6/Yd6ObWU
fROOwLM0k10qidiEf8OAIgO1btAoZyU6+TUR1ZbwSIA20wAvgfBPZQ3x3R+fcgDb
4BO9w/CrvkW85MKyqLryOi8LfHC8b5g8ysQhHYjAZQ03zIidquui8VVQey3ONyv7
N2wXYqIAK2Jro43gK1BgrNMM8AYRn/cDGg+G5YJ8lWBUMJU9vg5O/dEY80YxrV+K
iimauKInFK01jt/ezPY88e1h/1CFlau+4XFMd9iOhP7e7S3FHh2UXGeaFUWV+ceT
StOXr3uLpcs51LTXDD+QkXcOHHaEGo7epGR3+H4lGoGgTmclMxqDnk4vH24S79wm
UF9P5AGRQ1gJgdP+dDRmuj7HzNJ+I7EpDR+qzelcbiDQLKOjoc8x2f6xqiTexKu9
zTKoKODZIg6Nw+F3+llrsl+KrHjmxlFUDupDgoSg+nsfWAhpCR2X3yYw7B6w6tL/
SKjvz722D9MZu3mk32PWOmK9PmCdEym/e3cFrMTCYYzdSolYBjoGfOLuu1ARDqdl
IPfVw4LhUJeopa05HS4G4wdcPK85Bn5RolgSiAUym2LsQs8trGGgyh/FmmAVhZUE
wFokUoAStLHEeK0cQYuaEKfxZNCqviZ0eVIEvD6Xzh+NhR4WgjH8YHhlHJ/xGlAi
MEraIUkMO17Aj8Fye5MXTxuNn+FYc8qjs1b4gvjlxGOuZ6ZcWdHvUsRoqVLkyvdd
5WpGrjDWxbDQfbXofRzhu7uZSsOfIywTn0xtmhBtjKpCSz94Y1U+qoi+ZzJ+KTvz
xtQsiiLNv+fTAjHNzyM0noEnLQ8p2QDQiH3zYe+9QMS2fXkccrGy20irGHw1JIhb
bTjwxMMwbZCZtoaS47lVWzjsUvZpDD/LWMk6s1C8V/kIlvuuu6ueZ1db6ALTGZLy
01L858ntV5aAzadQroZCLyF4dRGk2aEjcoaNmdvmfFK3rd5hyh1XiRta5DNJaCzx
a2yNrwy0hGt6DlDd5fLzBLM14k1Eh6rioxdwE2cmyl9qI+jqsRhU+1rO3nabMWj+
HGmpSdRexpPG/YDUOrpFB1EaBepCt6flHZmcaO2HjLQQDl32brSMORqCmtvvsv8a
7Rye1a+mU6P1Yl9b+x6uGRYmtJfQkBEXM36lCMgK8Nunh2BYhDK34LY+q7IsMCIV
spv50dGCnJgfpc+8YGJ1FkXA/rZhOmNfPf/uYWtI2oWr50LoHWpl0fXVjv7O2OYG
ZKcPEomuBVE3UewK2Db1yKP5zpIIQ0kWCzyX8Mg2dS+3qNQru74OJPEIniGQI6OB
KLsf3OGDaV09i7MMkCmSamlCLZb/uHu8zIIkspfzzanNsWDXzEbLQgy1+T9302ii
aQt5KrZ5rqbQemlrfjzRdhLwPp66Stax5UeFfsOuSDIl6wzl9erQrE9evXbpiP9g
2VaSKEIuGoJ/tQMch1Zeef1r6qsv+ndh6t9+Nq10JcqQS1JcSQFVqMY07Yf5fC+V
tQrSTSaeDPKr6/iz7DDd2gtQ+wG5B1TYEQrAyZJpkjnqwmIB9hAmgUAipPYKM4Ln
MhhQyN93FmQC6gZ56cDaF+awfv7iAaFLZAKsyO1VWyh8VF9e84jU+fA+zIeYlPVi
X6G93LBwbI8glgbTzUmvdoEIhxf5cGlAxndPCEwKlr6k2PE3X+eOG9mlEQDoDvLa
JkCUCgMkYWwMXB294h9cfB/CIYdGOQZGd3/QL3qXohTJJJd74MpPr5e4W/DNtvc5
SEJCD5Lm5S2ookBvlX6jT9zQx8SM9T9IREhSK1ixuNwhocnDkpAW2HEAiiuoT7aA
5h1JKMBrg5/xhwzUFO8kfcyEsrEzh7lx6YBa/Gue8HLaOuKDixHqiMZaTozu6EKk
K1b0Ne8Nso1Lmn2mHGvvmRmWPFMrrnxa4oFyehLamGb/ETKU1DPqeqny1Bdiuhnl
grs8h+gvOQE/ujPYIf9PjxgDnfwtYoKOz2X6uSxiayEA+m7XlkVCTQvsB+ChY+Do
ZxIgVoe91k/BPGlEPbIOgMw3oX6qPs6VBFancvqaaA4+kD4qrePv8SQgR1Df598R
QN2zDoeW2BqjPZ2U++zcbShEDXtWOSw0JHoNEBzRpkuxkj5Un5Z+JYuiFbQhZie7
kuc3ujcdVc1OC4hrjbfWhhM+urfzW/p9NiIhfszmV4UzF1KstbdOREnIucraNZrP
AA2ArG+LyADsf6dqdm0LhB9YsqtqJ1kTa6U9iSUCU9RhlmhmYg0uk4bBJtc8INbR
B18jPrZqs75Jd4GpFmvqh4bjeG88cDAQg2uiRr6Qa3Y4N1xTbjne1jPpTV9q4ztN
2TuwhND8US0aLvowyqtM3Jy7RaVLgggmsOzPTf7wHAshyiD1ye9FPJ4n7pXjBY5I
GQ6y9i7CWqlv1I5w+JJ80tpeoCDkrdZ9Z6j/d2aF2JXP5hBwNbwOoJ2c9h+uulnP
P90ophP5plIjCIYE24g9Wfib9R5/ikEcIsbaBWgz2z5u/zvzpHNf9r27Y6VXJNmB
Rve1HgjgQzJhn/XAXqQ2VMzGsXF6I6yCkLa9yyOJn9Z4n5ic7o8T6UB5WS9HGff+
7UUJzXDafCcjx9mLNfL97/hu8FQnH2NueeT4v6I3W4pa/DMumBHKqVTI8A4GLCqJ
CnnM3H3qQZmYGpkl8Yb65JzYLS5fp84ez4ZsDplWlZvWcsNKYjFoCF7rk4wGmymV
LD3vIkKTSb91SYG355hBTeqWo8KNRkbz4rTj+zrXSS5aGaMrM5mPJ6iYgJi9/dbd
mhuYvfKHF2GiOYPlhp5gNjK3ndkTiTQ+wNtFx/o2zobTIcShPBpy0ACx+dig79v2
ec1xjnbUrR2LelEyR538jq3OKdAjMOkeCHDjrDAIkkDnuZ+e2WDJ8YBkppPNcQyQ
p5llaKLngCdJ3NaTLzCmVqPJWIAtVzLTV8u+BX1yqLut4ftBBG4bXz34smHOGoVI
VmvgNfS6Ky7cM5afmBSluGdAmGbegqJAiqyh6zQO6tqMVZwzUWaY+xTnqPejCqff
PMwU0C2nG1L6xDCDLTDLB3ODi6KRDX+n8jT7ZOgzBNGMPhbS7wm2XZzw0NwfgFyM
NmzqO3secaMkkw1EfXBwAVPU71mL8Pvle5HdiR+CAag7h5cgrnFpRQR9sBsNFKKX
skY7tJvFb2NaflruwZpJjEvFtN6EHnu9x28SvW7/SVxJgPy5WAqxoHApsb4J+uFw
lQYKfF7sDzXCe0MNa1G9qbneZnPgP+cy0ZrrGu6D2z2eOthLQQ9MVCxjmXCEq/O+
Bw+M4ztFiklufy8L4I2TG333wz4THI29hludsK2ue/EcBwVElFUY94b26WW+RGSM
D9dbz0zL0OCkLIZRdKSl7jXTm18T8k2QH8n9rkhVO1od0YUi/ChV6zDP5VK3sCEl
TosHv6zBoPL0GIEDBv5TUI8NOH9Oc+26f/h9nm40tulPseZn97Hkk9j3g19NOXBO
chCH0GJCbTXRRlG+QiCjdz14N92GunBt+3uVsKh3pmH14vWvdC6pGCh3iqd1Eak4
sbBR5B0Hyepdac1jdfZwV10yT8C7pyXJnmTbXs3SekG8+GGAlxSqflziHyAh/0Qh
fYRI/TeYzhCWxw7HStbtfBG2qGWbkB/kvIrIgFHa0ZZzWdttjNUsqv6ocrdU2pxS
HIjO0nJgDi6RMfO8Hvy6wStN5bZzMgMcVWWli8ej6hwtMBDYT01fckugr+QhiWv6
UDjAlQ7sXaNZrz+6AhYYnp8mZJr17Tk3kJyGhkc5I5nQSQEKaF2Xbd45LhC4nrP4
IHIt+dhDucZK9JoBatZp1xJ7OyHSGdrLEc0mqcj9q/AzYaxC1pUhWNK73ATw888D
alvpwqd6lBHho1z1zxJizn2Ri63QaD8nG6JKDm3jZpqONOhxeNQiCIU+arBkcoGu
MKV3ZME6lS7wZcJ+kfZVXJ44QcW5u+Bo+53yqeOfAF85KUYnVI6IUppkrbGpXVJd
opzU9JZ7SyQCjtrCOtfxM9Sj6VhvtjdEryu6RpeZt8ToCgaAoQAzo2uA3BcW/JSv
LtL25Qmf9OmxL4v4wmQRKjRWMQR/24/ZmEyc6cRuaw2w7u3Lu/4rAoYgNI02Vb7Y
Nj5crolnpoiFVdhqIiR7MGI6fAq7JPm1oC45U+Nvkt9eYEtmD93wScanEJvNacOh
gVztEbtg9xFG90dKuF8blCUHAdoCTtrC+qLQVk9c4kj4TUJZMphUr9syEg51yAfk
9ME+MmCbFQkhV1n0cM527zH71kwFcWXXI8fYQLnIDljJapjSrMl8Z8/zzMZr1nL1
69Z8WgHRmp8Q5jYgrZTZSI4QLa+ofmN0Hv9rdfc3t+t4XFEeZUxnWfbC0cj1dP1B
6f/IkjJoKOmJMsKddh/r98BQVD/dAqA4wCM700jkOzWtWYNmDegbCrsJVsNmwef9
feVoOzHpGjfT3bX3PnUKQPRP6+HxiMCVZlhYKzeE55ywEExNKhBA7IPcNXmCMbj3
KDAQwRG2WWpPKIp94jofn5h/lMc7FVjbxdyHegrrSJkWCModycz6E/rfQR/nUzZz
oOidBRQZoLS0GsZN7Tu/lYcMWxiTzNkOvp6aL6pnCTGg8DEv59MoFqYhOr+3Ji4f
uNZ8F59/HGKU/HzNKIGxEnp4SS/6iA12N1V7JMIKuPGuo0aYf1ZNuwl4+bGnooYc
rGo29fmKQcpMGXZG4gaAbDE7BTD5CLT1zapsa0fwtVw2MLb5QdYd6RLTER4/dCj9
0gIkgSzGXjiO0roo2KQGXiz9xIFbR7s/Z2W+RACFv2BiHCZI+HK4z79RRCxxOKad
fZYOYZFT52+AkV0+Ky1AKOScsX75i3dLROq8Vz7dN2yb80QL628PEqqERpWEtE5g
L4pQs3nXHtXRu9XBIRqxhRoFQ7jd4GqLtXpUEKfx3dbP1k1SP+bEQrTtsjiP1SB9
36ZaaboDnmf8MUx1Kc14Ow7DDwpZf7OE7rR1Xl6HuuJ+TdArX2cFWvejJo6MG3Ug
wI1BE2Bp++t7Bb4a3uBCVBa7gPwXAgNBC953YHK+Ahn/SnsCcnKDCPJ3mcsYLZU+
KEkpUVEDZarJ5SOLqXZSLRlhFyXcaYJUh6fZeOnkwGHZhFsgPz+ghIo+kYx0D38M
um/eYFdUA5EUvu/GKwqCvr6KMLz+mZ+ISNCkTbTy7Z19Xh531beVt1Gr3RAOgYL2
68jquMTvwUn8XYB19RocS/7w/rt/KLhiYSb/xiVSl9nFV8oMz1J9tm7vEmhlj3XH
whyaqsaOGpHtNLTjTs/9fps3ymNL7m10Q7OM6eHOwTIZaOOsblQCw7QK7+qFbIHk
bCHm7Tn7nrCxalK50kIlgHYgpks8bqOneRugGuADldsznUKi5OFqljcRXt02fTk6
arFxjafm3ZVTiH78tYhDWl6NwTwBJKDiQMpHJnswNBtz2+a3x0gS6sdu7MYsghWY
/eB2Djlk0mtIUCKO/Jg/hgNEYCMz2EgoH1559dv0wd7kK/GfGrdYXh1MjqR5J0Hg
BbxbdFeSH8OsC4kL/rK1yRT9e/VDSzdttX2ywHxHlUNE8xVhWLLgohK1GzSxrvfZ
KSWKjvDRII39VfN/Kt8EcndkSsqNKpySKYGrJ2MLvR7oZyde2cEdJjHVVyUxqHvE
sXnbSLIBzek8J//g5oYmHUWXPbcDDBiTcCN8QkBqJtthwnnix2gZe85g7mLjckCO
Zzqh7LYs2Oszq4Dj3M0rbVqTK8z7ptrOwHLv6VbmrChe+OVE9pYHi6t1TqvdIWvj
+mOT/ho+pcbPyvhftMWz9bI2Z7Vki5yvFB7GdHkdPQY9IscKc+FYtnjUkJ6aG+pR
uR5cmv4PXXJ+eFumVubKFtjbzpj8MxyY2Kae43DOt7HOe9Yleeg07lWlEaLYNawf
0g3YWp3fWTtUwsRT4ODVm6oWmUWk6x4itViQ52sRSeBfVtDbPOWu8TnAh7IkEovs
NG8tkWSIiJq3B28KTTHuopGp2g+3fwWJ+dvzQ8cyYkTZdHrFX7ZZEkJNpSAsTP6E
Kq6blKTfi3a5eq5QMKnNhJMN80GJziWBa9GYNZrtMlfIpsf+nNOo/Vd5X7eT6KAn
7GSjQ229z29lc79PEPAa0Wr3to7YAEAiBrU2wOzooVMttBnC57I11CsLDa3ZyQYn
UQ7yzZrNFn9FcMlxRvYHqmSj5bI5jQXy0m6LILX3QfmiR3gq0K02Fw+sRLWy1k+s
xXU8uRh8JGiXlPnrI79V1+zBys4iRMRirmbkyKARrDVNM2WGrBLNVhSZn9xfqUke
AYA1+N3Oij9OJ3MiqIrSwgC4+fASQLaZ+9kwPr/c2EmZxIcIBuDmkO/JhW+2h3xu
Trf3lzAKZh4MhbadAgNUMnX5Hy4wtbSCW877LivRY54235WWA0LhT+sJ03qmCYzQ
OubHfzrfPI+H9YEvEF5ckbZoAh+us+B5Fwqip8O/ZRneNwWmqgDVYko+WcX01TW3
N8Xs3jafnDssmGMnc70eCs+YEj1+Rf1sNQU9KhCigxK5hSui7qn2uGwfOq5cS3at
EVvfIgWU+vMc84EtAsFI3nRJAnDY6LE2Nna3RhQ13eZPETOsdNoDSZMIz3OnAFG4
C2B9Mpc8qNQUQ4BsN8nr0YKYVbmYQX3dm+eRhXlnnj7uaJMI2ahvTEHDpyyDgDKz
vDlq/odpnCPMK6yoAWVt8tmLboF71ZK2mVpIoetNQLxpRm84UbbBuRjiKvI9/sjM
2EJmwLnGLiTUZXSIXxsfZ2r21A30ElORh51Z98AhYZSKp7vTDPBIumRXlWrkvlEc
roIaNNrzYguy7JOXgO5/wSaHHfQJ8oFNDrRQxdIRyOOzRt6hWUu+w802ouQe/XoZ
Lu2+YlCuaS87P1rJhaJjmVwALGJzmmnyTbnUsANUJbqBWhtZlOpPkm7gh8c6hFWg
bCJtT/nlw2FqWbysyJvlSuEbC/5xdtqYvafFTLv09Yig6/RtB5pIShlza1DmsmHH
35sTFqpzgBaTq0p6gvwKnH68d0eCIF0fp5VumltIuJySffWKKf8/I+WOMDAGUt36
h578Sh6GBOM0jkfW28daEEngajlEtBBj9+J49xL+MkwpSW2YmfT9DE2P/0/3DXB0
xdxPyWaS54ocikHEQirLPyvCyn3Lk8RNlyZ5AbiIJjVz6wJmzxwTDp+nprSFAziC
uNMacAaqoNXE2zGgungjENj7ndX6A6PHZ2hecuDvMx///ILkTdixkW5EC2eV65mM
Tw2zsw9MEB7mtqEz2irG+ni9L/N7jNTBKNnC4KnhZBb/4BlmJJ3O5rxCz/Rqr1kl
YEv5B4WDkdpZBIczr9DaSxnPzqzN0cpSSYa/I6lZPI4mj1UFBeRw7TQb94eJV4YK
pZugh39f8++ZhCZkJEcX9ZsyTLeg/OhHq5e/Z4MNarMl2rm4oO+uXU96uYlDOkxt
0SDsyoji4XZCzS3Gkdfmp6h7u57o+S23s6E1NqZme7loW60STNzfzAddu822FZMX
cCtidoquOHxXRN4hsfIXih8pX/O0/AXM3Sv1XZzt9p1uEJisylDbcj52j8AR1XXo
G82E29NWS3FGg+7JGIT2vHoITbUgDhUUIOFyVpJI2ay15IqxXZMmg+9qIxL2Axlx
R8iFWwer1UFLOXbFDpAxGa7wtaNdMEgbrSjOQ7DcBPWv9HdKoByMKV2wriP5EXgb
r36ZzGOl8FZQIzY2nWjQJYIBr+VShA34WKziQxP6tH4VQOYXAoher6jEZfrKrVgZ
TogUcf7A1rzlAIA7TqU1TyU7Bqqwm/HY5cYjF66Y3Ne6O4brkoj0g8r6E3NKb2x6
d96l+9bhml+a/DPXdz+GlsagkJ3NmCVfr0RyJcgbVR4aVjcTWvKCNrRPpq89yhhG
sE6tP+R6PVUqcdAUsmCDH7qjh32cgec2+njCUQI0KFv6FWcVUqwhCfUU3GtRDiQH
BJwJQSwAoSYTMILfML5/Ztvt/LLyfKDzzwrTN1nRdc+bIwvEr529+RBflcd7PLJS
BML6QdnmNWGKfiwsemQHcccqdAMoF6Ng9f9BuJxUpq/TmcYsC2k3Dzx1M1j8JRtq
0tyujc6vEcD+fh/jOmjN4g6oCXHCN7IeQBrkeCWMWq7EtCoq+p/P4U8KzIhpXJg9
J3c7vfHxSD6yLDLGXYZ5c6q4fxgFtPTu63+p162g41cAz1iyJ77qaSFMPeq0UKSf
L6INaW+CUQGTS/tCquZAjT4QtA7EL750vlTCH2UGm961vxJ4XWA8AlwcAAC+WUkU
e472wUCnSBj84jtEnkuaG55M8+ClrPnGvF09Zh2mT61eIfFFIu0ni4U74VOKEJCo
HEaotr4CMxs2SQMPgWGDYzc7L7lTrGO1uYxSHCuPMCoCQ9Nv/RGpWnrjKGS6TJjZ
+a8XTJ55oo0Nr+5H5Lun2pQWpc9ILLpLs5Nd3cHsi9qaGtxjM+4sWr5nJXSqPYa4
h3wDfObHCGzFk1Lwijglvlh56B5dGpqDbgY/DEsQaMTOGP4ycprNebrehlWRUsi+
L0f3GGuqi6FpULeQU5N9n8SvYlfzr0UvRHWx9q/ELBNQCPP74+tm8h6BJ3iqpafJ
k+Bj7rh3iIpDRoyK1dsUn2qMgTsXCWc2NGlRKAOt1uJFZ8pRsz+JjwcsPYEO+pf5
YoQ5ztLI/hs1kVZ8fNHJ+p0wQ+a55tYmgpVTHerbJv673t+fm7SaeONfuY9DKEgZ
Jjg6Fr0aNQPSzp9QXbShRFNkzdx99HleETG0y6q9Fg9we+aCqGHzZH69NmL3EKG5
OR3X2EYuEYAsc/HdgPrXAB5zpAoqge0bGXhQMwtgHOlpIWR29Ky1tjFsQhiA1pV9
UTmaTakQbNnV7hO+uuzDgf55j5bpPKMBi5IgxWcOgHzAfhxVIhaoycN+EXSMz9VG
8CSWrgqeliLH9a/ZXOSobFnOzmpe4wCQO8eeSmMKjB/7uZ0gej28Uy9kPbCr5rtw
gHABLoP1nV+NJh3UtO2jAmkCeGOvcZWlPd25ow/pOfipQK38LB92XMLxW9qZqLXd
5ITV1Ta/P7Hfg9kD4pRhovMXT8Y00w/mjMeyWr9t7FTQL4jDO/Vi6cTHm5SCGrsa
ia+phTIpBl9aYX8xvz3yxtJuDSZ8nJEyakjRi6xl9f8M0apCR0f+D/r2nhY6lrR7
DsVE1Tq/NEAU/JYBVxVMB24tHLXO3SGefH981ku8AImwVMtO84VGkL25rbQYqHrg
4+LoraRwBsCacpvf1In76RzkNpjx1605JJ7yZZvYE2upgrd6Y/D+3GN2psyCUkLC
rhsxLqL7/kBlWY9De2QhDDFUwdiMrnf2BxOJeb93y8RvNoswzYD29MVJaJuDlYFN
1gCiYi3drWDGyaKuLiF1qnWLfW9aAvcgNHPMpjlIQKSXZFIN9EQ2Hi1zzewcFr55
Gly9yRJgVkzrJCibp5wHyoIgB9dUOI5BR5asd8oFUV8m3Z8TJlT5Sf34z7p0LRjk
GEBym8Eh7KieMzrTUYjZZznybm2V5XB0Qedi8N0ahPwXOlLITPxE4zdUjguD2kIE
NRPJxcPpu1hAyWntLJaYTnKMQasoN0peo0YogbFzeWh30O/xPemMM3y1E++WZhOU
L3UYWi6qjXKkFCU5alWGQLG8+IvNS9QWqg/Y2q0gGRdLyo0dL/PC0EKgYV6oLwYI
5nEjDYr/tDBfyILbyaWVoVCOeIDs7Y+A/00f+Rx3kY8qADQMLI40hNovVKCjRFc9
NSzhl4U/UsOJT0VhQeGSOx2fDEXoeRe4jt7it1VkOWz7CKeI86qgsm2G7fQ+GByw
Ob/mOhcoKSzJo3CZojavGenfUYXW7g54xNhUPRT8yEpCMxq0JVFuKP8G/elW4UIh
K8e4ENZvb0r6efegjiKxx0Vk1YeWVbBXVucTMWiZ9KF1CG8U9DX0r8GTtoaVu8yQ
OryiVEGAq8bmHag21zO/RRZQa1X5hwwLPRACqz+XnBjyqaF6sYIbT30N9Q/P/PDI
7VrO321BYkofslsTjC7KKaLjhc9qcpLJF6Ct4ad2Li/ksSki2Us2w1dUTf/Go1wU
Q6r0Hd2hRPOvUH01l/EYvyo2gW7JMMIVlUClEjIava05Ah8n5GeAcBJZmUIBj7Zo
8jLmRONfpm02ER82WVfr4UrKvU7FK/PcIHPbU9bFtvOF7HikJCOxz34hQFNlpK8l
BJo5h/lixNPCfyOKloQ9WGpnTX0Dmti7rJhrnnVkrfAzSYIdC1zrO4McHlP1anKd
jiXzDlcEf2Px14dGUqjupfeBUrfXF2EQX64xqF1F4ZC3u0yDKUXI5rC1kImH/o/d
2iOlxvx/MGVcc3/13y0q1YF4tPQHJdDNec3bFmBVulXvcK3/yZsTuecp1LIbiu2+
z+x1nex5R/E+U0H5xCKn8418PhD0FlF/jowY7NwJY9WAOLhjMlK8N9lyrEfPBqBB
91J6kTOYw+DVAx2Z6ssGB3YkKtzVp+2gQh9Kvvn19CZjhBSTz5CtO1ayb4zIQ3xy
5izRQ1O5nXLcw977+AYJXNF8kU9JzyZihSHup8pNLaWBRQqcfdqLRlWqkvDuXyer
cJV6nJzlzjTPztQ62O3eFt4DcoooonJJHfK5fiRCz85kvUinn2SlJQxFOi72GbLV
Q5yWjw6PZ8dwGOR3Ic5R3suXY4YqGFafYLKMXP9b5BzMxxwWw5axQz7em5T4LkQO
YRuqlNu83onV/54ceRmjzxXUYwcvXau/d5J9zvS0y3rOSoCdv/gJoDyLVNVA8Izu
IGrHgLGfQkbZGKwlekNUlkRdhymlQwxMtdynE5WFd9Pud6uVL6VBy/6doQUxIu3q
HqlThSyCBWRUraq77BuaSzflGe6s3DVdD9uEERaa9r7On2AAXfJShZPOhWGhVgfz
3m3+Xw+8SD3c+8rJFe7+DTqLCV8QPq6+5l/GwUtI5m0gWpXUWVIaDnmQwD+xh5AH
sMTGaeL3xK9i55g6Y4+YdwKI/1ABmTjA8w0Qg1eXm4hzUd1MKlrOBLfqKBw6LzWh
MKZ8fk7jABk9PF/cK2VCGReneWbsHvcqLhYZ74VRwQOR6V1X1UGNV1NWwgMNVn8q
cI/s9bH1z5mtC/BaUGyFsoqBIugBzDDpQqwCaK4Z0dDpFidIK1LS3UqHpmMzIe2a
P6Mg5HiAFAWs3o2qb0wy40T6SfGP0gXFAbWJiTFZ6bvFIhCVFEu0DfUo9xKvyPgX
9T6XVCg3OPa85V5DiFuFDt37rcTPsGzJBykRlBdU2OHGfjW+uaFdPoOURMxhN7Jo
qgw2zk5y+IpMtPQ6cWYG7ono3NoS9wwl7r03oYcU2dEypP5TF/GjPKr0CRxYU4uf
n0pkO0uzORRRQ19V3fIYkBy1v1fVO3SmQQxeV6T0Y/0yzCUmU54fowaHUkiOyfkD
BOFBmJkNIWkd6IBYrfgdZLD7z9aEVtiCfc99xvdAabOisEnvY8IRntF+DIynH4Op
KKrb+A2rCia0+REdBwrcRTI159KYvZBigr+vMOZHwLjfA4v5aXWvmXcfpayxBbD9
QkHi11J5pCADVp6nVxstvJYQLEKmhNqZXiwRlol5OXTQTX99LHlGXFKzt8J4fm8e
S1/GHg+tpqIIfXMtGswQykADRw7LSbIiWPG3TiyYRHGXxQwsgOLMZC2rkXFSDFeR
QfAUeCf4fUUL2bJJbgQl1wRcj/HGLWC0/nidRlW65+FVxO3m4T+Sqkf6GjfxsdqH
wl70jNLiNzP8F9AetO3vNHqJ4M+2GGJjGZPkjBz4lY5X0h/BCPRsV4RzfTcTWXi6
sKVZabio+AQwlGoinkkLpBjA3gQ//HGChIiTzRuvTgpdkYeUYf0BkYjfDTYwADJc
zubbV1sxxN3r/iIdY/riXXiFIUQRfayNF+kxQVEXt5utORsPKTc1ZFAHJnblevJb
tNsv+I23v/XeYNGf5gwmxWi8JV2zxh1Y2FlAopcsvwBxD5ViLN2yhHQIxlby2c9D
+bN/s3ZxUbQ9KubfkDNfZ6rrSrbS+mf5b16v2VT/Vgochqry7T+ZD6+VoCaQkrZW
ZYZJphYN/WX1yue4O/RUBJTAuSUFFCcPk9HUG35MB6WYWxjJVh0rOVAivM/1/mbp
9ybjactNAql7hZpXCSNwXZJWj1D8y6jqV32FqiPSvX5szqU0K+1807/rGfLKt/xy
MTb8c42qc6fmYN8ryBhiKcLAMiwFbICmlJjPf4E+p7uBvUSN55zc805SsaW9N58+
ZyeF5b7bdQZFWwF1MAa9eCEB0Tz6VrNEmYdRjPShtWzHrG4y+012WR07jB76aANN
SVLI3nrMgy3Dyi3xZKA9pznhv/RoS20COVYB9U7qPx7nZockQYKB/Ki9OwQQZ6mi
ckAR7zomUpWKO+V3lL5A/hCBmfZS3KW9RGWviUmso9lmVzQ8dsTFCaT9xGMwwjjC
zIpedGJZzLxOU22zwEpoaLc8uV/xeCqSIhtugXy+B0O2vZW5HuAJFipXwBLQuraH
E99ODqmhkNNP2i5o8BFxGrgAQmFPldrAZ3ZobQ/eaP265GIJ99Bse9t64+r95w3l
eTlJwuB/MjwjC+OmM+taqpL0dY231CNpnC1qV0GYTbGPPutqwaKq0dLxCIZHTI+9
/yNTLdZP6DdnJ+K7C8yrvCGrpDxue8HMGp1IloJSBhfXU79got+zknH5NA31YkpP
a9oWtlgDvgO8CeTk9Tdcme6uEnN7k0A0u5pYBk9QWHv8BGOlLj/gcsYjCyFZnbfO
SevAb9/YUkh8xBRWv+jmxR79PXsVsZ9ohxjGtcDU0mkm6OpP8ptK4UbeoXsCA9VL
ov6I3g5sTKMKMWF4X6vLTWScNS23Lai8ljwLWfawWH9AVZJKUaS9ZyfGm6lY/2L7
7g4MQ3eVInHLAbDs6G/9CidIB+9CfWWXj5QBXD2tJI3ykq3Rxt96iyNmi+CYo3/p
Qkwj24G9D0Nxc6ZzPUsi5HC7f04MiMgP2lECAS1oCaLT7wtShr44+X0bXnZLsDrT
+TyLXE02Wp9UT0BydOoCxjfOga2K2pOncAbuFsAPC9cRLolUZ+pb4mGvZqE87wVR
2QjQCx+xByqdmypVabMJwv7dsKEvCr0FZ+N1f6h2xhFXOAz0tlF6B39UTE1o2I2x
Ag012/Qb0xBjFjpZTyaQYEpcN2rl1xvLI7quWh+X70GrCd8OVXZY6WTmJ45KBRG+
T5+k3qGH7W14oPB8BYAfkYomXcRAYS6t0dk9jKCWJUiZYJfEjjKMqmW+zjNo5vO3
+e07UykTkJ1s2z15mgpxMpL4HF6Y8dzg7xXZQs1bAvH6RT3J3Y+K0E6fWdCWXZaF
sJUPywblarN7Ui+nvTi6xhMVbVqlZsm413sB1xRk6y0u5GCPXyL6R2lyh4+5YCKL
eYAvy/23EkJV8sFpspbkRc3hu0u1IKNs2rhoJrm9sQtI6pLgLSfV+o7soOWc8Jo/
95IUn2orGpU/ramJFlwBhFMf7LAkWNImqZ/gK1dHssKWqWyGDpYo3VkAiOHPRA4Z
EXtsRhCKdWcvUR7fy5xGk7jfcU9l2k3n5fxp6aDKhuBSTV3SovJ43tcO1T2Rxe2S
ynjRfCpWCMCm/jcUewFKwVC7XjnTLjrq/CRcN9TEKKbDntNpl+y9YA2MEvgEbPSq
bn2LmuVqYuwR4BZAs7YiZdt87rJ86eYpzPK3Fou+CbfZocUi5dPIHYKbPvqmpUBr
+NUitcNsRnyi2DzDpDHxkqMYiMxPmZFS3j+Mfs1xGcY9wf0jB1M2QdCVuJAFHRgA
CsOTb8t0euSglAQwdM5gRgCrHQfW+OC02iOtj5j/+59mjg2LqJVzNQi0GN3H3dxp
nlqrqw0ClCUVs/Yd0NRF2a4bqryvHTWLgvva6IRAEWNtpZrxn5LDneHffxcrJt4J
U2X/+KFK2iqTqclAaCrVUC5KorUGqXE5+M49mOkZLq0F33YHLw4vIChxoDxLMqdJ
vhG+CLJNvCByudIZK1xOOlNrUd7tytvvql+bhrJzOUtV1KgdE1BTxe7tOw2kTbYv
oqwk1JnZgV5tZTYodNxpkbCUh+P+u9dk5CZnSGeIAz+XgQaklGFq7g2YZB0bqfW4
45kfuh4I/bM+XAuQlIBdOAcK208Sl9IGhfr+UDw1tzXiPgiEroh2j7jl2Kqg00Jc
ldHXJCFC/B6BEgQzQnVnLNsUt5xQlC+4WIbwYKX76WUSO9/mJGVw6cGJnfdyaQIK
l0eC+6lf4y43VtP/kjrAJdKyf1H7fHNeNq/fKUM8Tsdepp0G6t6J1SGlxT7IsjFq
EEDG+/PG/SwtnNY8ZQzVxdGh3zRKqjhceu91IJ6ZimlyJQAb8nTAdxmsy7NwjTYZ
smIQh9KID0jkwb7ZuzBoxjIMeR+TiJLjNTtXjgV/cRDMmJjhDm+um6IwxLdNgjWD
ou2y02r4p3S9x4bN6+yLH6OAQaMntS1i1e1wKqWJIAR9T4vfZN8UXMJtd/S6f+ad
h+0SWEunAjP0NLEn/bT607Zr2V5jwSVPvbMrcIjeqR9/VWn0kBZTy7z45Y9hADF/
b/PRWZyMGWA/hrJoj4rAB2ckFWrxG0EJ3RpEh+MMfDXvi6bmtcylSdClN2F7wgPi
XREprGX7zOTfwSQ2Le7bYm8YSFjlOk/womgJlljNXt4KnBwqjizSiDqexKZuUJQT
+GgKEJ5U4TvtyESVD/kuk6emRC3oL8QCQDgWRqc66W6sdvAUslMV//4zEMeCyrFt
kNNySWEJ8uOQ78xbFG+fOXtToNYkz/YpM3oVBN/2SHiRc3aHyteNg+MV0BVIaTy7
ubBVFsSoAzCYbCtNALquPRu1gzOo4mcShS6OB1tBGveWziTNbpC+YblSsvsP5kXS
kjrgYrgU2t2bGjbgWdIW84G7ZeaUq54J+MJLkl5vJHWAzXycrW9cKK2HSq2hoyve
fCB7n95Y4TAR3+bnbrP/HiDpZr05JMH7wEYjA9HFhdC1/BvAH/CVPpxDu/xU0eCD
5XP6hHC6FZdKpf0eVEoJzgpJLhCQRaRR6GUkyDB2gHq42VmIt2VCdyvB5YxLyp4N
RN4TXRn3fXkYIrPpzPWtRrqBdJjm4r/Ikgk+bo6xriAW4cn6hmIoF4XDxaCxS8C2
vWtqAWukfrwHS0tDEzaTKks6du/gAqj4fsAjR2PRyyLmLfdDJ0T77kF2H/DQu/zS
ViycxELTYL6RuAsJmJxa8SUPG7t6NPUgs1nKuApnPsVFvKzPZ9GhPUCvyiLZ/8tg
xKXUZ0DAKG0Kr8pSLmqUDOMGhD44YDpa6eEQfqzR6BLK/x+Iq8oHFoUwRCWkbSQG
g5y6mVANDDmllRBi/T1KvpaAVP30PV264OUrw1G08jzzlxEqfnKVqn8DAjJdgDdc
jNsEExvpakuKSwMskBjuyoqXgl0QzAROOiPavSiyZ2EcAPPX0sVEB4asBscdtQO/
rbZoBWZpkIR9iKmYTMHbfKpw+IVsq6Rhg+KuSGd3LqHRkXQ9NMcyIUvxCWm45WJE
N8Pcaq8cSnMR2PtwACO0jkJjnSAZxEhmPW7I3Yt2QPUwcMRUEq3fMY+wb8VfLRtb
7wkHJe1eN9ix6NAlM8s29hLrAN/VRpRhBY2EeMP4wattHhcjTvZnlxQYtEvLRmIC
7nXjCS+F4pZ54ZSUmvUtB2S+mOSbQa3yjtF6lFOsnpLpzPqMpLBkfvP+477XXsrZ
UxFlR+2s//IT+GYpk91t4OTdHyj4RZFBWruKkQ8T8hP2UzBNKYXCSRrUuG5Hn2bk
ZBb5N+aFk1EqdfJ0+N/SQAU0FNtmHl6I4uShdYcc+4NITuvcrO7PX7ftYsUUZwst
oHYN/WF66UrMI9nDp/2kML0RBHRBydWVn5MgbgOyywmPUjeeK5RCqkg9vLdiyDtq
sxq61PLPIs73Q8wzH3YuIcvzlmAgrEsBgXJgHcS2uY1jUWeHmIH3agOohDoiN0yC
aFGleabfnTvHwnQ/zlCEqLAv9I3i+FOec8ey3bhV3bqR2o40g2k6sKQW9KYoZWdv
3HBzGY1lBCSEf+hP6c1+4Qkx4KmU8AES8L0OKr+PgyZf3Hrw9s52j3phpRwjoETx
5h2YN3X+Oojh8RBhsGRN2hbwonpjIpdqCW+DopJqDdRSs32TlAKNEybHpiHjw4Zx
gsZkzOti+ThMTZoZ7iTwwLR0Z4c3xWVdpEPqOdwcLKbR1b0ZkyCIGcCfY9oeYnn+
o+FEC0h7VPfqDTfnOsMzEK9x0g98W7GMrng0bCiD2cEv6nzdxWOVZoGxWju1iyW4
265PP5eDJsEgQ6zNT2n3KRO067O3MqK10u/jVw862MB5tefm272JqKGK3qRh6cOK
/o0EfEsnynyYudncA85VHSIt5/Lz0I7N9m6sd6b4xXKcQKDWtJK8Wk13UIuT/dMH
1SAZBvm3CXfuQlx3qN4pFcUaVp9WXqOPs93OGqXnKrc4xQU3WexFm2PqzIO4K/Vw
J7c5j/VXxx1WbhRjUP/OXJh/QKE9Q/P/ZyKfhDyF2Yvg37fb4oszG6HVultbYuqp
r5IY6ol1N9kAEHN3iWmMPxMk/eSB0yhaOnCCRJwSsws4EdSbqSKjw5QXUuYIZ2gQ
6XZojz8+RbM7EKiGdWaxfmbtiKC3pdBVMwgjtvQPdmfv0bCldI/BDQSzBs77U21E
TKM9DmxBZjBnZVAVVs/pKhgzkujVqWUpmr5icuQm/+N17THJwpdckAPdRiWhKpey
tQqj9+7qL6z8VTWFNfgxWjIVHybEcuD7nrTbp95gpQn8g3a1Co3Y6oHsBBbKMKCD
QGItXhm/NkqBnbwImCI2t63Tx+Hz0JJBSyeOqqX3XsSj3TtcFPoO9UzvO2ctfq0p
KzhiMvrEH1Rf2gs0k6MGqg7r6C0Bk5RV3pp8XNUpTWEmgs/efYA6d8UijTIzu6Zx
OA3eKIe5RjztO3uYHT1sMX53dVXaICpr8PuBwvgueY9wgkPJqNg0vfsYfEGKo/VZ
PmZ3nilNWLImfffFmmpdyZMECHYysw7k8EBQ9XR8m9nQ8vZ2XDXDzLZ8qroODFZ1
0VZmU1BcsHHyUOR3xsrSc5sI/n/Bn3wn/Gk8CyFN0aVvQzx+5NIXbSJnR8lK/6Lr
SXkgNs5VWwODHzpral7Pthfr3XiLn/aN7l0PxcLgwoi2aDgHjH4awf+Q8sAl/xSi
7KBmdzu1mKZGg1OX4UcRRGurIlvxfu6EnxxmOecYbo5oJhqBywBrVX8HRJLevEmu
47g3/p+hqs0ZOm83iDcja70tulGwE600FILkDsEgXNxn+CCNW3IbbR4OqaVuvxJq
WX9kW+kjd+YbEmj30zQfMshUQe9XEZWud8hgtpfx99FLllMYL+bN+d+etzlN3bJa
UPUkx5S4HL5iQjTiel5w2KxIgpS+CcHLBf74lBGcHZ9dvpULssIa3AZAAEsp/+cu
ml9QTLNGf8X5Bp8vCgE7JpqhdErvkRi1SYHidf3jQq25HKZt27xu/wCwekx8oz9a
g3i+45jaq8u0RU4PuVyvqTWBFzMhbglXfmNS0FdAVBc+pKlqqcuL/p4XuqoQb/JA
KC14Z0zOXwK8xIhJT+O2GzeuK54/9jveAdtZMTIQMzxQOdPmLh+ekoLbZbHyPgF8
qqBc5mejYoWuCdR4xxCj7dIBU0Qp6MgzPetiW61w9URbnDPbHxUOubTqIseGUF41
RUukT46jmMR0JLiQtPmw1TVnmvEkH5MVde6XuCUXgrpiqarTEjX1pGteLM6Ak6MC
JA5Rx5sQuYaGPsglSlQopth6MTJbTpdPhp3LpoG03C1x+WtOzZEny2FT402vUm//
oSAyVPy3fdiepe7G0+1w6WzpwaO3qVWuFdLKwYsphcsN4BQKxFw7ehFQgRY97cCs
lT4ME+KJmtfthNa0d+kPpdPFE8AjZKLyYB9Q7p8iTMMvwwEb0d0FWdwCZwOu8v3R
MthNfqIMi9Dtzly3/vOFVe3y+cIndrwGpS/KtVysW+dmdvdp1OcKqR3wUTf/4hud
eSpVPPkY1TjFpjEwAkXcDwaPojjlZyZxu3Kv/oWQjqbmxa+uMYExUJLVHPak4wzG
0rUmcwTC/5kGult/nGE24nPmHhaV+VBROBoImsWCzuS8eK/l41lYXAmDmPok8a2y
WhM3g/ixrIZy3gm5LDQQt4k+7tpDJFY0PIk+FyrQAEN0PiFPACqOLKPLoBYrCOvT
XE09HaBWgAYXOrJTB3n2wp6T1uxRZGpQJ2J/YHvlDmxElY8YS3S8yePPmnic98Ag
pUhac4rMf2G5Yn5MUP/xLbaUy8qiv5EpmDOjNnPmlpAfwApACmIyjS/5gUU1nbxU
3H7Oi0/M4SG+1PZVcxetV+HPa5ekMU/DGWYz75RL/SlQxVM64RywWNFFp5vqCYnq
Fl62pUzAy060G9ETQwMpOMXYl11yHk2okJBaBGy96QIPVFxjT1INI1mZdKP2HuRP
XPq+FJtz6smVahZo14TCq7dT8hL1A5vAaMwtNK828zygXNLyWMet4uJCFy9aLqjf
9xE8hurLkubTT00tCyqC+DUqo3tEoyVI8W2bCW/+mdiVmhmuNDWNXp+5Ulpi1xYN
ep0LwhmRDour9zdNRZ2BpmT1Vmb8RxMYYV/2UvrFE0lyPTbNg0UnaVn0pLwMf1RB
arb5vWGLHAfcl9SHCcuId9oxRZQQJc2EFKaW5orX1Wl6bFCFJ6rrwSQ/osarau/D
+7ZaShZKfPSnqUgswFvCZOeXPTW9DoadXvZpcg5jljAbXTxzn0VM2kGz3RUFuje9
jfJFoudAv0JZnbFMOdxdTMLB60pb3fG9RP3rNPFeVts8/Yz/xRJ9Y5qKGSoehOg7
J1NS4JguccjBklcceM0DQ9WFHFcN8lPPg2W1679zkl3beg2nhfaIlFALwzWu87iC
T7WmTGED/urbBjy5YTl/H3+m2fXo4ePURzkP0e2njj+x/Na2lPJs5phZSjSLQ2+E
M/c0TZgrReldc9x4GCdbjOMTEDgfbFDypuGaL5icrNp6BzmI3pwis+hM8F+Kx+V6
XvVoa8Q9g+/DQRwDbHVHH5w5fu13LJd9Zwnt2/MkabkSlFbI5HiR6qeClKwasb8f
IVOx0SBQzNV+4oZ3d23pqbDmInOQSSPiS2ObDvyvrKIlbQKteDFVt9SUxOXj8lCr
f2uZVINccbq4fLt9Ffo+bE8lLMnL2w3YzdNB6TFteZPyTOiK3Z6SLbsDyT39KyP/
o7jf58fjn0MEDF7Q5mvyXeHFLBDRsd6c1LRXfEnm8715wJyU+JsNZa/rODngUh12
yqKA73r1qLfup3ojwBYeJpEkkd4lE1skdwex2o1hQ0rkNYK2kYFVCY89ZmB4FNe8
qUiRneXpxA1B2TBX4WcBM98BnfPHv+EJ9daUZdEW402tWNOXzZ84O+W68CBr3Jxf
wH9RJ0eRq0U3IY24W2PZsQ6qCUnGCPIKYBWEiaAPVkvuVzHa3NHF6TNX4i2GkEdO
HOuEIL8vu+UF6kz2rzEoDKMfQsdZvdLevPxpfLbUiQQi7NXqcX2sU9GIj6TaJx5P
vykq8VOjGh2sCVRZQCKhMAtf9XhERKPspgKs6V8IZU2cZDtrvLWZsuNxJ1LmtH7Q
EjsxrrRenswXqk5uK4gTRC2u+3/nBDAmRQSzjcK15PWncV140M89HTcGx0lzdSle
2Xts7O/dJ21Y6kiRRNbdb4ioM53ihex1StnNtcYQSylE4umsBze7/BHzGTu0EIXJ
eWjAC1181JlUv5A/8rOwfnvoplsBLdmv8ygayfzo74scTLdH6TY5xCuFiK2Hm7Gz
nxJfdIkl9WJzcACS32++KQVeWQmtxJf7mEQxCY+YexacvnAJz+HdVsN/EOh42Dnm
yXVqjOAp3lBq74GSLIUeovdZuLhwriWT7aI3gvaghq6YoZyH3GbYuDTlJPpK+76Z
nWtRvKO4iZ8XMqhORq5VFgqBdqbYLi4PfRZstZBHwuOEs9/jBpNXj/pf1WzDdz0w
topJqr2s8me7XISZdOcZAfTPK+BamF8O7PPJeR9D9fG51GR1SIZSshgk5pM8NyHu
aSXjAav+y9NK7pHOq0NhfxILEXGjpDPqTzV5Cz+SNCH1bTWfu4lV8prGe+W6RB6m
b0vw6g1eEfvavFp94ZdnSadnZFe2LfQK81ZiDWFoFKvvHlfvWtdt3Wk4fX95bMzy
4rovv306e2dG98v9wDRaeFPLH+7rQI0LsdDJ9Xh4Mw9cNCNM8lk4ak9tSY29icVR
mXswZLalfA4SapqsCi01EwxbY8nAfjYInnCwGDOW6Zw81hT4GEe0E4vY/SmfhRyg
x3yPutQkOEHCOCig4Lg2ppBwfGibVlW8KUq5zW5DAOFJPNKkpJxDQYvxEmw5oEto
djTGqGy5MdBgv4SDZZEQbVpRzSExHIZzwg19Sz7w6o+3XE/ZzX2y5+fmF2wc6jzU
ndhRpUxc6kWo51fVIljRNUkEub4/0ESMCAuohXJl1SPQdtF4zhzhuewwHhcM1PyP
1nipwARlEjFUTUYfMV5iNaRx7DKBETnUDoM0Cvnk4UNaEuHhpo6WjH7MqvBdWP/J
WTxSiAsft6gllO6XyzELn5bn1INNThp/9MxUSPqcKGhZxRCZ8BTDAK9HHf8S9skZ
yYQOHPkzeJRWQmVTjdtw23Du/1QCYV8ThIJGoxnQYTNJPX7Jkk3/x1Eh69QLv8AL
0b4iurgqbHJeNrGZK4ZBOFLu6pKd+anaxObTy8kzG8Wn/IH0UdLWusCvFGTIsjR/
IXYiooSgNfwr//7KcJjdmRmqSTVJa3UWq3ClLw7J2B6ZV6JvhuWDhA3q9jCfofPz
e5VRyaxfNqzeJ1l8KhIEEPMOxrwitYCf+OqGAYeZ6syc0i6epIBLiCeKoqMuzGco
mfX9j5f4k2Zx85rhEYVtdehRIjd8KNpCj7HL9jaMvNcpriDPBObr4wVqkbX9i0Tz
JDKQjUVzofpmMPMIPRLnmZA2yzpOJsfgk7CjX1LJmpzNTxFmJemIizpOwD2qWCKk
S67RJdWv0q5dIWl0fJZuujvwPNdx73jWzkcxmNk53HiR1l9tJieTs9FgkYqCNiu9
BGlsnV9KIkwnoPVhK42ZKyk5RZ0gGJEc7cod13QBecnrBBA9inXam42wLr/RrjnV
T1F+LRo8AHJdbBNJITEmWn//lB2gxvb1ei3qb8ziCb6qinidUL+6ZTNZFp/El79S
uWgekW0awfHRSIEnEBHjqp589xaNzajawNFxkKSohQ+7vVem1o3xEH7/unsdcrlb
CCz/q5l9A85mBsW7HS1xbC9D7z9BOHpAyO+281ckZBmvPgOcB/N0Xg9gXQbn53N6
rVF/NavZz1QbvI83DS3dsd3xd/3wqTw/OCcaGhc4FIsXyVsWWYFMq5KWOmUhA9O4
ePMpzCffFyZu3ilZIDVwT5ITHya1XhCQ/97SjLgOOuUGbZ0i2Iu9D9TyD2Sf38PE
WLiRw878UYyGoFbZhkK6qX8hEKrMhBhFP5g2/BCH1eerhuD57sHNKG7T1zrl5NrW
M/fOUasFzwQaFcQ6idehB56eS6W9QOGG5qPWwCvylZFUmq38bXq7Tqow9ZHj1FzP
Rs0cpPY1J8w3PVt36p8qBes6ft5g2gdGBcaF1Iw3b3Rtghv6mAcwToMOPJeoPxF7
XiNoXcj1SkP9/SRPmOUq/0DYuUCtS+GPBawjwEUzOTaSrSfDhgj+A7YIB1Vh5js8
pFuLqZevKYlzV0ONPgHOls8ie1kcq5C7+aAO4haEpxluvViPm3jll7QabB2E0M0K
bV/eV4zBmRQs7nwA8enS8TYNArGd6Taci56lt74quQ2DKoSLFG72sPZ1rlR69fey
C9mvSNo9bOnHLHstljVEKMLH3uFYGQuG94u0rrKKPYWjX8ouTwSojFsEVv1d0jbl
Rfo0szWGP9KO7Zl9LfX2emzZWhoOuwtBeigq3LJ1FbVmLTujfhlSRiJsY2SKuyQZ
P4AUAkJKp/+AlkbsyWAnTljBoIri0jFvAzepU6tfx2icYZZwtibMzpiZQMkMCxgw
6ArWDMU8JX7T1dScR1MruyGm0kh/0xmhYJvtgZyXUYraoTIX5mXI+ZiQc9ZogLNc
cwWWp+dTuNB+U4RUgfSEl/BNJnb7WgNlklpL04k4NaKBstunCEZdWdp92qdyTCGW
V1WLhTk7tBGvjkLmalsh3QPSxuV3EO6h8dsOxP08MJYDnXmOsU1/FvLqI+EMIuHZ
zFK0lIamK3tAP2oHw9rnqidCWZMU/tLelheIsD5WJdEBiEzDiLU+0iaXF2oCxTnj
PVzrVw2St9SgOeMbe8gJ/cWvoZyAbkRWba3VH+n0IAbl0AKFc4ff+9zTQUydImQX
OQAdMCYcIFkvnS+JnaV0Ii1Byi/aP7mM2o5Ko9WZdyusYQqs93HANhqDrt0lAAsa
X0UwF2vHZjXTZAlPO5jAvMnRpkUnFy8OcmAyGD4ZBgfL8vtBU+zH3LDFSebksTg6
LyhO6nweFkQYaq2hNLB0R+EMqgiqYt/3MRkgISlLTLETNH003gwfzRI9gfoH6pwS
DB1lPW9pYec0Dolw6ZF3YKBvUVKrmRrndJrHTPEajf2dWhSNar9LcZEf6w8uOq/X
vZ5BEA8zJJIH+nQrDLbE7sfavpur4xOKtnJyJYwRVw91AVBkMm4x4I3aKhwiK2Oc
YLjFi3TilkdLh+8rEDqr3foRED3JPFVSZ7KT5lrqkFSxHNAlmXvdk4vABAGnVanO
7zosXscTApZJE1TlELZnxuuISbw8BCSQvHLflHN3xok1Uo8u/NLRlZ06cy9/AjIv
FoMnnWJ9BUOHjaYuxj2GO1UzO0HXiVo+pNrQDMGNKJtOOMBRaz3cszmwSPf1dnD2
IqtPmrtY/XpKu7J5CeVaJyQsGFchZz/8Eo9sdvLsTx+3Ul6PaMbeiD3TyZ2tj5ts
Z/XRF3geAQEj9LGy7JFHp4g83yH5IN47bibfbrD2R2xc9f0ZAUU+NPkT2teXyu4C
+K6J4PAI9ZciZYhl+wRlpr70l+9eL8CqzsRCi/Oh5opOn9fk9ayTd0HpBAxK34f3
VG3lveJu4UAOOQHsQtpCt/jWiPgd0FuJtbpLEI8ne0E7prGX9BrLl1qzZZtncvPb
csQWWL1RrYJeBDqwuyOsK4AKG6VDeZtWmgFf5WwhwrpmLF6d+/SSN+6AGz753P4V
o+yNrHouFXWXxNEjQDLb8NKCdxafRVA3PUXldSd74tfl32H2MhSaW+O4uUdHiA2s
Eg9qZ1gJAI6oz7qC2dy0q5g6gZzHPqYf1QyEqJ/QxzZ72i4+LR4Knu9T815xGT8Y
aslRjw/fmPw9drz7MkNBxavgopRdEMpP9J3DsQB6SiZnyzHcS7dR1iAlt526B0cX
pJD4sxc//O7IfF7b+6jBcAnnnXxkOxGdTemKzmKGylxFOUCuTxFJxkjqdrQzcO3O
B/SfANb8sGJ3XpQJkgVadyRsaip301eNKaDQOQjwuqY7K8jQYiCD12YuicsumAAE
xS/vxBZXjU+G0h/Uy+5uL8IYS3CAAyu4NIVIIKb8oK4nAo/wgGHDE6thxhS3/VAI
VRqH2WRUxPjGP2SoZ0ADW5+dAbxhoz+liu3RE0xTM8kelcvfSmQiUs+d2pHwPJu9
FORadtBMXlkkVoRIcgcgp8SnryQWjhoD2a4zQb6k2hpGuUgYMMluAiP0qtwH0/oM
GDcTfMwBnNqzdcnQnt9sGFpdPXaRG8IGqk8KeR5vORbrZMvh3Ww4GdJSHzVOgD0o
KaGshKZPPRmWp/j4x511OXHiXFOrpaAF87RRlE2/KxAIjJ474+4HS2hTnNxqVO9T
6mnjFTid6djMHBxzTw7vO9UpYr62sJsKL8CJry9w4Rr8LT9N/YyaK9fpB+janmgQ
74dLBCyvZqmsDuhjUFjFgfWJZTBGWOLbX5aecEMMOc7u+1Qkt5gMj6IhfD1pJCIL
KPVeTdjoH8JMaGERG0GVsHCgirh+tsHlqNvFHdjTXxAH0VoQ5e/ZN84QKSaD7QWx
AHa7nCq7obPsBXFLL85SbUJ4b4K1+7WFQ5d3O2KFMtsqxPZ7nTgmC12BK+0M4Fwc
ocCBAD80E7oAtGJf3mwwTVMHm2DZtkpJyGPIEedSFtDxsqbbIQsOKWjddqgMSWC1
fYznIoD4AxLTSdZiFZfVVQy+Pw32ugUeGoXIROZqg+ULNK0gg+LACT31WYE2/XXQ
SZtz5ySv1K2NJ+DGnMkiWVz27q+HZ9GAYUxaz+iY7+nT4o5dObDpKXWs9/L4xTQE
JpiyGuBJolye9ztmMCTT615XsfNpVhYd7hOFP5gAWGDPMqAPQJOLqZFn+8L5JjEb
O7M9kJoZc5YnnXrGObWBbaM5ZjhtgD4fgmVqucETU3hsaOtto3BnuS+A9SPr+XoB
Sjljexw88sWMrFkRALXVp7Kv/XVfgi2omk5Ga0Da8+vNUpdKR33K4ABRj9jVbN0+
4Rkspkr9b9ldmfL8dxh8aWkvowiOuyvqxdc7e/L7fd0lvN06HQQ4GyCw45wXBx0/
eS14aYy9aypUI8hV58D2Wc0RvcUVLxZIofn33D0lyrM51XPjdvRO8WK49GxCnk6C
2p++4n5R6qsc9IlJEvFFX4rwuESqXdKJMC3SFd5jRd9mSR/LXDcFlqdX7EuVg+An
L4j6A0jYM6659hvUfYVo2OkwBwWFlfShBkmQjKil34APdlkKf/qkfaomhzVprgin
1Hjk7nxgoNHqfaGYYCbOTowW8K6m4FhnQ6z4BvnlTIEw/BWio2Ftm0xJp1SJ2qfx
qxGzHE4u5dKPmGCm28/5RIdKpN8UN7CtVM0di+GLJR12NF9AtqSAacvVomLqhnZh
Dc3RY+rlLrHoUwRre1nME275KQiV1OT34J16Ohn+y36zIlpCPwncDa5nYemkDvDk
LNEYkmIt6Dt7xauYpcrJutj+rZdEyiWfFz44/suBnlUhSbV1eaOcHI+Nz+bIHeTl
u6dFQPCvUrBAHWzyoDEMvIJw6oDZ1eir7q8c9+M5glU7OZteb4H6HOi0yCIloDaT
tRvKoUTvrBHByTbevPbcb8VtgmoLtjS+iBHFYB7hHV0mE7juGwFCOiEomPJbrnpw
Up92Zw6Xu56Q0mDb3nTA52rfMcA8HCUBGOsFwr+OhPRTXUfnxljuJf+IxPFe9pJ8
t+hGbdSmyHly23L+365UEkKgtx10uWcDx4xVwLWimw8t1aNTlSRghjm7Divw8uCE
vSwwHpsm05m+55WGzMtijuObd8CO4DvHfXBgK6PY1Zud8ncKWDAVIKNvEzRUECDg
S4JdFm4xDC8PvaE8fedJ2rvPXbLDXLY8q30wE5tbpoiotGaZUq+k0ZlP29M7gNUS
3R4dmXwQ9opbivCBQn/MbZik4jWIpcmrCAndQJDq7K9Hz0injGLIv2uQe2xo5yiY
5+KJdKpJFrcB4cMWaOdjWwplf7+ZHteA66yzU7l+o99bBgfoSNIjhQj6fLls2ydd
l603g4VQcDQYb25W5Q3CHqWHSgIo9RaSZbzOxdLj8G8sgysw1A7sHXv7uF5iUSF4
nLK9uRKiNoEfCRAwkSfcP6AavBynEKROOTp1R6+GviTrdPFQh/jpxkiNu4NpR3cg
PlCErl8FrqbNgqjDIlINPttPgKnLranbFyD6IqsHAsllkwXddOIBJVZIzHiMFajP
MfokBKEYUcsCAy+jRyVFCoSRU/+apCrstr9FKAxwGyPFtFWo9d+r/9kEhdRVBOmU
9ttwSy/GA4gt/NFdkMXz+Ln/j2Rwgfrhr8i1LYkpFTiEJjvmNI6EHX2pp/OHXZi2
Sdx22c1o2nDclovJFbXefHC9lGrosOXWXrHyXOByeVMUNKRJ1ZwsBPBUOcf6UGiI
EI7TPAcCKOLMm+G3z0bRJc/mNzv2Xh6M7CV1wujULChpI3ryxEY9EY+f23aD9tqU
0tX43gVYTYxqg4s4JGZlC2vPiP9NHoaGtmgnScyzTiyuR/pKU8KmNrEmdmNWjiaE
LC+sUhKknmiewUeywjlmVbdac9DQaRk30FLUthrvOkBf4DDjRBVo0hPPAXP+LmCO
Yprw+RAFebKCplvJrQgDh53Evq9hPI7uiqUoxRIrB5cCSgOjWYHfLh8wrWOl56xT
Mxda1zecSyVUcCY0AJsRJoVRQde9gQoYYmjpsTB7EXb8hegIVfoUS2IttuW3TXkl
vyUWkTs4QaPJxObeh3Q17FEVjGdL1mKLrpz1gi+sVuTSNWaXzvQqKQwrL9T3cuLt
UixY4XUmnZJvZXncYcpqWkgo1IcZDBj/1EinpdSqWYzcBFfm45gDixjbQPHtDlQY
IZCnyrUt6/hBQnSwyGVdxE6cscmZZvANEOpJEn2uNS1Ea+BgJCXAs9q2K9yHp62X
Xnrt3l4X+b93OkkmKBUSlbYRdSfhY5st9XZEAlvKv9g4Zk6N6rPPrz3VsNabxKio
bKEHn0ht8GMAAy6tmWfMEtazC6pyWsP1Ew1QcZse3J4g7mWCmTKkVyGjOCUwBag8
AV1zKDMjry2dxqlC4ZGINn52MWBPef4ID745rlLDRp1UiDvuJ861fA0B+o7RQFCq
yPdoARbNE3IuTi7xjMQ5Z0nhLU5hIia4vaB2e6KAqZW92ZtZ4h+U59tq+LiCfxGF
CpoqAuLHA+CMHWUrmC3WqrJw+VXHrK/ZEXkBJS3bq35qQyK5PEqyC4VZt3dIky2l
HgMjn6CYUIFa7swvpXEP/2U1i6MNC6cROcmAvtCLW6rGCCn+jp2wB4ui11S5zEYR
TgGtPW/BSZtDROtdS9N2HLCrw+yRbXihNR1kDpLzki5JWWvrnP+4Cn8Gp1WuZtA8
6/F0W6ZueOyKyLAkbiMj3SA18t6D1d7ef3vPVZcvSSOyVXmXHdCyg/IOyFV5whR/
C3V18FMmMUAk2VvaAGgZ693rMJDvJf8Q36SyiTyZ5RP25oR2Yw1thoCSFzSfppWo
e9lPl1ijF2hSMDH9AGsczaM37C98vph9ORm/4uKTeQU4wOgNyYpAa4ygcZMeq3z8
7SRxqkujsaK/Z7wYm1acoS+I+rD/u/HPrseUhSf70z45ypDxEYvJqVwvZOD3JbYH
rYz2MraLqV0feLL6QB8YSZypTQgV+A2ZQ5L4P7d/zuL24AjJ3YtnyXsKeSusYLYM
kgUmC1meE13W2JyPVTEKUMJY5E+zgCfzITPmvXEokY2TU9637Ix31JYDda3+rgRu
fQlrRrPdNvyFQUJM6ukrvOZeA3hTylGb1tLfy39S5XtRo9I4xViRgEz6JZvraMRt
e1dA0ml+hJ5CY9Bdh7iSH8s9GWKFRy9hVCVe4HxXs1ZCKioAGnW5OavTEyiBrGAr
IgIV6g13YTYkpK1WaLANI7NoXlG5SM63dzP9xK8Dkz3ZZ+/+vlU+61la8V1Ct3iM
tLydSkqMyM3IJ7rNHz80YHH4orLEjOuhR1JXQqjUBbLLA5zXevD0m41LGw8wpFle
D3UBcRlbGJioKOWHg8RWO/p1Obydx4AyOqnFEyabsv0T8OKTtFtXH+iYfSKJk0ZC
SeGydfftt2ueLV7iMKghOyllWI3+2gyawFaxAQkSwccIc9VYlx792ZgAk4TNlJcv
rnzR4UDx0STDajEHq2GYHWCbOECq3pFPcgvV5o9e7mijiE4eGQaj00GnJp3kS1MW
SZpyrVkBS3jWtcaMgXTPdyJT9I2qlzpygsNsqBy07oajv4CimFe/JmBmvDmVlKwI
tbdDAErqLZkU+qyABLnK0WqAM+ByTih3B4pDwCtQ9miD2C+PnNMy1WLvDX4CTKp0
50Jnz2mROb1xjDwXdtZa+HLS5akfjEbdBuFai2RvAIz2dCPCVOlq85Wu/SP6t790
DlOyp4V9UJzSaIIp6cLzyApcpEWAQZ73u2u0zUeWmP7iV6pP5/LIy4CRniA0wiZV
QmPRgqM/rMdEJxdhU1bTLfcoYHXfDJhqRRr4EKq8K5iASXBm81g/VccgzdTjhsu2
FCQ/pICRyG0nVvbb/B+0p2wAZdM3Y9cBAP0WMUFMufsNkWhQuuJ5rb8x8QeDWtoX
WSlrp1al8TcU+KPZmHwk7Z8Rl+iG+bQfpCtwXpKQgwRRiFlgMSziq8DztW6HuxHt
RMjry4gZtIlsfJas+gdTXGO17T4T5u3OD9WhYXy7eIfLCZGMKgSFwtJSFuLvfIv/
Uyx9e4MLQzq4aYOQkXUOQGd4GHnE7EsvPtMdvKJHVLEC7b27OjytLS7DT5hexnZO
YSDXMGTLMkwTRQlJKy5iK+D/+EUBz+3Nj/B6twvkC04THuY5fuDjQMO1x5zkXYmE
aA6eU3JXgPjtUAVXNl8kIAYkRJsX7P84b0VFkg/TLXVO2zshGNtKAzFyasfJ9KG4
GrqbjBslSsTCrD02p39QVK+nS6mwNxun10lnvJf2lDwRcZ4Xn/F4TcOMPHiqzxJR
eD/gxajoAVFd8WHHAXYU4BOJ5Bt8eM8VZE5nDNO3Q8GHOAs+iJbN8X5eEF35A9Wl
Qm870eEe1jsBYcstHrOozvNUhI1wo97aT8I3GZgSizztL1/nT6vLATMDDVFRPJyn
s0zYTgvP3AsiGWriuflUrO7x7P1Zesu0vyp5KBtVwtoLIbMNF2eBKsOQpWVkoI5X
2X8Is2UnPs2lnlqX9+9ZBuZD1tY8/4bJm755FzeDopoYGEea83ZUj6orjobstqo+
fkDalN3Seey75nPB0lYoPUotj2DVxpf/fdKJsj+Nv5+D4SQHInok7D0GpAyWKGxN
MZKzOuDCwFL1i/AycXqhMueXzWLGqTOQ8e849TB+l5ioowlp2V3GPs2jqCWZZCrN
QAs2hG9moDntMCRLTSSy4hKPUiJhwUhAvi5D/PBtEDXbIU8Ir9ViGp8gAQAtomIX
uX8iLoznHxuYIGFQX1YZu3tLwMMYFvbEWvjIGVium4K11+uEkTsW29/6m80t6dWe
CQ5mclaA7PsfXXzu8LJQjlI+fmQhIOQ/IIzt1VnDY1OH1ORkFSEeMknm1inR/X8m
cwo+3Obh5g8bPKQX+GvxF7BaIO4XwxIuI6ME4oL/tqAdTvhVqgg0iyL8NFy5Apkx
qhC/RTe71tQwuZi9FeScW+00wTero/mm/3uiDK3SFgeLBCPe5zeWUzQESBu5cAV2
S61UwczvR2fqv8tgbvlzruMOXc4RijbqhQuZB2lUaHUNt9i7R83VFtmvhtrM5CLG
LGnQ4oTsZl+PrfaElVctCGH2fGnp4R1C8YBs42bRazc+gf3vORBLxFeiKKPDzWwx
lVWtZsMURrCG0L3pe5wY9OfYNc08t/5GYIJ1gqVOvFC2agNrYja09C/PnSDk7xKy
A/Di81jHosENjGK0yCBI6r+2qxHRlO6Fd6vuMwB6RNTcLAXa7sajdlNtBFyXBcm/
7ny2d+9pAwFn4pmCESG53pIs8Pytj2JtQWmr4Q7N54w+1n/TkKOEqyJHaWYdW7Ng
TaKITY1lLQCgIqc84xYugmNmIKaq08XqR9v5R78evmCvkKFxC3eabngD+ODL8gUu
GYnut5iVu2rHOSjXFIFJz+cMbV/rsf2wCvFZC0ckaS2rWoV+sWQycGXm7lZhI66f
BEhN75LPKBtdjIFPvXAhttL42wpd+7hJOadhkFasja5AsRWlbwZy6fcpRaozhS0m
xOi5szfw2NExp38hOSkfivRVY1+z5CQBXcHGL1/MZ4Rj/tmUx6MQOJXJixtX6PZN
djRnbf1xqTAq4XuK7gA95cFemy56rc8piQ4fwBsB7rGa0fTDmB0lVHEAHALvPPuh
hyfQh4bAvotqz8yz0UKLOH6ehlN9AVrJ7uPbqgZkQdGcZaMGdFsU6f62EvJEQxMZ
5DmbzGD1Ht5mBxGPRqdTd4xjtIJtCqyAAyGD+sScC8C4civvEkPtVztFYPdl5/vw
NPG2viIdf8yqavIV48OYMnm5nqqklXA2TSaDJavF/Yh5eMmt3ke5WR/i9N2UxlY5
cMuwaxdiW+YjeiLlUJRZhkiJw3O7H/84tvYJru+PgUfVPbXaMBRbW6ud22RhDHAF
TUhbJtunW2to3OQmORJ4gX3dH8u/R+PZInVzKQNVggxnEucfjzyj3xNK+2hBLpZD
Pbnvs1n6XheAJs7C3+Iec8/0sP5GCLRLegu9JGA5LAaTBmlUIk3aY4hPq0vP/J+J
KukY60PXNedC353YQ67Z5dexmxzFG1YQ3N4K/PAoESMZ7c7PhiNAI2HJKoGEiDyq
5dsvKefg6zJt8wFT28RehH2B5YCCsIZlmkchrv5ubaYPuuNOL04w47MUlVBxXpX2
T1xMHkRwree+4QnJWi+ZrxJZ5hLqHZYCHXlLLpaew2fJdt2D2L+3+yfwsVAGhnB+
EEKPSxpaD1TdTujGylxgtVXNToix4u1I8JmPPddZxbpsNYOv6/Dl8+q26X/tChtV
JasJOjl7gYpljpGIZO5FV3fAeH+i5boTBAwI2l2wjMTygFCuQSYiuz4uRf0pp98C
JHcCipgFeEbpX3SNmXIj5uQ89JixAYRGy7KnDIEm2dVDpbr2cod9kJZcudY0EPmB
3fNF9eLPF3jMVLBmZyU4Q/YytlfgvJGHmCK0dbnfi/n6ZSFNOQClTeUsCCvQPlMG
+kKc36RYusGoo9538p69irlL2dkYxoJh8Kx5gHHS4Lh2YUcHPdZVCfJ0MF0JiCIQ
kMMWROCBWKHoxkyo2k4UF/vf4o9+2gKgCnOJqc2kK0hBJMm7wwdtq0nUknFBulHi
a/IDVacfJoplO1a9daf7hbO854fLXEJNWm5Yi9wYHmnHlVDkew7i+eih8rWNNHrh
KlMz37dH3fmA3Z47GJ6aVWkn7NYvLu7ItZfI/y/3hjG+S8F2zmi+MfwP36HBWhld
C/j58fTArvnTK0/PLzkOR5kgrewqw3g4yXAfddezVxUNs7hIYI5qYjmQxJq/Qqtk
aGVwkBkUloxv9VfcLj8QwplemYRXkqiiFBmLEWwdudTypVYSAy4h+ASS+N/xPJB+
pO20F79f1YQ2KvOUMf6CYtzb8WAhfCUmVcJIUEkPRwxFurFLDxpxqj1HOroBSvoM
9R1VnGun3pEWQdVxBFBSvUygijAoKKKQEVCkxq9OQMsNPZknXjly0ejWo0k5L8mT
XYpWrny4uE8SIWSgMiCLvF6GBY9PIivklI5fLXNeih66Ed0uv7wjdMWbTxctMTvY
fiAJEjw8ZLMsJTl8lofbYXrbqzGRU2ptgRbbcymacqWbpagie6wQPk3kN7EwDgpi
uiGXuPwWOG1DM/Szx6GpwVT+V39rt6HHWyTLBRjPi1ut4VPPWkQ4RAWiEHVThYY3
IL+0RJ2ahQV4OKX/JhoK14EnVIuyq8NCPa3kZXLknP745Qj9zkdRWcRRIZlT92/9
++CubUfX72AFEe/atx5ddc10fSarGlrSXIkQVurBK8/VTBm96NYYMfcuiFbavznX
BZHOKQJviGg1N1QZ3ht0t7UPT9L+x2b7BeF2oo1d7POG3828H30Svs52c3pwdaZ6
uaeMFgNNagmmm2eADK03plkwkJ999Mq1AY2PI2pBsOmrXb0weyLD9ywVj0dX2fYU
YBsb83Fvinnno0zokMxZnZAQjbT5t4WD8fVBH9jMQMCZYmqcbQopYiX9p0jKib6+
SrwTYtnp2/3cOt/M9iJ57+1rnJmXeqXRgI3toidzP1tln7pXA1zPCNWNxLzi2oPh
b80zoGnPjB8IH1ee/XEQJ+dUKaNlg1CIP/41t5OVzvbuvaAlDCJZ6wprRZv56o1Q
fasZGaX1AOu8FpL6ezzLpI7Jr4ftx9By0t5PqqYnPN25FeUksdsBEmFkkEEFV1bl
e40sXjDnQMl5iUoD5xFL3NDDm6QuH6osI2eIzd982uwbNWKliWig1DySQNlqDRZR
WAPmgIpbYr+MUfRmc6T+fUr3Qd03IwgmFY3OnX+kl6WvdkPddoZPpwh7830L9z+l
9J3AOUFHzlSNpwR4Yi09J6nA1QyJz0ODiENnUOTGN0fMjjXh5slE4p4vv9DRi/lr
9HY4NQFRRQWPwrdX9z8QdVYBiQvmlu10GszS4myRLl78UUrNtZkkQDsQ8O/GbwxB
hfVBuXqZz+2fwHNLnSVycbG9V1sdw5gg+mpKH47pEIoM7uJhirLv93WXABuX783/
Iazinp5hvpKrAjzPGDbzE9i1UzXr9m5pULXEzIWbNMV0sCHLi6KFYIRe+bFTX7fL
dPrX5zhW3iJ/uKYNNtTUcPBCmCtDPFtRDaJzaaZQl45aqASXCprPCdB5SyLfxhdj
koIF+VZTTVcLrI5dNmQYBM538wpajcv2g7XK95+hHk68ku+VDLqlGOCZqoYWIJlM
5BzDh9ecmtJ9rHihQpNH6rFOGM9B74zoQTzuqQqJzOhsrpl4CZBo9RQ2rAGGIoQJ
yZX0qJuUFd+iV/zYt6z9t5oSdMtciYeR4o/9DeWQEnZQJD76JaaH+uMfnJvZSYxq
+r7MAD77q4o0vx9r+Gncurhm7zXEeZCfZMxY2aJPasMrL/tjcWAkbXYAxOVVIsZp
2zSttdyS37Gu1VzZtYnO/YW+NBcWkjDTz6Dllwd/eMH3GJTS1lc4TBNIDIXwEAUi
4ZGsTGlIYm4RJeh5Gu5+/1g9U6MhGDYnXzNlA/xLd7GIMdTXlfck99iuKSxYbdfy
exO2GInUyDBKypdr0sE1r4RHoMn9636X+9w00ozQ8LmV3GvYh//6wi5czs3GapVh
F2MCH3qSQsbHpVKQLpiiqoa+UTYVGo8uRH6MF6kGx+FWz7G+pDXegcC1rpoltAVM
V3RaIfJjxaFgBRA6HR7fMzwnc5UamOsCDoLazje7caIGnEy+tnGmq0EXlpB0tyR/
loTLQfGSJhhpKVF18PcOUTg61Rrm+jFHYSPz3PiAPUwG27Dti9/Uor9q3ec0k0i7
7vxlTavCRP3Rgq3omf3FeoSD6lTWv999xmJKh7q2JRf4co/c+akkJ75cIWizDDQU
nlEd+SOztZ50MJ4Tpqr3Z+mJOUCeAr01M14cw30K3184a7ybd8o2M7kYVHcvgZCe
uqb3ktpayoChyaHcYcnY8sS89JfxzJ0vBPdN7GC3dGCkd/6EmnQyzz5WGlTJU+Gp
nLzY1KL23+W9CC+cJ7l536kYNSMsmj87rngDHbddJriU3s4CEwxZRCcLa7dOCfd/
rwyWm2L8KfahUC5l+u4LvxGus/BoBrwHgOLDhL9lHmSLbwd8LZ4qAz7dcETRwepW
4xJT8gVcOaEx17F1MLHwLNAVqMFs0hTe8g3RN4vhBxK1NCXDqJbHGytyIbRgUfhc
kK6W2oNVEWq1U4RFRC5moe+ENH7ZCatbHrbigb0OewKawisCy+AsZzAXpYUBFkiY
JauQ9zkXwHJoMFIj0bbhIcuX9VtcALKZJUpxbrCN1GuPETu1OZ+H56C1cutbUN9d
C4bUd/oIQtfUvFn17zL6geLh1oXxcM2GZO7wSXreQSDFh0hLxK0oYXFXXmbnAKGj
7/pMPat1GgI0uuZPTeFX/EaG2vUKfSkZ6aMsWrDPYS7usHThXWCn5SoW9GaRPBKp
YDeO96qJgueHszGchhe6jAvH+Y60EAmtuW+6ioi2UcTEMYJDahlcO5uX/fZCFbmN
P3sePrAUcs16SCFuy0VYKQKq0aT+LDtjZbNrKCMgyMHIBPtNTq7aOoiyt96IpemL
3DePVtTjiy+JdE6KCg19N+mDAX4nhCF1nmwOiir2lAtalzhlfEvJY1+aXRAM9G+e
Dn+xDzyq1XNeWnLixgMWAUee1NpMSd5XOIQjltJqyt2390QuzQAzy2Ow2+xIfS26
KUNK48MkbFDhlgr2vJqBiCCMDCc7Sg6h6VNTrqJwMx4oBoSM2rwrEePJ5FKnf77z
gnq7qVNlQjOx7B7ARUmOTAu4gU8j8y/hEITJ/ogIR4P5lHegv3oFCQaPVL7laPiA
jPVkxvKUq4hxPPYuA/h3k36RwlYrjZwn6zTlm1q1AzOXKjQ+fPVC5qN0vuNLjk2T
hm6CQqYjjJdaaUmQpdqZpA2gKITQCbvRSI0gz8r/cjfXDrWBXfCKFHgo9ik/i23q
KJaarLPnBKxvFMyL97mo7H5tExs2g1ltia3KSynbHGgsNlnqWYnZWaX/p0ZwfMeW
ZrgNh5PoPpw4N+QK0SdWlbhXfnAi0oTwNfBIJFwM5nKHPLkV5h/EZeXXjfThCcaK
sp7Q3iKFYYi9r2cAqz/rNmpQ0Hl5pM2u1pVv23AFXPvaqg9vIW+OPae2OGvtGpLZ
YcqDXkK4yMJV2ffFpfRmycoeOqLB9XJgaKp7YzXg4YS2Um5DTLTGaV07BkTkxhAg
PTNHFk6TTItWyPcWUg8FD/h7M34pEl6cTNHfp1QL5BNlNrgdCC4scau+IxTNG0ES
k3z7vV+V8nrYajQGaFA0d952xrNQhClt70eyw/741UTuwTYphXdjvRwI9NH3P25c
gPqi4L/Y33s3lsh7MPqFE99x4bc0HHd7VeHOTlUB/OqxnNaUXr8c4LzAeWktRkWT
Y8WmA2mqzbF738dj7nXFI1JVV5kkTVvX25NdnxsjafebUJyi8L2nWzaC2+ylUAKL
wAN0i58rLcogXRS1DcQuvIxFYjr+/3OT5IV0rUbOwaD2x1onraQxSpxZt3tbZiLM
iY3q7QbQZQWYHEn+B46dLM1+RDPDA84j5RvxNozx2V3w0/UnKcJlsbiZMx1rGHSM
g0RQetusJ+lOrCqIUSzVSHC8TXxaed6BOc7YlMP8azup1UqJCuvwEiUOZuovrKPe
L555RtXI8TCrrJm7rELy8wtflb6vI5dL0Tg7I66W2n9H0SEe8VOkcUqTAoI6hz2+
ByVshm6iRd73IAd5VAJIeIaQYJSdzs90wS3jeQZOwEUY6qLALkUO/K9UgyL10ZUm
Lra44FVsn9OIC5TzbDNlHFUC4FjTUd3ZjUlbFksfchP/5uG6ZnMjpnNnrHbIxMkO
7E5umrxK5ArIq1MK+sw6+1qIRY8aFSo1lX7VXY5rNVO6XWcwagyb7FD/jOoGAhDg
cFGsB0PUOZWJayhTL1wF3qQxddr86PgcDqs8V2ZuDeZsM7lYzc9KP+dNKxQWAz96
WJUkZPFZrxvy8ESMHY+Xv7Pyt8AjoohQ3ypiiGv0mYwpbNCL/vg0goKl0tLL49Zu
j7Td62/6BEXhTdQW0fa+5ZyKPbnKpWC1EJwBD/qGFKDk8XhU41RO1bVDAwIanQxd
xNuIIZjWQBcwJl39+qcSIhERMBWFa3Mg3ZdNvepcLEWJ6w1P1YdPda3fpGA7hgM3
2t4BiuRn4uwOB9TLWAedmb7Oi4PsJb+adRQZld+8B3xeJgHkWofAACHlqcWFPg5x
PXdnue15zdl7QpPoy22ed9BWF06SD2GomgQT7y4UYHQ4wzLUczBs6LkMUOqQxX68
S+ti12ov7zKNHuBV7A+kRUAN+LYWI3CBqAcTuUq5eK1m9FcVuo2XouAfR7d3vcKs
U9AqU9ZqKQeNlvz5tAeqWCqF7YSBT44Ndy5yVcSwqA7KRj/pVf7lTSJRKyKYxTwW
kIsVJTUT3b0UbFHXi1ouTw5TVpP7Hz9AbgRomePhxVVGSZ73ojKB8Nq4eyUOqlLX
u093aRM4mCpsRe3qnB42AaEa4tFv8pzF8ZGmQRmIBph6XmXrxLBuI5GSxWfZw84k
l5WPqnuHqz106TaNablB1uZFUSQQnUvfBMe8hazo6QJmBx45v3YS/2pehYIUkzKh
W85tfJexg+HP7m15e8Q0FkvKHu0tCLVo2a340bfn+PGKfJeeO/3xhXEZtgXOjNP6
SsnG5bt6o23f4hzmRG2vmYL+1ZUVBNkXwD8ho8fGj/Eo62Dk/7F39qrLLl22r+Bf
14u7v6eiYXuLzZ13jC20uXpa39UWvAugvtkMTuhJzxAhku4xP7+AtxuqENKy+1I+
cELtb6nopeE3dkdF3rUhiOQ6TOGjjas22Wt04+V2+xMIy9MQ8E3rkbZchxZTO/uw
FRN8gIrTw+rHLs3NVX7+Iz4WRWwCtdAtFW9FlZQxpKD9bk4BXj2fGplHhsVC6CUc
5FwPnibj30ojqhe0jLK1za1geKK2FeSxPY7FWBRQFnSmVhS6GiV5dUyvKo2ww9nJ
t4ChIeL9JjgPsoGKvBEjy7li9IBafgL33UnIo8kYqzrWk3WG6kfN8B+l2IA/NJnv
IDAQsxBKOBq9COzm1b+0vY/vREnfvuC1awO65VyM1L2LdMemItALmn5CoDvLHqaD
DsK4oNpIihc409Fuaby18znEVlnVoUwDMSvZUkpRBKjnSo1aBke5UN6qOjRNijqA
pHa/yjJjnocJu90TX65qJMvPQwnBVp/5aGk4GUBm6sF++zWfUU+WVATJP58wxTDH
adOKbPN1yxP+si49FB/Px4jP+u6HAw91Y7YXYGhvsDOQaFctka+Ustkmc9Yv4Yun
aaaqlU5aKverf2dpXXNw+bElZVXy0PLjRIMnljXIQ3pVwgwLq24JoVqrxegZMDl6
awH/j2KlJMbckSS++OTAwRiG3voTxM5/CtExC839jzT8fsWOX+NRIKSeYOKbS1t/
guVLQnp6bxYX2WkKrtZmrkeqRDZO6FBClkpiY9AaCm/M5PmNUw33Kiwe814IkgIi
27KtdaVKo12Lsxo18/6A2XZnXXHzPlbA360V2In5GdIlepVJyIED8yUqgNCoVpUs
D/b4EuHpeMsrfFybbp2AHlFarpqHrfta+SLcFmTYfV4Q/phn0Nm9v+HJ87EYtZPv
Lx29V/C5HX4LB5k3VHEF2tDPCQVYmqknL+/2kPPWQ9J50CsGkRngz1yqYQqSwUtU
a5R6AAY/i8DyBVb5+73IB7v8M/7YkHoLulVD9TgoR5OfPn23aHHjIXTfTqDWvJE1
DXSJEiz11JEjwrn27KDJbmKf/v0N6l60siGOcUfsdVfmwLotnenCtHlGvDpooQyp
3GuJXQVJiSrLJsBUnvTZ9ZhuHw+NxAuJOP4gs9X3qyW+2Rzk6aB42YWp0JdLapVd
NBrtY/UgYS5QACuObS0MqDxSso4CJCmRISZ64Rbdw/DWlFDQVLcj+vvaXqJfUtBa
jbm9zeNqdtjJaXdxAQvW4+prJFLI/lQqeppddBWxqMG86DB8nwBoj37ZPM44f4G/
VeuOslrqJBSyWtdbP1TRf9oB4q3aif0kXzhzcaPnkihm0gxpYZFCm4OZukE9g3uX
hxIPLcdBFg+kUb2Tm/sQLKqEWNRR5P+sWeaANkIaD4GYFrxfRCpopXTSetaTvIVC
ji3w4HcQ241U9jw2XTPYG2Mvj8EDHQCjPorzkLzjOvb6IPlHFxzh2S9NxbpArhtd
6I6IMvxlqXtD4oyaY7Kai5ZCerqjPtklV0qBLYmdwlGZy1QdS/hhFQUA8k3IF6sI
yQ5CDEKlosrtHxk2pHX586/Gv3PGzjGhBMk/KFa0sW71Ucf3rS12dE38VeT9TuIl
gTVm7KXh9ro2VoWhQSHWK4RkVmZJ89bAx4GyZlMlsijIHqLDX+dGR29UgFcXeQH5
dUFy7h9SWEEjFXu25zFZ/VKBkjMPRRDczbA/rlhheh+kAD5TRhIhJjxGtK4HaT6Q
YcQvbnLjoUcETOajZnuOJvmta9Ha5b/c12V2+iyiaXdHVPRBtztVXG/V+IRzxymi
dqM+7lVXoZm+k9haasMyYfwb67m0bgCozGOs38SsyTngsFHkZXR8cceqw79UDxka
BlvaXfA9+2hlG7d4aD75rpsnmpr8DGbqlHMN71osgwe5xnLX9SowFvSe34y5SLEb
8d5pX4pLFP0jkELuNMN/BPi1erMgEg+I1qwXd/c0wFLANKRbl7MC1WYeRSD4qJI/
gnB4+xpPfK28uctLRapUNvc0GW+prDTTOWhnIZ2ZKm3/TNNEn9xjImyhcW3EbKWZ
PprmKicGcF1Bjqi3xFaiwfSTwWWENYu5ptljVpEixtdgh71MEjS7I+a5CK7Ft7vI
V4/IM8nMKZrSIkmMBi7VgSttQmUj9nOkjPWY4QAjrxKSBtKqxiw4YCsZDEzDFC0n
TAG1fghl87aRN0nHg9lm+urnRN+l/fLa8hTSYWPw0UHS4f4eB064+ky6dbvQ4PCm
5WJyHsjNUnO8a857RwLHJXADWef67e5ntIc2iFIFUP4rueSfGUuhPnVyfwQZ+uCf
UwBLBuszEgcXtpv7E73olKeiWNvDm6m/gtAO9EwgtpD8hVxVNpmxHAWhwTo8lYr6
8mqiTlPY0rTAA2UqM7tjyt/ZHFPpJxEZ6Gdq+d8yKhKyAEPH4PVioYfuMMBZVuXN
J/xcPogPuaFOOJyUsSwAd1NVgUdZayGmp18bbLal1A2WvbwpgggKOhXu3m6cI5KT
n4e//rBXojp3iNNK4KQkpuz0zbh4FniYuyfWQk49GROMXf+I1VCao23yZgL8JzdQ
6nBDwo67xOIG4JLBYM9x+TwKR0UaoKIfEa5pcZAATl1BvqEP+18u1pOwaNOLmwOS
x1gBDF8lchVAzDfhuiFVMlTTsjUhU/vnZ3mTbRJlAtA5NZbGV89Uq0o05H3xj2tT
6jBk0Femoi6O6HGCHDOY8jvQfpZoXAwjDI/L8a+IJWJ8uIQBdO5mzePWZGQ0ZyPa
vZzqELU7pYjy8ZM5TpV0vfTdpY4Avt3g2Dn/8tEtCwalOv1mXiYcF+mf/HSJ+LrQ
MVAUoa2TzPw6UqWY56hGNZk4wNpvraEqQfZvKZldWtlvRwlnbqBhqgltvRqAgaYT
QMOQ00wHPsQvTGdVosA5oomwyOOqJ9PhoMbtwGQ3lXeqNTgOUume1rgfYbCG5HCC
ioo2IOhbLp4pEBoXo5Ns6bfCx99P5/7Y4uvA0/3SqO1Aw0IiLvRYek392CyaUCU8
iSsduzJfkXQJblXtgMpFld7YtF483qjYA7YHWMqXzgunBzNh/I1L8LDZSTntTXvE
Xi7KNyxFApjOeWqTKQG1onfC2MTn2uQEJ7S7CgjLQOIEpxx0HIqf96Fgrt78MC8X
NwuzFAxrYRKPneChLnj+e1TmkgBFsr7n6Qw6zaKuaut1HHsOC3zvUN8MqNnr+zh9
QmYquw0JICcLwbL+1d4RdhoOyihiEyk7Lgbm/SbpCOKYN2j+1Rpf+LJdZDoimmP+
MPtzw8CT18UEFjpdFk7m8xOvrIlEGKEY6as/NefmwHm1gfqdluL8Cc2YEKV307Wt
dlOoswTsfa2VYaNSMPxmy2Wvfd5YgcNyzjaRCIUOJOu8zxIa+B/mfi8w2yiqbs1N
6yCoGwdrUwSktZThRYPRcOihrDhH+SvTqSI5XGfj5G+Tf0/BOwBFFvTIphVasNIz
OO3RiU5xZ2Cme77t0+XHOIh22itYobSa8xFEuqrBmCO6t22wpeS54jHV1S57pRC6
YTmAIoCt6+viCXrcernrQmUdWvXtvS6zkpWA7dfIvIhtBJOgHX3WIxzZ4+gPD5um
yC1Q+iLVARg4U81ODGxibgjilq+WI64r9X5K7M2k49IRKnWNpes5iU7HpjQyijtl
6/7Sq1X8xamOkbmnBqdxQJrmXCpeomzaQOc5yVtyzSdt8uZ42/JeF/tNu6rGiJn/
fzE7Ru8d5YNrLkzmtJ9/hjtwcrY8QOFg5VXzLThhDsncCPZy0amNoCbX9dXW+VsD
SHOiFW9bXys0GaoDYa13uia72/91RbPneWZcxFKu1iMOgCGrRlrRi9GtoxC+tKyi
l8X/2FJ04H7Tqhl0JuCc4fWZKmerOEeeGvLcUx9LFdZCRGfFLfwnfa5B6EpLhBkj
xzGMAptHpWdcS3o5WdLv9x+mhYwBrPMZC4ahSXT31vCcBimuCMKZcKf1rUO8YZhI
m2rZJGkYDXna/RYnF1qerioWz5baJ366h0XUOi8dmY+EVPZTt7HNa0wPzl7wP/YO
qHCqwnJYLld+N+/p8Irkz1iQOkwJqcTWGX2rnd+wJ3yWzQClS/QmAXy0Al5RHWmp
8wcI1UZhwCQ9rE+zeGt2+3n9NQJ1p9z75itZm1iEf4CQn8lSEKOVcMueiDGNmljx
vKJCeS9wlZMKNz5iaU0D0Q5BF9ux2wiT8lV1iiJ+gTT9wyqayJXpIcd0YlqJB+ym
IezuyHsSTEYaYQbqh3Jg6zNGzA2RTolurcVIykX/Z8Oz3IvfszjjsGtQvO8m9cyQ
KkZ6u5naSpbUBivReIzfMcElgRpzBCcZ4655S4ZGVsFgSm+2vMnxJdpaHfTHLy6g
mMrFVkWbkeQquYYOCaFnnAHyBf2D5UFb0x6PxdTem+PPF8K/XBZdO/CujGyXHY6J
Nshfz19sPCrx0wz5KVvMGXpAXYlbdhwfCUBBI97n4HmKkWW+kKe2R+lzk0zm9xDj
a3lMsgFDqEoQK4cC5xTUBQDlE9nOsOVptkFDy49cXNOzRyI9VZTRzJ1gQUR6UY0s
GSqpgbnQVnKbCO/ZiJOzM/T1O3IwfT4vUTTg2nHs0EEWqP0le1rbjZ3DxQ12Aed/
9ol985GT8R2lFasuTfrUSF8UGqeq01Mf8DAPjzyn0MmTaVrg2kFmg3nrh4+xtgaK
zDsYL7rlPX9N4vACv2o+MvkOgBy8TFbmrRpbVWi7jxuty/GSfCZuBw2+unTYsPjc
dGn51aS4BrHtWsgkmhCzq5e/2Oea3HCsS4BfL3hcOQNfsfcfb/7o4TORcJNjvDBX
AgJSKjC+SjrA2bdN4zuwzOVAXWMf1frZdSqWAIphbsqW9xe6EQH0XPN6+lmL5jIA
fZZXJEJfu5s1NK96HlCpdobhyiW3CJe+W9UeCVPeMqVXq+b0xDZpYlBkcVTHHH/7
9J/3p5uP9xrIRCKZ5xGBHAoWrLf2VOXEiI3O/SY7XG1MsR4pzlBLLZYUjcp0a9wW
cNhqCR7CLCS1IFPyyl0wMCxa6WPrd9gI8UR9DFYfHVXOBpCAuiOOv8gHRB5kano+
AOInp9LtRx/Vjav1AVJiy1nQ2Wp+xaNC8AOkff6xqHN16xYlCnq31AAldMQ/VLKP
GjRflmrWGEvWADWksbInmaW4Qw8J0YfTKrBYv299d9QKFgZGmy6NdhLBMP9Qoe0P
BqPLJRSXWCheTK4BM8Vci8c1SkwXXG7Z449S53UhtHzBroDBZ3RNt1QkD8DcY2WK
t5h9xx9cU6+Dq+oJ6cmyNZGN8iEWDta8yc53JgrK6FJIxHcuWOvbyhz84Gkzt7bk
/9gd011YUiiF8lxEwLcGuySdGkzZBGtrgw8AaRAXZkEllBYt7oBmZwhHigEpNpTY
EBY6hOmiSMPtWUF69nyax1fo1iZrNZey9rKdtmDV50iIj5PlYnI9evVjK/+mZ3p3
hCUR1OvsJVBzXyMC/HiRbRivHRZAmhi4SLKn63g2FiE4bbwUm07Jwxf/0cTUFnyP
jzHJswUzjL5TF5rIOOaaLkfJBHgwM7cyAmTuuL/Hfev5QzLhPo54/O6dL69MhxJc
752W9WfpNYT1UG/CzgdTWyb6quuUIIwqPL30CclPl7wwR8DJFOjtIrCpua+Jc3fO
MKr24921bfCCPamFXlL+Mc9eF3zVMOuc8Ws5pTmDW//dPTfNoDQxjj92q751phdv
49c/liB1o+yL4SqZLjSJMHlUb9y3784jdECvEwtd5J9SiWC+KQ55+fwWY+rhzISK
m+eGCX5unZaVrcPI8kl26VEpTWgcAyFc7j5H0g708IgmoljdUn+eflDCttquGPSX
lzQPyuwprg2nprsj6ZJzWiZLZ2ATCylsTVszvVbC6b6m87bDxScKKCvBbxTkToz1
pziexJ8x3EkQDOPnVFwdtMDVRpzqcec9OLtfZAVoP63X3+xA/aF1tp4lY/TGFPCh
BwbU/KaJdhJPWG0iHkXZlh0IHQbrKbJwlrRCo4Mf+Nn3nyJsA8yMZdIsJPCsHBMu
Crnaa07W8NuYT56pqyT4sreSU86N83vK0IPuBZu/c+lkVdkHmsF2IL4UOfkCR1Ku
j35VpZu+dtIrdv/LSDVMB222k9pEp/1DY7CccBET1BrCYArM26FjyWHx9846AB3y
I733UcDLmlJKi/dcQsTR+PoHOaaIOmb5doJwcdB1QWK5WG5tiTXh3sFVr1mF4XKj
iRXg51h2KbuGS5S5vU20wsldA/reG7cNfACvKEMJTlhT2KtOgh53lg5MWEmCHriK
5Kvyi0bPMByu9LDY+/hdDME3I87XXM5HCS5hXPWoO7P1sc0Ct53ob+C42lJRBCA/
ISd5RhNiMkfOeuNb1tsXZhX4KiGLYiFcTFqZ1JK5cuHCfFuWo/v3OoAHUfIgDsdN
AmQNDNxQSRCro04kTNtiopDg3DIWYqF94WGyEIKBGoaQ/O4eTwyzIEDMmIharP1C
YqRlaoTwGVrwZG2m9gWDJ/e5Ad3w65wRZgtSqp1Qq87ywj/cxnegQ13WsxyiBsif
cS4pXWH2GXL488br8EfEzsE01AqfqSw8gYIp9JIm6uO7MqD9rY1csqpXvGIPfoTa
x6kaKQOf27hK4/paU3fgVOAUPcTNAfN0WBHhzgQPgaVrc7KKg/QHM7Oy4JSj6b2A
94eAhLvoy0rQY47jhJGG6OSetD3F31ZLBQ0rMhjmeYflMIYFDUfEIQvQcAltc/i8
qmWnQs7TpW4jh1CLreWPW9pvv9HVOMQ+FeHCx4Hmks9Iq4i5TVn6aNNcyGBB6gne
zeQIGMdV6jNK48M2sxfF/QZqPhI6RpVAjDLWQE+5iKDU+vQGRPDZKkUZC7U7gefi
ClEATIXNSsTadnwh3BXJ9098i/dP1fWuqWfLDy+siCNjts4YIeSAzO5VPVgoiIEp
VYOij4zKbojH/qQs+Afx9IBTB9fe7NUa//PcekheHH35TN6y/OrX6LCNmjVOd2Hi
5E6aNIEbYH4ZN6f9jx/IoknxVcSSdkdrS53zktaHmV/3xHkTTAIrYSQU17kA2n+K
LbY4ZQloSPkhU8m5W/3miiBYjba/Oh45Ue7CSRzjzMqko9yHuvkytKldcI5PQ3bO
3d17J1X3rmRKgIOFD3Ir/NkStmnn8/ADV+G21480RHeqyw/HQJya018s5KUs2pZX
90jtB8bxTx6Ar4nY2pFvUzqfmVkOhhoyveGrfXS8OSZayS9TOrWLBh+tHuXvx4/c
U6fQKfnE07Mt2mDWiW8eYNidmaI72oWDE1MQTkqOPKFdE18UYe98wHTtEa+uLBXI
qmSLP74Biy/ehAYtdI3JcoBY6p6qw9MKj2TqY3Cm2bpUEei707Ml1j+AkuO8Ote2
fEuty+jw9DuBAApSXdgSasoCalOfmP2hHZUROjhYC7z8gvR2HkArRqljUSwfCczR
G1uEjm9zeQ0ArHrMUSx51szQIwaCNXYcwwEFwFnd4dFwjzzc1K/YYZMBL7Lc2hP/
ZgKHvXqG4DIcXH1D9WnlLa85djbuSqGpLM6qwjcq40GPCUWf29m7T0AEoCpM+ayX
D3VPBluZobi7cuHgTwpD4CbCbE7BWXtP60oeOdzJ7/yKOky3+JBcwUf50ZUt+lyl
W+vQtpullLIxiOUgBOHOuW5mmFZyOBissm5WazOXo6twV9IGoGZtvq3fXAmOZ5xa
Af6Ijq0BYm/sduomOiO2MjQxW3UIg7VmMfJRGw683Cm+A1xUu3+H3aMcz7fu7RSY
6Gp4+vUD9SJbmPwd9+zVGgYJSfhD0UOWCMOe+ZKbJ9cMTjrGdtGK11gm5D/VB36c
Ac6ZIYOEzLvjocPGVjnuyZclGJGHfJREyEal6FbIH9jOxUTPqxa8YoiBAQL6epUh
yd6CiBI6pk5U0ITjRhi3hiZkwHvUQ2m91frecGuqEIHK0lVqhQQWKIUwOK9BGueT
SCsGhwpIh4xM/iHB87op2Tix62zWpQdacOoY0ptE1vBiypRaUqDLYO0fpU+xv9ZQ
DuCrCy+k1s2OsZljv795TDB3Ksx/pVBPvtUR3joOR47/TX9WKqKXiI67Pxk4w75F
Urcf4XQbjMtPyAbI0+iYGAZWBkdlblxTyLQ466h33RV9qIifr2QZCXtAT7p4aFyZ
hL9ifSEpnH/QfjoYlJJ+rSI+fR+Xt/0wtS7Ke09a4ZAu+TP2uZFSHq3/EsgJQfKz
qtTM+aq/fxKcnY6UuBR587u4/9wW0eIb6C3ZTrZ1Oz2AdUB0c5o3mGV5ZlWQ7ptl
ewnp/l9Mtv01k5nd0lsChjwpDNTnSvXz+XsgD4KemRlMdOJhjbSzseUW+N2ka7iT
OVUe+iNbWKRRhrCAHYSpoGVqmkYo+hWku+8Cjn35PdTWKFgs2j1BQ1CxtUZItVT7
RHYzDmWfXKNCT3xi0NE1vJDqN7k824yE0HIyVXyJnGPF5cAm2eAp4yxvWBrh1QOQ
2CysjhgYZ5c6uSWa3pE2B1VD2VGQFbezeVK9W05iotG6Hsi5zUkVwGfFxXBw1TwW
5ChRBlNZD4mr7ragUCkO5GgWM8ViKzDknart2gRX9U1qlaBoRknChJpvglPosUcE
Em8Cj8T3SrJlU6NeuBvrPvTogTbHUgWrxJ87CEdJQ1T8MqDdlhm66MfqINmBiZeA
4GZfNOCWdkmPCo+E1QzxNmx9cAqj45dUwmDzZVLbbZc7dSF6y41ipyXXIKT2Qcgg
NZ2tIgEV+RHPvN1mnaYo30rBEQ+R1Ube5jZX3WE7hnp1qkT6ZM/xksCJHvN68kB/
Pm+eQUSXSeTVQUJPuYM4cFoRBHGhlKnvDRwJKQwxMCb9RANh6Q90R5Ywy1fyRmcE
CKyl+F+uSPMJNnye6GF2TsffT/qC81PftRAI4W4ABgTw6+R4SaHYsrfkMS91bU4o
aNCR0BDm0e5OiKSL8tiZVybcV8sDcjLlHm3H/6jUs9JHsn91nuU2dvz3c0sF/ZCb
7vku196pb4Q9kqfCiSXRk++HxW78PnS+G/bW88pB6yQuAZEbnmGRNcn/1GpyOhFU
BbfWLLvTtBdhTql9Nx0Iss6Pk4G72ixTyhnJxhFhXGUDmlaTYRioJt572AComKYd
jsFnL4Y6AtpDUcgML/9R31DwezZBO5tpuZMl/vPpodGXckVyEmyveAZKkKiU9Xo+
6EKT3hjKnA60dSOUTRoDe+lWQN8ZWxlkt140XALZFogTfg1zgPbVh++lh8pwte1k
8LGeKr7xKIvM3yreRVaOlr+fak5ineI0stKx+lMZlbF+R5YWEcz3YmVNRfxueYc3
EpTugmGgFN3w2F5j8+zL+4gMB8s3RC22+pehcrf8+Y73y4dhsfCPTbZ4KfsaCCvf
6TSioRFHGa/94Gsa0jj0dTK3xAjRi8d6HL0YgAAoF8aaA4fEt1z9u9+nQYlyT5tq
e3cTMmvN9GyLs48kPXUuZtC8nzxlnbeKzkwB+C5sLweL1AZKICJb2CmxAsuNv5aU
9UBVxReibM3YzZzzfyeS+ARNvHdkia/z2+xm3Nbs4K8fUxXcqDUX53C0BSl63wEk
i4JtcsH3CEN60gB2MuJafAYSQozv/b/bbunD8mCnd3n2FOHE8TXtFZRtnlYH3gkE
rzyPViYvVqjzMEjbQw1H7ONKb3DYl1ZqQElOYhMLcfZMT+F1gdOD4xOCiYxghOb1
LUdFRifRa+AuQMfH7Ma8bQBZ3226WBcuKBQhCzunb7ycUQ+ZCBqIkTI5Fg/DBAly
AwSZ/rWrIy9/+27kNbi8GWxX0W0KJhvzYJUmoJzNiZdL8DpU4CT5ithDJgTuVHv9
OeBCyc5q82437pTKaGSJ7tMaPAFouw/z1Y7UtibZfQKvpOgin/CzB6Ih5BlvPim/
vv6FWrkepgO/GwZ43Bk+/LltyAgfodN8ihnukSmn3MF6bsYakB1XyKLBkfbOUBKE
9sJR7J55dLc7ffGgDQKYYhQ1t3EUso8xksSWZ2m6Cy4fTbrL9cTm5C8/N3G2wLm8
G006XyPq5Ltu2ukdpDuDRVkCso06yxYr+yL3tvtY+INNgNKLu3S+Z/idjdZgcx1B
ZhthV7bU+qpLJmRjnRY/WutbAjwZk4qYWSbKiFpiH+KMe680RLOh/LFFyEnYl0KZ
8YOdtMUms9gFPTZjCroDSrdWQWlb/QkCX1XXKqaNnQRruwQOtTD0d3jMXmGPB/cf
yPYp2frAyD1AxM0g/YjbSYBkdbGdWgWT7UyrjTxnxicESwBxOv9A84lJvNYj72Lc
VcR4OmVufWfL9QpFudalm4thp1Qg6dX83A1inDUhP17uBNwRAtJ6bRHyUs3fTpBj
6dyBMeV1su2I3j6adC9pncvbrUCLA5hKy6BNbGhEHI6RirMKsaGWH6olOLcqSAFl
9w1PdQoCJVlRledUuaQ20S4cpcTIIeLoRBxMupfB6OVvh5qGXlmVeA6JUQFwBcCt
/YDsGiv/st54/HMpE0SHMpDTJbZAKEAgUbwcR18l8jv8fSEmNR4qNjA1i7cysHmb
uGX7imPj98aU/Mutg6HDiG9LTLFVoOoDEk+EMUBa+W3LBema6oSjiAmxpwSjYlHx
hng4MST5srXQ/ZCj8gycKRtTPty455dux4JpU93AMbZpr/CtyW1rZqv6ZrQZ1MUn
tPg7tzI5RillsEQ+CSi0GWW+Lwlnd31nvkSb3t622hYdCzwfwJ839JuPEKEZon16
XDr8jjqjHr4nJI5YpJDvIjvS6+aT6MwgLxxeR21XV4YKIxctP79JFaDWYzxbwAv4
EcpSaYVPFF+oSTIneXjFHUoU/k1FKruNqMO270X3nvMZm4wbz8qSmINZC3/5gPLk
p/O9Y0+d4ASFQsOYjUda3ojbEm/E1vPYd7YD/f340Dz8oli6f8eNFNUYn2dhcLQJ
OkX3URiI55vqQs8u+uII7YptF3quQCr6wncVDJqKsaT0DnaNJIruYGs8SKRLk5T5
87qb4xpycwe4nk7XMXjsIHiJD8w9BaDadrtYvxv2E1YY3CwjXvvnHLdAWMH6IN0h
3hRtA+XTFwI4rgpHYg5AUZx2ggZEtaQvDIzHydc0gnksXUE0YKL51xEtwsXvxDkT
9glDxY6jC4/iz4Nz6LS3boIFLAFiwtWd0VObeHxt/JyX/+9qt3XsBkRGJ30PELZw
Lq40zbKkmRoK61vZOMjgXaIdGLHD9HEbv/N+oEBspotwYU+u0pD6miFbGGeFQq6L
WG4rD3ad3YGw82qfvE6WRzXLtq3efF9jKN9sIj5c+/COZpOF8FAvJrUf/0jBMNNW
fh6sTsvUXXMuXbokGkFcN1adRiiPpWTq4CVIBPaALlChGMNff8OLR0OUsGpetAw8
eNQBVj9Th6NNitdJ8kUNQCKVcm3m7FkfGHM14goeXrrQh76WJ4w97E4rLQIXxGUk
EmIK+DR67eC6DjGcMgCB2Z5zghpHUbQyBhOT4Yoq4A76u7L+8UT1h812tL2DMAPu
MqVuoXHhsAQNyIw69MgywnMk7DLL+wLde4ut7N/Y3+h0aekw5wluxwE0GIl1mfkZ
yFv/hrLx/XUaMZuHTz9q6mQp+0yWpQxuB7ip910kyXCtbl0JtYSXzSD5d523kwL0
f0OF4VKHahq+S6ley54zDOxCNT7pYlaizICL3uTQp6uYK14fDm8qlbaVlrlslxnl
//ZT00wv2Y9D1lR732G0oeZr7o4zaMzEpVMxuNrb8sinCPT+ncWJqp/6eyTCFDzB
94LtEC0s1z3MFC1SQwMPC/Lf0CufWJgaBOOeD6P0hAlLNMh8zoBwObrqTaATtGJl
ad+OgiEdUmcqJvvljesjFE04LA6BOn9AGPwkYve5u3TnqHwVYESryMVAvr5IWj2M
9EiqwfUBvKm56jD6fIz148xRrxcWeur1zoXflR8PupbBoS87giKBmh55IM9J1UM1
CZJwF9w6c+rB4Ezqc6OqxOfSqNqMD4TUwyPyDLcikZ0oik2vIdtFSRFzZtemUlEw
/ClvBlEJnbaLM93kkTZMmhW0/HbpntHhXZI+bCT2AYax+bDy/C/3mFE7641n6OhF
0TOkDiBCAYgQ3LH1qQy6xxCsftszNE8teUqgY0M9zUnMDg8w3eRK4vVUio9TDTiq
tapHcEt1A/8zJA81Sm8xRvDu5wWggqJXyKf9tIMD9Y4oOFfAo+gzbGJ56AsR7TiO
A8glOKj1RhKqf60G0799mre715voxLKgGIP5oYp77VQDTGI7Cvb/IghCjvktQnLq
yqrttYwfipBm06eTd/LpmkmJMMkvaRjlWi2oE0mtbvQy6y8+y0mTyXHpJHYDiRLb
nPW9+Bpz9wTSh0ryzzIuFWFlOceIy7fwem/izLozFEMlNv96nuZQkyHHQkJMczh8
NFLKUgM9dGnFR9ZPOTdhcyyziH3ZX8Phx65AWire1g9vkU38UbIt6ZdpPjQkShvT
/sM6jEQHtsZYz4QgRI9pYAOLPeQJkdmpRTCD3+ba58HicVLaxjsEBNGTTbps0j4s
9OlNuWfqQkQeve5IwyxYalwpYWeYoyT4frzbfidj7hyXlpCov8ntXoqaAaj2XcS7
oIccMYx8UD/F6DdvR2aSWbwhKaREk+AtjQYluLHhBcdeV01kXxQdYx0RA/OC8GQE
0Oa3+EyWCIhM167esOXHU2S5ApiiU7gApLctpngEPwBPAr4PUMSRF2HPB2Ek6lcP
ukEeTrWb3A4zw9F8SyUw5K0suu4Z8VhPfhjtab0/TL9mUhaeKmBKed0nDPWzGcpp
4XYf/Ro17UE0GyoPB3+D5/Jq5wI1h/s+P8GH1DzEhsHh9SiaNc/exAoUjJBUZO+U
Fy109dpGwwMlv6mcEV+Nm+CnZhzSC9n8o5kj/Zz/rFFKcXYSUCUmhy5ZfV3cU+t4
dmwhtdVhdjauHXUZ6d0mv9k2UCwC4a/ATSRk0Ww8DLku9/XCytlxPk254Rv3z45G
MgWS0j37bS+IBeZc8icVL4+wvzz2CAl6uhuGMTO3xaiTrprCtYReHJO+wutlsa3m
MurGAhHN1qk1bRjp0I/VfrXP0LwukyYjysNtpv/sGrwGL8DmY8/5Yq8WCOZdTkoi
efiEgGknAguxNJvou2yqIbydVdttP8hUwk/GexwOoskh1cDnkky+ZD4B2ySyEgzA
kZ2Xo9hDoFVZ0pFyPn9PArjU5fggzZbrKdmFUCrkBKTktAa/xVxi8ZAceLKqcEoK
dq8vkGLxaq4/3ISuJ6cKnTaqbOqZJvDjCim66rQdb1+pCzXVlq8NhwWY2GLqf0g2
e7ztQI+9J+aYVURpIgauA2w9O7NJfZUGNdt2GcHs7SfzHDzW5OD3bcoNJOaPrJV9
m8cX3eVcKkpm1xaFbqOW4OwTZdwtK37Vmv0JdL8ZlPogZ4n9TLCRKMk1JjQKH9yz
+okbAxfDSi37IDoVZWh9I3Uq9X4zO2pkUft75R/PgO4hwast+fJ0vm5r3ei6ydnH
Ca2z7DRJI1671DzREnNN2/FKxq9KpckgS2TrlnDKEqQadpRk79DvtfZkVtEw7iJq
WmsYLTIV2jmyyjcjRmLE56Nj7xP5e5VCaTtkNJWQbfLmiQAEin5PTG7HCqSFh8ax
hD5tk0Yhlazb4w8fMimW4kHV4haIXky2+0Lp6mab8vqgkflA9tJ4cpmclEPr6kZg
9QjHCxZV9ftIqUkzWchbtFW5Qc+zeIcUWRKw168k0AB//FHX46N2eIwaekzV53Op
hB8WB8Iqbl3ojkcVDfwiK+560V9bJSPrQTlaDhDNR2BGPSaR4bfqOTy9O9yY/Rct
3/myoPnIEWNsOfUfFe1MCDYGZtIu5ezmdaPIljGEFEVt4oDJo8XDCx9JgXdMZomJ
PaV30Dayyc4DKo2Fq5irR8JRPiGCBg1LEs8YqT719RF6SRf2kSZleRtTOvJ0AjRz
BVo/lSxzEptnFm3AMrGvx+AKiEZ8+XxgwsQjR7cfqgS85cYwvzEzBaDnFFCLSw7w
Q4My6G5Bw2uJhAuT+ggNUEbwTLRqwg/QbdzXq1r0CWcWudZmuIWOzA/TiK0zN8/V
6epDr6QUOHUOzRkgFEOaMHb2lkPJo4CuEPd1Bwg1swtJYgkI8JihhlfIl2iy+RKH
0/kvCnKS8md7h0KctEHj7dTCZIxYl16y/OGZgxUuMpsPet6ibI+smTaHxkyfWAGV
Ei75rAN3g+0TiIjiD5Zyuc4mA4svK8JB5KYxjw10bN9cJSx9WHUOPvCNubc2ymAs
GmaTBbCDNES5ZkWxzYKGM6wacgmqgQD2llj9qeIPJadIdReh9H24wqoHwswFA3sg
7oWq2DNiVYnSQoSVWwfzgWZ6/W/9EmD0svheH5QKBaSEo7Vx3wAJf1mhz8UIt8VR
7uX2HjFDh83vQX+/4XYZBzK66argWMIEr3FjVvceojn22+/hd1/SBFxojIVKi1xN
y2W5H4rrct5i3iVRmrHqKHLiD1p9MrE5wfGxaMsNGtJP7qJfwwN594kN3Zt2F68f
nUychdXBfGyo3dekAPrPdVKgaHxuez6zK6aJzsjmYyjlFPVkLm0bhyAyQdu8Uila
hfOKLDaNjypKHQlwA7yZ6arf0obIGAdGmBnvry/3kBWPu5cd431bKVsAuTyLb5dJ
ZJ1JFMNvOm05qfk9dfU4vaSyXuBpaAO/nodCfJ8QShirnDiCZhAA+porufwX9fBd
nYFKgXE/OTX2CM/lcl+XiehCsJKuW1fg46mMb0/BOnE2HHlhPknvJvgK7gq2fdgB
CNb5pL7PVvdxIc85lyyb99ARWe1mo1YQdCbRxuQIgnxFpSkh3VOFbQsJYTcdAiBA
r/ClOZH96c8PQMrabEhy5eNgFq9PdPC1p+lkBSGV7DJebMKQxyRH/ooKFkJ2M6QI
Be0UclZi0s2qwhaWFqTy5RNFOOj4vkLXOrhS0Lxu9xJ/V/G0Ll29kMUOzpbnRaLh
qebD9FVPzSSOhok1pi2lLGAidDvfWbNjZWcTby8QkFJu2vWS1kCwoZBqEbW2a087
59tcUW90OZaQog3mpCW9us/fCtl5cE8fa2V2cbFTeZ0luFuTZ/DF1+0yXwPkq0Fp
tAPFbO6slcyPQyx6WiWVFEnNB/fxN5GYQYe6mZGoynLyiWRLX3q4SLic4N7btawM
QrgCAelUWzwa0d2GmcQUVwV85C+svFNSBGIA0uHCaVRaK289Y3glZmWjXMdZ5n9s
5CzP2GaZa0owh0CEeBhBtLVKYJPM3DV5mErCTo2vTyULkeOCGQPDqOhpSmkr6st9
iS4bF/VTkIqWcC/04yuU2mIymXoMgqPSuYBlfRYw7Xvy+Gz0uIQvRGSUIIRBzp4x
6pAhGioUlfrVBVAzk6AA5IJbspAi/mEEYOSDp/MW2BSwjMWldE9iNiRpXu2EI8a2
c+fYmXWiDgJI966/pN3waL02sEYowc07RIfyzOMJhJoPhdwWEkgL+u2xdpw1wqb0
jAMM8bkC5sWAeyQ41gdxId2g0Q4ZP2cbg1rYJNRN+jkDckSUC1a4QRLfZ9kIJkZp
7c40N7VwsBDqwcCcjNWoH9Fa78gxHfKpOa8E6Hoo5EwPykUglZZ4gvGutVsmKHEf
pf2Gt/TYsDBMQXbUs0JC736gsOCSvH9wV6kv4WuxOP3wDE1CxZCUzPupRIR4f0dR
N6ixuLR4Az0tVbBmmLw98TWXpxfVRATtjsrupAqyEBmag9Dp+xgd10+6ef1A/rE+
tuVA5AmAzK4UX3hJ+F9yeXlN2+uMlLi/Y9DojJElq6tyjUk93p5bJ1XCjE4dA1zU
+D5clRVHsMp+jnsDpne3Buo5saolUbg5s7Ja34D3oRUhuMNuDHxfNIFtQO0py/I3
hpGyeoNBEKnvccrK3/Y/FGri/XdT1OHvzs9tw5AyBg80Jf1zluUUwlUaxVuEQ3L4
3VVfbVCC771DglNiiEMg/giR5kbYWQKkCbFhKNzLc8P2dZMxKnACglfFgzQ/hw7n
mF47vDUQLYabKpWHvkxi5/pl3GMCuGeeDdPCh53aYMjmFmWVCltUWxaOC/1EdGaE
QQ2UbO4/AYkTGJ4BS3tHA5BDxVpI0AuoMERJ59I07drDgUXZb8sIxZCdnkCyn2eM
m/SfD5MmEQaf5CJ0fCn1CqutaWWlJbwVw/PXlNoolalV62OZziNPKbz3d1/okQ9I
QIU/WoHhdtF+RYb3HbIZqzsld7zMiCW7mYnExN4vlD9yzgRjrpbyZ9Ijcsyq9nXZ
h/4qvhdrZ0156Zl/hnRdo+h2t5JXmTzvG74vZB1VvtIz1q/x3OWCyTeIpP1DJmtv
O+vwfc/WHTjfM+w26Wf4lovvcWY94303AJVyn5Ic0hV5yHZnT+kB+dQdr51Iho9I
3LZGUzBV8XL0VZKB6IovGYzBogo48rPI3TwveDzvZqv3lhKUCHZztt0EyzaojDty
f9nVlIDeIYUculB/MemJEk49G3LJtG3jqAh4yjRDDCjUsbfHc5zvZjF1CAeXierF
BxH1B6cAgYfqMUj4FOurRPHQPAQtGp1IK4jxPddQ3hW75SCpyE0KzITJyX8TcuAE
lZYVn9LCMar8VnpE0y56iMySMuQQJjccuJ7bOI6iIOY2DqWq0JWd/amtShMw+HHk
cULEKo5c7B4j4/OmzTjQVTKf4Mxf1zuxp7izfIkZJYyZ6iAhPeQmLCDvHYoXoEM7
AzxxP6UWnPuun5M09XmjWThcR0fiRW9OWLlyT1BFVEwAq0nzce4AClGM29dSLqtI
4DpcV0HyLKFztkud4UamxJq18sujQrP/K3iZtikAfJJix5ldxvPYF49+F9+ayzAn
cONrxv8PduZvj46+kguQHSPBuncyoHDDJmRQUnPOsNWp2FYrZ7bHBDtq32K4IEof
53t+7KQ9A8rlAA0bQDTF+2iOTJydrUSKpteJ22kh/sD3NzU1Vc21Nvckn8gfRhCq
8pGB/Yhhl/+Iefg5fm4kU7xN04HlmpB24jnco628r+QPTibFLxtSQ19kWLpmBY6I
cW4eRS0fDk+iV4mX97eCLfDst4312xO1hHveMpfbHKjzwOhFSkLk3xJsRCroqHCe
WiBaG34gx+id/W4mI2eVol+KZcv2ZFEZ6ITjqXW9YL7X1WLSEtUZGvglKwbCE0ls
KyTzF+y6sO91U3h4y4XrPFLvj17o9A7yGSDHQ7PYGlR6HEh5C4+GoeJo3MIJzG3e
KI3qCKr8Q2kiXan0peiPhaQfVxcxWkBlW4mmOGJQCNcojMdUmQnPpv9IGaR4OvDs
Xo4ku3BI4WTX3f6B0HYV9wGO/SLRAd6gI+cy3Dk2y9GNaOR6jor5WHgpms2SbWgH
j0frQYyuk8jGAJTCO04lQDpH3aor/VqJ64mstHJfPHhlOXbihUoX5Qbjfq2SGCiI
N/6NtGklKfPu1mFQxHuICqMtolbQ2d2uDJoi8234my4t/AximpkoOIPDkjvicpNB
sJiCmdubRtmDTwyWQGMSBw0fu1+pK+KyDJ9ZMQR0wJ5bVvKYMBz1Kq990tAWCDka
TXL+Ht3J3c9ADX4DaAZt60mp6yV+K+XOuIGp42PQvNtJMT0s6lWCm75nBGN9AlQq
P/mAb1HXzj11QHdh23i//6lK0OC/PYGIJkAcEOA4M5UghM2YdnfLH8QnL1Muh2v1
b0osRVQOlMnsIygA5WVdkoyoe3prtamJfT5GudvWyenpbYNS/y3tM6TZLUrUKkTp
Q91tqBldZsVnkB2YkTLZL2dKKv3Kkh56DuSKQvSJXdOF6E5gLhGYf2YslEhIXfb/
pZsJb4oXZWRmj2eThueHPHAsHo4ZuT2MFvU8hANREOCpmhCNJVLDMMYrw1D3x0b0
eTBQ2hPx9zoI9TemUzXFHJjG9GdK0rOnRPBIsLmSOOmG7OMJ1nnrCbZtRwA+LHm6
39XZ2t/Eimmi5T2WaAsxwViL7ngaTkkP17yeVjBAbmr0CyIacwcZymRspEF1Ccmy
AIHuNU0xuwXJzfG3Wql6zP6gkADVzziXB+ZirBVMoDhpEznQGE/Ik9WbKq4QJ1rU
wTw/X7GfTv8y2qJSdaxkTpk+q8qd95jPfHBkV00xVSLANTeqDheoXURgjG2dRI3k
1kmPYPLuml/0kVTc9INVrSADe8iIC03/W3d39vdIe9t/qoumpV1taznv6rPTg3Bm
sxNZhj8PMTZMQ+CjlgukLjwfJTgN3aUN8803E3jdjAF3dzo/SZKPY9YSCQ8U7lJc
togJFqe0JN5x9Kyt7o8fm+OS6yiYqArZREFozGZUHfTewpr162LhoGwAO0lfUm7r
tb42y07Nkn3PYzsQPSqpbiIQgmkhM+EEBjyB+GhGcJsRuaAC08Z1zJaE81kH9uFY
c8Cq22ZBxLdEeJSTttxukResNGqBteM3M+b1/JpLvM+gvH07aTsrzp+yoKgTkeRC
wXBELE/1iWkiK3Y8+17VF3Xz97Kq1P2DRNBu9swmRPAsMjExUdGy9SP4VdQLgpXC
j44N/Nn6h63rW2GXhX1vlDlUyt38gKUtmiDFwdJ2/C4RcAntvpKPhBRefHPfFlMf
EZu+YHQSaYAUx+ZqEAwlI17dj48JCVXlZ2TvuPdmkxNmRcQSRXHtfbK2UInGnR6o
+z83QaGYHqG6YOohh/vRboBI/GRrCAIjK/XY5RnOTLfWMeRFwXlviPbmhLlptLMg
FgzVkMs/UPfnuAyYr0FyWexjT11YKgAuX/zzau+I8UhcE4XYVh58Ovtdcdv3e3pa
aacrh3My2uYz/xOtYE8w8olJmJ65eOrFFr+Z+GykcovGya4j6ENrtmwiWc9/P1an
L9fbRvO3/ToSWSHD5DZ7lZD5O2uU0pJOEIk42y4hWHwOpC2aX1hfEWG04x+uuk3P
T5v6WG07rGEEfI+Liq2GmImVsShY0owGDYqQ0sAFK41+Zj3voD5csRidT+CgyyPx
p0hEvUKj2mGwIiZxquoibdENvg0tubANzQkzY+MmwWbUbTYCqhHFjUv2Jc7yD83k
d6UIklr4sOg/R1Hgtaa1inQ6BQ0D2ycE997sNaCRg0pVr6OJiGWaB38TciynSICJ
Ea+6KiwqW0qncBs+vnnkQx42NMWXLBO3RV566XUY4TlZpGVY3nzBUB98egifDQQ8
2PZbBAeg3px3/FJXp7taWpGcG4hVDrp7Dsp+DkOsVhcHZc/ubYTIBUkV0P+MKnpC
EVdY/4BtoOqXj2m38qqBOhuRBgyD7NNiE/guEwdq6BjnwoiH2kKP4mv+4ANGQupa
NcfSpOFF/gFMg2tBOtAMuwAuHi+o6Z7AME3WpPoHduhyyta6wZ0dklN2XZj241I8
PaPJ8xzP9rvxHamt3OGDon9RB/DAZ3BPyLjMnibdTv7//1s6zGfRP9VGb7d2lYc8
LUwZekypl0yaZ4FoAcOZBniIWZMY8Cm1PTNkamvmkbkxydckm7CSfxPt9SRvuFNN
YB011lULUrQErGTQSNY7EYQOfqjYhMoVuGIqTJ+QpTfaNs47B8CxcMLrN/LJQBmj
nki5JKyoCS/b3V8cwr6OgOs+o3MeXA+/jJlbtiYRTe3sa24Vc4xCYQRYQFKgwMI1
dNSjiP03/sgMHSRoTxN2Y+CAhj6A6PJXVPjmAPDojr+zuWsZvDJhWwL64F/ONHuW
Qzh2DbCbcZkDUuaSqk0Iu3uL8YVPBcBndsEFFGlNv2sVXi2PuAXl+3MuGP9zEtXJ
YQePW/u0cb2dEtrPCaC6cBPSk1GNq8DF8a1lKX5GWc7RMj1glRKgHKqhiP3NBeVH
ZOKaTQWVTdmNG5R9wQIK4ulaiSOUJN56e2MpzxWs3dj/Jso5z534uGj69mx4n4ye
lBDS3h9Iq8GscRaB2bECesJrNDWbWisF9668Q3Z2pEUin0eLN0WedlBxpRb0xSgW
gTTWChyuW2wRiIRhG+Du0xlVv02RFodPjk6rTGNNx21jcGYt+Yr/87AufuqM8Xt1
azG8aI47RdcjV0xCg7uKG9RhVHu5IkMuRbSJ8gjBjYJqlUn/jbCgaCLtq8aqRXKs
i2Lvqx0NparM2wrigSSpElbZbT2aFIqFG7jjw8KUNE0Nc9CpAVwhLahfPDWeNLHa
K6gCq+ehxI5jFqBp6i/yj0mM6fneMidqR4qzy2hpB0cPLyg0FWl3hkLwyaJaCfrj
3J2wxoP7vN+RAMlWFNs63+mS7NXqirGlZAPJ36tcqoJ2Ym34xRuAjtYYEz7Q2Pk8
Jv3EmhpcmA8Rv64ZxO1I/qD1Ut/t8IvovkGPSQ/rWurL543wlJsrsDSNIyYMaO8L
+1OzYFR6wyc7tq/HddFkun0X096XEHbpwG/pQjcU05xBSlhtwvasiaduMMVG3/ZO
iNolKrIywcxwadiBvUrvZQ0aOGNTSfDJoMH4gZWOEGkuGWOAKxrbEoeSc3P2Rjwg
pCMmQ9UI5qCjYGl0Eou3fw/G8XMMDHtVJixowCgRCCMXR41L0vJ5rye9wBEsONzn
0QDn0aw8XiVlZB/aP9RyS+7fO1qQsoTsmIqRc97/QFJxeu322atYnhV8NsyymV36
BL2MEDgT9R7NS7siFAK2FM2YRb3aAin5Cl0txxdaoUaEuc0cR6lPUwhOvh9XDr+d
CO0CztWBe1eXo9mhzgBfGRtrsQ6K0AhoWHjsMUa+6VeBID3g5Wdw/rHNYBFbwSGJ
ttnjlI7M3XJvg0AVF3XuCxL+p3w8HQDRNDGYP+M99zqVqvA1ov9K/2CXuf0kMJwK
QDvltMpNHwR2/ptmjvO90ac6WQkkrBhKkhet0TyUQCG4KHDL0GQmAkGeBieWa+vQ
uxfhNoMr8LF6Mjoas6WXabr/7Jr39dxPPiZjthcb3bzpvbksmVhJpJYj0aOQkKzO
qQfb6DNPBEBMKzIz/rFqK6GzGg2ezTDLE6bSlzEHrFEI8gx2P9j8YDvm+a/0uTfT
6p1zBbk9+rV/wQEP/eQ/U7sqEE+t3Qv2UtiPZVHdfT6xaE/1YjqW1Cy7Im40+zOU
S1mojsVlSqLuAZs0KMngI3hKFqQfNf7kq1+2vvkYb9Dx8kH2oUl90mTSYzf9q+7+
AYY6oiig2aAqslvRFjSLO0CZffKFsuuLGRwTBIWPxCgXpU1n6NJ7B8s/fNe2qci2
7+woCxp9bDPzh6Jz390v9vel19OJJU4NX2D371PoKDggKLGRxLqubYjSMv+6WJBM
6dXmP+X5kV9nrLdgZtFg8ZGErMh8MqXH9d1o+k3y3JjIFwhMk7UVheO8ayr/e32f
t9nvW5UAxWRSWIVF+I5gYY83PacfP7BmnHoUrK/PFBUkJUdecm9n7zeAv8BIw+ob
UvIB/gHmjnApYkSPYJvbGJKsXM8w8h5bORi18SXHMWj/avan20goQGLQuPzt36lQ
+AlHfbo5Sed4i1bUlp8AAYz54/yybqrQFE2TMef2GzWcS8zuv0nlHTYAtaURvxqH
j+CDEcVRfJihxpodIOFYVdzyqxFzn4SmPIV5dymDcbwWgESJy56vMR+wzfBWfYOr
gc5J9ImkPFGWKbqaXW2BzDQ+FkjdQLmHsIosmgb915BhzYj4hYMYuSQS0JECuFni
1wk/s/4FolrGmQO/dZsahk6tVzQoPoTEu3uu9QKlLgO5tR8TcpeZ+fUbg9uvIIbh
9U9U2NwOtfe0HylNeEoj8ALuH6MbjgQCVRo9x9LFn0Q0/8RuJrajCjAu7KsDs2bq
PlBe6EJoGPof6pKs0dEIvfr/Wf9Q1ysbWUcLGNkOe91avfCU8bysNS5lXF5G94Wc
1voBWC/Rc2XnjY5GYU25UB/Cn4vY1iF5bdElz2dQ8IE92z7FFdXGjTp8WXNNS/jU
5IBDPg9jYIPOdZy96PXLHC2s4pVLn3RbC2qoqy1pQo1DY8Wl0xs6RZilDXNiRlAg
5YLHFBDeHqgInyqRGPLm3JwkkU3mSvFVtE8ZrYEEBD3gK4pyJ1s1rssO2weURlQp
WLwg9JziwPoKdfvOQ3rwVIgwQL5ANYJJ4aw75Hp64fA2LenKbxKDUrjtD5I5mjXx
gCJz/XEydpuBtqhgoR0cqEjgS33ErAM/6iOBjAPLvJcSnoObsy/6BtycfDfG9aSs
1zKckB5TlE1NE51i8vHaoYQnmQELnt+sfQZXDT+yKovViorFx+mM5L1X6/wcQObd
qDIxyYdFmSwg9CWXPIC9lHGefNWfscVUjJjsjp/v7qLJgVjJutXYaec3AyleVZM2
NZik+8xa+pUuX0XzeQB2OyYO+dHiJ0+74qlrkQduIttp6pf0njFPNZqJx7aBbp+q
dgC5R4L4Rbo8Gmh04f1ZIbuYoaf8lvp/NoYj5Qrx2AERx1zP7epMc4srdchmuAgD
7XUe+LSGBtBjns+qM+GHsELyV1VhNZCZwWEss+HW2k8gzPwH2TNKgO1Pb8sx2HTC
Q6Q+H9oFo/tkiBo12G0CDC38gRK0OFyWChteOjXmohyTr2NlA7+snrBN7vwAacGR
7ydEkHMXiwy9fcBVCytBv+SRT3CRlXt3ONRWfDtmZIHpVXy2B50On+3m9g3IzHMt
GqpxnGolJonBRnx+INn7lxmhTJSwVSgPTgBeGySY0KmsjDAer+4uVamyzZYZx1Tb
bMVySrFWIFTIpPjjoIXsivkuOGl5nJl6K+nRms6niiM8V8/P28EO81Gjfhs4y+TI
jA1aJhLsnmu+OLggpyqJkUq2j4soaqXM+wDaq+GIMngiN2NhFj81tKDV/eOd9W5e
tCAQUpot1UEY6SKynHWw9BS3RPxIACzYYi2CArHb0DqiTmanX6iP6v/xgC7pUQU3
4gV7QBQJwGoZ5bEmKl7GYDm0SOG0Bmd02yzM2DxGa1R3bFhB0MK5GrjqBAC/gmZ+
yQ7woPNk7FXB2TJIpjc1p6cZU/d8xhae0KPbfpMSLr08D5Rm8GWLEecuXPyNLLkJ
fpNX+PW+eM3/0bmPVPqHGULtEFmID1df8wnmM1SA2fyogETBosB88tA6btsz3RCQ
rJjZVfE0Ttn25qawbsvktllGN3aTmwgM1A8iC1fDFNFUDijhXOkCZI69JWYgIeEW
7Q9kMP7+Kxn24rTZV3D3Qfp0l+OYQOBZmd3fsCevHvu5XZaXNY7MX3YLu/tWYji8
m/BcLRNLy4GlkEVOl1NEo4JpPslLkTfrzLxnGoMUmp1U/kDfcYecl/YtHYGHaF++
Hpb8uV+VXC8e5mqDEDxAGa0t2YLVn6RH+1fb2e2Kyov7Ywl2D0GM3siENGWn7dMx
wuWSor/WBKg11zkZuTglNKsY7MVc9eI09onQgT7GuDe4ajxssDtUvP5Zvj8miK0n
LVSDsOI4EQ6VoDw+LPRX50XeS4Bz8uhCk/LjHvTtbSSytHPt2fp7abGVBdYwn1VK
K2rmSgE2WQtbWk3wkh66F04MLiaB0MAgZ9Bv0L/QiHxm0cgw7alPkL3cUztrnXWZ
ffusxnaFbexuDwd7NXJhxIDfw6hY/0v8lCc7x236qQ9RvU/GUSV6q1y+7sOrWz1y
5D2PCGReUjC5ZLxj995jwKYSKic65tNjUkWUP5tltdkUDvseigIleLEP8htBlTGm
5c2B49vvG3TIpyZzdZEnZQfoa+vSvFZ02PZlZcj/rKq80kjFfEAOAW5P9r/OG8BL
qOO39Jxopcz4oyaQ1evQHf298T7MOCCW0JruR2HOp6TdynQeOEvgs3vjmsyKx+gZ
IheFMuK8HL6Aw/IMnHwrwqKdfulqpvTuq4ptfE0y52x0xysVTU8QQO1LpGLuWwjP
a4Zpo5cq/XmKTZ15gp4s08Oct3ZPHbN4PpkhMkk34YP4A64hLkE7Ja6n9ImWaoaM
Nv5NsBS2VzDTDFvfAwBp6u7f+mb8I/B5lGNoRyAu/VZKG2+Po9KZioFxiP3LR8dL
CjgXeUXMplENT8y4FDsxeEu2RVQh2SGHb7DJR4XfHkoDRCtEDfG2b0pcmI/D+A/t
OjrPxHHbuhHWUs+hG3JV8RwrhVBTNMy/V/JejxZGgOf7t3oHUBurznKlioqvCtXE
fEWcL3oOyuKAG3bDt+Qg4LxTn2yxhfcr8SQARSZO3R+k5fCSTuIDVDUVQS3Alfe3
IIDpePHEborwJN80iGUJSZ9jiuYX06WqIN5S5GJ0OpiySkqs3QHC5iHA0HFRLm8R
9oO8vbrGt91nAulquBFbvDnMK3I1m0YMLRXQUmY7EoIuqCNUB3BlXEkDC6XWhwAp
KPhAapo/V0nmt8MrlnAJmVkgx1CmgL/2Bc1AWcpqlqIMh9ZCTjvSCxujvZ5j+Dob
pnVFdtv5IUsQ7RZp/KedNKKkOZpxUObN+vtVSpMlbCqdb5AvTgmvMU+fXWoENgAY
SVl4/QeA1XMSD5zmwggZZ8k77Ksvpj1HVGtP+ENaQogn203nuNmkClWBkRoXdbfd
cTNp68QauDrt1hBaJGQqlynfCT5wJ1bhfZVY1NooNzrYbKSh3w2lxZikrCcgSOWX
l54hlP42yHpdzvJDEyPrEVv1jwmN2FLj76DeqzsWQ1b8uVp3MtH+NKo3J3QtNygi
XcdwS+hslZP5QuXNaTeCvpm7cllo9plJcRN1J6IeBEfpsd3R6hoxkPcTs81SgPj3
x3E15S0JGgZ8yi5V4SixeYqTCzWBbBnpbomdkq8FFo+32r/eoWd5vdOW0xzmqWzM
9UhfHR6Vfq/DXfjOloAZjXeXY24JHm0qyOd4WUCnCoPIqzsrFP67xAka+zIq7eyT
l3Jp1PsOMRixTZjYgEnWeINTXLw4p7ybU9LlbSE7J8lGxVmZ/vtFnTDPN6zDykJU
Ri8XMmll2iygIOPddm50XxFpK3TYHa77IPhQ7mtgsDa9msBDPA/84dxds1NhzvzJ
oAd7BNl5bmGaV4xj2Drbg8ldZ/mTlRBmRG1qVF7JDsXWQScb8auF7j4fKeMweE/U
wQ+K/NywW1Cz/BdtrtDz3gh7YRjIzvO0HWvFmpEjH8dWfzH6Z1ed9Pi80IizTr67
nyn40sBFagqLK/Zum6GL9Sg8OuKSe4tbuHmjny3D1+gwuZKo8+rHKh+2Xz14wJR6
jJ5VuYHltPTiV+dS/tWCee8C8ht9w2NmMvvNtR+VMwj80YJSyBA3y237Z7RsuIBF
7XuMDk/nSlqMMaEz6K0ZyOL7eOm28CPsj2MKuKd8ZMjXO+vMtNQvaSXLn/iUeW2R
L4JKDkRVBf6T3tNJmHkpWKPd4mqsQC46Y0XRoYayb/01lSYN8nXLWgmXAUFcMFDC
EXgIDlQfYN8ps58PBxC8gAanSJ9BM8iMyQ31PuVWo734FbpSBUk+z67Hy2GhwsDa
UwphGNj+sIE2hauRtAcya0dNnr2SHOWACUUySf8N5d6zgUZsKGQLrFG62DCw+ilb
pb70tmyLRHhviltxpduzV5y9sgSDPLUabqp0frDzp70/3Ct4oafGXWF6V8ARPr1r
qqM5+mYmFLppjQvP5XpcdaQTS16Yqn4HXInzxJ0ZnJQpgFwiMeyGDwdWC+EA8Yl3
Uel/VDA23yibHj9iHVJPEDWhaJIUqcKvuAJzmtDYBB8tXN82fzfZY1W+KxzvseJE
PlKh9WumCCVcjopDdq+xQQ+GDN1B/bTBQe+2sHozqGol3NMlk+aOwpEaBsYSiJRR
cKQ9nHN4YVjsU9KKVPEO6Zos1D5/PPli/Wc2GIrsCPjATHmn9zveydMy6GwYpHjl
dTbRmTH8nPMMRRiOVWVju3+MaIMSE9268fK6ZX4d7Zs244H1779qzRWb0vg2DK5Z
lfYNLPkJjD6Mm9SnjWDvYVvD11YKimqFb0g51uyY98zCIolXfiyHll4aWZKxa5ui
aM62r/7x3qPSp+yryb9SFFF3VOoXaRVg4/pPe8ydPb2tyFezi/HFPW6LjqkEJwCQ
KI7yntNC28S3MGT/gYO1haGBJNBMmgmgaEGjdwKkaq+3QdnoNZb8990YWkiMzjfE
KbUP5r2jcM6sKks1EX+WuzMzPTozN2O2FOfFnPByT624MT49ct5huyVbf146gFf9
hB5IXRobwfGx4j+gMIzHq15Zka0cQJdIYgLW5Hvyx6D9pggY0ZoNfxh+XmO8AzKm
qYr1j5ZdadO079jfo0j0eGxPn/yJ1gdCybl0ptD9rAVTBvLroXW5fZ7A74fkFN/S
kmcA+ehG4/JCQtwW2fr+IWNYNNcDa+aABwsNTrFHk6ichyaz1JfZP3FBbebSLpf+
UUsWy67SNeXCegUb18A+EwEFg5opc15Apg8/TwYjSA0VCRiM9BZ0A8A7PLM2apZg
p7Iex6noFgnsnpK2BXxGcmekm08WZnzkma3Q5Z0JntQES+BNufGV1VVVA9PaPtHP
p8TXCPjtCkRuejcldilxeG9U666QHXwJBTTK9R20JzsKKiIwB9W+5XEtOKD9DSha
LhTvZz/kUyAbd8SFX5aZLgpt7EjsS+RDtkI9MIAyvlr5kcTvzRNic7Xj2lo8FT2c
pbx4K5ZtXpBXVPrt4ACq6BDz0ktg6gNg3fV2INS60BRcxswgVDcsKgxMR2+4h9k/
4Ew8B2edEzQ9JIyiC2HL4jDVF3+PvPX70DrwySi1jwr+Z45SY0e5WlLgOx4VUYSN
cBd12K/Nun6Lelbg5z+BkVdqDzfi47rNyy3GoCEwGyISKjkIsIy0txVoHpfSkxBv
ub6ilwX7qFtueZtYrHe0VONAkF8nU1UmxehL8PQ6VkKt5eTzVq4bZO5ICpxs9Rim
7nUG5bjKOxmVI9aGQdBwhFp3aZhNBZz/egM6zIEbxqJKaJDH9/MvaNf/DF4xfT/7
UFxe4ip0Hhtl6kwIXCSFlCmNAs2EMv6URYFII+M/oQKHh1EQ+VpryuCw5J2LegXR
CzSdYXeeQyyWsAVe4pQkI5uMYsmjn38epcTYECBFdJCm3/km8OwbvLB7iugW0/s9
IsE1fTJ9uf4lzbFaVAGXi1Ztmkyi5EKiwwZbB1F3rb0Lo7YERG6EXrmcrbnMoGvl
MuoCSx/4zcuBxSuoazXJbVpw1KAzJl3kYHLAH4VmLTqxJt2EPfuWVZjFX7JFD/iM
P09SkbsVDcBGuWActebU0JJkhWfueDrkxi//m/cJDNDwDp8bunjKoOxrKOp79QCn
5XpUa2LGYCJUlCJP6jGjYWEnUbOTzI3ypcbRlB3c2i4PfzUsZBgoDtF8ykKouQ8i
be5dP5JTUUtvQe4UlJ6JC/70WVpf1dKkf5JXAY24omAL5XN4cToqj33f2dQ6/uCm
gH8TeSICXQ+C/S+wq12WblZZHtnDIgDRO5L9T0AAjmFO15vdCflHFsrhEHHTHosN
PuXczhAMDiZkmTNdZdOkVNMeZkMytCYNl8hKgtK2fSFsrRRE3Sdn7k4EgjSrzzRr
UUm6ff7EOi5dNOm8uKNu54twJRtSxUS26kVdFNuunKMhR6tC1vvMg/ikMrN1LP3C
P81CTESzEZkQUfQ2bM9TKNv7TLphM9+OhqHC0kZs6NIabWWTo7SMNXcJETxbflxB
pRL9pFdn0L8cb5K+rHVgMUEzdRQZq3HB/Map8y1V7aQhF7QEaE6SD+w4BhrvjBjQ
EI9nzXmquEdZBK06aLAZ5EzAwAoQvBJcc83g96TRplVjjNeOnGqwyHv4tQaZ6ssc
OwZpEsLhI3N/loaWobVYdtb83gXHcKslWQaz+X69BVOPxwt+oV+KELDpjyI8HJ4d
HmEtq++aGojGOX+MVqdDJ3NJwVfA9cda0ktryfwAkB+jJKhxPIhzwaF0vamWk4xE
Pd4HMuKhuyv8dbka4DFSHycdtHpe6+50n+XF8QHOis46rkP11PmxXl1ITzDLw8U1
xg+jLMH8cHP/rM9aDI2zu52QnWtvLlcYXMXpqkZ81xwooofnuS6gKHEF12zdxu5F
qN20VJlJxdhGaFZ9jfiaKjoZjwK7kEO6rrwXcV0aXujiFZNXRpWNHlPPzKZW4rSI
x+geZUHHZeHp1z2a5B6exCBsp14JCIqqZzrhvYLwmIpKwp9MJa48u76kls00s4hr
nVQPtvcSG2JHlznK/bXtnUK0E6k1Vec+UIXSIEPyZG4yrA6qfQf2c+kzpEI8DUb7
ktCL6tO46crknzJPXrNOoqSg5URJ/tTOK4icSzSn2hW/+KzQXySHaxmKYrMJP3PS
oD1c8RymyYcbHeNXFUzl4QH1DzbpvV4ZVuxdJ+2HWbwAsaOpVQIpx04zoGaSWEDP
2BxIsRW2KKSVgbqm/tKVJ8EcUFVQZYaBd/qfVGZZKbnvRNJ7ywwAGqsV8/R8bs0Y
WzowEnBVAj7Rlp/teUSSF0OUISd9iB/6vPpuVOAdNGSbdAvvSrB+uBExbJWLbks5
mF8AMKVvCkxBs1qq5f/Obr2IxGLmgJ411gysTgEOFnBQY2Q8pLSUXHj3tRlyOeIY
9MkJ55ez28inwqLOiz6PoTEyi28Gi+YcmnSFhR0RBlVHAdZOrjeHssBbPaBzDB5j
8NgQrMiQYAV+Xvtuy8NGQaLMAMfALqLimSqqY38HOjsuQv0CYwPQ5N4jpoUXoOQZ
Ta8zQQNUXfkZXJvYY/AzshYxVHKNg8NzAyDcP+SWafc9YXoXVNDP6tGfWQ7nJBBy
zNFe3UCtuUjSPan9RfF3QwMaZksxhZYPS7ZxBMs13ATAFfyzWlvl37D9MNbdIhNJ
7hJc17BS/1tVtUct8Ry3NGNHUUdbG2v2W9zKg+AnSewIvVzuwrFPTGH/vtgiPSy0
6f8LTAfY9Xft/x4hMK6hZIQr5PtIlA+5bNd74iWN9NXAX5A+Y8pOFHNJxh/Res8m
vohCyPWW/gCBw/tnizoFwHgzQtC0fJ0rzeMgjVS+Ezvo8hLlKsvTHRLzoMGuJj06
EYmst2P0tGUNvn9sK6TPLG9OOMiPJY3Ks3j9ShPwEgx6fhbf4XsiB4HD/MIQRiv6
k6Havqb83s+8Bc1UaNbmn4r7cIVcjv4TbZCapxVZRDrqzzwYtHh7QQjjSOQIY4Em
LYPKrfynx9c7i8ix/H/N5jkRAEhavSFktiN1zO0FtVQhjgqo1+v1+JxGjMX9N3ZD
4BzCtHHoH07QTB57XM4mEy8XlwZkn1OltrV/k9NJYN0pAtddy98wLX7CDvRIApUP
NOkQ0IGoso3fEFUTT8GocJTgjYKMxAHtcSBnmb4dXeQ3P3t71pfeJjunV9iladwo
Kg6hjrC+ysF/sElaeeDGqZKsHnTXOQ0mMzTFLvUUtcSChbF5ONFdYtg2jwKMrYU3
7OYE5DXZE9dpkutJFUHLFFwtMTlSVzRjEi3IW3Au7gFU12fHg5/gxDb7kV+eR/qR
ZUukZFKVvF4hyIv5iuw3Y5gSL4AKsqahNVP3InagE+LJMfEm2HibxFpcLIEri/WF
eijn0U91ievF/ggN2vkOaAI+NsUGFWoTUBxGX3vAeBZJMy/suPRxUCIpIEZRIed4
AJCMRRERXowRhxlxm0KexA2qhCetRqtrTLrxFGIy9wjaWgGhgyJ8DyGBgyi3fKLY
AQaGc6ufIYOrvRqGfU41kt1WJ0xe+rtWmDKKxclyg0UOZM08yQfw6fGP0UisDuR0
09JNrAbAvjyZa/cpC29aO5xq5lkXv3ymxYxXu6nbxsgt3YJP6hj2dxFAMDe6nUSb
mKbjW8XvSSWSu6pZfzFKRwe+HwPei7LRO9Svu1p+9XhUBF3Mvdl0H4tK6dsGmcI4
QMf+Cl4TdZvtfNRnyr6hF4wtGXp+QFqL3pGZielOyPDDzDTXREmHtVGSuZAuBmpV
0mMrkfYEdQWKJ4D0NeYsJVTh4Rk02sv7DFwGA5hXS6L8pSt1oTAJNatKv4J/Mpex
Ala/5wl1NyvqhwsviA0Iw2DPISVuJaFtINFS8ZHZ7TVaPEnYlowC+BQgX6iHNWIz
TUQmte66lL7EJSmev5dOi3pWZh8p3HlxnyjvoY3Ip86f9xi6lHYRrlUOSIkyYf9U
UOs44N7FyaRJQsROyfFG6HQ6fUmq4rJyAZLVYKwqfF4DdBzH/zimHChhxPTwJJnO
L9Ve7n0/xEOUJf1+gNolU4iOl/igaYxGgVYc8LIdbWSsVQ/iRFpHpA/s3Wyqj47g
b9n5eHC2l7m3Q/A3cOrcJvRholrMqdb0VhS5uJ4GAzjZGvPWDOi8dfY7eaDo3NLk
S339l1vddgfQcvesa7+QDU3D2DdcbUKB18qkVc2PJGa9cnKzACCTFVVL25XyTj91
HH/1wJEYKp6BU5f4NUlCfyBXJjpukgXlptB0r9rV4tq0rkNqZed6fkKrU4CiLnbh
ypzM01SNCqsj/7NYJtnudoPRhNDy7ijM5En9iirTiTuMOuyfB+aNmckWFBfTnHkm
n8ij41ltcElhGGlK0rChdcECWV8YPD/SJefFy4tJ1r+elcnx2Ln11J6SxZ9OSqpn
xlDvB5WrZqQimCJqRFqlh/dQtjwj1/4yyAWBRVH4JsBga0zXOWcXnuNBolU5JvXx
/Kqfjh0SZeRGWigsanEJY5OsVGKrznBytVk+TwYKUmJD26p7WeX1OZkd3u4TGLdf
7K4mjGJUYuv+20gYJ50/MVd3Xkzr4jk184NiTzxgq23aGLXVRNQZwwgXmpI7GWxB
k2sMSq7EML2e4E60MaqK25K1le/RcnMWIrhUVmVzMlReh7EwkIKpwRJ4NiBRgoqO
gKflDjhLYySXJ5buTuv+Cam+WaiTzYAqXPiIInphaqrdu4/DIACZpTx5vvwk4pXd
H9fFImUWli2KYcACFkDWpRKguxKgY4YRbGiUvDI95IirDknkZNAPtGhphun8E7CH
jsbd7kddh71tkOjUA8NKxeAj197O7WYTZDuhUgf3MfYW5pMT4EuFWBav5UhW5SDr
HvptoV372lLyoijPA0Tjjh1HSWK2vKGSdl283bj2NQoES96vPaK6FbWE1xSgCn93
+ofB2RKuvt3ORGz77x/7Gny0dkDfCa6g9yQM+UwGHOrnem+dNSSKkxIk+knbny9h
isOe1pzXgIkz1hqruKAugzvjfM56MpqhD9AIjLX2f/bqN+zCe97jnVVRD8YeCxiu
6d+rCSl84VQEhgZchBik6rmLQCMM98tAPdanmPMseoYMhLfSj43fLxGEuvfz9uvk
WJBNN5m7r+UZuiaW+YTE5DCkY8EmTSsyqFpQvg87+E4bI41trjBLwazX4MXbVkvX
zJNp9U+oj7LymATJ3dWBML/gNFDKV7yyEPGmKkMr4ke6gg5hGARaPQTZ7vO/cz7T
/+cFvg06zZgB41jdyfyXTqWHIXnnq4idB7Aq4IGfTyQ1QMCgB+aMw4rpJP/0NlcT
O4z6iJTa6YukwOAQSCUai078d1vIIP46hfMQROuzelAXQG4GKVBdUo/T+0Vd42MJ
QuVJtgqYyCvWhxZ40eI45FYZfzhheFpMM5xCUXW8ISpakcsiAgoQw+un+UyIlgTR
rZqukNXtPwh8IQUcziWSvi5zC4hkzkmlW+xPu06c8rgwIFx8z13Dw0fNnuL5mOcT
IpFoRcX8ypeiheq6pO8OcB+C+P68TH+My28hf8a9Hgy30GndW4505s1gTF1KZMPj
xEWTzEItFLQzVfS5PP930tYFCvGvSI+pDsIvFVqlYutQuhh/w3TbBtV3/cq0WLha
OfwaDRoo7ByqvDgTMYmypeJfDMxVmJa50YAATdKVUV+8LyLq5QdIKpDEZv1JuyjG
T/ZSf7m046UbC7XQR2j2aY6+RmPrnXlJELF3QeIPErh534E2amRHpP8b3lwP8yP+
KpALcYsoN1dFrPcxrQIwnOgOrHdGOJTl9OrAKqIOlQv6Wa32RKganq8C/4WUi0Cx
iljZfLNu2VhX9kvwFk59kTnhisyzpyPTwKjMUsZsMc8UQC3m9H81rf/opinrqcCC
NVFXOX8QWvXdNQSmAosZrTQgI2Btp1YEBMOPet67BGPiJwJFJ42yg/LJavAloR9q
JFPOjLPaFn5O9Yv1g1ZeAtzvA1ej5VYtqoTrNAZGSUf5AAb0hAMUuAxFc9AT1uTG
G+FVYyne2ZFDySqHnr1Opl4CYRKLCKp4k1pQWY4fcJsZvewE0VxcVSVMLW6zJCtO
qbvw3jOPO298uBqvIvfCvok6bEN5eN3gZtNESMM4d33KoPD3RRdxb0pNXJVdQBuX
K/XsPOU8sqojN1Lo6Tu6+iEKVJhC2G7Qj6dO1zDvOh3VgkAH+Gi/pKli/yzFHXqo
ba17jW43R+W7KCacSvlZFoPgTHoPDlnYeDu1X1PdszQ/eTfrN0KLbkk9pyVubT0H
F9RkCsHyacOyTBju0hdix/B/t+DRffc1ymxk7JBqw3iJ5AabYY1/XKbnOir4Y3TP
zVmMcQV7+S2WWPeqXJhm6mnz8vxOBEipPb5DMlYd5tSCKUySPX2qqub+ltR36cno
jWEM3lPgZs6q5a6WBB76dRavXUOx/6MTXAfZ1hdpkYHbneQA15f0Tml6zTT/Giej
kktXIRk1BFlropkkV/v2C/cCxEP0U6ChOm6Bbl6XKUhVGj4a1RsSW1+KtwwMOgW3
soDsCu4/PwqEi8NT33pvweeCZPDZe1beUjgRebaHCynl+BTxlEZQ8XeOVexsexVC
NuPGnRt32Tt8sZTIIWp2F/j2rhoiTpINFFX6FZscAlN66JuQImk0j4kujUbd1jMf
1Yw3gsHvao7rhKBjk9aSch8tO/1ABaF0aC01GKbAOyzjr1vQbDlk51TLc38LLGKL
6A0TVEUzn3CKc/YF319HUxB7tqTAui7yGIdWJ8YUO0VPq2huKz2K77eVdKuTmHBn
qNI8Bs58/jzCfoRhX5NlkxY3yf1AfILNLPwyJLlWFuMPleE5GbofyUKJUAjCjygy
/zAnHE/mwiQwsqHS5/XgXJ2CDhD2VxGxM9DfCPMN3f+sfnfbnkPrCOqddqOodhaM
NoroJ2XajH5wjIaVzIEiDAMK7QFwRAOAw3e6jcZ71KbzLSD3aSDs56wqPWICuz9P
lAlLif1FkJ0H6OV/sjwdMMrbLe/OhxOW4ENDPxwTolNo8OCYYUHqlvP2bTCihBQ+
Hl3T2z/a3PKjsobsoIGsf3ZkGbidkzn01vA7Y4/jhskQrMIImys0p5q6UVoLYBKr
GA3q5czWHilVuZ/lbpgzPk3vhEXVd+KelmuWl74E/6kWJXkbBrH0/SGQ6YuDHQyp
bRjCBE4ji1wcvnBVqbcHVgN3wj56+eniVrbFheh7EMVeJTxEBEk89ql/+qrMcE5b
98D9y1D2jJ0HPCnYUzST6qwbZx67Jwxm90ml/BlfI0d4aAwh8v2aFJN77bAugmf7
eG+NSBGH9bnpwMoqE5PZiabQcH8PEoWDe5Eue0VVQdbqBtISaF5/7jfaae1Dx4xZ
ZDLtchWzMk+VLpt+z4fxVXgEUtCamQrXdTR0h0bwxlePI4riatHNbnHpb0/lRjrr
ttPr2Ig8zHKPqzQBGurPFCyLtp6SwrvffkOJ+aN32KFtlJOiC04ZlImFVG1L6anA
RxELvvy8N5GyeedOadpVug2HEixuFRMUzIqlTZ5VQ4BtP/M7ygY9QFqOp/hCPhTB
5kk3P49ps9gIhxLaS5V4SR/nBEGYU0O4okzfrxcTXB3E3HtgDiKPbC5Ef9hFXacY
9fMiDLgqV4IhU9zTMSlYe6ZLvjDatRKO/3yIWzDv21ImAxe65sg1OBqg4VLSMU3j
fIg0x8hhdKvImcbPjhe0R9i3P0Q8PsYr0yS2g5gW5O568pO+H8EA5CXbnmS6M3gI
4apaDQPSnahOtM5nxjUGs5bPDT1EDEtXG1/etmR4gv9hri8tyBywtR/CPuvM3sFb
R9mSKdraN3s2FfoM4my9ztGD3+F4Ni/mzWdbyklzdS58ote4Xdw2YqX/pUy7Vnz6
iPHVnm6Rzru1MW09MUfZbKDg5cb69o6hPo0Y3GUhA5786GpcxxLp0uBNnLYvmARD
di9m1qdop0363LJK4CG5BklC7J5aIsQK0n9TiVrMmgIghZ8TDUgDMLaUzdyb0F4F
JJqCy3tfq23UWnyIK1T4lFK61gsFJbinomlcwu+YzmlsCAAy5Xs6XbciEQ2emcfS
tFjeIUbPzSvizjr5w4TVdQfQnOxRyyf3Droj9soge1l4Wkfx/im8zEdnGgBRF9pY
l3hm3ZJ+b23XvgJqwIhY7D0VDiiKK5mWDBP7yPbuKI8zGOFdHu7CHAspbQWuV7fS
YKhk7LQsxeGWtsDwFKhfZeAFx6qmFGUiepAOpJYgLOesc1QBW91ZeibLq0mQU3tw
mmpk9Qwmvg/mghWqX0+vam9oD0UZnb/uGeDcas++5Kzim7dgHmk/+seEibUt+tq0
d6YVAAYv5RJ2kFZ+kRARFu+MbilwnUNge3Zm45gO3Qr0sHOpVDAUzOvR+vQTpo5q
UvaPmJM30u1kmfJoekFb9/wRUfKupPQMGLZ02pVHaEN+gspP+WhcrHHBFqfSGw8k
t5ldYFvXaZlZPkR4WXvU3oqI6/TlZBRUpwXcdoh6ShJDXWc+AoCcYB7en3choJZz
myll77As1GOVYOXlWIqU67mrxpg1QI6tv9yxMYzARB7Dqi4rdKcfp2Hnj1i4Gp/j
o2UmHxbpJWY0UKpE71u4Qg41YUKl36U8LGquNv2qQemXleHnF9xAXg47qpgEItUg
R/RL+G0xN2coBhcF4h5dVKhV27uojLD5mOvvUTkFRDpsqsIAGXxYjLI16FbWOlna
ZvYlEA6CQ9CT0Jinq9QniTpdZ1a9HkoEayN8/vAcb/YOzS28abRGW3CYW2KZIxQw
mcMNRvktorfsMiLrzwNxb2Kv7VBuIVj8hfuf6Tz63xuK2pvbsQDrcFx5TxqCtDHQ
1TM5oTY/fUgawWNqsBuSL5cy3c4NlfHeUCL/hdBu6tv07VJzB7FDNAyB0w1G7mky
848gB1+xQvhzMdmid2hpqfygj6J0qzjgJYAQEbvNRc/aQVchzhN++S1h/SAsGiT7
670q4JHsKlYKVLO5torYQJ50zAnyuVYamakvN6C57rDN2CX5kd2XMLhfFgWAfcYa
ExOyf04gogX/Wmr7sewKkTR/3mM/sgcaYEB4D8Z6yESWWMOt68Y/36RrlGz4f1Tv
OysRnY+HmEvJA4Oe3K2dX9kty06OKs6Z0ShJhsYmaExZsvtPfui3FztLOIoevkvY
AltCxBASohiTVoPbTfa35c2obcbMt3ek1ZKaxaDnENOOqtr2x8aeSo/cMIl1ezQc
Qe+9dDzAXGNvmz+8o9X2CRlpGUCIjr9cgz0uibXMhxkLq7R+Z2Je7ANPSJIstpdu
MsGOgc18nxcMup7Kd8uhGWbvR98mAcrR2CUzaVbHZJKwZOKDTO06xJvK46NAdWiF
3y0sjHryI81gIIv/q/tC92dpV4s+JIUEBpYhqLtxL9m5waHeXxMC+8HRHMB81BLC
YDWgLa5VMzNiNVGmwAE1sz1WsPgGBjj9XcCIOanZ+JM8KDjgcQ9hYrX0QOmnENWh
KLT8Jly/Rg2FcWOEHBUq5TNY0iUjV7mbkaw3FSf0PIxzWQTqs+2840W4zXc/pxWV
pKmSACk8GqK53TkuHtUH4hr1Ubm1irISiQGJsdPkfmXVrP4FW/Wcg4zHXYqOoXGz
UbgRK1yMNC0C1/JkDWZzFNdhiObzxQN5AqIpd9VKq1k52L0vmJ7tzyVPzxadt9rA
bKyi2Tnl++NNmsM5KCCqRgmIHEfXe0+asnM0biw4h5DX81wIo6BfM535n02Bfk6V
nngrnq/xQ2TijLnVNCyxUnJceMOAkey9cP+CoyM1kUSqqjPedx34JkzN6ZjcKTON
gnSnqUvDjfIl3Dc3B6Ejrd/SoLag7Oc631WvDuivF5CdvD7GetoxHfvp4JC1bJX3
oCIKcBoJhlyCWY8Ww5oc+mif6VwlA7s7FLl2XGQMXOpnLf6LB0T0yknlHvpnVL6Z
KNwqunqOyRPP5P9tHZPvmy6NSI21CsF9FYZFStUxj3KvO0Oewwk20L+Dp8f+rfCy
2R4QXas51NYfbqv76m0xiS2kJOna/Gmf0dhooN8/yBAWJjo6uPlH1x9m7TIRUDfg
3k9atfnX96JF+diMdy7q8H785asESiNHqACaz+BGf0Ii7eFoVh0c7MoFrkawKVAB
W2m8EcypixloYA4YML/RA3bIDJcoQOKhNlTOl4cKV7Upk7Wwi6MTO2EzewiDirN5
VS3XgZFdNAYGRp53q2h1hkadEsofDXmaa7aT+QPK+41gJlkt0/peCGl3W3aCVYa3
lkG3n8dD8jsbYnyHCeWA3t9/RYVgOI6fGAAkpxEWeH5nFshfQxWaw02dg0JT0FjG
tMdhuTbzeGQ8TZHMW5ou6zzlJDfSiS+y3KjBiyHdYBl4sHlEVEhuEn+gt7QAGy1H
uH48V1hZvP8kJv8BADOhKLP2hRTBj45TlV9cqvxsG3ruCGsbN3FdjpSdNzrdC13+
m0WbGAk2ehQ0Qc7au9zJcYgffeWj4E7rjraNHXmDgByGRQp3ARYgB7iAPOxPD1bm
6f4IMzxOWLb9MTiabsHugqh9mFgO3oI4/86wpslBG19DejcBtA8Zh2l9ynd35g6O
nceufQgxchP6ZAOUBitynM9lN8IyCcgVnWi8LmP9Hk1itV/J0xq7YjvwSYaLaCSP
l99ykEeiFpESL/Usi4vxTBNmdp074UIryBaGgLXwJ+q3Xvvc8KDdsXOvdrbxUoTJ
wa9URpSRnf69h7pSViRJAvIkxnaD7E00wNiaqCno48oAY2/bfHmsf42khhhKJxKe
p8DjWFn4VRuFhUMLffBvMklf4Yh0qr3mD31yYpBmPXH0HXt+AP7XMXgUh4fAaD8B
j29qctcD86qEkLHLSM0vCmTs36WkCzGLqi7La9PGtlGxSbhNieTa+d9SNo+43c+D
7gkNKb8bYDuYCrwG3BJFfc5Rj2lfvGqMDy53z0s5BbmSssxKma2m1I6RMZ3cVG73
I5X3HFVQY9C8FuACSmuWDw69y+DFzJmIY0qigioh767Z8sfgiqPtBv/EXNf27w55
2oDOR2twiCe/OEhgaiq/geeYB9HArQ6bclA2noT3jNvaaXRPHLo0XLcuxGVcHyF8
0gt+87/FfnWGvuMvYWp4wt3k82KthRJaCKIa53Z8glwnyz5fsQaxmgZLy+sZ4CMn
s/HJeF6LKBB6BFTMIsGe3cQqdLQDbHnNHoe7VkUtEfEB7p51OxRpdtCbiP49Kij7
Ok151f5uenvxt3hCEsbUmmHsaX2EtZGM6f8g+IKz3X41z6FOcaGLl1654O4eG4A7
OXMQYi7LPT0fcdU/p29tiY+pR1w7V0n1W0N4vEPxQ58yNnKkq8cmJD9P6PbIS4dd
0CNfitmXJzyAT3fCxc1ory1djd7CXFAPneykn4US81RxbrSWenTFA7fCf5QGbv1W
KvVbSmiTtm3M+p0/Yr/39J1scAj0uMrT7eYV/w26uJk3rGayEZNID53PuzcnTyMf
8bN5L1/2MrSXlsQ5/FsSn/0LhbjF5v8jzck//RJfsYc3NOSxABuyJoNRtji1fEOA
06S7yCONfugKqQHBYGxug3fb/QrSLpF8vYwQIPrSp7Zn+J4j/nDbk9SKlNtwXYf4
ar+tERRycCnqNiGsC0wqGak/C2KrWLw57g+N5/Us/qMcwEt3B12kQ5OrjlW2ynar
ytGBeLjZS18iShVocbMmSUhf24xma+mBbRUIuI/uSM2ErKt+DNHWRryZdl3mPFtP
23k1j3NgRZqxXXaoXbn0SfoG+iwrfggfaDOBEMV0/1EolO7lWr/ECA7Hed9xKq7Y
2+yBdFQnZxHPo3R2JJvSs0g3wlQutRJyOvrtbL0yw40qcHB8+JIMlO5F5gO46kNr
lFPEy07sOlP+BF/ZZvoIG+iV99fk4+YCf8fUK1HPaFK+cclxrXfYiq+q6LHcNAeF
DDWY+HH9x0pKz/anAKviBeYn8WyEx9/XI8PTIPnbH0Whuv772TH1/veIXaEN+Omb
oCsaPqNEJeS9qw7WdFLkzD6Tf2a1H50yx+UeoSzVdvuYZzLMOMe/YVHYaUjznWcy
xAH/9tUoHiQH6PtqScVY3+DMtVkxTdUTwsK5jn2qD0zi5qwnhIy7cMngZr84eC5n
0ubV5aVt6OCWG05sDQQZv2FAEP89Ut7l4/4nRppT/sTUIy7hQ+QEpLl/LsFMmOdz
UKZ9F2jpFph7MiIA5Mia32n4tkoxcWPpe/mpacs7M89cDlbT1r+r5xlSBvfMiumz
0+tFfZ3dFMqk9WDfHSYugHVfmARLmOtHhYoslzslzmt3BH6J+vVNVVAkxf9Y8BNv
BgqbEpIW5jNaGiKy2c4QDCcCXvB+FaAYlqoeYhRYNAjz19AccTrygrSs4HX1qNy7
IVnantu0dBtcg7XTxScW4NSMxWqpgavqBdt4pono6f11fbuWHepzSMdKnI4KbcTI
/v4VyrwTuXWRFaAbzy4FpzABLeQHgfwVLZPWd+4Gq3yPxZkgrpFS6FkeyK1+Eh2i
p4ijj4m3ieiD3ylAMGYEbmkV+aoCvHdfU+IflK3EIyxJ26aP51+wN0S22CGL/ei9
bZn4ZUIBt/AImJZpdtyOF15lJJ+34WHAQ6q3w2VcYWuAmFo3kBjgWsLiATVOOPfs
SdK/On/Uf/KkaT63X4GmRUpBZP1JWRYuhnlPVTmy9lWBX5Du0T7i4JVNuJUH8xSw
y2Fr+LP60yk8/430w8iqqeT7PE9Ql4joDIQl2n77UoSr/E+3vJ2DFUVEz6vHZrkD
5mZt5e45IH8+eP/nx4gu+3WkA3YuBjK6mj3OazXNxHvlegN9n0GtT4knGgHfwRsg
CKv/zaZP3lKQOjmY/r9VXlGN112mV3fEYus0j5G41oma2tzvuGKdHh4pZOPd+Bwe
71o6OsVI0s41qJDjKb5b7oPNzqFmx5nA81erzX+QyihvIviX3aw5P4D863b89a+6
V4nXEsU+5SE62fiRlqPJMDywcXfZATnBuE65Q2CqKdM9e8polmpMlMAVkkPVKCbh
9+5yamwL3CLEDXcDohmbPZo/Kqd5L/9TcvtDW+nbe/Sc03wsTahF6XZpi9g8P3SR
Fui+6beR9qAOZ5OJVTBgdvmAz5PZAGjFIZeEdQfl5bBtOVyDN5brJ+b9v/V2sYwV
jpjAThqJXqsjjKyRWpwPzN9SOtQS8IudWUjIHXgCVqqDcKGdzhqoAEh/yt8/zN8a
XkY/ygUm14/eJBmUI4Fg6G5oSlIrLFrW3u2/6/sQxwfvpUXeOxsu+sjyBgQIZh7r
ahb5l/Azq6qbbFzv1pvgv5VGnn7k/cvte0tRCJPLaAmM3I8QAF+AWb+0OpDWiOgD
zj7cfGv17bHnDdWidHEV/mLY8NS0s0ER/NUfTiBQq9mIfKKWF9wfBowbPt1SZ2JW
3WH+6ThHtZcbt4ISBWAhbzEXMB7Mx3btYPDkER/P2jYgLuffq/5la8+FDguc+e3+
DTbgjxJAhw6NzH0QC5r28BEXgL4+x56HaM8Tuz335gQ23p5mHn/A+fNMJ7ttpCNo
IpoVvd7a4vci1G2YZEIhjs47LXeJDbu3+ydDp4cpj4ITtrQG5njubYr+LYJREbqz
gTMwLZguN6Uk+MvHNmYhuHeciOFR/Yu3uXhnfeknOliZby15DwJV+qkvoHhFliXe
qjsUnUek5pMqswQ+Kglo41+g+YMqoGDKg9uWMItywJ4cvV6gqq/PqQe3JcyeOeed
yVCSG1lRoS7WXKVuKBYl5BsnQ8Y0MHGB9DioxzyajZkf02pg+DBdW8u94Rl40Z3O
W8+pmVH2BUNjhHDf2JXemGxK/CGOvB63mHAcZpZWwIr+aQ6fkWtMzT17uc4TddIe
RhXRu5eszrpXePS3fxoBHGHjQCCxPKiaY6yO2R7R6x7WSjqoJzSA0Mgq/TYIRvWI
gVCsbMuoh7JxKSqOOAD9WH2eiYdTSVn6hQVE9XDRp+Z8nnwDamJMo52wuYEcXOAK
TBYYcR+f/vTHk5pt+iwk+pQrldCn/sqg4l5inH9+3gXMIX60sLq9N1iHhM8GNjGh
tdIqEj4lLT0AP/n1GittoLFFvHvK2QygVEYdEzoR6DuBFQgsLkCuyE5EhQLzURk3
TJjS55deZvovtll6vPmaDlc/jXGAloNecHjASQtQMvZxydMNX3u+YmNDsJ1B9ULe
pF9k8j108Fblc/EIh4slNpubd20kH5EHIX86UILc2BPfQ2K0Vketf85ViV1FG/fO
uD32cDcSw5akPgFLQWid+KKln8meGlk541hUUmeVsEt2l8CR2rXzUQOnKFxgVSaE
h2dG/s76Zc+ZeVoNkdKWZfraksxlaqtqEtXiTgXqHFIYAcNSUHjjt0fqU0FJhDQq
z4qFDvRGwMMtAecANrcPbT+PGmwE5sEnAqsh+SZ8/DweAJPaWM4fwJk34Qx3E0jY
JtmYhi2neHDRzIlsYEL8yqI+lR8Y5AZqEDqwMPeFox4IZcUUMoR/H+inULw8EYms
tB9hUBrmITLVl+kBSQl1B2Jgt/84n00NwWVX0v9rv6EJ1iTeBIpyKQCxiWMEPSPi
6DiL4qiufZ9Yz8DczGwedk8yaTFNbEL19trEWzB5VQ9g1IKsiTsbAOWVV1YwEtRB
Nk7aNgd3aTpoJUzgKcZEeskQGcRzmld2mKdoyGP6EwY9+Y2cTc9EkhYnk6mT/nfw
wm2UlgPBJbmxh+Yd9lfmnmHUEr1BeHtlvGO2U6jlptih77TGBLjLxMLHN6vj735W
ZrvHDOVQYO0Hak62bD34L6cQGDSovHhl7FX3jetRF+QtoqtHVK9o4TCFx+WQn5Qq
2EZ+XRVxSedweZNbMth0BQpsBIP8BYf1TJXXDKwJLLLebp6gvbleb7ZGr7/bloTT
9NZEuH9uixiEuIcf2q7lwtNG3HBy803TncBOg7B6MvPg1YNovDuqRRRHuwVtpA3E
ick7QKHPUIaiO6jkJ8a87Yg7ZMV8NqjSVCsf3Thml1GJHUSrfqBVqhkZuQglGBp9
bXbGGv3EbxKyYRZw3MYa3E/a1TNevcKkUwx5npiGmE+6tX2EFPJT6X6wTDBSMXF3
bZiJbJ9fFsefHzmKtS9yIdCOJgp9+Xx8fsGGdk7zsuu3bat/tkBESbeWRH+Kciwu
9nHbXRj2ol2qymS3WgrSySDvXd8Q4d3KMUXrFPJCyNjE5zyqghG6PNoHbB6qnPIA
Yr2Pfvs1cUQep4JtwdgRSqshJ18uTh8lF1H6BLEWllF7FaAAMI2K0HAWqOJp7ebm
XLAzfG38sgtiR6qCZ4Q+9m00PBiFgbZXV//tP3gY2O8cdaTf0Cl0CIafwvK2mWLQ
yMvPx5wGXkQRe6n0SAZPy4fjPstdZdurHCshRvhHX2Nev5uoSkRIz1JtIgxkYNQT
nhZu68TSZASg1OsecK9QjTNfWoa/gaYg9b8F9Q6nAjjpKhZdkERUCGmBmuhNWq5m
HLNq/jOdzzvGynDI7bKt014euHZdNvtwn+h8VG5m+rH6dP0fursR2QuYEMhj8AD5
7ngel00k5+X3HvwrjohtB6tHIkeXJ12rmE/mJvRaOeOJnn/cm7enISiF4lWT9HtO
3XkL2dPkOFordP+a23PY6PQnJ5IrGKWKjKyy8EPTQnRfbRGi9L24qqTtLex/hZ5R
VGLGuuHY+qzdNSC4xarcY39mlGohUukXpfipXwLNRNOcZzXqi+NRljZv2WeblAVZ
OUN5FhNqTx+arw8Y2IcfzSom5gIJeLZsQpar00Wz0HOSwJo7PQFG4S4dEmi5eBqz
471IWBVzrx3wVbrKOtwoE3Y3diPM8T0LPwa5JX8hHx+BFPl7jNIzHNKZ5CAD7xgR
kKk/SLDLxzqHkIlLQu3gF4cgzM7FVSqHc1RPJaOyX182XvqAyq0Au9U09AaWAtXu
2BSxgbdZASnbBLYoAb3SVVave7Wzkc0/4Zyqp7cuXUj/8gnW2dJE93EvjB+9/aSB
G1eUZ3xpIXIJGJeObAvJpda3qi1JEnlvhWQlIZP1fA9Sz/mDzTASqVQ24Xut29P4
lrLFWoxKw/ALpyIbS2mo2DPaugJTh79mNdFzjvTdRfhSlzuAcyng3zH3ZyMSXAu7
qP7iXiHpWo47bJ793tVBm66gQinFEnqKx794CdvlLBLE7lqVx+3b1SXRw/pTEG3d
tT6BTbp2/oMMggeAllfhn3f8UNgm6iwDii6pOAxkmLkVOOJx8/UffaRN0VK74ptX
hjw1a60hzVEK0EjpuFZXh0viGiH6OG/51L+dpGH/YiWU/4/Dt11MHwbP3BSfe9eq
nbP4ChuRgrktccuuJQZUpTQYjsKRqdgXT4bCiMskm47qk7RKe8k0ofDgC+7IlBmc
W+oJhlKH1rvznthbtAJv9ZO71rHn9G+luxc3Bxw3EOxln3dsUCbX1IKHwNypWajC
OWHH51ZqgMkhNuyuiT6ZaxFOpUSaNLoOIVttOcuFpkqK6AIcTqE1v4UGwv3e9IId
BfuV48whByyutqgV3Ch7J0Ogf8WDyU2L1GtJ763lSxyYfpFF8nj/koHpM0rw265d
8Aq3dCjllg3WvgALdaAsiE1sNyxESr0I3442QlkD7FiusILJ/ga6nrVDRveOZazc
VCpPFWw+S9xFvfE1jA9K82qX6cFWAUZc8g4Q/SOsCxKrvV3u/cEzyIFb49nsDDFp
OgF/i9eMlurzP7pPJi0LHO52sm0m9FskNLYHIidTI8aUrQsU5QOjHraY7Q1fOWvD
6X/p9fjGiYn1l8XTjdZAH+Zi2bB7+zrO5/7Eq6hEIuwFrHV1TfZrXJLzrQAyZXzw
nKu+yqim7pEvlnhTxVFP1dvv7ZW9FP1jpHmB22gO57mGsBpd/wawdzMCG2t189GZ
nLMhNeRc1Stb4jwFf8GOy1bw6d2YHq7E3bEYjl2vrslZW+VRGRJupxCDN8iLAY4h
UEAW0dAkJUvFHPiScteF/YiubG+I9WEsy6JuMfDNPkL3hz0fPjVW4Fw0ekuIIweY
QJchT16X/Gj+0Xe5OZ6WMHhxEFk6D9mOEKbNce6AyCl71CrxA3fqZjU/LIJFCQWL
p1KtSmSSktQpvblThHJh7rJ6c1CfxpMib8HUMdW1RalgAKte0m3PSIZCfCZa+DVK
g/ci0xN3g2pXoJxC0mYjH+a5KuW74oHCOTgIQGPr522/WVKnnciWCGTpqf0p2Emh
Lb4n9OTcZx5IFzDIAp9RuCJSA9JNdMGF2yXzDd6W49CjtergolMpJpKcsxnHh1Yc
j1KBjnUB3sheWrV4h/bYt6VRgkhc6dobf9aLuCa0usPG41rT63VuvMbRS1IJ+OAT
KTfdOlo4SS741lMkMiRT/k1R3UoFkzuZSiASdpf81IBRxfLHP36hx1CRXTg8iwkO
7+tJSJa/IA4F7RRUV9xAFrIdYqGYLhAIUwhh5TGmenU9CkxKsdGUYcndaiBhfyvM
7nBipz6qC6uyqdiRF26I6OUWFusNQuNQUKDHOTo8jWaIqaTAU8y37cN0MjZ/XBXZ
2tlbR2ejN4dveZ+c6ATLYRgDzlhfNWjtwoAFLWVca7HT3a75mxRTZPrOAesdAqGx
mD4SYm/0peu7klRimw0baNlDpmMUFP7POFcxYxScRpTOmoDPgI6aJzPJuPTE6g5w
X3zvw2xvXZd8MqVQRjei7A0CnPzu5gi1+r8YZQv1ZXHLwlPPHA7dQtF/pM2ElieG
n6Gtqp33nkap13fvcpDPjabELrcbQD3EeXytSWxHNRZ35FSJ6TQCxT04HFTxxfUY
9zlVpZgHdI14oCLJIZVkxXj47lhWJBVaKkWrk9k343B7t7p1Z1H8/d4Chi3jx+eX
kn0xvrqBadnBx7OystBCLY+lLwgkkaRb/vYuS6iZJwhu6Ljpw+R2BxkFjM/Ujaew
aUoY9dDhB0SG0ZaKztHBZr1agPZyHPn9v9+ouM9OP59mG3lClCJxCheSplGsa9OD
yEsPYFFdQegqdP6LRM1AuRO8kJJRiwu7qLNJYPeFqM8hyQ4fODPnF8cDhzBpXQkg
IVmZgrwTjLPeRdt3HFkQ9bPA3sHF/mJenAN9ouRqOruW5myWwaJjA5SNRjJCoMbG
dKIiPrL/o5GnkRJYfcS/DuqI1lgeerEx9JEnlk0cAum23YtU/dSEffee3ITj1FR/
L3IX58wh0O697KCy1SjBhDcd+J/WWN3dR1D6g3rqZUwJ/0CVv/2fFxXu8Ovqlfj4
S1Tsd3e4skggCLF3BzXFrRwlkXjiphEXX6OSRlcREJFl28ddQVNMz6DaeQvggCW1
6WGYr/pPMS2npxH7qO5v2EtXD8Kd90rmg0g1fQc4/yjQmT9u2Y0SEkqVI+vBoruB
LrTal/6QtYteygIWeGXLR32/ohUVlk6BBc97TVVrmpC+E9ZIYl04C5HRz8sDW3a5
OK7+M04GFMcU78nIo6+G3L0OFmkJCudRxOfzTY9zPJ9VBfAgr7+mbIqLbuZW5orC
3ClhhDxBDzIHB78RrvBP2HnDs3pUAxlfB/1rb2MgF8TwcB5BUiLxOWeKxd30pdnX
Wu4IoLtbWnEBEn8XMh53EmcVz97qnX3W0XWJZGZcidqXRLevBHn1tCe0B2QvccNg
4rAQnrx0hYyhs71Oh0LnaLX5LiI3Q+Zim9OpVN4s0NIA12w0qEoXYt1dVnWFa5w1
x0+oO8CRu1QAmvU1zx/AYfnzh6YVOcCSx40bpslU0FVbWc+Qqujjp4YdnKTU4GCh
UdjMq55iTUS4B1AoSCu5MfkRzyTDZreXM42KdYnvsnbN3bClGaniMaS+oV8B1LRl
BzMswtwuHKJ8AxwHFEFaXU/Q+nAz06MH/zhRmFt2kZg2NMO1drwX2ULtTlb+d9pA
DpCO3PHE13KlzCQ2XzJjOgpvbQqcVTlYkzRExu5icHZXMCMlX4beTJp2gC+iEGiu
v6jMrEQHOltzh+JiJ1GLQe1BOlw67T6a3N3Vdz2mTAllk4nZ4Y41L1uHydjL3iuf
nmhIII84AJ3qm35ReV7/kgLltjOmUFRj/Kv0+wP33jNyq8EmSPfDwqMA/eCkgvvj
VQdvBXxRkz/Gf41yEGl6PAj4Ms9sWLCCPfVNNK8UvYUOuH6IyoLce0/R3TsWZqzg
5d2kULnKJwQ2z+yZe2ULIcLMZmDu5+BoE2ARRJOyH4LZ1wYYyL9T2JnTKZEj7KFB
SN1jwvF5FFiQEOhKLWVYPunnYGwUXPxdcZY50XawtEJgy6ZdB7XZi0LH4XJEIHso
NKlTcVt4HKYSlnJjWSBuxqeyWQ2Ab2/AxHXwifeOYqnLlMdJov/YWd4a/B45Yx7x
AsrGtRYtRhjAFWITBuj3H4is7GdW74D99ffQ9oJx12L7GzpwC41h9raGO+YAWkxe
+WPhOXy5YLJK4ehtpBQvNcJdJugOQIVP2AS+owF30ewvG3NoO8zNKrDDsliLWIB4
1gOtm4InYSq3dhbNGwktxRGjUZuG6a8hIoy3dBKMGYDWoisSyom3+E4HgPZhLOLT
GYgtzV/Il66GH2q1+A68UsFFNLAuhVm0TyC/9mLcfwNpq+m1iNK1/b7F6eDPM6mA
5oBTVsZyIMOxgL/y+86qHCTJjHVIG8ooF1dxu7KDpOhJbccPPkDekBrWN3CwOL5x
r6rC+5+MzhKafLPgk+ssS88yhZnh+U3iGmcWgY4jnCqYkL5dpXBlWCnDU5+j5SH8
/M7nrO4XWOUBHzKvmv8XPklWYfCa60GcJLOJjUZc/Qeoye4vMglDjl9phS/4/lRC
SxW1ikrbWbwdk6zqZUvlg9YssaFoh/PI/HGMNU8J+9jy21O4TF3Y7TmCB9ZxeQ1B
1jYHEgOfcDNOXbt3weJ7wgswtkolOPsjAVXB85dUrwiROMkrBUrKE5Eor7Ybak7m
CkR5aSKxBee2ycA3W1RZtN9S9HgJWYvub2m5h5NC62KpLjwmVjv3ila0cmVIzR6l
0W7jh2zOc2Dda4QH8NQ6LlcRZiXiw9fSWEPYy+tDrP6/nCFGkXANQxIdaq0f40Qm
QvGZ+YLa8tUZmongQgTcpwfIX8BxQNcitnmAuRggGjXufHy0IDmJoL3qacmL1NH1
Z1BvYcj1xPgsEqJTJcBdcVzCCNBI4d9nnxfakimKDHpVhOZebdC12FUE9+x4K2uk
doPu/tO5X4vMLwpk9ViV3+Tnukhc1twS456/TDVWFttaBWRct0o0wyHESZug7qxp
mHa1E74ihMbbQf5rfeEpVU2AC8Drmf4y9TmSADDa3CEa9v/rTHiFocte0Jelicc2
c5RXVSkb+EIPbD3O6RUFU+7vEgWJoMSYuTeQQqQfm6B/w6M0Yzgjgyozf6wo1mJQ
ovZMQU58oTCTuUtltTCBgAIXmifMtLvt3OMLjsJSZZPIr5ppxtU5feQa6+qK+wOS
iAcF21YDqY6l6ZtsnjGFydjxsicnd1otEvRU8ckUJbM1f4zdt1VMyfS98JG/CdeO
pb8d8cIUPCKc/afx8CLhzI0KgSHAoonJlHHeoxMb6Fs+6eSN32EcLtcw6/mziIUR
DETpih5f1qYfLHr5CscQjv8VkZJq5BG2ZNxxm2kKbPP2LEqLwFgPaRYMoQW80/Ha
Eklqexzz7EJ5I6KieWpbxjYrSuHdX28mD4i0hhvn1QAVNgV5BsaXL2vB92TdOjUV
PWhGzHa38cvx0J5tlKIil9aYqTXZ02gCCapCsyv/RkKoA/o6Sm3wgSUBWeWbCWgE
eeaW1Jpt0R191dTw41/xnIc9yxWyxIHRCA/fnUBfwgDa0qy7cADPGjBkjSwEVE05
K/ozFI0yuSLQ0WaGvTvL9vfflYF2gSG9GK1d+td910KZe2zgY/TDm9MBcq3dBiF7
sanxXSGi7Q9Flz7Xaw89MaWtVD/acXod5CELDJvEedIadcvlkFVk0alBN/M1107p
w2bUO+MlpfUWFY/pX+C1+sqMnxuY4ZcPNxjn5NRX/0hhL4yn+GpWyLTU/A0v6kSV
L67UjDjox9GGH4EUToyjs+z/bBVMCqYqZAjQBa1Td7iAwPIS6aedp16ku5vm1O8/
f+NLdSXJYCPQoEAcuu6Pga7vFuImlbN0vTKj10S5q6cYRrZwhB0sVw5LCibuyNa6
6GplQ2Xl0xfQlIBNUSugsga19nR1P3zExJoXCOzGvA+uhzBZgf976by8yYELF/YL
7x7jifIZ8rDtmkAPm19lRbyBW3WiW0hA6WxPBlsiRQKxxfgBlWM5i6/y2BmvR4DJ
BrWStX0oHUVAPTYe4DmhV7Qm+nPYRQ91KcaXy2NFESsCsuz23EgxOV4ibhlg0QEL
wVjaiqtOofpMxc8Xe499Az8+Fpgvl0dMfWP/iBddAp4lzLTHYQjR582oA2bowTlm
2X3LppyLt4KnqQmEJJrLePeCfL8DU5MvKsgZ8QawBQ09NIci4mhEGt1ALr4DbBGT
H6Y7rzA9k+ec0FC0YsXxctUirTi3j8brKxXkIbUUgeE1c/24CuXMGIJV1aA3xG0i
SiXWlaPkPblOrH7jjRi8DXju9En3sUROAoCAxaKou/5WZ4E9bt5bwYu9Zl+6Oo4p
BulCwueDDWCFEmzPFJGEqhzKY9S+l+WjgSDe4BXmC10I7Xrc8QXMVNRsHN2INU2+
BMZQsKCUCCFTXhF6QQedv0hKCjhwux5kw1sylBAminN8k+BjzzvmunDtVm9B3MRa
e8OuBJYpLQdBKwOH1kEsP0T3YKNtOGQQvX5CW+yoWWz4FGyFy+4+gGSgLtVpPt49
DxLK5mqtO07cUi1mzJpMs9q7y/7giezD6JUmUchC2TcweY+h+/PuW/tnDARw7SvJ
QiJ/0wbSFrgY7MD2MWSJ/uGZRMbXdUcPoPyeMliibN2Og+xS7flI11ic8oZ3tjfq
JrwsaDliwjkUH6yXHaRqMnkh/mpj0mxrHemnH4acMXIAVHL+y4eSlr6iaykcb+OR
WhhlRNJxeA+ozM/NGkW8bSWlm1uHvKQbZ56LMxmnw2Fjm569QBIRd9L52m0rd/nL
EuD2KF2BQMLAPawEERpqsz01er+uA+ZpTczVr2S+7EGcxs+/GamQJ9zCuTKukPQj
S8WBOa2+OLJnpL/MV8WWSo+DPd9k823Ivdlq8pfkqRXn/Px9pUYNJg1qygorWjcK
NmIPZq+7C2PaUHnA1mpokC/7fYEXV18m5VqAAkupbjU7MY7bwBay8nW3jIe+g4f3
4bK6BPGkpQkBUf8yUSfR/ukXfgQeocIWIld1hBL9HG67h/YJDlDVhZ+UskFBS9kx
SyiMxxfSu7SygCqU4WDrdJxPHIN7Msa6htjN2gBlV0A1TPR3vAz/oELGbkcZ2ISM
0ebD9Rh/moRTHDOl/Vl4roKj9CCNqcFPu4EnIf+PsYiOgMBuBP5WByRki/VVfh3e
Jw2gc6epviy+mfZzv2iK0m50jH5JwDOCq/ZWeA2RWsx/+Kq1Ifd8JOKwvvm9v0Mi
v1gX8twXVh226YyCop6eiA7AFgBD8V5wiJQDx9cW6aJvBlO32CMZ44Dc7Ge3t+/H
hlvQ4Q7RtsBhWOzvvswzcSgwx9UL1XvE8ntQta9e3j3ObCiFuRZLpgXWTpL9paol
J3wmPVy1mFUyhMIYuwVDC97caMXyAGMGxJlyvNRLWQUXEcR+lcExqV1PfQ1KLu/7
hCPBQISs7nrG2Z1hGVemBKdvOZPXxZTgLPzCGgXsL4Qn7LFDoW27hYeZXA6zlemI
q4BN1MVzvy0FEtYCbR7VqVpFkgzg0XI5ESHp1WCLCQT7PTGHX9v0p7PH/5HvfrLp
xnAiHCtz1m1mo02cpX1FPLC7T2rHKYnuJWepcx05vXmzk5d89QaojygPDZUdX2ud
T1hVGpftH7+ar/dWF4tnojt01KM8P4vA7VVO2MJSO2m20JUzBwEtSqS7wUuBpJJe
UG6jTb27xnpCOXn8u1jcXmHLjbfTJMjRERED0ut2OwxOHXbQqeCQRf3k8B5AqQIQ
nYxFi1ZBz/0RrCujI7m8OknnBYLWMtHlOIi8A6l1C3LG3yftrjhWNOnDHLycVN6u
HBmg6+MBuEzLnHo8uH91uREBsvwXFe3M8qx5rCJCe/861W3QVOyGmt6HqEpFcgar
7fb4DMH9wSD/7oX3C8KTKl88yOCbI109IXwz/lmypn4s3ruTxIMptNCLV/mNXJ79
JnhTuSMmtIVvwj3qqQ/7lHKexn3qIcmG7IQUkuQwFhZJdBVZrR4843WgMfhAYHoA
Nw6f4DX/qS2eQRMkjTrKduaGqw2h0xa3WtSWru2g5Ik1uDcWoN43P/cr80CK0Pdw
ju3NdU5e4qa2KaNFN0WSoKb7Ls0OYsHh93q7j79J7S2RJItrawUOfWDWSyBgHrnh
/SNTCpFhLNgc+pMUwmzXQmBRr+7YXp2jBrsM0Coj51VYGDM3uEfagzkAAMB4Z7OH
6v6qzjWrpXeLhE5hjwNJ2/XaHXZC1+2bfxhfVmuc6wNfgNq58UoJGtBrO5fpgrnC
qB7GtXOEp8p3INA+6UMl3JgOp8QFsWmhT9JZSQRIYClgRRSUANQU3JqilRnzeQLz
V80pp7xhKVjvWRHQmpszHI9H9GkUeNl1psiZkb75PzO9Eyj2hgi1KwYEFetdcImk
itc6G49GoMZgmSg0JEzTqk48LtkVmgq3doFBNvG90tBhTwao/L1V6daAK7ntSnij
+ywj/kHJy3Ypbfjj3Gqy4a6KKdrWe/cDIRkoZzEFgqJTevKIq13WIVytyBLqN8fV
aUKxV+dyWsbUzidDNEdGDQN7T44f6Fu2rz7/WeD28X500AQF4QOaiLBhgqfUjnEw
MEpfj4+Iy4VHvt3ZW1iTN7Q77qPRP1+T+NAISACe8k1VPCzE+hjNuWZrxqeDCLOf
naFnHbqwSyvlxcaqAiW4XHbUmJnVX7iTtsABsvSq/Eksk7kPX2FPOEdzqhjpwI8A
s0KzEi7g0hfYOwXzCZFlwSBwzrWgN1MqnpHZ7AI0m40OaRKYUJFIZdvtl4iwRhTD
ylIMdLF1yPpvJB3TBaH7nnJTG4PjixNvqVOBu0YJBn3mUboMD2X5LgIxga3avQFk
c7uBIszZu5uQpax22HkZzMKPIx17mWaWeVyKg95O5OQqMmIJ7Fm2W0rAQNUUhHye
CABtHAnjh3PC9sWj7GCW6wYonoPI8WIBHMTEdt+pCPhH8gito7+kPzCynzbMjE+M
lxpqqGaKKEo9+0Ht4YFZGirUa2SVWMlfVdOIl1gKh2IsA8mP9ZSKH3av05CVUuXZ
eLFI8Hhw42YLTPlhWltXnfytswBorYXs4Xu4oJlMwRv6dRFe9mR3/vdNSGT4QLRu
HZTtFt+1Co0xrPNPD78XyKue83ed/FvsHFlm9uWX4xg0BDa1zKIqL1ov0PLdw2dO
C83FLlQGVsNG5N/eAF/TTmwvTJP5ZzSajCr3HEt0o+S+o90vtUGu1zyblBmTF6mr
6Im7STZpI6quXVTRPPPE/wCuQCisnq5qb+LqLe+qRJ1g7kWo98kjtvTonG/kjsby
PIH2658llCeMPkT9+NTrmyJzuNfLeYcuVHEAbtw7U5cUCc2K1wA1zJ+i80nf+8Qv
xJSsWUhxlYWJ9jUbmSMvcXUzZP1gg/1JfUVoP/3BobeoyRq8zdDfoD3RvRWKNnUw
FJ7yaG83fghe1himwNTmL5cafbnL7BHHpJDppNWFi08P6bgVLUNPDleYALHbG0uS
cMaKNs7m0shOZ/Uwx4/008WSyI0gHGYZezaDC3cgSy48fjOwi5OuvLJOmvlcjVl7
A9nZ/u6fCcSxMCJSXu9zwsor5xHIfflkK8/GpfpTvm1hIVoPpC3kyq2eCi4YytMd
UcxHGgLFyhtgLLEGUIxlb0u8ktQwhu032w5LS/xdSD+rWc9hHXCg2S4CksLw5P2A
38emfGe79OX9J1GT2+o4PWopvkoVV6oeSK+o5wrIaKnQgpX26Q5Kp6ThwjAXWOw2
bx0Hrv0oQ5xyLai8LBoiLz+OeV6OctZ2sM6+n+G6dlHjyVyZ/3O3tykXCCocu/bu
ujOotknAW1NBcMhUiLM+Kb1/I+RqsaxppF3fSTjexyaOs+3mPKjKfRiJTYSUihQF
Zl68f3Y/rg9r57yI4EpqoYFr6hLHrsc1HGwCru4WlOsB42du9edPCMOIi7sYGFqr
Y7SMW1d2jsTT5+5iPLeJz9mGkfjhAb5nFyhYZXQNCnnlTMt1fTSej4dO2yWSfJ45
qTqOmvFyusIHFQT8ql+2uYd9X0MrcpGc0ian04Sj18KFOrRZvBvbkZsBaXljhPfN
Krh5pMHIEGbbvk14VhzPRgBwK3O5yQhS6wgvMFerY/KDoRz/0nuuNtWuUb9gwqDU
SfO/NQzyc/u9FejOF1ytxcVu7tryyoSjqSWGEMveiM8i8F0kbIyXv/oJaTFUd5xc
ljF7ecaN8O5w45TDCJ8aavys2qlt7pkcOfhwGMJXoN1M6hFWgQzVfS7TS1s7WQel
vli1rs5IO6blb6xBCHZMzzmU4VZpvhvGuErMOvcZAOIebRtmEPzG+aGx2lk99Xax
1dRaK+JNicDiiOMDUZ7J2/NNQVPNy4Ts3OEcRXg7+Kb0mGsjCRvTWyCL384330bs
NAS/4kF94rRza5fc2LpO26UFbG31gTsEisKZCcmymLYzasBsizHgrvQwHVgIkxTY
Gm3MvfijCIe3CVqn3DDjY4LQkwkx9Cd15zL8vqWODBYBNc8e7CS+QAz211NLev+F
RBjJ0+lx+TgaZxaTxXUXpX1xMbNaVbqzyF20DGrSwvjAx31EpsucpQbIGWPlPxR5
Fev0vVIZcuF5o47VSKLD4KlATBN4pM45OLCIUh2rFKz3X/wMKOM+RskDMJXRo1rY
uY6s4W64ss1SYr35JlSC54Wj/oaFiLrBPRD5XfOB7o7rT2jC2F5fstaCjYoVsobn
ONOMaw4rGYzDWMU0J87HzVtX2WDRXzNdNs4hDyKXjNYOGEKus4dVUUo8QLOJ4kGd
Bvhz+CrQ0dADcGLdlIUeGnXJvz3qonKY7fl89A8gJ7N20SmOmWmkYSZmeUe3DOWN
GJdpX5Qu/AfSMLQvugoLi93mlZXSN2YxkKqAnK944LuQhz5ndfIeBgol4/kpc8Er
8XrAb5HYUS4CefAYVHq9V7ldMUeQ6DgGvlgh889uddGJYt59G+JGByEZ6RjsUDQ2
MMUut51Tz74o+bnDINsKf9TE6L4fHkR5MQRDtPdwFkEAe/1xi0pooU6MiarRzf8s
rtMJwlhz6r+qK0r5ZF5Irr4rFnV+UIrwAu88cCb3DlyEE0lrlnkXmPBrAoH7Bbwm
jtDclOVAkVWQaCVKLng2ymF8uIIthA6vDte9RR/GTCwqJZGbw2gTUuCK6Ba0I+bG
ur6LZJAbL4lyhqDB7qfNGqpLcUOGaoLG4zLJateKxjbOCmpCtq0Hgn34PMqaRWvn
EH6A+7ZyOeKEQRccAycrAOn1O5hlVnSoM8JYvcSa8YgoVbH2KQ1S5O36WW0DZPpX
DiT58eMS4XfsldaUliKlIEjelfkzdxQQTuXlhbkxTJZzLlsZ0AkLBBXrzMHdcOqp
OCQ6amnAlb8J7A5GWM/9rrAp/RZCJnANDGAg4Q+SQe07VqjYvQNI01Rj3XGVxuX3
rC30KXYx9oBfiwvKXkDCoImcr0wnrEuhAX/iHkCgo3i9qHz+LUaUOtod1MqC372d
ukRzCBs8WO6TIxPNFIBnp236Beqt0qxX/YT7FTqUIS98c9kYaSNj7i7bww73VljV
wX5eoa/zEWzt66rGKZzu8FOQks5tWumzVz60MmuyxZyy2NgcvqHXca/XVWY+lGFg
DR3w1cKVoQjDcwqmwpFxPCnX1QmoH50y9ww3UIPC4G/HOudQiHQqcq3LgMKl779A
T5Lmn2galLqR9C0mKJLHA8Np6+Sqpo2G8g9H/+6J9sI6WkVxfX9TBXWDt5Vjhzqk
AbbOpjRmj3HAaOjMG7O5snk0gAJuxCCO3yMLt9LyXGfGCAUJTfa/MllZ5O+lp1Bi
pK/3xplIB6rJyJC5cAoSd/3soMF1XpZKBZcYvXQXDC5+Cw0adGZnJqv2XQCU1UHO
4/BgQgqRtUbb7YPY5lvTt+XX9/slK8Z0lBo7B8oYT8M7GY/qikKqDq4lvnZOJy0b
s1rksav/e422pU71G7rg1Mb08I8XwxdRUzkkdLk33IY7UOgGU45LwbZ8f5vJXHG4
JbBD4p+BjZvAIOgBcVhIUMZGpGB90HBQreiemmIF65BAJRTucaDGGneOUW8FKEuk
Zz7nA2o5Ai4xM+fRzQM6H58WVuha1sk+or3GMwUpUkubo8Cat/3AKsKgqyez9QbG
K2If64w6KnbNeAYRvBlN9mNDDf54NEBzWJCPVX6Y2Js4eu3MCVQ6h7y3j/NblG72
x4xZ3k3USJJtFaxm7dREvOmaB/Cg5kaUdHHZVQMiao8n9TENoOQj4XyDnI4/C4zi
glCZ4U3qRR1ZxqMA0VWGufG2gVh9oKRkkNL6NDiF9J8XHCJwytlm4u5EkawOttEC
LfOscVvighZ88tOHefCntPrH/VeCFpIpuVcYR6JeQMeas2FUyPDMXCseB7V1p5YA
zR24x5nsJVQ9nMKHJdcOiVBlLUmNbDCW9AVBu/bCyav5iaVejbxsarYTAxI0DK1O
UqqfAAWUiygQcVQmMOj3Q9lc8wp6bcTWG9bp3wT6W3HWF7nKii5V/5kNITkYrYiJ
NmKP/SaUsYPdPVpPTewY7M45OsUvUgJBdNOE4fqRLDmQq0laBU0Pa1/nB2vsQxs/
xtkIal6RzpXIMx7V3L4tBX7L85FJ+i7HS7x0YuSJmdYZmnWDA2fEcnjR3xmP+7Yp
adrGva5P6qrcS9XgwX9PnPr9nUjUwM71ui1otDOnIHFpO28bVwcYx9AHVH/2FpBh
SMdcE7Qhpa8X7R0LcdNqJZ4tzKexttClQ5Iw62x8hocXVx3wPSCjSyZWShFEGATK
mUKO1SlFS7yuhTUQOsXHT4GeDLAnY+zkK7gRblrH6ce335g9NCUQsrp33z+4ch/8
YCj4fO2SKXp1HF3jxNhc4VwHy+U32pkKvc14Sa8ncpVoMBDwo7PmcEfuqeaFb+Vy
kiGhpFSv8rXkODiNVMvaR+ViZeMxgagWpXEV4iYkvn1vQRdV7oer0+0XgNNiHrji
/D2rKwqG9NvaQNQ5h/59S89umKPcuMymG5jyQtfu0f43a83fdSC+oYeme9NzdVW2
jmmfR3ZxIdVLkCPV2tMCF4LWRn7kxngRAdLJq3nNnBnqPe5zV8BK9wOUrMvor+zI
/ETVCgRUI6pnGPMYnEbNclbS66VMAmtsSCbTRR2dRXRBLZwyj+5x3a3Kx9kGeDOk
0I+1YXF9KrJJHHFwcWvSCU0migdEsIUlql5OzSyvp8v1pByq4vNs+b+vLVYgTRBz
GRVLtLokTxztbGT4B0n4sy1nhBumw4WjJkHxWS55nIIjfUOD1LMckovyat+8N5Qu
SY1wSyi8BgLdONxqm56po+xfGsCk8qrmGirq9ab8gS1ordFzhX7at5cqSstIZ1tR
tGWVEQxGEgJ13n2VoClkOPJuCj2iWA2YTf7+mBRXA95F8nQtHJnONYaE/KlbYy2E
xk+Qx7zXf7LurdhC/QBMfX32OJag6MsDuLM13d8t/LE2yQEmrHtcm9R2EltEvdTA
QmPBVZNop08nrldtm6mCBdybuQzQPPj9BNI2d8MqEu8G19mGbTTxqcvYatPF/h3G
ERLefJ4Mv8gQI3lfI8RBZVzevWzYNZjgn2bbPMlv1bfx/AuazU6V+JkBLoVH78xV
Fun5sYrJeaNvEcZwR/VXwWiWjFj+IczfB0lEMrMTibQ0iooIOLoVb4u8s/5lSIoD
+PJs4bDTTqn+y2vt//l4g3Mf++/EQOtaLRFApEIGRU9ZlNGaNXTGqfiEuCvZOgB+
3A1BGrYLz/5xfLF2TZcYD5/6j/r4y09HjDLq6c5g2proao2HqJg6ccZ+tbDZ2vje
A86C6fX0a1sl9koKMDkYHVpZ2XrigvrvfiUn2xPk2QBs4Z9HrIms/yUIS9AiuNaI
Jitio7uh4mp4tDlY0HFAoa0f7SEx14qnwBKGZypf0h/kk4T+9hpxZf/rNIh/Yz7S
ASHzm4ScCoY+9JD+TyAbC/Hkms8vU6k00LwwRb3nRwtgBIO36JFbX4KLOdUnG4ma
XuN2BD6jcWBfOL41mb8VJKbh0R83PvEln5Puk5sncAJ3xV4ShiDHLHK2WzIdaqpw
VUFCU2QLagiT2sS9ygLvmU8io4WPFWEO60JtZ9NWa81e8vWwkI1PCcvCjycyPSG7
yYtZ61Ej0XLl6cXsNP2HThz97g+s8Hw1hGAZs+RacdYwinr+ov/1LOkU5NhIVO9i
l29GTvWkuhjf6oBs4Qu3GsdZc+TtkNrgY1XE39Ev8gdb+pS0HrmD6E9wQblo4PuL
IjLXiVP6PMLKgNnIhphocGu+32xxaT8JbZnISIM0ywVKCjL4ELLSq0K/A6F9dY4D
i2SxJ4rrEPh9evTb6NDNPIiVSmoR47+mUn9Obv10Q1tY/03vWOQ2CsMiDDWDxRUT
ak/QV6UAC5NlvrX3d5eBbQIupxQUV63T1AvcHWhtv2snqO4cRE3cdRDOvrTBVMq9
jVb1Nm7cSsbCOv/wQncFRMAIlm4wEvHTXQ646KU+nMTJMI0cSi1KEpPvgJSgTQhH
6QnpGii5pSrKoNx3WingUdhlnqYxE88gg7zOIiuWOoOyALDFIlW9+M/FLcVvrO7n
3FdudqztRqaiY2jUb6YJJEbK6FUvksjbpQY/b9eWZbf/0nDhkLWy1Nz0AF0lZY+D
xYE6gGvnzYPh1IlthEFPgqGuAbIX4z6CLOl7XaWZx7gDVIEGREMpN9u8qmZZdIqZ
LnGpaEb2s9ggDEvrG/BSgA2dG0TINo4ean2mMpM9UhvoFWT0vQkk73FfMh6bOt/U
SDmvdua0DzB0lZGOVuZCbRfUlfjniUIQAY/LksKfcGLaVFUdX0qgAgJrk0qqPsKN
44+tOMN74ysI4Rab04Zz4WsNV/5LY0Vl33r//6/P/XijAALJvw0KD2T6p53WIor0
JcP9oZiSHiC64cCq6DQ0zYlTP/S2k8wkg+kJfoSvts6lizFe8b7LvExxpXm/j2qq
20Q68z7bqvwWDLPwV1n8HmDfJsonFnJAIx9bBAeRmslRHVmamoz8siMbv+gjKJtW
fRviBLRtCHPPCr2ZMLrmKvduceOIoPqIackZdHibKkKbQ50kfeFRrUJuUEQSz09g
eEQ0GQe/kHsg9+I8j9X1iBPYpBQHduV4podHa47rWUvbOIEoy9UGfCiOfzs09IaV
8fil48qr8aUeEO7X4EBJZ5p0AtcX62bLj511PGhlN+Qi2KFnmOTVJzZHtBJypAyp
dxjh10W7HI2CEn0zNddMOlM5wqOX5Y2/A5BxApSLSqCMH+zp5LsG+7aDrzm0r4Uh
fIA2ysTo6DuQUnjc7ie84xU24yB/iGdsTI0otfuMa9nM4OPg93I2dl9QECE7o46J
GMXG43xSfBFORJztijA1AROHI8nZFextJlfSzjQp/mbOsFKsgC9LY6BJKzaWzB5/
Jhs8iVG0joKRBWVvmq6EsDW5ODg+CgSKSu/xWGYWyCnqdgOozNOPP5zA12x5rGYU
lAJLAAD76h6qeJ/jfrE5Psw2qxtgHsSDDp9/I57rCVdtZaf0yVrcrjT7z5Y9xUC1
abz+YT1/qFocPzX7uUtGWDrM/REjI1KubC6ocuTbvdoAWH2a2G1lz+1jfPx4VvSS
FuPpPQVzRQOi+LFg4ZdrEldlTKl9As3emlcbD0bqtLfI1fyLMEMMZTRcFM7cvBXA
XMNgCHpEvj3rdRcINkgu8Un3Nn26YM/jZ5urVrmeA0XH3PrilYcK+K1KWkV/JF0J
thG4LEm7ZPqWMP4DHaCfpzji2o6E4sEI3TEZPQotCk7AqK/qFwW7K+auQ5XmcDkx
A/fpeNm7sGScNZ7JKIg5CZZ/NlmncCy8N0xdB7VhYdw/rUn80Qerlo9L/oLPOWJ5
BPQu+iHKNQQu4n9KAB0D13qUCI63MlIvGI8AJn/vr3LBg7pkyUOZuM7GUlfNwW+0
VzygXpRM0CA707uw3YXZGKPNa523o5FtL8+IVIIEO1PfgiRZ3fCPZqnLaR6HY/pw
mKtJX9yUKfjqvl+PrL9OQVQyO4Tqw9XNRGffiMLQKqWnVQx3VRoiFiEKqIlmG1gC
7LVAz8ZfR2HgevtkniSX5SBECJ4qI3JoYkNNASGhKT7SdozRTh2UcUAf2jO4tylg
IIEXVHJptdogJYqb0cBGs5AsVBFhIWsW3OCs5lbKRQD/cYmB9XJrHx6HuyVAdP81
0tj/rY8F2sy+rEGXpXKFrpqZU+mwoRr67nS8/YnGK0s9ipnD/+e7i0vthruIP0cY
IBCTda27fLjqsPSOah+cjp2fiZ8rwSaaeTQaLzdO8UJD4TrZkH6PnXJJhRSp8NE1
AN150uDKlGrdzVKtXD+JkI/BZYUErf3/hOdeG81Fvz4T6x2hbcuf9uAziNk7Fn0S
O0llgs+4YZB/EXb9ZDKQ+JArNjLJ1z2NmtaM3Ga5xf/B605Lc5LIN2Ot7fY4XsTK
U3y+54wGjfsw/JQXKEOuJYwNReHJK+zNdXyoaZcIbUSk9SRUofcR/5OHL1h5NUXY
tXtcwJIvzrruJD0ncVXjzzxCIAykEtWLnDYLNBCGgdsp5t/LOKmIgm/JTWlH+HFh
kS3UDRWtJ2+wspQs4gLGJD2yxG1F5zTGpzJFZf06MtTD5Yu/gNB2UiQftZKOkUIA
sfmZv5UycK6nP0uVqpaPXke/QC8InfXwMnNWjXCDCQs1KUKz2/uvpHS5svn2JrBY
GDamc5mqYqqhEPoarWWz/FQDSGAp00Xnj3SwEGgTNDxyPhkkG2Y13lio0iL38tdG
o7NBFfESb4LSAv5fJxhrg6p7lAI7GlUJJqBj6iwjUbRfmzCPSrcI6BEtRKDhUYue
IPgGb2oniWz1C0jJGp9zG+ZmytGrYCVJIuEHFljIVT4jcqBZYX6vJ5vMw6DQ9zON
840WYbk/QdOoeAAflkyp8o9LgI0xs5kHP2nykeFKG9txMgA7yjmaRXMuxZkTGecn
sTbNLEDX/0+kXQctaYFYYVjO2HLr88V6XGnUUe+dojfxfMtYefelcgEQID3jxV08
9UaQzWPIAuysiGsRMnT+mrfXtsIbXxT5NcEbyFQJGFojBka8SU5EN67PKEngOdUo
nqk9z2rvXA9JpFKQnOohcfDrCWOfqiAoOM+ch/X3zlRnV5Mv9+J45/sPbsk0/G6V
burjQtSqSGFmrVet5x6knW+Ahy6iLY6dGuSMZIfSO8EqZh3/4OIWCwR7DKZ6skdm
/wJ2upGI3uNYTH5qcz+wMnrAciWwP9qe5XYWhOXx3bXwPG3Xk3KY+VB50yTIzCn4
h0J93V1JhukYhY9soOj38lnJlGJkejlVCCPSlsZl+f1ZvFIyhM80YLyAexoljEg9
64EuKv7wb9KYZz57EaRDFRlmjzj5OjmNpdiO5RfQdkYq4pzUG6LSsK6PY9Nn3HIM
vN8HFLDEBg3NVilF2eGarpih9/XqyPDkgX8YhbWCBPTuMLko3/nOuBr+N7AiY/ED
oan9bHUOjadBofOZW1oD9uHSFOOjSU4Aa4W+WbTUxyvIQMHUITjYtXxB3Kn9dZ+p
gWo+pTHTVSB32G/l0dJmR93bbDrpa7jyzdCtwVw3O+rNHPBoPVcoQ2tbwWafbjHC
FA8pJlawdinOb55u4iTWxoNW0MkioTg1vcGJfvPAJT+Tz0sBU8OfXVBNSXYR1APN
0S7jTRjTDyOEk1Z5G8J4bdlz7tfp6s5VWUUENhBniDqzNq9wLiIIqX4CvIcyjAVe
bEzNyJcbgm+Jhid1UzuSB1GCH1onorbBHrw9j5t5BpyX7G2zUAJRBrzW4Zub2MEK
LSL7z3Y+MMRFW8Z9S0lg4F+LlZhcu3dIdolqV8UFNtZJEH91C9Secvk8yCe6Fu9O
9PByfwIiQwNbxB/SeCD1eC1DTaLsGLfU+8UEg5y19he22fA5Sq6vtTvYQwWEPOEL
gmvqyc7vObIKZ5VH/RC2JYHGuuSMf5TZ/re7tS4sbU2KQ1aydLN2SqwM/vvjlhpX
/2vp3VLg3Fjb1Janc1KjNwgMIYnCWwN1HpBCvLKqGQdsClkPBuO2ocMniXpZJkVm
6mYGnxhkVBEJTBGPUIvAtaK4UKPVznJxriiCYc0izSuhZvVLFCzdvGMgCQLfCtat
b+nxxBla9qIsEjX9J/znAR9LV5OrHdU+hdJJSbBXmO5bWC0HNVC35o7kftKo/5Lc
ZgfY8pqQD07F5mzGYHi0VWLobvqGCSSdd3J6J/IRpuRWGpCycPpHcThz6s+66iDh
b5OfNpCVw6dGIs5xM/ES8m7WuN9JVPNPDJIh13NS9iOmgSQJTNor+5rRSoB+Iac1
n0jvWo9MobPEz1JrZbB8cydWx6JybYTe4tFyPZtIo8xXwxL0CN80GTnTnmhbF1eR
e4S4IwTNaWIt52xeXwvkOgkzAiSc98kIDXBuQKgOwskKyJoyxM2vQsmrGmMecU7U
RpN9e5/DJWTMw2nrBUfFERiS6xUOBCPUQBepTDI9pj7Dpsg00lfRAjGbbThglTor
dAe+r0wLf6TQEiHXezkcN+TGR9CbTYishApj4BnZIkDD6WJ0VI48cqHTKVLhNzRf
PPexP+2e3lsYw0bE8pIMIM0xdoQrexPMKJMMfVfbfxtwvAtr5YWJUEK95R55D3vq
4r2QK8zx5tcqTQkP8Ct7gBJY/V6HnDBGbcZhjnzCLmLHaJVx5t+eWxOCL9HcZFZd
xRO2CzsU5rM4hUho3T8iHK6v9Hble/FL4KXU91qmpxjR38q8gLDKSmXIzEANTfcK
pIW2J9iRhhM1O0elKG9oWHu9axGJd3FYo6ZewZeq6ATAE/xIw11o7x9M4lfsFHw8
7mDeKl8/1jau7VZbK5yfB/yCroLeOG5EI5SiVLN9+9qgEX7o8N1wEgc+Esbo+rh8
XT4PtpIngZOExErIIhi0OKSuHMxxeQDpRnk6f/c4aT/MaEjpvFEmY/9edgVQlSvC
r+aOoKeopklSNOiK7CgCK9rqTtqEDnxZz5K7uC8dmfP84uCMZOk9tf+cTLicmPX0
hfp3jCS4GHiLfkEuCQyMp979qs4F3MEJGUcR4JpJQZp+ghOXDasNoife0LE9mbpQ
tcaNq0j130FO02/9h2EvK+tnSBUJpDhF+AXt/j5riE+9nI6c2jHLtfN3/yBv89fr
+qrQYk8zZ3jNiWrwiiD16fNM+EWsUR7nsc8LvmWWJV01ePuJgg3RELlncykgIGRO
2v7s6/lPlA1SCWq1h3qZDFfLNd272tHy0QXpFohDOT/5hE0AqmFSNLuntqh2UpjJ
JKgWx+vJWFeTJd3oRzRdZwdDh2/OWgWzxp28+iI6Rbk3CyaZRc6rHYR+GRIkbx9b
LLYeGzXkRYrXGOGyoiz/QEdKas+szw91jv3nWRhZpsUyy6/II884boi3PD0bAWFh
R8Z5JA4wlZleMWBXnA1R0nQB7Tm/S5qSnGcFL+S7Mwr4jIOfLxkgb/+FgAfVfiVN
MVmV8fIX3g57Np3xKsS3ZcqBryp0dArT67ox/4yz0v6vndj1y/5ZNYPCz8yr3FVx
Pqfi5QpHSUuuadut/F4e8CUckMSkmUt5sdlxMp0eJYnjWpA5WP0QO/WgKr1dFbN4
K3EgN9NLBJdS1l8rlJuxpmNSCBvMy67OlyAccHVTmPwu+SH9Gi5xi/BiXRbGFs78
rw9xrGB8mMvDBMioEnqLui9JY3lfdN3LYpK5QsOWSCzptUD9deaQUopRWA1mqPXp
Sem8yO30LyHs01G89tiHkTrLCOWo8yrC91W61KAE3bgOE6U5sG743d+WptgIjsp7
qFIS9iYU8inTcQ7CDdpztEZskRsbn2NAyGgpZB0EV36sfwgzPHbyY2+xXUCGn7Na
Tt4jlfH5cZiwmU1MheuFKqvlk4eGAqREVp9YAlIJcJqqdsMJ7z0BZb8fqCj9NQVt
jmyWSESnLLha+DY7ghcYTjLVRtL09O1vjGC+I+CS9pS/VH8oDqJbQKz/V6wq6Wqn
HKz2kAsLxhwNnsXRcMLdrXKuSd1X8XkcB2voM3lcq5THWP6AEaMsmb1cbf+BU2L/
oFXyx5f8j+iPxHlJ2InlE2KA2fvNv3x12ukKSQjWrXB0BSqorTUnFHIFN1hA+rPX
eDqtKcqEzm7JQ/3WdSf8RAxkzl80zs9Q4E0pzK2uvXsfq7Z+6PjnpWTrzHK3Wy8u
HRQ/xxJrLkqyXEJ3C+z1O/EvI/GWhQAfk54EOsV1uduD+ziJaTyEGo1ZgveFUHZD
zEx0+hpUd+loAjrMbnCRrW3DIsAZ2cET56oqxbC8AlD+IyG6NsDmsPPZyNWkxIBB
xv4aWCYoqoKt4Q5E5ep6aG9SBPWy3BUKWJbN/ZGekT9auRbjKwIdRCn2cXyWRE/S
n6eb2ftQDvZ4LZ539sgRPlJHHrgGLwWAI6PY9ekExotNfvXMP0uZgDNtWNuOZVs4
1E6iYswhBqpwkmjUvWyd43l5Vg/4bYxkpqNr6S0cdl7yFZ6if7xOkmJFWHbofgIR
r5Qgi8kMKI9pKms/71IrjlzLNjVVTNJDuitZKHD00tkalHvph1psF8ROQ+s4AKLV
GVYC/4b84aoBBsBsovnSTVb+wB0+ZdNqlYytlCSA9SmRlxOnJ8GlghsmprAgjVfO
VSUm9E8hox9nv5Z+3Dowk2kxLJFIhGBn81ehlRPzaQvAT343l7yIyuCxaPGHde/y
Ps/ATFyLOyYyjHOfzFEHUa0emtKKA43zuepYqKnknaauxzabfT18KxsEZbz8IyJj
QTW5W8oWP7pLDkq0frPr57Q0F4j8+ArJuqhUwgAR3S2jKEqNKpb6BWHjbqwc2gvG
gw/kbD9/Z70sYFJEdnrGTibdRVzljW8rZQOVsYb+RZATcuUbnbQ6BiKFFkKlAGeI
jKHaguNKrj5OOoapA/pOw5GCDSWO+Kp/KRG0CMBbqSMb+AKlji0J4q3nCp8DWQRp
Q9EaTcryLN/zGXPaxNZLfjIi/hUdMUyEuQB1z2zEgupKoBJ9O2HRePoYIDBP+KBV
OQ0X9nc/QBYKfRImUvrhbMVeot7UN6NXHRl97VczlS2ZYMiHNSS43rEqI7It6D5y
qYy/io33skbNiphNn2zZNhT0BWxqLXSOxt2OQPusuGG0Twwpo7h9Yxfi5MZvissM
+Sz0y/PX0Q+1ONLI1Cghwc9Jipl9sha8FeatzxKIP4imKRLXGeWS+lFloHoXH6Vn
M6kDtX0VvItKK3bmwg19F+X8aqO1vjuZAOJntyAW6WdyEFoh+nmYQ8nXcSYP+Mpd
foDzYrQ2Rpc5M5NzxnMUx2nillebXhQRy7r2+8eI+ezGVA36ZdBa8z+vODTFflBB
KmYOFM2NK2J4na/v09uIKH30UIm+q2/S0yy7MznNdYif434AgZRfjfwNXXShpGS5
Tr8GX8Uiy7sabFO09i/MtTctpCT8OqIerKpcQ2FFGYnGRTxQmWJyCZR0jIkFG+uW
4QIFEblzWrRxsCWo9n4za6B8LHIQkpQHnv4uscJpA6D2uZ8wL6WaKwo6F6FtMi9Y
nQjyBRseO1UaGr04QuU68zSk4KYBwAnrNghxPkxpVo5iosRw3T+EK8GZZNHNKc86
3ZhTwvt65mPN/6y9n4n9geRFyRmcWsHbBO+sr6IPC7GRQ2PCd/6Nlr+4mlRfnl+z
byBe4JyaGBWPXfgeOqdKHCwywPvFXj05rPWrQXrf904fO4ZekfWgLolhz4yL5pt/
AqAqLRCoPNr89zHB9bX2WzojtAk+oJ/ahhM6WcQY68EbLyOivygF1vLUO8JtKwbO
QYoTB2+r1e5UQJIRth5IDzlH1rLAYNBUcFUfpfWGFgrjrwwlmtOaKJl1Q8E2gmZ5
jQ5VsC2tRkB6hsZyWJDsOtu0emv0upTUXObGfBUFRgAnj0fqdhdc3oQRaRoSEb2P
oL0Hmi83Gn7dvD5/ScCE02xWYDVm++YOZFbiIK4AoL1zTtaj1ti9n0NBYYXBhVta
/ywTzNQJ5K7vJQ6vh+OE4aQlUDUSfKNAGEFhpdAcpPgsg7kVZd+6WvpFdJai9Mgf
qWbAe8SB+g4C3SN7NKXtF/wdwo3Gtv4Q0qZMQdmfC+dkfiwQjybDmKotMNanXP0z
d4jgcULzxfqiGeyKBh14qqv9nip+o4RmIhFc+a77+fBg2/gCibAAPupUya4jVM6t
ptIRGARoOOMvOhyQkECcDnPoQJvY+7E2PJFUPSx4g73PZhWi+BLb7c/XHDZJvumK
/ytl+53z3hJGgZ2Bn6RpiP7ad08ZjijrPQfqs/YLx3Ao3RGIPNGBjTJlqg7EK84/
7yF7GdKrjZc5dfOPraPRMo2VLWwdW+y0uTJGzo6kxGupeBZwFj5dGrOcHv5zSCWk
mpIJk7w/Zf5yD3B8Fp/Wa1vUkTTfU7nuM8swhJTVOPCa6nlk9Bw43faxlPQ5eNWH
+kywdwh0krP4RK3hWzZGDWwt1CE9/Iww0itxBWErzO11F3gRgrTHWUCJeQVgwBh5
Ys5qkTQvshxQ5nyhJSFmvcrm8VJu8/45IvmZ42jSwWrZNFKsb1sg4+iW2LQYMrq4
Ww9LHeiLryhTo3J2/l4+pUbeK2stZmKu1FEHBU4SXClrwRq54aUzSDF+wTN+OpEt
R8KlBIsNn5D+w+ZP0ha5pFqwijAnqq7I8zO7dv1ostkFOJbY9C0HfIcQPsgttMWn
e9Lyt67uh2TuXTpO0O/AYaolTge+98R0nwi/Kdu9d5lYjh89ZT8XhCUx3tFavBN3
9HqmbT5D95HSoExAWjbhnDvndJgKGdHLNO6+ZF3oPBsn40MtOPtfPmaoSkLORJeN
e7eCErlTf3/ExW5qyH6Aim3ywt8Z1HTXvqz4y9xKoqsMD61TzoiSneutcNZN53K2
tkQiV2eYtHScs/c5NKINmlWD3O3pv0EABW3Xff/1BRWVoj9EKONBJtbwg1A1pd4z
JEdXWqsOgo6UNAwKItidNdj026hFx9XCgbGIDH9rhyW1OauozEZxxPB/1jq18ilr
cdV7sX2EsAELxEZsw7z2zHPNbQAmJ59bxHdhPIgtkpXlS7nr2BuZ2J6FksQLnqWQ
ZMW4Mg4OBlWmbtPZempBucQdFdBf7tonhvALiiyQkupvt2x1SKUdJP6uNsZlL3lm
cAYuE1eSGCSTgZAJWD4G2Up1v6w/GMtznHzlt2zwA3u40tAuPqpEZmt8cZdswcHd
pcz1bo1eWn6GEY9e6hknwjglAfsURY07Gmn796i/pG1946zWsoFEHmWwAfgl4FBA
BZ0+FhkFaRSbPQFSTfqM5IVabl28I4wTFBzsoJn7EcO1riBpaDsQiEQNhnRQ6lhI
BH7KWssNtpjSlR6H3998X8Ju4O0Y/pFg776SH304XvJC31FM9LQZAooGF7o2V0/0
PBCaue9j/xKb213YLVq5NmpBviws/I+EUdE8iv7tY4WhlfdDC6afWQGz9JC6nBAN
juApyylLWVWdaxRiJIvhwiB9oQGyElU+fSC5DoNs9V8P0ZSVtkB78AcDOBK9ETCZ
QzDOyadvFdf91uph1v2B9knc6cNUPCQ2QPn26bcLFG45wcF3W91avx5J3PomBOmR
cV94Jpih1fGXGkuGUt6aIUav//buo/ql4igbgkOF18/y+26MSOJOonVu/djO70Rx
cWZ33bGNxpyubmI1TBX6CD8uQE+AziGreLcw4H7tbHHTkM7RnAgxSgsMaBEpW3dl
5R0eSAHTHZLC2+nzh4FkIPqvP5WdeJn4yCr0y64h397WNvHSYG8EdOdtoc9VfAF2
1XIhD+A3TLvXLkkoNDM8icH4wzAUnN+mWVKxSMKnbCyQwFQtAK/oRIlco4av80WM
q1+VwGdeqhLrFBrTzFnRd+XR9Q9Ex9ya79FsUBMia99m1jdLXgAZMxwXi/idrkIk
vWGHb4J3wCX0SWBWAZivN/X745UZlWC95i5OaiSZYcBy0rMU621CXdZTmZoHbYWx
o73osZf4V4tAfhr4VWFu21bowLyYnQowIQCQ671SwI3mVesyK06utMP3vCBJpuOZ
dHy2KWEQLDW5UgxPZ0f4fny5pbiQoG8bLb/gkox9clIo2sr7IfvFNAaBL+YdMo6m
SGhFq34EeMZ8YjzVvJ9QOc0jbIG7uRfZlrfHGQElHm79FjzQMbEnK/NCNg1xEIty
wV1a6ZlOQYCt5d1vrl+19Em7/nQsP+KQMS+bUFkUaAQCnpRM0MGh7oSLq+ueWygR
2mOTPguwbl+lT35/F2jsJ6nOcGD1jMQtsF7leZzXu0Lw9jf5dy0HYMwb/7ZTEjnK
spfD7HnWzcKEuxT02qsJUKi5HItM2u/ldyCtqO9DlOMg3RUNLK7oSF38/XMqZLR5
lhPWps3TbFEhHWyD4Zt/obm+stel3W5sSN/nlB9J+LCwggmucAykPREcVfAmw8t8
cPjdXCvlbL71ufteMMZ0SOPSAVOOwwoHknllm6MpHnPz1SEZHhLK/7176emLuBN4
hITf3rkJ8nq2WAYX1sgFh/L6phR1ieCdve79RDG1EM6DZ1/9Bii1Q4S/4oBKF3ru
OQbJLXfU9tcrZlqyMmscj87UMKdi+Mc890VakAP00ugywoDKD0Y1RIgkMupetUj3
OGjYDVNao4YamYrUawqbfeUEYeVYiH8tRU4r73IQ7PkwajhjChgbz+zB/0aLO19H
FNLlzCiMx114TXQ3Gn32f6nsMenCW67eiu8UYEFk/TBxjb+Okx4+2+0uZr9qpi9s
HoyauDhXhsIpZpyNhbS1+nVc1Nsh8Y/9f2n1+eR3RWDQ5419K1sM/zRjHiWh7Z/I
Lnf6P1kG7TlC2fCaOCt1Eo+P196VFAw1kEITJFFqlxu8LL7wt6luh0KezYT707RH
KmE70QjrVcxTiR4pCB/BTyxhxbFQplPrZjw4S9C7IRM8QKoYWqhGTWVT7+7Nw00/
KR0jLOIerD0CbzCBjrMiSGj0qP9Bi54a19O9aba7mLMbHJudHxLK36j/ff7myQUR
8Nz8ijZ8f2CSLKKvd5e8zFNwP+EB0/bUOwjph9y4C5wleztgWQq0Kq8KPExt0t6d
CSYTbrFsN02vvlh73BPSGeozveKiBREzjEaPTLSn/4lbheXFvug9iWYSn1biqkkp
2PDksvLfF4KcQadyPWWkBZ+/0qhusuG6XFPnorf9To2Q53Q5x/VyPMwOEbs/A5uY
OSsKbMRooSOT5BciLBmZnDcOJ0aRerqIj2Cpajn+7OfVBNtuEuUVMg1RRx3EsoUj
sicpZnpfsxbc9ZcnR6C2KfTBELJedMF7j9cLY3fgZGftqSxw/RQWBBbDiUz8/SqM
6kIvhgQWrAJ4MmuwTcUhtQK+Zc+XGcwkQgLhkX2kH1bZPJRk7zzBkLg57JlcpQLM
oO6RASC00bpNbSOdIbpcIr5dLZeEdHOIjr3x9e9O6JlUwfIm6H6AhGGL+SfaK5d5
sUBI0xna9U6c4TDAV6bHhC7GYxsEvVnkAiIZGj5Zc6vTXszNUgKlmSwjmnVEIu1L
30tKbEE0QFGtIbzy1l0/+LFFaAebdtFqNgURDjNwQKbqfsB46r98ACfrrpaxbl7h
zu+Vp48HEBjlKBWxxBR8hXD7Cpp2S/N5JEN6TRzk7YOVBZ6jEzClzc2MWK+pF51W
RMd5UQ2NbSPBNoA2LiXUOuGkPT8N4s5vO/c6t+RY9tvTynMIdUfZ8LB9puT48ZKR
iWIagoSLgOyj9Lk7rQPuSGKuERjOR8OscFtaTBsp83MOdY83/VcskujvSt+G+AoP
XtQcNcrCis/vTewR63MKhe2WcMAZuHh1WJK0w6zEhKidMqfip2pyAR+7ttXtI7dO
JfG3RuYgyMb+4BWoZVaUsyIDtampVJ1nLxPOUr7EdfLIZPOtHo7r/KwnFi8R+d9Y
xMG1u/is7uP5OJWj/Erp1zDMB9HlyepjaA+I9cym2i3yjNlScVoZkYs3mlYluWKS
RdF3i7Ls1gVcRwalUPR+MFztitR/jMumdnyyXirJMU9njL+UJFfV6I0kIAqzN92O
rvKCZ9m9uQjppx2r7LHBk7c0USy2yrx6obX7sMZp5ulAOWC55xORZcfm7BJ1RmZH
MZYofmDLRyqmQEiDWZByYfn3+gZMrXK3INd6JyodCEwvdnucao/6YtkwX2TBKsSw
APOLHx/GyhthK4plN0JJMMZrR80aPWe5MrhyXWKgGdyfQz2Yw2Gb1ElFdFQasfU0
GkRckDM9N8RiXAyPKvrb1VPaB2ov/1rX4hWoapvy7rzSIV270/YQolBUwijiH13D
zOItGLszZen61R2TZ97F6VZ0YI/JUTX0Dw4x/eKvLOJds04ahtszRslmgR84iCEW
ryXxFddHtQKbuV62d2jDUdaX9cTs2THqx96YMr9jPs+Px0A7D4HhYaZEUrA0NQnP
CZt6A1Px3CM6WPUN0nlQiZguAxJBlm0APTdpgmTAGbYxugfKkIJm6Fn6wvwMoYZL
PF50oF9VkU271mJmYw81ztwmDgEtnTmfNUDU/MB+I7LLcG9P2tqqQ6oRbhql0MHA
T0pc7EXwgy2Eb16wkD20595YXzkCMR/0f76qZmwciUf6SZ57ajdv47TlyQndLnaj
FHf6rTXvcMs1GmwTJf89mExTgTVjrgq1CLtNg429XVxvHR2VBiA7JFcbc8bETwNJ
OiPSTs37RT7VVp+7NTLASDRa+FAB0JdX6jT85hMoHQGciWoxPeX+rW7F3i3r8yb6
mCGCMK6VP1rSp+h5s8vU+HZL9crvjeXEi4ldsMwkcJoh/apR8ASp+osz1AaldfCn
y30Ky4F3Q61qBtI+It1j974X8qD1zLWVXrqwcMLbM/oJzeVYaiM3sCxQRBODHtFo
datmR+pDiD2H4wqtSLFxhL7Pyvxwx/uNCOvY2h9Y0Soy6pbRnn8QqeCxyTwbCJh9
9frd5vjTZooRTSVfi/N/yC5+ZxRIDE5zbnw2PIA05ESErVVf7Ghht2tNcobmdyhI
OUapBojUfXwzM9KMNxC8Ln8k44DpUsQVwpxiqbLLnduGPLBvC7Z9nrvJLPUQnQoJ
WF1kUjwqeyL9i7K9VWAk+xAEHs0sYakJdp/v37arIh9dTSCxJlfGW59GSD3cVbMg
/DoiFPNEKQuGlJSn/YLoEftwM8PwbzRscOe75kkMfhO993Nn2E8LyS564V9hTXwT
sbR3B0aDpbTO0/4EQg2hPRM7BJrAxQu1IOeuSJV807/vaP5Upu+6RkjRjUWZJTmu
cMBr5TliIiGjLYXd3UTCgyfmdSA0GUhgdPBvqiwKVnxNgTIYJVM7TL5iSebEIT3Q
oVkT/9tY90/RqPFiK/eRPhJZ+ymbcX5Ydw6l4nAw5lZiwkSgrI2ojQXxz/lZzH1k
6iLggpT7LL+iLP4L6SjyxQTFMY2JuiJcIUAzlYnf/TWOF7qEyIJequYn3w+FWd/g
PpKQTafmX3Y7YzYZ/RWbrXMjPWXoN+TMsbNxetnBecklhR/sv2W161q+ZWIMDzLw
jMEMa6iFe2O22i0pvnkeAk2Nd9ILEO4ca60SDiXwj4bcjNvhIi5MfzI7NVIY/kg9
aO2uJj3cbGm8hTnHktFaQUfB/V0bA3fZnaLnSuCTzDEm+35IXoJEyHmVwt78cnWK
Hw7ix0EEqzwBhGjiub6ZFfFUnhHj/WgDDzp5PB0Q7tKAw7pQg27RLNdUWrL7MbpC
sB+6pdizfj+8PWQYEiq+J+mu9+ivEO3fqLAS81vHSd1hTS0vOuN2nEpGBUOC1Xa1
jNONH+PvaZiT3tLAVEcWKOziM6qw0nwdKuLNdcU1GQqlNkr/WYYSV9MHAjLXhmE0
90uPwcnWOM92K0Jo/m6ztfyD4t9ekubXRk5XIfZtFVY89gwNlppJYGTyFhFn2kpQ
P4qMh3U1oqWoLuwIGAMUIuDW3YTTQSn/OOWbeIVfHGsBxdEU2glyqXVa4dJR2RyT
VhzMX0OQOB6wzQy5EHKSHNndPoTjhM5KlMrlKA3FKKOmdk/udFPpfWXMS1+PlWHB
uSJaEzu6GavqllgDSK5WthXtgLc0LEwBZkuGFvj1xma3Ml36MKpxJTQ/kL+6IquY
RCGe3Wy+WrtCpEQY/iLeM/e/6i/8C5jTU24VTXD1D1qaROMn0hQRnHQSNIsjGQoH
ZqyeV2iZU6iXQIgYlB8njOw+O/V+cdRE7qUZhPYSbv4fzIlGAdQ092M3kObVh2lL
GSw2spT9OdCRYjGIgT7d/bARPRl+i6PzdhNC3UKyjrBWRxVD7Lqe0qV4W0s6B3l4
2p1okBrYfX3S4BFGHnqMmDpVDlg4s14L6IwqQRrkekX08HNFQk8A2RvKzcHzSqUI
etb4CjdsGmOtxfyAYAnmwxUKB/K9M4bvzoCr3gfPgmb18ey/sPFG0yuRITlnmOAT
qDbrMRJglGKGGKVIPWXZgxYVT+4UFXzfocvwb3MU+K5HTU4DVfU/VUhgp+Dzmt1e
rgDDt4Ar2oGVlHb5DpJhEtS4Djp5Gsqq5oiEkTswGUfi0hOf0wvLA+HfSRSReY6D
9vXwUQK19BMBOkjmLFlHma7buZKXoanNBgk/hWBdJQ9dWIzHaRN7klzh77QZ4j3H
adImtephJ6mLlyuO9Pn7V3Y3skK411lfx3kswq7W7SkTedJwQNcbmsFhIwKDA4zb
PtP8oiE+dOP3etzM4EP9inO4ygj53nRya8rLunuuJZjJfAHESRftNbuRszpgOXUv
EtUAaLRxXH4FcH9N/KD1fBMXO/siojJsstUkq/5pXkSwbOs4SxMbFVotbV/91aHT
ZXd6swLB5yy9O61y/OGdG0qnIH+tEQFA7P5DCFBuA2VldlWFa9+AxLrQt1nztin0
SMQafUf6noSabYlqHuwQ7/yTssD0/F3Hfn6h6IWlOYYr0MSiJLWF8lYY+3bcFBlh
gin1sVbad6uJ2DyCuiBI/6s7h40NN3zUC9eH5Ha06MNMSB6GJGzVKUXN3GMK90+s
oPNsvrAAH71EebJ0t72uGoh75wnM1btIpuIT7tOvL2LGsw1J6z80dPhxw7uiX4HS
Nkeg3yOxyX2VjMwVq38zQPMKVzUMLszgTGEI5WGHaKl7NQvN0An7itxi0dhFNR6o
YtnrpAaw/ou0VytaOCv/YRBv0QnKruJrlVImPsXwqZhwwzFcaBLc8VW8w/wpGrs0
4sqtuwnH4X50igyuvQdJ72NmppK00dJvtMV1j+aVNvTAIb0MEmgYS7FE+Oe5vbDH
ye7aaxr5j5FH7XT37QN6AX0nc0k9DOLTn6YjLz23sWSDOhaHHHA7At6xoFOaHIAq
U/sIDTMuwWrgsxtQ2IA1IeJh/eN50mYWpa6URLS1kFmume6tZn43cB7CvSR+CfIW
NILehStigrLidcLz1UUJqih4iZqEHiNJgRfLVDAv1htTWVZ9jP8+7HGHgwmAkUCB
xdlybO59NvkRCIica82z0aXjHW1bMfrbB0PJiylKxzT9H46t6SzFYHtnQ3/0bjAt
dIR6inoPSRGSe4fj6DYo0BwhO4Y21jj6d8N/T5di1QAr2KYusER1yH2DH7cHRMGh
1C34Zbo3d8u6lHGR9Ce5myeJy8OSK7ed0AW2e+FdiNjxfg9LXDK1db8CneXsr/yl
xCsoe6ROxvJ77Lk0eXbYPaZds+i0gSBAFXbEmji3cQY0PHwzK/HjjrpGAczQT3dV
cl+tvIyEawIAn6Rr5B8rEfMdgxyyEnFUfHxs2TZ16QdxjfwT+nCPqxSaohTADXWg
E3Xr2nCDcb+Kzpvza6JTi88PilTP39OQZTORkyxTYUVtGvry2k23ScUFhbKxVx4H
Y3KkODB1peUO8+1ydQ62+m/pHgeeMECCf832kU5kMqIGcgbKi3UHsy1aFV5VYS7y
6KvqEEHF/wlDNThKMaGUjrZWj4n36skEz6IAxVNPNcuguPdIFcxRBzd8Vcu/GU2P
+1S9Z9CdKaQBk49PXUHmYBKYOjamxXYU7plptlEkM3IxkvA2RrpGRPOHEFEdtIr6
Mfn9U8BcTm7ABPEboQi7UqoQSpRkZUVEVdUEFTstIoxdiWxHAbMZYA1fYOawL1vK
HrFOoU5Lt3FL8fHqeZnlbwfVLipU/ipuWOwsi86SZo6ol4RzryMi/jNLbkaVEfix
4zemtqtt+0RFq/7dagXkyfBa/Kyfu7SKi2Yiat/6xetTe/0WG1+LU+vxtF2WR1XK
abb58Ci958bbXQ/eAEtb034mVZGtPanIclzaWNElsk+VOPqOVDTHeVvte8+Prv4L
fIau3Nwao6M/3fvd7+8MxkDyj9pi6SszVZmi46kAmbqwrZpL6ZgYgwIXgytl3vlf
OI5lofidcvzh8pvYoGWcgCnpDD7qgmD2FxKoAlOkUALIVR6q662C5nl0cn+iphoj
FiQ/lCQ9Wi5dJen1xT+OdeOS6rCjhWuVsEVCrILCgZ/HfeZ3WXW+GxZzPj1oaXvZ
pgx/WaPM5tooBtyuwsvjj8H/0BH53joeTLooMc9vGH/lREteexSD97aO8FSpteJ5
EeONiQjYN7s9VjVMeI1JUN62OgCNTHlu3fwWfR6bOTtf5E0/IsVYgWjahDW+jZuX
IweM8kwkUwn1T70S1CFD6PIoJ2TZ9ppX/uRAKLCQSJep9URZRoW8BblVj4O/tu5C
cmpj7w8knp5EApaW+TKvIn/oo4QiXIXHzOeG3xh5jNEBq8OHTxBO3jdeocE4Qj3O
QnoUL1y9c24o2iZ0cwvALaxrgzTiZ+2Le1WDXPNDvFRSgFGklrRnDeb81GGem0sN
m6E5hvea4CXNR2GpsB3YU6lQE5TKLryZbTpPFLh9ZJXgp2jjfmkB3A80BkICV8aL
D4AEcPhzeDD/pQiMhQhq7A0mdbmyKocFfjZjUaz2BRkgUzLQAieHa4LG2qQdYMgE
ALPB0R88gqv2EsaXg72kijoQ3PA6sJmoV/8SKgj5vtA8TecoTZa4CCIpbK4GFpJl
DQcBgbRGMGNmkcgIZ7GxH7unSC0ooazZojMqELck4AzbpP+uggOf75joZvrh89OZ
mYhI0JGsXLhjEJxTFMYJfHruyhRJDlFzp4D/1nATiw5XjiLsm5arOOO1TB1h1JSV
qQbSKSeFF+Lc5JUWs/jr5+rDfAHnCFR+6FjrL2BWf2+y3u+gr3lfKav5tKWreyR6
29nFPlZ9aUOQFJth+I4xvxJMWusAgHwZNmczFueyX1eLdnaX4+FF0E/fzBEoudCp
HyMVCE5nQS9MdmsNlszEN/xMHUI58DOEF2hvjYiLHs3GaGlVU9SG7Z8CeXa6wugH
vXUJvcLmrfzrhPGKyHxZbqdiuStwvl+7kdWjBMjaSOCB5lSKkJ7OM7H6jEI2uoi6
wXUpBQHpsIocsx6/Nrowc7wgJ/UhD95w9o9hcGDXtRoiyFD+V+fksjtigwaCxn9E
o98CU7WdQOY/Gu9JOz+UZSGg4wZj+u8REoWaPscjYVce4BS1Wo+5Yvb9/CfQVAln
ZHucDObq2zCCLwQI9Mcap67TN0ha2DlQJHMz8A/or8yYWwssWMXt6Bc2OrcTCmDD
sVipFdTdj4DHU5X/FViRx+m4edG/PVGYnfC1fERFS5YQLKdPlzNdasaxzrKrGOEG
+5v4qsyYoKpbSFD1/q/REGsk69BlElxtU5futiYjC1TwPthQGwezY1lUHu8pHqlD
i+yQauhdPfzzJMunf4yodraNhrWnEa8FpakRADab0va3Iqs/uw2bNhl/yrV3YUib
Ru/1+0BBskItHAOcq6vjBt5a4LCPAOe+anYoeaoulJ9UbXalD5g9lSa5VRXkTBf4
1VbJB75IfWbmusVTTyktRN7JDUK6w+8jX3AkogNBEhGWkWMqylnUh+4bCyKhYO1c
Yes/n/+rbpX/c/ASa76/kIFsinJDsvkkHVSwf47Eb8zpY5AQ0CHeoyp+FmiLRB+B
TWs60JiZviC729AnopjB5vteWN0w0JJMMEg2XGHPnCPKaNmY+k2qEscgHpkEURwv
p9WjHrxvr8UwtOgrd8mNzxjS0TOB5vz4dgIvek9zmYMe1eXu2J7yZvSZRtu9w7Iu
ipTad1pTfNrGA99vF/nu+IlLgUjDLY7rN/Umi88JSpZpO7rhXgz+3e7IubisKH2q
LPVC/Ss+mVuBOFtC9c/5pK6p6dP6rJrq4dQppRHjKnfo6dolr6TWCUB82jAwlvul
1aANw6W1mQX6tbU65rWX2H0uVFVzDL4nF5alf81EEdhlKytftSbWS5qtkF6RxYv+
hyFxqSpHuLthK8BYzpOuE9i4zGOBMA63Btli39QeVPw0xlQflPgJLzjaLcMk/Fzw
Ix2ZGRXjDgIJaseyqfaD2lKXA5dAgBFqg36Lrmkf9LZlA6fpB9CPi6LnXSRfilCC
4e9bEz7gilvfy6c5CWPV9kLFtYqeVbQJCAofGO2AQScs4h9GkWZXSPXsO25Rnz6M
QAe6TRjcNsG8gQOK4UvNxgPP9/FNsvOJBRQHkSNGZX+DxXm/7XlxLOp1FTffxpwV
5vWacs85ectlRLXDf8zZ4kqAHh+ZWcBCvuuYtm1kEu/VNjOePCa33hmF2lMkFLGz
cj2FXNpLKVcQpX8GBOFOIRoh2/pU+zI8bawl6RyPSoYBLCxxACLNo5ZZ26NaLV5U
KzHa9+mAExy2vYFM+3b5hyIIWbcAdMRsOI6WdeZB8hw82dap54J1Sz4nYlD0ZVDK
9b7t+Z1AuO3fENhY7DNQ33HLZMhFOHq7Z29nKaaOFbiMLw3/ewFEkaGyG4gM9kbI
sZ50/CCmTNXe7mRB/xSA1x9Kvwj1vWmFgc3tYr/R67RAE86riNVyA77nlmqh+0v5
OtYSg2aPW0P07T14ZXCstZv9/2v3vK7MJHnyHwwC/d5mDfbmTqATwv9/sTgwSFy+
Dqv3Vm+qU29ylFPQ9dgJVsQ+i/2xXX/VmVrUxjJrsmsJ5CfIIQcv9GVK0UT9wgEA
jADCv02dMy/wckZKdXh5f+l4FG0aSGQmtXlVpERoJ1FXWL4fwecZf8W7e6QqZPrC
9nB6oSx8oMGjswp65gHWHdqg779dJ2Y171DlPzxXHsBRXLEs3mdh7A6w4vm/IlUF
i4PeQinJWe4QsWvTUlV/U00R+ls4SQZ7JWVROD5OzNXv9ls+lR0ynRk0vYux3zpq
Pf9SXn41RIVUIDHAB2zC2cvPI5YvHmiOVD49hI2+zp+bMM58tzj/QYReZCkhdf0S
edn2L1RDLXth2lMsoaKBiW+2C5UlkJtbVnr8SMqmxuiHlQqaDLS+wV4zSEmgHtqR
eGLUWFaWFUmnIGJJmQirC+N6zIR2dMIkNDA/NfivFHD+bfL+62Q/70/PGT7E1BwN
buvP9lrtyC8pIZoWXXwBWJBtr96VsBIii1yxxuCI4Rkt+ALN5SzKjYE7g75cNG+v
IRwgh3WExGEUExbwX3LzDkSZf5S7OSckJh+Ix+wtcVIBMXjZLBYv/5XDZm0Bb6z/
etfbRPEnH2MWSbi4yK8yPHikmGEqwcYK2KqQ0XvgzEV06dLofIvmnmVdyOmXiLx9
0p1OG3Fku/n9hYw48+qqhpBlb49lBw/P6clhU+JlvEu8SVxE7hWJ4DJ2JWW2f7mR
WSHekkL0kP2DfouBL0h7DCHIRJIGkIxh6kylFqTEBegZO2Kr8gyal2Xqk0E8ERKr
Q9L8fOpeiXtxRZ68Y5lGcp2taX5IKWtQk02dIN9Qg271OsLUCQe9BhhQKM0MmmB/
a8Ducb8cbzW2kh4NTnWo0qSB0gchH51H8qs/HS78my2n4P5cAHpSGpVcMYpUimPt
xmAOnBSC+hOOYm1+VEceMOJPQS26tqSEXvYDXo0Kpe5fNtYbJDmmkwiE4X6IfwfO
WzUCE1+05rU6MHH2+kyD3MRBoJUOY0jIS5t6VsTM21SxiVDWEpJALQxbSdU7oO5P
pUc430drlzo0kqzALEKu+4PVdiGRbQiUYXa+vUMmGoi5pwyqPwBJzVxXbwk1GwUd
afRWgp0QqxErMrX0zxHoNpoHynZr3QHBiGB1Z+uCGnN2Ha7DyiNIgIpPnIWe4ldN
Mt58LLEChneMVM6BDrZH3LQe8lUINDkcPadHghMQjaWjMMofopfBgH0aCwfvAln4
oEbqCJGjkpjt8EatXk51mmDA8fP7ynKBLaEpsGzBLCrd4H1xcoaZpTLJM0vF8RHI
xweysWzk5Mcg4AkQpR0v+lpuuoJmSN3OY6TVdNmBhXtg3/gyvb1gDj/mw9h2pzoF
7fNjsac23c2EPNKlocddcvofI+XJdRGtP5tB7y5T/bfNN2LfvlyOnT68glisvLuk
B2kToup9ZJAKaEWvTlozzq69YFYRqwP9bNRlYRO07tLUyIeHCFZftwhFQmsqRhRP
Pp4cOWBEyB/Dur27zeVmDcAuZqDxF7ivSUQ4IJOQJTvLm85q8XdBahQi7eooRFvW
Bn0kwd6AzkD3360Db9z4wf5Oc6/76Q3z+ntLoxxPo2Q1qHxQ5xxigXWMBdeChYK5
Sy5oX6M7YjCnBwMq1yZT2aGns9zrhwCBjbKXp8Wmz1tqVywWWAqKJ5sqP4G8IWZC
MR/6/uqzWFykp5Q5J5m00u/hXsnyJRbJCV6As8Owlc+En69Veo+fP9FwF/wIb9l0
fxQyAJO8LYt6Y+SRDsfq7DZqqAHDWCNagQ3KJX2PDwbn5jWNc6eklYZ/3+zTDEqa
KRPQZozr5Wjf5qEJnpumgJ9hFoxKh9uZaRwWOs9rIzoXo5hW0JY0el4nGIzhj28V
2Fxlnn4O2fsa7IA8suE2PetcNaBXIoIGBZc70yRaRcb0Uos65H54ljhk3e0+qoiJ
RGNSTFQppL9IpTyKI+X3HNxKHM3z7q5sdSAZvSdn+Nq9J7qQF4WGAYFy3sgLK7lo
p80MJGVFhQpcDPETUy6OWnTZmc5BNiHa2crh1Bg7ur17gKTLodfG1MRz1IjZd63K
lhgTJfBWhMPhcx6ClnyO4KLNooTU302BOR9Q4cK7CsMkjkaom9cR7LS1DfWwWIA+
K2fc3UB34HxuBK8dcQ1jsl57fVa9nkBKyzSpAule96Dz3akdJmqOE86Jvnx5VNzB
emNnCNCY0kcyr8KM+K8pgUj+zkMb/oq97SNOoIUXc2UwC7l8/gZkOBXHWgRJ307O
vT5+Q0Xf3ynFnFlJ0G0BkFpKxJ5LAZ7qq58CA0ObgE5Oy587qN9YVLEnHCeac8d7
3hJx82SlzcGDxB62vJZKbpvP4+z8sXJk/cSxxhqSdAY6Bko0rNeU9FvIMlh57CIY
0l7mtFOfRWpA7vjvt5gORnIh8a+7Qv4p/++LbXjSQvZcYZhiVOvMGmeB/EAa+yUU
6j0GsHr4FTlQwWxyi6ah4FPiNQ0PCy2DYbGkr1lCXjo8IhWNPbGZygFsaHqmXYkz
owFn7WGP3hoSPSn9lTKxsohccmnuRSaNLTbbZng+KS4HL60N2v0pFNtDAC2D1WVp
vCpfHs5jDp17go/rYlERa4hpSbx8Fb+RBBoDDfIIs0n2LQJq69MwDyTrGA/biSjk
Qyu8TcrJUMP8qE+FOROhA85fsQVoSP9b2MdB9+T7kGKOFASOyyEwJGW2ZNm/zjcJ
AkjDyncD5lac0bv+OvmiQ226dVmETdLaeLbV0KxtjHvElKXr73NVYz9exHLK6tBn
ITBN7PsM8qB311GOEupopMPERb1jnKMYpf3eUg2vuD97+FqXOcNQHxCiV216B3dh
vEhg16wO2d5nIIKv3AbmFFbGLmKhqAKvzA+CJoy6MWAnehDKWNZq5BrbKpAzezoP
nNm+hIXcesS1MVSJcdJT1nFCRXcIrXsD4/TClHnNuX+cd3dZhiXqLyMDdVS52NY6
ZVtsCZxIm3en5ujronOrf8pFOwyuMt/nHSNCLkVa/HUnLaayI/BpOIXklMtmdnae
TDgl7BM8XwVmSNOENj2yaEG3RyyC5sJ22RLLe6+BSp5Qu449gsDcbuZkUzWgt+Se
zFpl44+NpGuhWXmv+20GN4Uw1rOMnm7rqVY7Vqh95oWmsv0rIDOmNdzmh9rb4MYX
+aY0c/M3/d719lJ2zP08K159ddM2xjdJMcT6FTysFw2KseqfvbfX/Bxr/oAb7YRs
gOh+5CeBEFzEDUy/CjRKWyEhVikIP5+YEGAFNr+Hrb0jv/lTaSesejtJjXcwhruG
Aam47stEPA6ujk1QU7WdNRZbWqbTcibcUxtwLeZpEsacP8bC+lBlg6NVQSVPUTnf
XS6/QEZO7aBt4hTGQ4BVL1trDLd6glzzCbyQQrbuVpdKBkbX3Zf8NHi0PJmlNEG0
T5ywY8zMkO6W5NPSHtknf3UzPlK12bsdoadflhUMzcseAzW2vDA4tc1hkPNin5DI
Td4uOrVqIMMxO7hvXtLKZsKDeC2AS9mWq+SUwG7r8LwT4XNFYJ6UkxQnfJ1Iq2+D
PE+zIWwY8H+ULfpUUp1qGmKguDCFouTqjztx9UgxOb+QftZRrjbDgAj+jzg4GrAH
O226a7efAcEY+d9zP8QRywvkCMKRo4typmcX9iiMyk7lnWNcUwmt1vldeMDApRTf
HBZCKHWjUy6wgSCuA2glmoGAHAaUnZUe/kZNqGTEKN7IX0Hgn6LgQ4rejtClvlUf
TbFo6kBgdPHLWO2gVcMxcXiLjytEBlJVK0WYeU5N6kMgxSJmdv+lkwhbsgTnROO7
MTxuwYhp8VAZYv1Dtw/309rkalvt6QPNxe1HIj/sblux2lei7fxBWlzn6FhSbDuc
GIJNlcz0dccabCjs+L+NJ7RmC22101K/J60uS8JpIUPbmi1BJK6gYYVlCOMV1Hr7
RSlRoWwRz4P0b6RdgoUTkIerRQGo8Sth+IG9m2em6SAO9VPWCGpYcx+kNBE3g2vb
PPi+BnesUhrZvVCJUO3tJX6S+WGm4RW/iqw50Uv93DLrE3gLqxBQD07k0GtMQS6g
WdAa3uM/ESD/WOsK2FDcJLn2no2dKbukhFBZ9MWAd4gTzGwijxRPA2fdlCUvjGsj
pB0O3AAW8Y72fvLuiIXq+G+WTB7WjRVc2lK3E8NWx0fT3rpnkMI/OMKeoZlBvpBp
0l/W6c6bCgyyW2DPuTxwGgL+jCZrl8/Lrixnpi1Sv6GP897fp5+67zSpYEz+avjH
qLFXyUBuEzrMioY52xq9IsbekZ/ySqD9gojaaq/EL0hjW1esovy/mr54U3ewaB6/
ndyhBjdoSTQK+kRjOYKfiZYc3Rxw06M7Sdxd4wfewIe+tyUuymMdQ/YD4FsCAStg
lHWQKUKm3I012UQGhS6rgKmD2CaI9Q9oToxJGouhKt7DY++8W4ZQm5y+fLIOz0zT
tdzPZVADH8lt3UT8ohR+fNFc3c0KKSCs8PQPAM/v/f+Rsy5GZyaX9AlINKcW3ae7
cuwdG57Icrv5joJBYR4iFNWnIdIPla+q3VeRMB9RkBfI/OqnKb3qmyHNG68L10Du
imDmnnMKopIk4EsPntugQBYl7aH0rbYVnvB9xVeTcO+rCzYSiMwNFE6kZ9PHWH+q
0Gqp081jhMuIRcagBu22HCfPjUkVCSvKdNHhS/ag75StAOof71apRYMzLKcFQF1S
agA+LsHRA7mHMyKYEDDzvUOWta2eTzmXXp/jH/z448CR8DGrk55TN89OTAxBD86D
1RMzcJtornbgsNTlGLYu+vCDXzfPnq0CpmzHdMqkC+WrvraoJlbGblglrotzVfZS
p4nWuyHdeWZ+zVdr9L+wPiMwTIvn06hxAf3Ceb0gpC4qSHzV3uPRQzXtAlQnqdgK
hcDcsT3z+jx+JM7uOH4Tki4lmy/kTCG5L3ln8kdqaWfHBfTx28VIgPImqzBWi4f4
HuKga1T4Ll9b4gCaKqcCyk8E2AYXrLLSNcoOCDn+JBsKaqoZnxxQz7VBtscR79q2
igdwUAdQVgbGm7SvrR2Nxo0v/etDxCIu5Lgefl+++TwDrrZf9uJ4NR9Y39A7QTsB
i/s5oamPgPbDzswaDg761J7Qib+HhOTTzi8eNhC2LQVATgXn3Jz7IAlX3ox7uAMu
yhi8ONT2TaArrGTvIIbOj4mwjCFNfg+s0FD2yFKQvD8+8PoDc0cjhDFmNApFYkZr
SCZSyUQ4QfIV5focaWInOAQ3EnV/p4oi18IyA0f0PaG3yvw19qmLBheWv2hnbnD5
KGMKCstp6JxOfeDf+EeScdxV33R+7rpNQRnXTdirkzJxc9udxyXSgC7lguVg7LPX
TuvWK3s24iH52K/nmdRyxAycmqcPqaeaq0JPUzLMc8elgz9CAQViHWyVoF8EFobF
TDOVDfBoTA95/budlxMECnN3J/lFQj4QPIYcIssJe6JBmvUD00LDHu+mK4cNp3W+
2tjZHRnghH8eU7F95URO2V7FINGEVgGqLKqQZ9RuIYpIKWRfuPSH0WVidszSGT9c
TpRj7QW5F3UFdgJ9t2hniL9dAdH/7AXYr2/lyS+6FgBv/1dIefpt/8lhBmYYr+Fl
LBW+05O2UL7nBI3ysE1cxfaJNsEni0Xyr41l/Bb4EbO16IYpx5UeTNfQsJZ6GBhg
rVy25AsbODn/KepZoPhKxGx2xDnudFQdq4vlv6vMvmYeO15UaReGh6/1IlaU/E8V
Fh8zgS91mb7am4AX+RI1ZcfFtd2DV36tTbVw+fBd0HbxqpVMwCIVoaSq3gtp6giU
W10PYCu3CifhzzeqpmuOZi58MLW+4ePnTFYwTE7+Cy6VfWs7bM3E2tZSqr4gu4gj
BzCZixslQJzWUGrRST95hVkDYix+nTjAruEiNV/Hpvp3abhbwvud0ScTE+n+mP4q
WkpfCpYUWq7y2lI34cefgwFroXHPH7gvwCR7we8G1Fj3JGJmhFQwt+G9wXQEWjnX
W8Lym6XWDYNP4p1/WjBgzC/6dCc0ZkQnoaXH2Uq5rAKR33SlJWzhHdOGoE3l21mf
pgSCPvmsgNU3WPs/xYEIsSv1VNcUeW0WTT0wjiciomovlB9bU9FDEd3RY9wX+YRs
7QSApboCaSFecE+1gT/EeecypIDOOY7JK6nfwgKXN4/MwEEmcIIjMhfrgRqTRKcA
qKDOfSXgVpmXwdKWG8OzZx4rAzafu9EyIHz4ZWf16qjeOVcEpruQ3m3XfshjoJlJ
5wlEhZz5vQxVLw/GRvpHYHiWrAy+1oGcXSOamZ4a//eKbsgnup/FDCKH2EDIf8tc
CxXjeK6Kwk6Zzp0HMPQG15Mt8KHpz3SN5/tbHgVzkSbOc0RJE4MMJZKFll4fZecH
9SdlET19TxaVjG2CowgQIJ6axymVen6ArJcOtW8JpZicjpSKOuLdoGqkS4Peojvm
Q7ZijLEQt7F8Vs+KaVkWXXjemj4lGgUMAuNdkc/2u0tRHGi0PJg0Od2OO1hABRM0
hcPFAz8OcgWwtRULE3VuTaK3h04365vdHrS43+datkmg+uMu4arw2zrZ3HVG93Xw
45ia7mUm220eNQsi7INJ5xQcKeM7Gzd/j+3imSlaSyDBokpLbnGKnW2h9FoF9VPe
kpH2g5L9K4kXhqdggEav6UAwQxgeJaDNI+vNaycOJSmR+2QN/yRssZznt3I4vqMH
5ozqFW8JJ6vrPDsiEYwMqhVeI0/q6yDD1y3gc5bTr0NzDF1lpGpuGTObIoyGzP5A
HysVAHmzW9/x93/NfBxXRn68HjbFMbozDCcKwL2skQJWzfMFarh5B5pMpNfYoOA1
M5z1H/Geut+5l9qcSiWLcoV6nYvwzXEn6CAHUUwW5WIPlhQtbuBWvhbax7+7nEEh
OH8LIhiJKWO241cE53TswphuY4DjYXdZQCqelE5PxG7z6c9FpBTfwsYFvi+mTA2N
TuN6wezhf971TMZeeDHLrswOPg5lCzBKturz6iuSp/fD01KCAv0+7KJGSVlsK4OM
ZhmXLeW1n16F9NbQTTpIu6wVtShxb6GgQVBn3tEAg0nxPUKVbzIFJsFSM52vS/TO
OsE4+MhUU5BiIobYZSmHgB//r1LdL3PuirpgSS/6kbQTl6kW5DFMJlzGnG9bejhg
DShgYKGd+LuP9hQXaqgf44Nu1iFl1+V+ioz2ossbItFj/TAEB47r+W7ThWDTiEHw
5/yYx+Ecm0Sef8RK7JxS0fnz1WxaWX1LiChd4L4Y9HzoGEkIvMgLaYt3tOTbIDDu
frAo4eTn88cgX9rq1WtgfGaypXxSJNeH8sMBwbqM+B7KWJVOlijbjySsG2rIU9h2
iBkdUXPGMLjS73mVWVkVteKwvMBSES1XHzmrE5yPsg54Y0BIZ+Wlwk1iqRiOQS7J
hVA2ybYO3x9pSP8eOb3Zeo7X7tVMRugm/IUj6ycwHuBwyvPMMk+FSCUkGnj2aOaU
wdESaS6/dBfWCU6vwsKEzoX26y7z1Gn8TONfr/Oe3vnFvCS4I3JfYbFY9O0U8k2t
A0agBbkbLGXUwpudYQ47lU4UiJq0ZnueGmTZrge/6dUkV83msTzH9n50QUhvDF8w
g2P+Jsh6lx/9vzHaUcGonS6wWWbMt+BUER6FDoAfwq0RzP6Qt6DjcnpbFA3AFitD
1dOHLL5edXZ1avXDf6q2yrylj7OFqLtS/jKj/TJdKtYEJ9Oso3ze6LpvpjGCaP3J
rfMIp12ihd2WkwrwmnMlk00Ixzu8ktwgkXwPyF2PhWDaPjg12Wx9nWMc7FVIczkI
SpchyH0qW/vu/x37IsqLgKqnnZP2vvGTxbXs/or0PYGB2LGT3JxvYSA4gKvrwA7u
kUcpx192zQbu6XBeZQpcVp9e3ynDlqwk+V8Mja3Wf4RzMeuJoJv4jPI9Fv7xXWFG
qXl6Q6t9Xmm2diU4IS9VwP58LPD5w4TVdMkw0wx2hbbu+q6mscV2zcdM5CI6MY7d
JwgtyYJ5fW58U/CyBpV3TMVvRavYuBJM1bjhq0W3l97BwR0ZX9vUACBi8kmM8iwT
mOeeTa5ZPogl2OTsSI7F773oKdp+9dkrfDkZCj9a5TBUs3C4YM6FMixoNHhBP9tc
uOLlu3CL7r6RNFdi+BZJsyT8il5kbGAjEUpdViQ7oar7Fhbz0UkoFaWWUIcFd/ql
vvZRc0w5/Sgg9+FysJ+QfZuekMsLC3fBYvJ13yKTGAcCAiCewILRGd6iSJruN4wP
jjBQ/oJ2ee1/x9c2gZGiLoaM1lMhwwLz/PiuB02Ks6faKCUB2lgZZDxWWfs0Oqr9
PPT1+2ADG3DZ2e9a5S/DJSTITawghR22TdpLxKe/UXxc4ifL6H5o1ko/tpHT3Pu6
zizXEVcYg5aLtYk3RH9FTC8Csb4IrMwJCQorhsiJzU4TH8By5kmGnT8kE0aZKhaM
BO1C4ATYGAmerjwZSrQyTWEfkZWcCLFU+SV6i7TwWuyYVDnjuwcfsvdjNUyug6MY
OJ2/DOW4D12HQ60glJCRSWIxvKDjEbmRh6XKK4sTbRxeLPUsnVQzJmr+Ry7hdVoj
0tCGPw0YMHEiZET9VQXlchb0I9TGfoYDzWCrcl/cTjgoGcxE+5h6e5LrpnPExRN1
NIThQq+vU3yJ+DtprgixHrVAPpw6LlgaO2Ukl+e2ZZ56YDDNqKCUAYTI5M0EN9Bg
TI9b91AJ6thf+0wgaPRYaqRbyz8qFtRFYr5lbkH9/QasB57HxQLj8ro5N5xlOrcS
2IfuIRw3d/AXXdS3W2IdSA+IFY6WPsJcff5hT2WP50EYhsyfNrP/uEQB9MzOUPJJ
/gfVHSLX1lcXJP/UtQsZxBesCvMXtZQdrCE6IboWMCx2ISmDKV0RQjk/kH79JeLm
kOX7G2wGzJRlDtDd8mtJ+sstHV0S+WVc+LpjVDCf4gBX8rfuw/AdjMxMya9IN6Jl
LHYmAOduyjyDoONHlflMcHQNwmgbTzwsOV5Ud3JBWBs=
`pragma protect end_protected
