// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:27 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aaQ2sn9HLeVhQcwjiONXCUHXN8sOwDvw9N3fT9OnNvA2SZpYiVlVnDXDl1DQpI1n
Umbvg65jsS0TbU5d9CVwvWnwvL9RMmQb9wnJVTCj86e0WS/1QbSjj7WLpT741dGZ
G3vNbYtsOLtaBuUglib1zHPL27omjpzZnkomB5BJChk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7696)
vPD/m47Yr9xEDk5HYFzr8B/URTWY2KateJKyMc2CvA4PN6uQOymYVKivBlDAeQMr
lWLuC6D2NztoFCepGZpSA6oZYmlgEi51dVi1q2M9d5EbVaEqw0f3FkpM9u0lrJNB
WeEsI10J41mvnYOCUp5UEyCol6J5CHGU8HVo5ZgPIvBlskidKuCvr1FU8BrlNUHS
zqSgIDOiWKP5idtSpmDofGOwu8Lg9Agz03V8I2FnU9/eItJyjAIDmhK8tu86c0mb
0COeZRSg6pXS2bRE7dygcXG7ftH0yvNHmtpOX6thFstV37CAYkLwLMugYxhhVBsk
y1WOAjBmQkGUs0J6iv0BjzDwDqNgpimUgvdC8HDCxIlHr9W+XYMUsRsYwVWvFEFG
TF3RxbZgxLw3Pgz41W29MEvMR/xPatTXiahwNhqXpUzkfcRLqohL7M1NWRmx1Ujt
gghO2a2azkaMep68AbJbC+OqMYlFGtlqSaKRp3SvIdUz3dSNdb1vkyWPjeR0p5c2
NHD+UBluIq6WZ4wSoYt9NiL0mucBaskoF7z39/1sCxTeIx5MpjhMEC4iqAzVud2H
9fnwgNulaOta/bFjMjMDT2LIQHEampVyN3LpC/eDFo8mAksPW+NI28eigoEIViw+
x5VQ86aBd/x5Y/M5iwdLW4oJpjlaMqmyAHSD2pThBTeB+8tHXgtQFld2AeF7WLOe
cPYaq7TnZg0cWSVmI8UBWf7mR/CXJRxRS8EU9QlMDqZyqXuLoXreQT8QA3m9FDJP
ttgklDS0YCreaW4fcZpKhCq+zJcYu71IOk9voSCN25rXqyka3HwtO1K68CifZBES
kvBsHlsa01QadqIKUVAcuIk9E0XMrOVzz+X91V3gsKKqbc+ZBl+aKIsRsjleej/B
rFw78fBNXor6zMI4StsSds/mAsBojarlaTft8yObix/gbbq2BM/0m8UwvpZnBmXj
WgWHDpjwE41Sj9mJ+5aj37BLpcmoZfwQG9lG4OtjeXy+rcN9NgRcXG0SkGnIxvmF
i+Q4fz8U8A9eV2LRpQz72ClNoHfcNbS4Bw/bizd61eI9ewYANrNSBnQlyyRi4Z4g
MEfbqwQdBYMdebs00dktoOMtvQB9cX8brntqOgvRQLhE8ZH3SFJGhJEfw1v4cpoV
PD197z6u1ZZ+raRe3qI0cX3k4XdUd+4sSeO7KW8c1kGnQXa8yyadpneaDQy0pBhc
9abSpqkFm+Csf4fcaUjvr/e9USKsJ7AuJx4pKwo0NyjHN+RY3Y/4bmr3J/vHM700
rQaTUfqrkQVa3ZyMIDo64bp54kkdbpJOOc9uCmSKdpk92PXVwM/bfjdWcKuWxxTJ
DhbodRS+s8nx031TeQDGnsBrAYJGwAdU95vD/pEkewBAHSgY6eIKe7+2l8rYbZof
iX1qqt8wdzB+dD9Jn8Mh+DB70FQhKv+KaEpjRhILsZO2I5IKe9WQrk3x+DyjoON4
w+5wZDeD3Z7KkCPBetIqkTuBTTRLQTeTis25njDPkn0e89obq1NeylMmwUnABqLK
lpzrRLpfIkknYjrsTlJQNc1S6Ud/CNxx3A+ZwthgxsUUDwPj6rkDVwE+Cjqun9AL
hS+swIOy6jio8bdDwN8pPK+TIKJmOUK6qa5kFMAwU3GUNh/TCIYu7AfMwJTA4pSZ
FafAwIlCEk48FpEqpRhC6WF/ta5lkwaJOxShJH+cIOrmtXE9sQ++VcZZ1jtOg5+t
DEmUk1gFIzHVidcOCVJNoszgq3oRS7F5zMkLPcOiiIbmuQ5bLgl8W9a3ERaaM0jh
VbE4niJzwU+myFwkxABRDBVvWj4v5tm7m93gqJG2payuwdCUxF8DdH5PkGI+BLta
SUvl4haQKEUz6eZuC0hVrUvxA4xxrAbA4mr8oM1WDSpxClZ6ciJc496N4XY0bLJP
i1RNSIrf3ndAyS7XOAIKEFcU2L6vd5TYkEO+Wow7iwU8noWOCV9HkVm3I50hC/+7
1j7cKjmGaVgKF4Kb3XYi8fZhXLbgpLXJZRNAMV8W8bsBNm9uodgYeJlCmqKJBJ00
9Yc04avourZMKcT+ziIPUG22lBBXCMfb9p3ZPEFKtMNptzXlMhzlZUyLxLVjp56e
Zxa+g4hbD8ygrfXtiinAb8XfvKVnr8rkC1UGTMbPdAQ/zCqusZTN/7/GNRABCoGL
65nsWNen3J4C4vNASUVl5t2hhSIuEi9dkfbDvuria9adcS9WzQpO9OgQGEyBdz0a
4zdauBLzEXrYOTsrmAuWBTh5fYjpIRTAwuYVVZsj7kZCa5WeXXiyDNjPjPbY0uxw
EW87xX+qicaX7jB7Pt81a89KA+A9HottvxK15maR9DFGgtTdRY4OJ5ToHA3KIVKd
/AuxC7y7ZLP1TlBaauDaL/psem4d07Wtqnn4jLuncrzdWjXSDB0U92/cD+s8mLGm
VJMFtJ1XYz3MekSNRG/3+ag1vCXc0SmDdjXbSLPhl2zr0ORSDvKuNZLQv0hl+Y45
t4PlFPcOLod0mLwnNiTCpHUXXa9YOCOu+zLicXVvqrXQVi7YVGLeGdcwCNlCvOIj
w1OyjMba6my55WJPGptFhiD4BGPaB/S/G71sEZM8zc/hG/yOwnBvz1Yc+IJXFeSn
EgnSF3+PTe1XQGWkw3GICejbKWW1Es3ygL95Igz0Pf49t/8qY0uTt04JI9WTukVL
hb+EtK2jRM4hs9PiC12gfB5ITW6xTyFPevRttOp/YoAXKOXvr4/ch/gBGqwh2sft
eyNKaMN/XEkIqXWaEzpEgK0CABQGCRNvIV++pPaCQCv926J0M+Rqo6NkUaKy6tt/
h4pKLXcd4eleyJAP0v7P6t35N8fbhKvmjtd16rzchIz4XahMW9wQSPHG7IJqa8E1
htvVvOSBANRYfnZymaRp4zDWPLPPisuVeNCuJ8Uht2PluSFC8qrvxcK0SbBEoX6N
hiVeuhXs1GBtYNC3WtkwNQuuAaeGK4E2zyJhkjKNvcMB3I184kMo5VC0LPwppEtO
oZj2cau5lFTFVHKAZfybQ4dyUxqOJc/mopJXPMNw2UH2B0JyMWqqxblRSPH1wOxu
qGbbudctzhaDtYHA9W0vYELmiU/CgrFc9tC+UmYX5NmtaCIypGuHuI0/Fhat07NC
L170htKKTPbF9/Ckl2sIps2Ds7o4MOe9YJF88Lz9ZmKEVJINIebZAdM8b6PCZceK
8IfOAjK86P64PILfK/EDY4bQ4La5V7KmLc/kVzTx9/Lp5J/1TH6zEi1eA6Axbo+V
bnf5VJ2BjDhfCQrXi3AC0XDoqw/wACkWoyClZGa8uzvRo9plbyBKBe8rpFzitHiw
F+ijibOrU2eGOKh/7uSwL/D455rBicdpERqsBr05+rC+yFH2IKkGQkWKA5HyjbEy
j6fBL823HCuD22UmSIYugOfyiX8H/ndF13Hs5d2VdXGTYzBRmJY2rwk5vFxXgcta
JBMQuZpgKm9/0pv1NHzKck/EaYwC6g7wKV1y6g3sHxFMCxytmtf6X6syyCRkzRh+
1C5QLo3Rk6AY+NsCqnBJSeSxlCEjKSWm4dDTzY2stIVCircrp8zVnhZItQhP15Fv
oRzgOAEqeUnLELdK99TPjBDik1eDLGqGf7+2Ck5rdhKlpgEY18uu5sBDRkue7UDQ
7ail+jgiPaCQfjZOC+SAZQyKorF9gOAQwYPCu0mA0FD6Y7wNpgB8s2oUnKMcDK4y
woE6lyST/7RPGmEi5GeUmTjD2M//jOLL7xELiS6tp+zyC15Txws0FH2IpKNLyX/v
UpFqcOCyIf5YyIBL6HMtEChj30GpnjN0ljq68aw4zNZSJWQvQjfDtj89Gt5KCZsO
QAWLx03KcjBjC5s2ZOmbHHIaTK9i+7x8gjjKyyiRKFTXuOfxH3LX4VGX/9HUqwNf
+540855C3A2vItd4gb3dvSRIY3em/TQO6oyz12vaN9sqLaKZPUHV65aZB5cOBgl3
4zOuACJPXPI4cP96f3hyBH6H4VC8MLOppfRTsDQkNvm2o9uNn6vGVbe5c2dbn0KX
PZziWoSdQAs9dwmznkcp/UJpjGOHkHadQHi7qsNgtxqj6oyijFQ/dTSRLrXOE3Um
gqOaZ0CYuD8FWNI78q892qjBbGFU31te7EkA9onSmc/jTgy8N02pFLXAW5ho31a1
R0rNQVoeARO7+hWadp+ifuZyfQMqMwlK+58QSr5SlDPo2UUS6xKOjUXVuZyDj9x5
4Neh+PcAbw++0Oh+GqPwXWRxnpyscUVPWIhn3UINLEkBeN0OnIDhOq5IlaDbxCco
Sfv1hECz7aQe8/VYDbVMldoAYQXTngoB48pH76ywTUxpozeyf0HAwjq61AgUi/r+
74eN0N/LxE4LncdWvC5Y/myz/xu4ifQYKtk8dx4DjvwL9BOP+gDj6d7V/HG4v0dm
9YYNDOyW2WjX9e1bMv8iP8o4kH7lFIXrl9pDWy1js7yxV/CvmnLeA6E9fQG529jS
KWVxmb2DU/PppOev/TMYEBs3fqc6mvVYOThyDcJ5AVm2DL5rhEJbK4U2oV1AASsV
fh7egxSCGDrysFQ2pU1HIG3CfK5Ksy3fdB41VrzBVKi1dZWXMyRi6r1RNgGndMNM
039miUm1H9MxXeQLLnTQBP36P2zZ5kovPHFyw701o4Qh5nLCbsw6mBFNRsg+MCtp
B1LEgCtvj0RQBfB6VHCy0GFCiM53Y6fguqH2L6C5bL7Qvk4zMTCdB0epaqG9w/pu
NfTSJEISJPVh6eDR5aOxSkI/z1HukhB+wZm1yZ0DJCiSkE3VowYaGDY7jgHddd43
HL0xAza2EYlFXaflXAcVsv8p8x7lXS1iThfT9dJjjrU5PJIhGYskKNkqEw+yn/St
ROdmvn8D2tmEh/Iffa/kIxPNf66/JesH64n3MfSS9Nhiy8D6COtdJ3QFUTNqHt3T
JHr8ZqXiRJOQ4aCLLUrddPpp4z30sjZrsZhPDPx18w0uQ3PJnhG2nv6bhFT1l8vv
MaLTsKDwlJGud39LZ5tOdjimR5JfDrOiDvpKfbkYcdTBIFpxeMQMZcewhWDk+9N2
ypfQCdT+EQfHohGuyc0AdjT9Yzhhl9oSC9Stkmsmiq2fGaZ4RsK2I0cZPrHAJeCQ
gDJ6jNoebV9G/nQusiJGLNjxryk/J+buwgNEr9xX62lu71UTS+979Rm7O4XglJi8
/+Jp6QnXyJowBghGLj6MrY3tYgRUswmdQKOf0DmaiyWJ51lfoRN78+Sqzii7MAWp
zt8lCb7RGrPeeIVMImhWR91g9Gk5uDO8UeavD9aHSOPx6AKxYYZU5HBLikz0b25R
3ht1n3xMxLR3pblZV1qZvkDzoGsg7ETuWltbTcgLJmAr8jD8CjCLhA63iUFW8wtb
Iu6uBMACphBuQJs7W3tvqesL8fhkM0Q8ph1rOuRcoJovPtCRB+o12tdHEGVz/Jxt
j0TGLo8IbaIA/dstZW5qRcNEEIFG8ZxE50VJIU09BFCGc6YwUfImkM0HT/nnYwWG
j7tTd5HLHswYCCXtBn9tCiH17p8SXfdKv53MlD/Chka9S5NhSZIfdQolb42VQEjm
2rbsVmFfdMo5QBvkRjW3Q/GnEsOp7UJJlY4mMfqBx61zpavQ6nQDxxCIA1gcBmKL
uEGWqo7rDnGyYenoyXn5riliDrmahZU2O1nGYpHqVUHsgA2AUWmCjqcWizz54Pcj
7SQKzm1QUwVItrWS2BzbI0dzWZj1hDdESHfhxz4CCWIFYawUPbQsPSO8RpU/7Fdi
mUrf791tmE4oEE9lMse1/eyRYD4nkF7C4wmvMrVhihGd+W1/MT2cla9CiTeI+PJm
3NnQ+uuEsGzv0Ukr+MRcer9sWU34DjulnAyd/utI/EhCdDGZnRnmj0puyMfJHc+F
R2Lbc2yBcJ0Npwc2wjrrW7G3GFgaEdZTNxH62FxVhvydQGVsn5cBH1ARxtfz2Jci
6k3K/nTzqjU6Zrsj3mW68xfZEcjDEKDg3c/JOt4GzqN8Gacp51ww4zTUAj8iARdt
cV/CrMvBp4Ksn7JutyxVcs6Z3RBc46ek4qlLRLnH2juolAxdQ7ntGpzYoFbUFCC8
RlFZe5kdaEim4Vd4dpMrcjB6Owi9c8omz/mut0Z5TI/MLxsiDA7l1NZHggr2cCAD
Vha/PmK6zHmRX98pEM/KQ0Qb89IaBGbKzQKLMIw7czfz0pJZUQxYd9iZ1MoAMVWw
gI8pwQUdcSA/flP07WRH9f+U0my15cWENOvEuujkmOYZOVZmu8+NQ5E278DeYBgL
uztaa60Cw+hNbTtcqRVXkitSv7MmVrZIvqixy13YCAL2yd5RQMlVplQbHaH4JGK4
CacnZl8J5O92iKzJ6NP3dkmwghhZZZ4hXHRhRybbVuhxsUPgFr8ZOfYbgij25u2/
a4+3x2wkGCWbP6J6/KCWuK5q9sd5hmVUeZ6/AWbpdzBLHvmfsWOOA/6RsGfeQvs8
Nt1ilBIO1Fhcbng1nWDrI+WtMwEUxzqi3hB3NLabbq+dn291lnc4CJULqBSyMlPM
Hljli7HzGCukL8bhg/qF4MPTb+C4mYdRAvfNVmVuslDlo50QdtVx3p6b3d5ntf4y
Y76X75ZaqSD4yYeCvjBUFKJmMKhwYWOv5TBu1DwYAF/wMUgXtAqFOov5Dt/TAga6
Z5SAf4WWbkvkbQVEB7f3Q1835UhxMO3gZLVntC0UEz58u9Yf5zrDptNO5DAzY//+
DRwmGdz0f476ZQq0T0l1mczKFUTbDbdunEfkVjg36lJ+M1PdAdFm+W8LQ1KI/I97
qqz88zgecZkUosJxSzWd1egfHgxmdZRyEEmpSPsapAjW/UoO2nOUOc29K1gufeJc
cYddEr8/9I1xwZmw2Bx8601WepCYjrQdZLP/4yZvsv00ZuPPsHbzINXukFRQr7vs
Ugf/3U0x6hsKfNOFfgcjWp0bwsixHZNzIAxfsviCfgMZU0aTgZe+TMiUXv1HYzVB
zN1KWJl5qrMFHm/DithVEcSQbiKfRsezr+qSJ0C5Jlnn5Mu6iuCZ5hNQoC2C0qQ0
0JYRFH+rVf3o8pzKXmbCoJXPJGIgRS7leIHhbnkd6Ls2ARAoaeXIVuavUNUZttGJ
qRv2yD+7ZHiz4BomWzVvqA892/bfQtkWe52wO87HHjhKFtFQ9pG6UG/LA/P9WVez
tsptVtpicKhtI7NpFg/QcrX9spVVnVC6tXxRlaVyqOhD2boRi+kaH+txoU1pRGoS
Ge2bAOL3+jR7EeoAGCJ/FPPS5mx+Fj5EOF3nbRohDbcBiSgmYv4ksF40UnWPuJLx
sJxjkxOw1IjK7mWFWuPC1MiIlF8Ed1mYR6REQR1kdbwIDiqzAz1bYfbux3wPZapu
7iTU3zZ3/esoJpSQP5hS3aMGncl8rh+Wb0d47DNemEvj3hVAtgNgEHTXL9s69ezg
5UjcpzTY6rqCVT+mjA0RVOUfT/xNBWL9VNjEBen1n7aC7q4LqqkiTV71360zQnVq
My8Z4Hm6X8x3NuJDGxgMGntFBECijgqUqahOEwEWQgMokq0m1enzOYfivWkFVtF9
itmpWw15JWr5Bcg7iPtpBn9KQghYcPzna9cK6LhCRg0lX5KshrPN1NEb4UFMomCZ
WhrVhDKoQKyJmct3oWGLDTp2EQ+Y515jGyH2a6V6ApeLVkQITs1sdXi/S0jxaPTE
R0wsW5FFrvRHphl1rP/45rbbvC18otXu4N2BWuLYX3wHJeBEQIVHBkJX/BQeU30J
6Xv7Bn/Nq7IDBLHFJHDW3deCY2KgQYnM8+8PpUQbJT9w0BrrQMxYd1k7cXqwF9Nn
0RZ3NtjD8T4+Eo4CmazlLqtHtI+3fbTl7wwaPknwha7LY4UHU+84V1zk03Ihhpto
FEyswjm/Mz5bYYERPtxMvcN1btOFATG0GdPo1vaJfygl/syrdjHkYJaSL3WtPNAu
GXlLp5n8YexdRc5cu4HCYE0VCAOIqJyw17ACW7p1xqb3wMtmvHpR1mxloALGEFYl
h4s0UNlQvodDqoYMvEq23+UeuDRo1lKFsctwCCk6IT+hqP/eFpnNKEjl/tzeUwet
GWyNH862Ta0bBUlFgjt9aT88bxtQkiE/QQmrKVuIlPn3c9Zs5hFQuJ2V+gi691wu
D5RzTfZBBWc/EV2MrjFeTTmp6Rm4A4r0IJEoZDQ/ngMz68bZjJ463c2DhfhwX5Yu
9BRTapMJyQrJPoxYjASjB7Qseu/UdvslL19CrDi/cnYHr/Z12MRjvU0GhrmSARtm
zgCsXtj5JbfTYFBFwktWp7gxDH4Vumezs42QymD3FATqPfidXjvtwk9WoGFYjIpL
xNzytAJFHwv02UpB/+vShsdDOC4Ww6WshpUFCG9KWKBDfurX5gmpUBvhHtPp1im1
gA1m6vOHdBr5nXwtjlbLFGbm7ZQpSCmxn06LEsXIJ4ldKniL37Hl39Zd1/0XRcnu
KAR/cVfGOlCdFgZagArHgnoqMiNfzCV4CQNNFYcFi9fluPeiaNr0b61j0o89SQMr
IGlXFxprMQthE6bBK/wj86c63CF0htBlfvxDRGxGGwcPqsEtO8X3akV0psl169JC
G7t+Q8WqbHbcuHnpw1+nPHNLrrcpn5nck1+P+x7MzHK2dbpzNLGzBCIIN3uj+Cax
Gkz1fGThRhIOXZjzlLPn3ffDag5w4Ey70FZudH7FejiSuAH+DcpD2TQpqmhu+2Sk
KJgTrqASeVLXPUcCHFZ4LMBplittG69BB4wnYh1+92ZME4AK0wGsLlLY92pefZ1g
y7XzoP0pqloRb9UD4eMtEx3XxRC6/myWaX9w8fdhmUkPzP0g4dydfg3tA+mkmwHK
1gWPcU9ivC7juNhyvqv7myvd4z69e+5DsBKSFt0Sxf/YkJeJANKFKVu4YefluWpi
zOY74fOHI45K+qt+4mBY8tligTkIkB9vaQc0Cc+GfJqEZXgvoGw+XOG6GbLOlMGS
qAdLe5Q7kDdoooPF3dMTU8+922yAQmoNCtLTIrNGVT3KQy9QVh9Z69isi+Uiva0J
Wi9/iP6oeqhntx7K8ZPKS2OElxhj25grw1vRgCYv6zj+Al72pE+VlDm0T2uL9D0w
bJfL0gWWCn+oFAHn4Hmf+8em0DPqiLF1lMLdRcJHHNM4NhWE0uPkz4CF4vbtSSSc
c9zhe4cGUI+v7N8D220LJAI+XDb59ndvdNc10EsZKfIM5mORa4Jwjvi671fhJR9x
LOuzozJZMg8WwNEhvodHfljkNe1peVx1CKJ63oprE9cOADGNvvm2kVHYKT5hwWt7
krn504qQzYFu1iFLbOsrk+9kXgnosZFyfDonh5BQxduXgPOq/v8BMe30VOtd0zZM
0Z5bovJ9LE39v8wh7PAtXPNvTYBjKDLirLxlm1IvLHdZ5xXIFgBy9o4i2qBGXSNm
1UjoyD/Tk4/zM9bDrSs+fZF9ZWxgWstLK65S9rtrXtFrQouza+rEJwz6RBRGcL3D
8c0Vb1HzS5MXXhY9RdUN/XEDF6m6rlfpfEWOrIJ8DpELYiOP0DY3l9HBZVLX/X1F
6YbRL/hW8ozwMceuxOdJnvNveucI49LDzg3nb32rE8840ghLas7W1uKmcLz8eVgv
95YMQm9T5QUc6R+Ebal86Nd1LwhZJoIZb3xRBIwVBluyvjnxloSJpBs/WWgOa8iZ
lmG/mHZPxQhpUeh7QP691Omjbc0RvIMp/P4jjBjLnTfWfPYGS4WT64ro08sK/lh6
kpxW2/4HPjzcyf6/14XedakOJWcXwQaI+D2CkdMWszGampJgYt1GgxxE88LpXKBo
k8jmBCMI9IIfbe4rgWac5qE4e2XEFCNapDB5Zd0W14wZTi8s3iHn3M/iB+0fYQ/0
2KoFYuowyrtZ4BwYW2ate1Y5ZRP1c0I86WvLJOSfQ0fbJj0+5QOx6QmTsFkny4Kq
b/mHhHTHvoIzOcmPePEpUdrVQQIpgwniGlrFpNhyY03DNiW5iV1qzzKwIa1OSZPe
6jIDLUBHOKBuQXrYpHHU09xblPN1UpFw4ZBecCqb+QqjdT2oPGZahFrro9vbpCG3
QFajuujybC3+hN0NVI9HLOfYf0RbGGNbI0R8F79vQXHaEOxS70VvYlwtB7dC1MKO
1Ny6DHkyBt8WRu9pSHHYGQ2JhjloE9H44SWB746FmR1IDrhSJHv+/6DbttQ2vFdT
7idrO1mjTLGnTrOqOOCXpPsqIMcfMEZxOpguOb1PhywF9uAyeQLwzQPlI7RLDS0S
vYR0peoNAUik1GtftXTueg==
`pragma protect end_protected
