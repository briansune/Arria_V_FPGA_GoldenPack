// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:20 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LaYx2r++q/rzuKj6HpmkEzTSEydqzFPztXD7IOuRKPLiyFL/vu5hYr0TYAnjWjTM
OheRi0mrYqQbXrnmXXrQ46EGOyDifnXhQDiHRU8b2907Uso3ONwDWv/uIk2ZSTZv
bX6vZ60kDC2/ELVi4LlkpulSqK/rvgFwe9dW5ZvNRkM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26016)
qyOidhusG/Mu2fQHROj8cRCFA2B0S6Uifhk/Typ8qH9vbXZBRCgD4WF29ha01Mvt
faTHL5TbslH6Z9kl/7LYYFYv+BLLJ80pkoZeSNhZ8vNFwQoxYfSN7Simq95pQC0J
hTTivixkYGoPiy9QoAjPz1bf/N+zZmjn4ZEiiKpd+Uc3orwf3HffM4pFOKXybpmB
GWaaSfKU7CSAf3Db5aPQPXHTgSnFDu8xwaHDUZI7oNxOeUcrRycVZpp+oL+H8tb4
GjvzJRsOmvAm4J7OPVbuy4EDOlD6TkgAA9L+iXJp3N4aYgqVS5InLP1Ib0pVfs5J
bnW8GjkyGeR3KotBx8NgY3G6FHqo6uv1FIeKnEqlu0iA/BgML2/2X6Cwqu1c7iO1
cTaIYZKODT3ib7SyCBNKMrzmhTlQOAdSFsh8iHINznKqF+ziiLJ6IY3Yeg59fras
P1VAQflp2vH7Vg33dlxy6b3ESnJSi4zGuYM4WepRS3FCXV5g9FQa5wxWOamdV73+
c6ydOMMg2dLs08BgDqkodroTfG1LBi04sM1ASGnQVmwn1RGYqLMIhFN6PNU4Z9xE
V4V08PPRTKhUxOmPbn/CAKJuORycfDqBhMd3Ujbg21HYI7BpL8145shvrI1rYabn
5IH+03dA3qBLrUtkooxHYZOwi/PVYhjQKSAPxmkQKJlt09haXKmsYMthOuOC8Vrx
5mTc//UBpovQeumIewVKCFgjuBwltnUNcJ/x2LWnQhx7iXIeHN343uDXtsm1s7gI
apWaxIU9Ec8TKY808pDx5jVBw/mHBuZNFK0u9QdL8+FHeUJXZ+eeEO0PNJs9rWUn
0hPgnV7ggKwBRgen+F7yeuTo/2/AQSx7O/NIp2hQDfrGTHvcGQxWReTbYsNw4vmC
slqj4wGihM2klvo2drqodCLVN2/unyQIymDfLTIDYvWAzabUOx0jINnyVu2BgF2H
c/u2pKTdMv2+xb8Y8XGFDlrxSxEnc1fgxLMUw+qerQ+dSP432WAvqTneDtT0XfGF
XQMdv//67EirOipKwx9fSNuFDtSP+ceUzYd1C0/iFWoc14R2WB8dryZSYKFW+rbS
UQUrNxCWGaKqgSzfB04R400rUezYNdCMahbrIC/x3dHbqWxEo6NSnUbFpKx++t+a
Rv9c5topkxkLoTY8IZwoAgWcQkXubHRU7LSs4YXGzWfOFLaLI6QNf7ECD46j5BHZ
5Dq8nXP6JjEmvoeWVHKuk0TMn+hXyRTXwDQur/SPHkOhNzBANmR/tftoj0acOMaJ
HCg9MmrXTg6n05wni5aFoU8TUOi7MJ3CTUm048JtNTlT5Ca84ELLIRWw5qRlFLbc
a3mjKZ9P5iu0F1GUqXC/UTMF2qLUh1ipgSEH79DkU1lG8SxDNJt7WqgoZxUPPbv0
IsxdTHCAxXgaR38FU9A0kejAc9mYtk+xl9Kp2irRudithmxJZL0oAXfN0GDwpwx+
ZkEBFnVXQ1bJiR8nD5XkJ+hAv8vbQcrUsMoQarrrqF8rrNM+SKiJyjOYqS8dSfnU
DESAA1ScJBb1ARu20cJhZ48O4fNIB+3PBwNhB0q9MkGl2TUn4fNdEKNdQoOAg4ij
uNGz0LActLMo/4hLAkgBgkuZuz3BhZE0lPWoEHZqPGlMBfGdIMXRlRkBVYjvSfC/
QAiFYIcwiMKD+IUULvWmZs/rQAajThlSqtPtYPLCduirGNCQBGpdqN3VN8bzitkb
ivjvR+5IvomQrTN8tafNu26hKLyG4XiMAUKFYvvVJED56RSXu1+o3wr+wq+CCgDK
aV6Y6NKkn+1Ah/Gkh7AqRPdeGqZ5Y72GUHHBKGXRME3aOOykx6C9zBXLgnGJyUT5
baVlETobK/PY4bbLqZsJ6U+X7vc0J0OcS/jr1EtaUsX4Pwke9KQ/MesYZgnJS2vp
kzjWu/+hIl3RfCelTbrOyufcXl38oI9WXe2JuN6aryqF9JGkRgpZQmAjvZ/MT9SD
1nfKZdWBxF16/zHEIb5lfdx/gKqZSBQNcgTDZATl5c2o5hoYzFnSlfe0ZUPd1pa6
jcbGFcevto4noS/U8gmMBAyTkT1p3m858PZr+hqZq/UAxmzPz56NeslcYQpCfrvW
flqeF8K2BPAQuYkuQl52nw10HOHaI99/L6LjCIw6pTvmGCrQQt/uR5NgxvEF2h6K
LQgxvL8904LY7cQBWDO8TbdivOKn9Ak3v01tDer+dAGv6RXAsk4HZV9wTlm2l65Z
jK8XBbh0e4gVMXZQEy6c718MStMggnJA3e3AgkWrzwNIdxJrbzJintgmhhtkGejc
iBDF6N4xqjFaoLc2cfZhrWzrVpULdgZHu/wYgFIwXyOQ9jZNy0Hx5iK3nX69X7eN
Y5uei7PtsRHSGuDVJt4IPfdVYLsbu9WXQ0sVa/Dlsn2lPV0Fc1l9E74pZfp/6QOy
zeJz4+09ct7wPXDDrQBI0fQNHKS5IucbukwqzG6YlfltkShCr+wy9vv7eqCY21wP
vo+w/tvxPxrFpOzz6d5x9UV7hWLhKPjc8GK6TmKdXjVcP2f9VVOxvCWVMLnKfiPU
K73i5c7gSeiU4CL7ta4L6L8ibNBE1CfY4FFIOLcyBDe+avRawczsqwEOx6qVAEhR
41lzPQLev3dX7G7aKPeTic5wGl/OKDFsRnd1losVRzkJa6ftBPDRfvhwyMtISqLK
T8xezXTU5UNohdBGWbeE0XCNM92iue1mnevYiwspw00WtUXnb2gwUWAik0q5zmaW
AFqEAZFEIJR7N6zGuoAYJmKScP+7NpdoK279TI8Ms/kgD5a3NFp8KDn6HzJcLzZ/
5hbeu41uprDE5NjJiNTD3PHxUQT9/uQVaY0ino7ESA9AT7jJu/axA+yuArssQwU+
QCg7bYAIa51GvMMdCnW16Pfkhx7Zjrce4JpUcST+UA304Ps6diccqYnQeegcfbXG
UD6+G2dPAACEqTdJWcF6yM01Y+rSGwmR6DCGbas6xJeUX3/P05QBVCcQLmVGgtyK
vn52exr8o0x7oh2HEo7kJsutHfW3544E4Z8NpKFRlaykmCFE0IuYyW1jOB6ASMB5
UJubvkIBFnnDik/e5Gr2Q283H6KMp1mOULA64OURmrqi0MSnzxHGAQ5sIe2aQzc7
6rk0/CZPecbBAEggC4aSdfrsq8DY1G5N9atqLL1ouvvIo7k4p6DC99dnkUJogUCl
l84t1kOYifzZj6VzMbeDFMlLSHc76K1laYC3CIViVi0YARROnlqWBPklEAMThMrM
uTCkh+31TbR36o8bIR03s4us1WAXzpiKiULx79vHhxdd8WwL8A1coxsy/K8BEAZc
X1Lp7jZ9BrylxCr+wGLv0xIDyv5cgDnU3v2EIJvwMjCQ7ZesYWdHEtLmM63DhQms
wrSTiFsOfr71AbeHWjdmnwYbqqTYUtcbBxBEh9pmygYTVy/1QkJuqASRJBq598ol
gnO7S9NIYMU+m/zsZcFU0IO0xMmK9NFq3M0dpTe3NcaE443w1rPaTqF9Ppne8Jd0
S3h/HGfSzTJUhlkcdW9VQ6FuofGvOxEmB2i411dKB7vZJXcCUzERBtMOElHpo6/F
QgjzEebaVKJXEuhrgRJNYzMQozs6gQ8dCDuWCTC8H+eyFwgmbxjCJFYQLPHq8UXC
3zdlStmmqIQUZLak6CgBRkRFUN0AMGw+g54ziyUwvkwP5l1sO5patl3xBaOeSG79
/WqJUf2s3mQa//FL3QZ80q+Hwy+TPzy7TZKa0zYRH4iE4rMEvCL+aYR9LKxooFY2
4lBKUIgQ41LCcOmUL03G+lo3rWaEQXtZBWNXg2VVbMIIRWDQqcXTNZPLlFuSa58f
njqryAPLALj0l9qZoYupEpBDrxuIzWnaa7tIxo8uV89c3QHxGTnXAUv+5sM/lF+F
oK5qy58Vv+XiQZplF/gvr6t1r6nNaj060TV8hufnX3Ph872RUB18Od42gt7JUMTp
3Dnt9QEX78NEC9rC/5yGXqHEWW/Bsp9LcXBSUmPvy1BSNJwiarlBKVE26EvuP1rQ
/Bj2o7J5VWTHCQnF/lT5DUoiihY9PKK7mXNudNkyG5acH7ngpyKb+51kj4MxH215
j8M5vI+cZFZ4aXIz8oygeSKHpPvv8yaCmx2lWI2wOfaxyMhl1VQlUb/xNoREO5Na
j/WDtFNv+inqaETvmbg7T41FJlCX0PoMyX3bG5nWoB/46d8YWbVIRsVVbsX2yuiR
zD0bFk9MQaRoJXkT2d9xtqRGm3NLBi7wVnUXmlN2W7zScz1qX20TeKo8ewNZYPTT
F6QebQHRsuomMoMSuYIxS3inGVHn/3pcg69PJ5PwYAYEdH/ypvAigiqcJg1F4iog
0LjsaAtjCXyZPiwF1JzNZ249eI6H4srtnfD+e3xLIUQcMHUZcb+eg/hSbHurIq7l
aCVCdQJPU0V+nx5oyo32oKTwiJDM3XY4f1xejvDHzHeQoCP86DqoXs3v7trLFfb7
HGCHxzPHb8+UXNwYd7s0dRo92Vt/PcUV+pzuvAUoHVcKdnJPwX7J+sX02flavfd4
X15upEMnY7yTDq/fbE+g0YnGJJlSFBL1k66fQXxs9aZsbxM6p77VItbAabPLH9IH
sZiXCdFvSC+ZPW3Dr1eoqtoPwmHXrQiqlPA9U+jzZhWdSXEI83c40xyjMESmFvVb
F50pbA9pwkJWZggMNafCLLLGfA2PuQ+50y4v0/OrVZ8ODIYxzLDttNZ539Lvs7MS
qqlNm9H61LoQvi1L6CgvnFtE4tVPtcGsU8r4PS/J70CtxWSH51H5J8TtEM+7YVv6
If1H923n6KlNys7BnKyrlLx7N7uOqeyP4OWvYeRrX6g8euTFXY0bHMkkOBQLnAql
gi8eJWVWym7yqsOs2dglykNyA+BDLGrudTXyc8FbmV2OSEWDf3IP6UiJ1jcho6DJ
iV45NU46Oxmbf77TWT1ovFlPz6lxu64yKqEM6+PB8DcnJcRU3OfqN0+fmzDhifi6
4GTnsZfj9e0OltVQfoUnW5aCbp9B98K65npg1Y4Bai7oXwMnwhgc/XgKiQhA5W1V
KX1pZQruNlan3jNxjJAx7zpRJ3xXe7ol24J0feU5UNLfrMvo8x4+lYoR3O2uJ72l
6MZkvDW4nqv7vFKhYGRmDKiyyaAlEQSEcq5gyNPjh2acHN6i+G8ECJtCStqxIu/5
9XlxyFQIpRPcLrAmBzIdcpkq/BngItzzL/BXJsZovtmNBgUiyes5SV3GffJ49IvW
GrJYPRDddmZzNYfTdmHC+rrl/3A0+ymJCuTRIuKtFA05B3ZC9gQDrDXaIeC5Z0oe
/ZUgMhArxvVpo+dfk2zGw30SfWL3PFEIU7FspKjqSB9o/5cY6JF+n17Of+0bmES3
mmf58glUzB4CpZ8if07wB5f1ZkX4PX4hLF+IiJNmGmGESMlz7aLXt8ELRUs6wXAg
8/CPkXmsTXQozoVKGbjq7mC87UgQBupENdHZosSAHY4xi8Z0FWfeDeJDcD1WIBo6
jUstP3+tCsgM1bmcvqXLxxZygkzJ+LADw1S2OLAEOjPJuDubLQhTix3+jGsu87sq
iSObBZSnyA4bk75Jj2WfsVC2kizg8C+kK9Mp8ExdzyKu/eHxNLCvrA6+0ob3jn7Y
wn2Gr+mAevZwAEutCXrHLDlEbydKa5DzVVRc2f0cxbVcvtytSwOR5iAG0APdSi4G
iOq6GE2CvTWhf2VT6VGMfvGudeSAhj/TLt+pi0iwPnFDJjxrVT1vDYKvuMpqsf3Y
0XqdMj4ZmyBrBaECgGygq8be84q2e2DIFJ/fMi3Gz950M6q1Wu0OxLbPSN0wkCFc
A7sbawlaMRGzqlBJIF3a57+vgRTwOD0Ry+jnsv7F803s++TmTDl3qocue7ZXmiku
PMNoFxqylqX8AHRIQal3++n4Kj4y0ro4Osc1IjZYi3NvV2vuTU0kVz9O5stcrojU
WtMqZPvH5tXQg/bsZCPqvuEwtY6odCSzFJZY9Yztz2AatgzCV5kUzRLYc1F+iwew
+gaKQaUSqoXtTaKJsSTYlhtmzSlrJWnymyanarqohyvWvoCAzEKw75wc7oJctqoX
74DrjYQAO/t1it7Yitla0HC+1A2kvGFmOiHeodbr+dR/NWQUiKqlSNb0gYx8m+2D
P+0UVST18PMxbm5hX7ifM8MXlspfYLEUq/WnGMebqWwAiMd2aHHR4E8zHjKSFFjk
Pv3W7Zy+bunqSGi4NMYDD6LxEd2gP2ryndCvqpBffRo14kZZTA2bu7EMrZK8+Lvr
4iR1u9dkylwAmHWkE5menFq6vWQU5d91lK20MqgbkLe3zxZHJRZxQm6ZVuXoRTKK
PqjBPysscKKoKV++1wGVcZHgSMdelyFEdGYtsUuzFAvktZZeWKspcNZ5vD8RvgOa
5eX0zqFrrSD/vJhocF1Q68t4oFdg+p7DFcf2FBqOdXtgVK51W1XjsqrrZw5+h6ax
2LMQn4mzeozayLx5murS3G3HVr6Gt99AaQr3uUE7ODnM2STVKlgA+aSbeN0kVaVd
pcj2XhThorHnisoHH4i5+0Nqlu0p/dyJ9JZNPNFAoqfZvw/HdOsyR5Obwq+wTSqV
E9IHQtZlMboECBVrAOo7MMrY4I8RWJ+Jh5sis+qUJi0pO45ftM1WhrVS1J9Ssm1p
butuhik6brRmvUYBNoi61IgMMhMEMmtspzmj1auc6HaupLXhbIvZljZuPERBiaXn
zOS7u3j0UgqySVM6ndWcqkc7jXP0VQcFvnJMmv2s+8KzLekxgXoTo4HQes4N6sXj
GgKLSqVpvffL4QhccX6D3rXsko7alD/t8pwEqTWuGe8lhOZBKP8Zbbp9+7WKEU06
kkGQyDHmD2cb+ABeIGuiRyHOp6Zohq+M6X6Lo9Xi5zng3Ld1oM9CE0KBJpX/hPCj
//WvjqRM4vwxtcYKhm6h8pS6MLpG4eTYidWi9y+KjbNXm+YtGacBxYSBo2JWMWc9
9ajv+9Vy98johMG/c3uRGWt2OoED97goOD4/DtvmxZM9C+iQQw2nox08PHNrGpZU
Wz/4XDXHMOYtINwWLxuakCxe3VxrjAzUwQEk00FAvWKewjBcBOGZULcSImMMRtxo
sHvoBCDHxGRRn6fszQiw5PJKSME2iWjcrS9mHypcLrFEfq6yZLn60g3binb8/IS7
GhxxkRvxRt5cyZyu8I05qzKRChHPy+3MKPDwBgNEuCtnQbc9DrQhF3fnnnA4ChHw
Pe6y2VsoJzz8kfY9BKRJK8clmdy1gVhtMZBqSvyrzRCsqat//6Nsl9iXa0t2bR0W
MUTEPMMq3CDs7ePSf1TQqgqMVt9dsO4bGO5rxUec6vbzQVzFEzeLxSWzIDx94hVM
5Y0nppSNeTuwdPw40ldfJfH7X829swLWqiYLasTsgdD/ftI9IrSE11CXxD+EMpvZ
EtU0/Z4oyTy2zuqlUn5AnYifvHUvbzYrecxL8JHEBzriN3cgfQOGTw6gFWVYnqnS
Q0bjBqNBcDG2awHAg3x5BjJB5y2xyp+9t4rleLH8Pl62DXOavA7y6DzxXNl3/gc0
6VV5wShYhwxlbGJHHQhyrPEW40jEFtDqwhCI0sgBon4CvQ35fAeuHRG/TkLFiTj9
X0TRpj9bFYzsKT3Q76h11SdU2Bl1d+JBX43lDJTG0V8eYzTdTlFjr0FGCCHekUvj
GTvk4C0MA7NDtJRdtf35ChtMrLlOtL6mqDMnRONLS+/qwJGpCFc106lzC+ncXicz
C9tEmD/wqrZkxqWJcBid6JIZxuw21Qiv7xxFiPVlkhut46tZtakhAKZpKcRVUpac
3bVrZ4oF0dKr8DzS7R1duOkrUlMqdhC9yRXT5amalLic3TL2miy5c8K8KlDmXdQI
GNlntPaoA/WoT9G3LYAFzfbUZT4q1yA+m4j1bALwB6Dl6tvFHWv/qGh2P791nSih
9/pZyK5oG8ypARY89sz4K+MiBghYBI9mS4qMJ1lPr5EB45CFr6aIAlWa2WAa0jCX
w2t1TCvb8fhVr5yHeyaAwbff8ithilSBCwRHN0tqKjDHLok5qXFgrzsJsvrJnap3
d1Nioc+6o4VCQgnxJ8HD+LCCiDTi1Z6uW8YkuTHmHctyNQQrE1SmspUk39BHAP/a
IZXr/KRn0zvt46xC/r966x3og6QWSSVONUYykvPuhAA/YtWfJHsYVON8bGJG8NYF
Ya8HJCT7jCsWLEJ8UVuDs2KpSZiNx+Hm1/MYc4BIHjVOOJZICaB/QX/kCp9LgER7
BjJKwLhBoBfjfsPlC7B+qZs9ePTy0K4pTfL4NjPFhTra2goVULtbvl08hXHcGvN6
bgswcy3kdAlArYhy12zlR50Xfopp0eearqGpv33XTswJgmvXzcxe0oHnnUekvkvQ
g5mP40bnEZQL0KGcXu31HuwARfmq3lT2OtqcIuxWsnlQuMDspygX48VenXTKnxwF
QYAEh6G+GlRZqnr6x2twlvtDyvXQgiXJuEmpr5GrGGGLzvluaxIp2T/GwPi5HtsL
4glsdvoVUEmdZWLZscYb6W3Wr+crhSX1auU2fCJO1/ac0axMG9VOKnskTeVAmjRU
NkUphjM3QJ/xoiKdx3+yzMY/ZF41gJL57SdqeIHxCM+T8w/cPfuTn6FUVsbQCefr
mMlCt/mZQ5Mjj27kkFvW4T8aU3ye/sMDicnOn5z1RxehcTPs+Dy4W+TFWu3OvK9G
I9Lq9ilfieUFWqoKbHlGX9DqpSSZpCfjdA8MGhiR5DV73A6eszmWEeSg2gnDlhVp
Cr/17M1GSIfBFafrjezkB+hKbjMXrqnPFkmcWdhT0oASTT1FtoJ1tn324T0LPe84
Sv4QunWBVUDqaA0J+OB/oIHW6rdiRlVPeE6invr0VSnBPHsY6PEI5KcmfAcpvGwy
/Syykp2U+pGqgegut2sUUjAmrp9aImqi4gwzk1BnDd2w1+YAxR+G/pDAyb9PlaTt
2+kvJIrwXym8CdgzIzi4p1IA4ZJIHwCaP2b2ExLCKM1Rq0daq805XvBMADuEFt2v
CnQZPXUoGW9AsE1ETou+w3ISHEELtOTJUh2YpCpSH0JhIfdPYmSCK9d9pH88EIws
f2emALWDYsM1XsLjME0aZYBwFDF2uFXhoH876laSQbaLTi08Kr/PfKvKT+FG0Iu0
BXFnVQEODx7V1ko/ur/LelpbZYKlSVJfHj5ENYcw9sj+7fX+ZGnFk6+H0EeArFkT
J56Xv1Y+EuGUdOxiOdufafIiZYyvJgmCDzFiJjhao2td0WjNBsvQFmq1vHfG/I5r
qdfw+7qdD9SWdnYxM5dZONugE9nbbs9cLbhN0FECsn2UrqtYnPHEOh4+GTh2Sibc
P/kgLMvbkysBIV5UwP4WnNvu27qVobOmDzvNm67SaB2KRAzuVv6bZ4DjEPS/k7Sp
qBo5Uxi+mKxrOAUVpKJfKuwsnBa970AvrkcF8KZlaynRTQTJViO9L+iaDK4e6uSn
LWMfFyHfUWycWoLYAYImveqvbBUF38ChhnQsdHXgZzTu8p94MxWspEvHLWM78AR+
5bLMtW4cxHk9OfIgEBnBZNbdeR2KE+Zs7rY5iMXbtqrsmlo8tltSiJc76aD116X2
R2ddMsKx6QEYLs86/vAUEKTGgmYH1IKpq8bbEp2368BzbjYNHxP9onJaLyyc4kd0
yPUuodHUQGVkLwIYhruPwTEpfub+X2uEqjmy1tfDLJdVhNFqGcVF7euqtfaEhibl
v8Oa+OU4j10Ru4OzshFN2nP1Tzc48q7I0H1oYtrWRSSWP0HLp8YdOxzJvP0zWXoM
6PV30uucBRQvk1a2l8nwwqva+/MxCX1RwAIBJSKq8jPfnryEfg3znEUltmKRvChG
rvlYSXsa3qZr8O6RQOQe30pKUf6LSoatrTP1MAqwlCMHAFFR1qdPgqdtpAiKKySG
Z9/LGNTh/PxWO2Yx9R0wTVnvM0wVOILCdogllYkd3Ig6gySwcw9B6mH7hOKrJHZw
gnDBmUR96qiV8/cHnoe7GBZnqEcq2Z5Po7jYe7dIAnN/AYbAyNteHmWWg/l7GHFH
zFyUEF8IPTvFrRq6BsAik3MXzLOTRiUQaEq2YNnT3/Ur3LM6JORcF7Y1oVmmvCur
o2T0g7hRsgRI4NysytHoYynH/x957kfm6jl1d9eL+839jh1e5Nz9OnNWsL0KgbRc
YOshUBcFrINNJIE1GRnjVNLJbduWjsgRsDKH+WS3oSLQNs6p5Knel+7k0LmzksyA
XowqZRx+7CURJHnDTQ/sZ2vsiZNRCmYavMyVAZUVqY8yy4pjxQZCmWZ03bjqoPet
tqTNfBUdXATx6lrtK8VT4FLRzK+XOq5Ouqb69jrwd2lRzuoV97zLzx6jxfPafm1E
TNr+jjfm8qBaGBUlk6nADOl18HxiZoZZ7af+Wp1mKyawguvdhKVyiTNPh6aWXIBU
oGccwx8hQa3GkU6frFIksWaVjqJgp1zjjbOFcVpugFG4CzLUWkne4pWjgqUZJDXq
qvWeOQtFQrlEYzDN1aSHpI4wyM7NzksPU9UVksmmsnm/nieOh2vcxY8vUTXlNEHw
OljZmynzzJ5qpc1qBrYo+aPAgtghQW2SQrPbW9HS7a2IWnN+B8b/uf80Yio5R0xw
tDVueGvm3i9SXjHAtYIEYXuNr8/kQum3NQSrfb1i6Ev63dKLrrrxtYWZoZbacm8B
YCWZ/+gBFUvaoZnL6p/7Rp204cp8rTXUeZo3uvSRziDRvxCYK2DJ1A3YWiC4XAYW
825ci+MaGETp7ESG9bke7PPWUzFj+H7JdcfNre+RuFs824NHd5pXdlXg0NzRwbtt
hi+qYj4vX3W4O50NkVGkm+n2ZrIwdP+JdNPNSwjjJ7AXpJDjvWnEdUjlDOrwCJft
ZWnY5B3jNI3/cvPcV1SDUzBOfsP90Vx3il381IQaKKdA9QSQNCpxtXNeo1smkHOS
nTR6VNDqF+QoKlmJoIe8V+1lB7PlxVHJagJ5v1qPIhG6qJ9e8hDFHC6cKRFfatof
BZd10DqoEnuDb0A4MI4wvLrJok3O8VNBDDWuNqN9Zhn5RvOscQ6//s3tTNqtNsdq
ZSyivbsj7KSHJZ1jpHr039y+8D0KK3aSQBYE9+24ovtgmSHJpWDHgC950DzBV+vk
2eiY7ifFmbIz+fxQELQEe+B2hja2F6oYPEucfE/Qq+ORcIYvptMM2CM72GwmOYKt
pDHEaKGHd+M4X+Uohs5fpqKKOC71aMXM3Q+tSHBtoWMQTuLKHkRSRejKseEugMp4
/Wpjon9n9gnLjVhBrs8G3mfAJmgx15NQPRMTFlufqDulfbQRKpfyE1zszoIPifky
b+pGKSzE0oIxlA9XzhT3OzrxgppYW2JXlUKtAuj6z9QwMJ3eM7TjK8Qx9kQwUR+v
iFmbFG/6xVsGO/Aeai+X08jicyAwHBwtBmNV4iWaQjcFHO45cGUTVpyJrerUID8h
qYjDB+nWSD5Twzr+IF8cgCUoAF3GIQWMwzAKNOVrXsSSCkk9kds0AhrOYbSwswIx
loNRcbHW8SiqlQA8VXdyCGZ3yed41FCiDZ9wJ/I7+KKstN8tAuB3z/3CuJxlRiCZ
0KWP7YkhZw7ykR4d1pMiWMCZ4I4i5zMMWAt/F6M34EF+zdHvVX1QO3IJbcPFXmBp
OqO7dsNVMJyEHKFkQdBHMEcZt0LmbLBPtsTTkkphDwWD4tTmbx9UdjKCKbN7eVtI
x0RwI6kQAeeZvtWQ4hH3MpVznLXXEp7mrdC/UP1cErD5AUs7aTjLe8ojYy0jewcc
K6HWvP0IkkXsbHgY9YSB2XLDer2perGTetCzEJZ3T2yyo9CVYSjq4TnsDgEkYPPX
1wPVJUsUY0/chUay7A3c0j0La+l+HRff2k61rg1u/y1lBr1NbsuRfUFdm/GhPNEh
eIwUrb4/w1tqXpUowhHaunyFse35mVbnFT3O31ROXqV729U5lDvNaIGqUAVbjlI9
BKm2psH9pNe8MLR1aobf9Ete8z2bswEc2/9tGHPeeVxxU3pF1yCrQROouqoA7q4C
amxFnhKvqDrntM3gsztX2tSvLM0+ajBh59Q3X7PY0dv+TOXubNyWjeF3/AiokKmN
BgXKFO2wx9mowjegD/3SJHVGZGE3LBTROSfK3O+ilnaKJj4KNyk7s44FC0lwFr7a
5O8bktuba+igxeVk9c1tqnPrE7admIqMBXg079FlvVngVN78NYg9SLqYaw34flCk
hF9PHF6ebGLrxeea9xlGdJvqC9mCGHeHF6GDUOw9W2+HX3hyoZ7fnPG/BEWQH9EK
nYnSlZp8vndyaFaVvyTgRUF1RlXFTCNHcnijsNJ58qlQiNaTbOvk2emopSUZjA80
E/SNF+UVkdO8kX6Y0uTQEA+YqWnvGYOq/2Bmmrf1d6tf+jG3+IsqP5Zfqx3q0iAy
kWiHNVNxkCkwLIiK8pjixTe7Bc3Ykz7uhV9YiXrFwINbUEWczRnAgdT2Tn4WCE1Z
LbZt6Te3JborygbWd9Z3qApoy3I9KsUp5qhCCYhNpeHDt0WLwViFbaDJ32uLY/A+
AXayfmoF4ia/6zmsbpgO9Qm5QGJKwy9Ve+Ls5K1w1dgfsTTtE6vIqVV9yZ1pJlMA
CX4Zz8P/87IoRMKEJxTAUAD9VEk4tnsDSKr1kzShp7DiGsIzHIpkcDzWjXX7hynn
eB0bIhq1n3ieKJrI8D7UtCo6ybSMwtctwuwQvFnC4jHzy1z8Nr9bv9vbr5GW5bbQ
kluhw/YDukcadyOG32P7ou3SI4+hqBNbhXD9fwj+xrw8PMzc9gu+z1GCfENLbE/n
suuFoIQklurGHXdW4C2XONxXiZ4rGpcRKXt0UdEF3FnJsayvdxSqqZnZLXZXtuPJ
I+oRB/FLV/o6BH9q1T4ascNHEC3aHbJj1wDUyqAlhxYIkQUJxbzhhCV3IRHZZMnW
j5++LKMAmwS/gqy6sFfsBtvU8hhA+Om0f+Fc9isca3VuVoEB69lpPlL0ec7YZSSV
p/bXk2q/FBOu6G9L/SOrSC/mVvSwRUrP31EoNix8hQ6I7b+ng4e3vzR74hngda1K
EHl2F0UQK9F+k/yQWEVPJNZ5kXdM+WgWInB8y/ccAZMe1jpeH0N5fzL4YBuSc1gb
aALINeB56plAHKd4sgKZnx2gjexdlPFMWHdGNeGoheUacFxema+AfARwJTuLALWN
DqTimWtYOkrWqgqdsMdhUHe73fEHxwFKWJVtI27cVGcvYVeovDrlZvVMqtaQy/Ch
X94NFCjvVpGviulXp45HtRFtBM2f3xCBAZ9cjUtJfQUoJRpxuJez7PY8XCyrjL3l
FkaMUcngUMIOp7jWOcSU3Fu7tVywXwp/BNxyZzS9E3o2s9QT18mBcNOZ8nJuuA7d
B8nBaotmBMLbPJ1+SUnOqg+GNCquyWDM5/VIoaDb1rEfuHH3rUak1bmdj+/d2Rtz
miE7K6uCC0WU8eg7NsaexCz3eURoxvs4WTucadkG17avGLNnSOQ85yujk3NkPvEW
8+w1BgwBbPdkBh+tqWUPkQZsYyW2G4RAeqDiq96NXvYmqLGxk0d03zG7R4TsjxG5
QUVrPGtMe/jl9/b2x8UcO8dBAj7b6d9nkYQrmUfXuBPJyrjtyBWvA7APxF95CASn
4UCF2SC61TwBzKePEc/mJBqlKWMyzM7QDh1kyjVd1PQQwQ9gcjs321O5/0F8/XsF
aHWInlzqV5/KZ8wh/xxkK72cpez6t2fqFbTQFNoqceW1Ybk/uSe0VZ49K6QPFmOt
ICJ26nQAJFH/aRAV1M2pxUE8HS5RsTsonbcQLNlm6GVjzDS3pvFdYXRoY3rP6rxo
S413IG3/E87Fud4r2jegpmsATUHqm54lWU48YPan7srHZTFa/cbXPJORQeypnYTW
kmtgKoel29Hj4C8PQHTIMZKwLPfxEdszCWEnHODCWd872yC7cwgepcjmLl0j0Gq+
s+cVUCTAuQcD0qHr+prF9bNfh8uoyAvaAFr/o7OKIA8yret0fAxNLZzLHM46lVps
aCFZiAsRclK8254fh2bO/0a0TSr3Qfm/FahRIPUIoGI0RHJIuxY4cMh3b371Sq4d
8oCCovYO0kdvY4HjOcc9njWPwcar4CTyMK3Hh89DGGSnlgNF/9OTu+F8ctDnB2h9
n0dnozpdp1XJwIDy9pBtEbwx4vDalML3wiHMF29Q2yCXyzMnWZ08bPbXwiE9Iow2
tT4ilVjbfaocJHQ9X3wXhAOqYHmbJzXXtNSnJwBPHoc1hjr97XV2NAx2YubbTr0V
TKgKtKaFD0TbIXawydK8T+IW9GRk8TkTBxCYS055cwSODzm68Y4QDYUxV9PMTnwM
eM29Eh+kE1ug1/sc7fRQTU4MJqFLMGyEcE0rW0ZxA8S0v+pJGyXldGZtACGibVmJ
fia/r81Bv71LOEsNxJHoSvXf0KciAimGN6uLoXask7FXJEpmrfkGQC/GE26WoxH/
+59CO9kZKUwGciokMJiBJte7JDGQwB5k4tbG5cTkQcuWazjMeB3UAnf9bu9ubrlZ
z2Schb1glqRg3YGvEKVet/BmvHc18IpsFWjjZieF29Zh/ZLUnCVluLoBXqNDGj7K
CeJFDLa/UJI7we+3aMXJnzqF9KJLsnR+63iUoDLDWalVSril3Ie5IZl94FSrYpmT
PzHPQc1Mg3MRP+CvIrxMYco3eWE6vf0tJxW6qOfQ3pSpDWUY4jI/K6esodiJackW
dzh9qRCdkBHWbDCH8Yl+WmCrcB+5euNEWXgiaKESO+myG9eWm5cpqKVImL5UA8Xe
SWhuwJ6dQzE05AhegwxNQQJpcYxUGSoKgWt3j7/N4MI0MG+ztkGtL8RvCHv9p2ri
f6ScUBcuFOX/l8PHMjsDDdJ7E/yTva+6pJ32Toqc0fmdSK5wCDYwbI5NTElWZuB7
8Xv5JEAxubLbLHCz+GW3UBSP7ke+J5jyaCoxWqiA0J7NAlcwrEpBpI61XzvTz6PM
xdQw1M8dTSXK/iG8n/hxI08k2CiiryC3VQqZmtkZaVzGi3nXt36BRvM3dUidaLbD
DsrRF/sHOfuwWiQV9X+dctrpoR1OcJkl3DuhYseXZ+HyyruycXJ7dJFHnLe50++X
ZM+c0gshxkMHhOPsTSFm8DcuNB11lqVbQIs5EexCqAhiB30iIF83j9QnJpOXQqk3
2Kkk3jKBz52RtnM+PArrasi76qpeuima8LzvKRNkblL1kqmsN1/do83C+jD664uW
GP4xDCst0iJ/CeEMkI6onsxZm/aVvvV8W7iHg+I/qPCKmtm8rxOZy2L4klr51Db0
3ec9FQi80a6Ng0RakokwKs7gzWAd45VKj7EpOaeZlNmZQBfQN72/fwlu4Yl0zgj+
SIMCcLXhWD98Zn+fDgLE+wKzDyc0/zUfPPlBNNtaTbQAPxOBfEtOjI9U19ds2FIF
eLHa/ZH4GEjfEzRTQs9/nXYvTWXVm39u28/4rgAxL+lnorr0OwC5MBqDo01I70F2
Axn5rJikVqllCSssMKMvIntmC+M4TL1uNQ25i/x9bN1Rm9+XAi4RDEUZdffhNniC
+NHAfx9Rb8kkrUUtTW5HZV/3IiyeGa5p5hzny9lYPIjC7RnHkEmNj2Uej5ByUaFo
Yne+GZC1C2x+fX4PIxuZi8T/Xo31kr9X/oPChOmEfbMIf/pwcghZpo4BCvx8nuPn
dnYW6jAnvu7RGXIzvfdMSPGDq0I21ssdSVFEif2ia5nsUXrrr5ae8RQ5o1afqXdQ
Z4k03cPLSk/16y6AxHwGg+XBYrOuTaMfG7MDjo8OcITW6SFF75MKobpWKwLrdTeo
FbLSyd9HJW0J2lto614ZyCaM5EYPupUoUzyr8CtFPPEGumw0rtWyvNRtKwE8WU6M
yi+SFT94nkRqc6tzkQ85lYywNamiU5IHR+D0SWFHuqEWzmcOOFf+7RJhYyNvB15J
aUoK7kcEFkjYS7mL0fKjSSlG9y00RhNP5veGMAPNIOGTMcYU5E4vyR4W/yh1lphl
szUZSNTTd3fsbRyuDn2yeU98lAB9xWVlGIf7DL8Rh2I2E/rWYOHQ14UROg6tp6Ix
HuYQUFZ5QTuT/oA8+eeL/M8O8S5Mdv3bRLR9RY8DIsF2EMB8l+VnVAAz5rP242Hq
uAJk5pdYVEQald/YzqNWqL65Yoj5K1gphIueyoEnfVk/x9D1IrG01mC5QZLc3gCB
3HkDZ7Kb/44MWjwtIfDZXtsYjpVxPF5+1JUNABv1e/pGIMFEPYMmo4rvvojvqD3+
AdNq8UTGzd+ThxLhqeFAC7dWHCjrg/cBKfUU9QIkuUFtBggBp1/Te/RY7+wCj64N
ddrz05iTGvtKewWRseM1w+CC0WJN3QiUvpNBXg8cusCAk+ByDDsuk1rRZ/6PONbE
hmlFRZEoHX65l0h5p63UXgprXwuel4DeEkdxMtWQxD+Q//CMZpfSFGwdqtcdKXjS
m+N9sbtegcZx/wqIEOC5rr/u3glVx/aLTk+3AhWAj30dKjuOBY6b2+7eHfocxgVJ
ndzeMgSZ85u3tB7XsZ+rOO7BOo7lnz71gaauI1ESMSejp8P+jJHFmesvaMByIgwE
sN/PlubVDb6L9r2HRpqn/HvdTSTU0GXPmi2mOWOmEF7okAJXptWtSBC4hcJ5Do06
YAzkbgdXjiu+Nockh7zxjQYxIsl1qEvCKE3QocidgzriuDkUp3k6pyOlboM3dZgg
98zLLMq8L/y22/m1tsu685H4cQtNM34S6B651miEIFMiW0AIX7tplHBuRpGsRODA
WKl9yosEhX9z3JR2NtXgDhmVqIUreTjfeahPOzYzsAeXcQ12bEo4+mPjdRHIMtUd
OE8ZrxCN808O6sA8Jl7jEAX5ENVRiP/rUKMVUZ6V7nVBNo9NhP+fSeEQER+Vw6CK
qLq89ePk0IxVJdHXVGCGqUT9X0JRaNW5DskteONGY41qi96QNttGs2+2KX+X4G25
iO4xSoHEoCXexdjjcvY8tiZ0Ng5wXeJyLaHDUSv3Jzo5hCSpkINDOMIG2Ph4N1Dd
MgaAwfGo3ecWDp206Qv7AC1XXElIoRXn+nTbZ+BEU++o2vOlvxihvCoZ9/xUFtJ1
fj5I0jpebu3FMTg46uIR8FiFKBp//G3xkrImSchfdJzAWNlWJUHlr1PrpUMCbYFz
gz2qqF8BW0utiZsDw1r7aN7pJZG+uRLf+Iq8HIBX83m/DzIJPX9Q3zgovY61vcOf
JTA/HgSq5QfegRi6uI/Zfj+Aa4Qm/4gA6s6ztLN9XrpgylP1/bey5NNne2AWSXLD
jRktCcBEfHiKlAv2+0IdkzjDS/mvFs8No6zF6T5GGsflySiyvrdeVqcwaalQcBIw
RENNtyM6baiQJMdYS2e0jx6TUErnLt/jQQT7PF8xRxnEH9dfpiKPCBgjamnCvdWv
bVBQbYJoHYOYXPQyAcbnAmti9LxaoYCzEaBvLGs9pGNsuGuShGFIZ8Da0vIUoCGl
ccNzAcQVYMn0JdPHXc1qTNkPZp0TvMcz/SHOGPLPsbjTeBjgpeZgotIJr+kzQYKN
no83uhHGSKKlc+oIn8s7lanAZ68brcQhPUhU4tksvUZMy+QIZ0fiLolFJfdWCgvY
Y1YKdMe2nZpb3kFV5Qa1szEGsxqsMptY6D96iFFU8voaunVMnPBseXifr9LljB1F
wxmAlcwGjaD7zEKP5stY0SsjQxkc7H5BOAL/0SxYZMi4xSmsBESDjDupdbT1eIXA
zmuQe9kPy/B14dS8N1eJYPgwPx10SOX0vJ5jUUwl5/oytlDcK+OF+ziRDZgAHeum
2n38V+5jqvg2QM+Uy3ABMaZ6D3kSdP24eCEyOVFsydtmMgqfQu0c1qE8h2E9V/RS
j4bbtNNDJyid2teUiCY5pJaT9V7/mSmXHAf2nhgqMY6pTmb8qb2jE21NeQyDFP6x
PBQIIl0AYbF7fjg3DJsWWZyz9evcw8UhWC1GkoAOxrJgpRqb/fRX3Dg9dahbHpEf
1p+ZBp6qUmt4rRb/hHt5BAHZZB8ob35BkvHa2+dxodjdWk04C2XQHGuDlMgQnkB8
KhgMpCRXs5AXi6nmunflmhGo2d164MQXGdj2aAAVgUPnGW1IA0AvH3QzBTttk+ur
fpbTuQDcS21kLdCucBEn7rX00soIlhlpq7DNcyO1Q5g8elnG9Wn3Nmhs/K5gh/y1
kmQkKGAhp0i3vbD3zZaNh2NreJcp6spVnOJdVxRMIPBRHlfwbwZwQ7k82QwXekyi
CGQgPiKAMAzfVWFrL3Zz/DmIUgvJolb4mGTjzyak1uFdzgrJYrM9vMR992KESbXz
UpA6u3Mr3nK0vR/jZ47RRIf0SdkToJmsC2qFPyGnSaPDSRFvfJEvf5axvemdg93V
zLQ3XDi7jWCaXvt2jfxErBAcZQM/SgBYpZMdGzbZfs9UQGBrLNZLVLBtU7MijWN9
jTcw+Yc9cF38UDrTqNExw73UCSRYxmlkJu3n839zLyyt+obHRhe2/gQUY21IdmC2
VwNoxOccs3OjV/6HaugqzSrn0162NwoJptPsBQDePLCBAtCKNa8zghuZY7dA/ON3
3J2wU/IFQmipKoeSbJsp6oLJ7NRjz7moRM+fuv9Rekq0ql74M5upLnt8ocMmSbgt
2ZsJErv9zliXLHSuMNP9Jz5KJIMvpVpq3WZ0sFlwhALqN2Ko3G6KjL4t4tSPM+ud
2XpgRv0JRu9ijH7n0bPODHGqDO93c2yMaXXMS0DF7XBG1lCfWB0uF9qHuuyVlOLl
OwYEc9fv+6ijCIghIZLArh9MfDG19rDJPAw1OH9BLwHlsrR5vIZ7aPzffJP5XX4V
vomHwCMqyboQVBfaqRRTciIiaYgonAUa/6VTQi4ekzs3DnG9gxMlZ6elZChXZ4pz
lga0q8+T68yap719MRVyr8t9aCR/6AlREsY5tdykD4SQVGVJpLceT2yJR2wUzuey
UhkiuONjTqpBRMz+w/mDtACaQMO80aaoGzLyvG5pWfzqk0tNuUYjPf1VoilZc7DM
CPqJRWA79V4JklCRzie+e3NsugrosvwY5rsn9TLgxV8FWFVaRf+cETKHf2/5CIVi
lPYCt9VbuzeAjlQn1aDZR0IaxREbM3F1YpBxUTKOlWpyPHeDL0kkrVfa8B32vUBV
tjthVlfvCt8apa99ZUuKuq9NvuveTaf+CUduQCAG2bpWU2PBb7sBdYCgh89R2cd5
Kqs535eOGkdmNDvfWWOEMM2shPot0zr8BIsMwMSVXT/uGB7isshQiU7UHjOpBNNz
92yUq1wePs+tWvWnRIX14KfS8Yu4cpZhWOF6uQ/vGbg0fLxExEXe7zzIraXUa1mC
GaPFL638moquV4X4/h2p1WXUwHBVzdkCy07MTsnI4N4WDkuD0DnQecYE26D1Z5rB
M7R3CnhhZ2jtBw4/3QfDL3JLNhPMTyYqyMLkzIQUCeM4D3jBPz0Lj2JiHclIYoM5
XRFFOoky3X5Sbeh6LNEaQ4OR+P+9o5UYt7xLnxORuqQPsB2iKdIum2ia/q79hCOI
cV1w6wriAm0f/rd/uA2lK6T4Ehm1EYdW8yeTtWF/i9he1C0o0xCXdI3NXP5cQd/a
ToRT+PFjTzZ1QD2SP/9b2t69i3yQELjtE53nvHjaWg/6v1D3Sim2LnDV9pUQvPIZ
jbpcwcuuDXU7BtQdVUcQ7ZEzP6Qi9QR/o664kPqsnconv6iEtGytHUygY1SzSSpS
z5qlnXqpWceEz99iSzWNIuxUE6ehHvUdiymNkiTvF1StpFTcMh24IRQibxHPsrke
/RjZPPd4TiNWdRVSfRYMYq6ZSEsb5A/pxdCen4FwYGW9/rF/B5O/DE0BNVTd2ysc
YYKJTQwYVbgIynZ2qiGQHM9EQ4LXQ3HqQw6eOjtnV9JDR1QHcRP7K0JqS8I9j8hu
hGGbTZNzKRYVMBgRqByGGt4qOQ2JysDQPEydqgZ2bxOQb27wsERf93WPtFVXBN0K
HNo0wkYuXvkvfJUU6PDKTbwlEOwlx4r4fQt7JQJAQ+E0oqijr7v/Ax8w1fiFUi1s
6NsghptGOhfZHZvRB7sJFKT7eYiCFtu1y1aQsSpcuFBXoAXi2SHdtZAFEezcpmMR
RMBNWeiOBuTz7s6U/73XJqnTWDYA4zW0cgjV5C2n45UspwmQr2NDsdZT15Hx2P2v
l0JYJFgjv+8pM+9QM4DePk0X8X6iMzySS0ZvZE31bH6wWpoH9CoAw6R1QMN89/Y1
UpgyChcSfntcqktYEvKObGz+JxRhz1MxeoJCcwiDnD+pGfIvEGJfj386Y3tm8unw
ileaBxNthU9HRajvQX7bu2L0QnPmuJVMK1wY6o4eJtGk6e/0Xfj8GoRg/JOYkK55
44BNBiJ61Wfn9eYWX2/+KP3Uzcyk6kqWa5Bpyng8iRKOJC/hVM90JTHLuD2R2w+v
IjRPcO0kA7V8ii31zf7mS2OUQaTj1pgoel7eoms6OAHmABq91cXZIniRIdKOuXbF
oVRhV9nizgGjZuvCcMg5WHxmz0CO29kf73/XXgf3Lz7cSJOoO/VchFHf3vJbHhR6
2vUYE6RB6W6L8pIIcBf1k/ZKPVIh/ys9wDhRtYfnj/APTj5q0aZYpxoqhxrzO/2f
dhhhutOA/lBASQ1X0fijg2KHocVl8/mLqj1t2z80wT2++rjfUBG0IyIhU02q3s9l
0NBG3s8/mpaHut6g6bTE/EOBoJ6gPZq3D1D3WT56pmDMhVK8OS6lsXQ6S1Pq/B25
aMzxonnxoKsSzPA4JJt/I6JQt+dHRW2IGmvTwctuBu9eGStywhAoyHfe7Xt243ds
p5pTwrChdIL0LJtvVSTEvPSX20+RMP7n+inrliWiww5FaroybgYT1bECoLp6gfs3
7qyereFrI2n2AfwJll13lyW/JdZJ1ZyIQK9C69xrUN6WnLa5QEGxgfHiG83C7S+O
0/zGReghpn69mrcdz7VXKU/cJUh7usn4evlAAylh/qfUgOf65ySKSnnI+8X6eSvN
cNxqEhx4MOjodwrUGjua8Tg8eyAfClS9SYXCT+l6DipdN3kL0MaStxxoXV+f8nJ8
bKEx8+jkBtcvtczMchHFfnrD5AC0V653csMzy4K90ku0uqHAyKR46o4pTjwB3Ra8
Tsfv3iIu4T/ecLVWJrCpe5gVJErFLLCb2lSeWExKYIHIN+ogrXnUiGUXLvWv8Cd/
35gHXzRtaaiSuIKSDReGkzoJr3R85/05/RL7HFxE5EFVrNH1Cn7KPKy98U876+R+
2Dd7/NAZX7syrRr84+7XAZMWCTtVR3YkBSoFIdykNicoX7z6YRMRerOoCzbOdSz1
bhuI0Kzs06odGpxAK0GTEBJHH31nvjePAT9W+RfWFrjyYNln4iHnJzVVzDDcraQ1
HvzBqBMp3KfaI2tdA/gdy6O4cua/E0Hp4eg0pO1i/ViFWLBha42jMSYNdkCvxwVH
mjJTLJ1zq2MJmBkFsCRW8ij4seLqfFql4H23J02SZMNJqeRNq0wrNOckjl5JYIUA
cK80OIC/SaVqhU60hcPlhuNIVpsf8XtIlXQ/h7garmnllpypZfInHzN3GSY94sfp
3mLU+tsEG7W4fyACMw+IvPLE3WC6y3AbBsJAouUkPRBfdqOdDJ8lF330/epn3kzL
ce9XB2gFbiLtAZ8XugwzI/hHwKxgHb8o+uYwyEfFYR2j2ZH5ejucrojjDXuqlYmb
G0y3nuDU+Cq1EmWI+XBlle++xFsUPd0BUblqSJlZCUpV+1VHuelPJ7/oWfUgCNbN
0V+p+Ej7b3kyro2R1Kbvnc5WVKIIpSh39TuYaQpjx3vjLV7sm373rqsp4hMx+mmq
q5R/fGKuyxFkPJ7Fkra3s/7Ujiehy1ExzrvTS1t8+VuQedKlQylVL2+7Tv77nvYZ
QSRUlD8++8uJDZQLwcNUxAwcljsNhl3mO2a7p8aAzqa5J35CHXl2sdMQeeUasPEZ
4byiWTsbUYic2oIDGOBrXlYO3aILybkI1W75IzpWFiupKQpSDXaqOpiWZsESkSc+
j+m4d9nrPDQ6kHU6ymhQXzK5unB2KAqhSHmgiHqeba67bsWq53ZeBPugP9359tFf
gnGgFe2jai7ZyI/GqvXCwoAtQi4mwQRj3HtfqrpC+cE58Jrx8+4kPJ4e34bPQtvJ
T/751bunHsUg+I3pdXyQ/xZeZb1qm4nKW7wil7/LGIXMG3a0cIDngT20tkMbzFcI
jMQ/sXGe9DHSoXGhIxkfK1TbECeuu5OAoAp8NGhsV2sVM/CsymVOFyftuvWWvCAp
OEoQxGz7jPyv3hwA+YllJcokn0lnSVgqxH6yB2WK7ts98fWA8HyjWdbpepECbJ39
GtiCLC2vgNUdErA7IIuzGauBHZa2MTOaa1S/S3ZwAn3yXWEJJXjSMZrP9PLApC4B
cge52UrYueqTmCWnZ5BaVarHbqRdEq1/LERZPTlremlZQdOoCHGg9NEU6BRdMbZi
VCxpPSD5I1bbSRxSe9Te8EpM+lhZPEeMPi/RF+Uz0dQebrazBHK9/b0ac1VpOCXz
y3yjo7irmF7/fm+T16EddQwDLSEous1U3lKdz9uSWkBCJ9TCd2NS00TyyDnnxSx0
CY6/LMO7XvlUYgO08kVdN0ToQYqTvxfD2wsaIVnG3Mctq3rQxxx6+njTThHy7JOo
X8QOnOVjTpg01+rjKEbhBcF46XsyGpkjw/TX2mgpZdLnB4Rwp2PMI6Z2Kt/tSC5t
RhupAf2GpYd92+8REKgRkYFiovm+ytMVvuPpCMXGFM/XSUNTTVuEJOx3gQjXEegI
LE+NvIakxCtIlyMsc2RC0It1qGkgvt6EATiMRTKdyMHrUgkNAoG3GFaW22cvyBY0
C9MbkwIfrnLKuJYulT0SMznzGo5qX0F6j9Y4ibWtPY32+I6R1kLlH0cY92i1ncdZ
7yF4iKeP9LTVPeJUQ2n6VWLA1rBcpdCG6SpVtwfpyznJYKE0XlFbvuyDA+5/vaMM
1MrxVB48ibs1A7PEuEXDiM4CCRr5XQ2LGOhH5S0GkXmPEjHKvt7MccnHqwHZ4GBA
JEHHsrYCu6COOih1sUDJdrsXQW1/M2Dy4+7Id3g6/zhUtXEzjE9tpj0WQLeDjfBj
CglVWcidJfkzSTjlQ5t/LgMLR4AQtCG2hYW2n5SUEDz6gFyBxm0rLhBg8RIM6PwR
t2ffop0JjVAOqyPho7EOg79jd5ZrbVBIvWdEGBG7id3ZKn/LdCFDpuqySM+Q+p6n
1Y7THx5KkPzpC1bcPSe0cCC0YHr6ffUl8tIYrZBvvtuIvFx1zZz4Ckg6k/isP5Tr
yjx2rOYMblIc9Gbr9ouGOVCy5wgIUXnZavd/CUllx/zUvDbVJsQgy2NxlILcB9T6
fKAyZXxUwCDXFjJaDbNXm9D5VmPk3QJj2s1SH8X679SJ5KwcAAMVj6xI9jEgKrtn
bafdvIgd4OihGb+VSdKepxwuWALh9zNN0LgPm6hhE8lqKJE7RH3W1g8k9cvL0HXP
Xni30mvf4TFqs4Aa+q/U8aqwaBQVmrVIGxYNJRXfgt5Dl4v5J2uxl0KWLxOFRWu3
u5M2b2R/2zq9DNoCpG9HxI8HF2Q5XATXUkSN4x8DERrmj5+nn+wX94nlq35GIB1u
R0tXanndTX+HC5U3wLDJlAXAn7gJjadJ/rov11WSeFcGurecZ4T9qaDojAhC348j
5VPp5JSvvT4TbejVtUyOaIGOcxYkwJojEhhFjEbON7eEwUpmdbkw+/liV3b5OH/5
psFoJBwmVZW8Hs8H1tljrMwbUqMqu3AVXPVR1KJk9plqlO0lYhUMKw2rIPAPJLm0
3nQ25q9I5VAVSuvsMqhIj02vpJ03ZPegWS3tZD4TR3htQ8D/9wbSJDJjmfhWfftk
BX293pdi9gQ8a+cHOCJ5RMw543BmdbK2Kyx5oyDfVx054XuevwwJSXNMyaN36SEC
ykPY7/cLtnBDCpybzySJEKbeQj93s0F2tpJU+3Qtc56AvzW8OhCx7a01OTiex9/k
hTiUL/RU/AlYBPqY2Rdw3zKJr5pmB/xe+9H7n/L+P9Q6TdX30mlTaLrk64peaXMf
6pvh9yyO0fKXJ82PlAD2QQ5QwWy7OmzXV4oWtajg6BB8dD9Vc94uEYwO0Wwitnaz
rpiTkEtYmm1rgxzzOGSShoVvHMm+3pKaL5GFp5ar9K6EuUbxqLzmov+k0yNNAlpF
oqsrWc0Ooyyafu1sz1TRai2yk18Ygoat0T36nOxVd6r7W9RCGSOUSTmZU8/l8IOl
hkIlzzTh02ApFrFUG8h0Lqhkns7k2mpRT3HqE3XQaZ6kjPCvq5Fp8lCo5bsygyMd
rrEkhaW37LtCb3kvmLs4ktd3G5O+FKqmzyyoVScs9mem+zMEE1tqN23UqeAde9b8
ES+yCQcmVDZw8i1ZkXx3AHSvaZLqvLsbL5cJlZQuamvx4FRm19lsDE2AzvswNGRA
QRq9uyXVxOCwH/eLLVZesmBo98jRaBwxqmMjBzmh/KSR0bNNOieH5BeprC+h/RIq
xMBsZiCCjQKj+17f+ptTYa5RbWPm7KouZrV7QvqTcNzocAOJhRGSfDtU8YuevRA9
G2sXjoXR3sYMg5FcrQE7waKoXuHHNA8KQnp+/C1i3lgNs51pbUQWIA7AM7S8UE9x
PBsx0HbbIGP/tgosvtP+eHcM3GNBdEL1aJXAQWF3/L6BRM2miDfUZBCRc+Anbxq6
30+vLbtr67/30y74Cm4te6SQZtwPkHreQnZCRipbSllbmS7gz2tW5Gv7GVunYqQE
veh5qXNvnrUPPur4KQVKI24BLnrKXqLDtMf1Wavv9jdvdbe4I3XUor4myqRasvQs
gNsOK0XAaR6Z0T3R7km9OFfdrEgjmGsw6tu7OV2FqTcQdtAzwTXMmuocPorNNPXT
mKdPwENNMpubEHz6cw/hnSD8vjfyel0/P8LEQxB8wgk4Ld82ucO2U9ci0QhkM9Li
NUGokzsYVbofosTfyj2wbUGJdxX7qshJdWPDdXMB2S1o+EvgfJ7DTGecgZk7GJw+
cDi1772l6WpYJY0d3/WDgL6pBO+vzlT90GkxqSNRvmJUCPItQ9NHOeFm0UrQ6v0v
oye+HDGgun/KGhlPpXr4JaBX17qKC0AY7/MlEIYTtxQesD2iFQjsbF2KYRuLXhf0
P1noZV8nxbjFTVkGXYIMQfsum36G9ZOXKbidbR+2qgUnCu8D6/M/giLweCYvOHtU
geLOxi/irKYCWVt1PENviH1wYTVZyHcfgwuonhe/lx8tLwobMz4N+2XnDF/SDXS3
LpOCV6Ipi2VS6tBhXgE5YNUKGSyIZDGH5TzZkbBO0SAec+Gh1k1rGbyj8srqAUqp
5J6d7OTo1pPLCixHnYpnQhZdrwAzSJy+RdNWnliRfjGrK/tHSaEInZQ8WitfmkUV
m2lKiU+O3+gAYhmA0QTuP4ys99jq1ncD0h5XsA9n18Zo4bCg4pfJTPyFgEtGGDcc
rbghVWLMBTCrP9rzecjNwRp8G3vW6oQKTYlBE464wAi3z2NgDC0D6ROT882Wwz2W
SrZwdudAjF4kaXSdIw3P6rQ3OxixP4r0kMdoOXp/g7K1FQV44w2OL93rGGzZVe1+
wqiJ7cWMM3jaJZPpfd6hzZ7NnJUT2qfo6XFypfGlY80xy8JB3dXdQgWShgSiwGE4
BwSj6VYtX7+DYgp4XU7GvQSEnt0wgBQPdDfaF27faVOf3AaZHiDKDrry/0n7tR0P
vAH7J4uMb0i+/8VDsuJCzpD/pWFJw6jNjaZtYDGQU4zguC+KKH7aaBPn2lxggNJc
OesgrbSDRvxH3GvKvHjZqjhDii7H1eG+B/tks4Omg2Zp2bZ6nLby1Go0jEHwLsj+
BEuLnw+bMwe/WsBI85vivl3b/uyDn0BAH0n1QIIHoNLtpcmUH4Xlq8gGnmLtuG3O
w4vUcBb3ps563Pv8U2gTJO5p5veHXBGWED4C70heoeMpHET+TdsWMt1+4+fBEFvk
62jr6O2mC46nCGIlG92+TMyJLGnNgAratVifG/Ale2HA5zlvsm9qFq3IJwxQW53V
ci8wvRnYPLFevSCBCnD7o9Ck10NGyitF2+Ta82VPxSNuT2eGhlhIE2SBZDIsQXBj
KHcK6i1x74iWc0hg9P9gSzQc1loaKD13ZDIZFxhhrevHo8oJd6pPm9oFEjzIrEtV
yYCGB3rY5PseLyCilhSWGqPDSbMR+weymhKG+c+jtzz4IX1jssaXyVVxG8XlKwRX
MbpbUrWLgFJM+HCoaDoW+clZftyPr3+JdmhecP+hxafxMRExdqk20Nt8LJrB5B/a
UaOk+kQOc8sd9t9Xgtsu9YSmUeKYyy3TscXlwfNkvMzhtCyMcz4PkdhjFFYnijYF
cV79EWPlScjrhT/74CZ4Yx4lfRBdLgknnehWxtS3O8LRaSEG0Vyu0FrTJ9CzcbLl
WLmfpaRwxm237VXZrYxHEVKDzV4ASgOS589lIxSqMd+NQq5BNOYEN61W0PEA/2pI
pB76HO15gK46kyvrODnK382KMqJbWTsl6cBPVeyraRSj58JrLn5EQXPGjb/02bJa
a1juoIAerkNd1HqClzV9q4h+ScR/pIBh25OSbWTaEmACqeN1MFVmuXHXbg+1sKUP
3C86SOucSlHZOMBZgSc6rF1AXs/I8790eXwoqp2jmV0JGskxAGjtkplGqPAfsgJ/
PNxbTymOpz9Eyh9t/4GTQaKpDcmpZyDNe8KcAR4bvpJ5Lhb2x7H4V83HGNWz0206
gWNvv/bOfadN7vhUix8TraNg618x+XUsqMnR7JNW4aww5ty5bx/o/RHqX7w5tcGQ
sbxmNNZAwjFwLQJzFcu7JqtCUbrTnMAPj7Diw6ikIOadBvpPxoMOGfbkU4pTzg2p
SXGT8zb47crwtLHzSI/s/s78PH5vnG0T+08i20pVGvy0MGWWkmFEUxnMAw1S0vae
BLtF78JJq6bBiG54T6W1qSMe+fiCt2cOR8ZB2FY7eRGEqRZcp3AS1CgjPaOkKsP7
lGp6d9XYiEF1w8TBM6FpmkE0ClUaJ7Hjd20Xzy+hM3peeyoEeIP6sjpr6GUVqYw/
14UH08xHucgNAIvshr2HBKM4PJrqkyt5RHwzFL34HOIEJ+b6sEwiXiBthMeGDVOZ
KNjCfZm8mVVzpFDlgBCdxC1gKYVmneUIlpl+sjseu0UoikpKlwnof/Rbwszin21p
TyEKgrj+d6Jh2WmWRUkOwEaGyuRk0n7lA01Klb3cGKyX6aSaHvmSrHRDrupj/yWl
AWq1RK6ddCVIZ+f1pVKqVI7X2tA1aC4zMtEmOiSP7w/rlJSSf8auPUu2HY68/KyG
gkF97gDnEY280okjP0bFevE41AAeCrxsxtuj0dXQgOxRgbNOVUXBc9SMrAv6lcvt
c+AXniGxpjUGnw1cQJKq31cYghkctTu1D4PqN0yW+AISVn2pmrkjT/YqRA/BpK0J
84uBEj6STK5AXcJ0HswxwJrTNALWj5XiE+Y8iqYQtwASmZ/WQrID4NiaDwv+swDv
Akt9a0r0xnZ7X47JXLAKDsAVG85NFT+DRaScEvTi9LPUV3r82Wt2uZS4EKGn8YCa
IdY7NS7TZMlOnuVM44xuTVMmMkZSapKoys0nPdBtTZ3MLS7/nFCcWE+UkiN6IgcM
miqd2KWsnFOICE7Y2NXFfSAU0MuE0ePugr3PBkW+UMTfamamktNWWWTYGxzwb07f
+8EDhRLK5WbAg1SgIWGtLR5SYYRNF3aeUk3LNmqPk+7sFD34nenb7TmzIDPxJIYH
xjAHpeZmwdqJICcPNns8Gpi0uvj2F8Z057OAJ6Adf2orHOLLGE2Jcc+dQ/LlHwEb
OvYtkWdvkyQOrojBi6r60E1/tu0494Aa/OAhV17wdgzYI6cwOKypzogH2GM2RE6/
eWEkwrqA8rQZjo8GvNOu96UoOMWnZ6ls/GH/mgoTauo4kC801i465qjqxMo48Xn4
PwPj38rPlUAx3MQz3DDTOupAjidGTTSehcnJAKHxqrgsK4Jfpb1+Pr6Wly7RBNe6
tWS6Fzzstn3OJB51lIJPZTFx7nE0X96oYJ71Svs7icHEmpUv2sTNpy9tUa9FPg2B
1L7+smc6pNBHLO1cc41qAEGuRAQyV6PPhMgILCLIw/RsI1DpSTfmbidBhVsaH2rY
FB+Eja6JPEmf8qjly1WbKhpEQVnm7e/nQz7V4VWmHBNH+roVYzi8Shy6lm8PdSkZ
pGpZ1n6UykVNXIbz1OmMFJowveHgeDtfcEyYikysp66bXHjhp74YPbcPkHgoS53L
gIcc6i+NXP3bOJtsC+1ptCAbguq4idT+sGgMeX3HdsQyopFAVa5menFtp/y+hxfn
IbBlEYAORqFKssVJIMf4ctVplFhGge4HXejLM/+G/xmOfNd8hfJLrS5ri8sm+Ffm
Id2SIKMctvNgHAyasaAWu8P2A3s64cOxIFuqgXC9eNfu5yHFZobzhgZY3RuUGgH0
ZStIkNi3tMLu165QqYNa6JPokSBOvi98M9ze5WRPkNTeWoz6SkaMi80OAG1+aZ3C
AZRTfd2hpXq/DEN7zapJ2jUU2viRF1yCQHqDJRDq3yFwwiEcN+AlF5LtbPSn80iJ
cJFMBPQ97Me6FaCSQsVzTJLiIYpr+uOybOZsjZFDgrs7Xqxnfs5sJuUOi2eR6WOR
tSOFzQvl9I/QL60WS7QiqPEg1HF2tbVbr2bA4L0DWphZga5055VVi49sYslE4bGx
8tESGfVHqiQ4I7jfH1Zgv08UGHtRsaOutQYLfTbiiHXLkIB8U78A7iLRSejhXALb
3AAESCVOr1+8zuumFimd0PIs+pUasEUV4SIxIrX9M37DGP0md5UdXf6qK5dUy0pk
AgWz+qNItF/A2bWOJmosa4UUJWTjPDgiERalk6LqXFHfhzDew/yxagXfCgk7N9z9
5/uiY9+3dZVsgszU53RQNX85g5o5XMyYoDc1ChYibir3RiOtpPdgr+nVaKGcXakZ
q4uZFc+iN9dkyRgVNLx5l3NidpOY3EDXtj8p8oq7AyA1naohDB2j6snWcMkK6cMU
O+mhRvU3U233xJPKqZM+/vzQXtrkmcLqbE4lNBGAozPIiIJnvN6WaNeA2Qp3po9g
Djn+EfDP+js2fLprv3xWTwkqp1hwYqWEAocO1uaXN3BGDWnYbt9XmUVLU1KIhOc4
RkKaPPZNiNz3ChZA0J0bbFDeSIX6chjbRiwFB8XzX8OuopSOIxd7oSZMrhpYvUu4
wZJ6E1nA5+kbD9+tVoix9tHfjJdKyAy+/EuMTQtC9cgNZ02AhJwfbQL3am6cIUX+
GU8Oj1+sdpHoZV8UIbYprmy1XmM1KHnaKp9zbCDScJjc6dksg7iymCwCfcbFGhSZ
r7gqlVJpB0HI8cL8XvlZpg4KKpRN6tbtqCQfRUbKlsbeFFzrdZ8US6tlxfYAlI25
+Rl6fOMcb4Df8sLgKaXwSja4JG1U4J499hky4DssVu0DDtGCf5SYZ/6P4yjmv2/J
h2fe7BtMf7UxoheSdfmAXcMFTO755ZF/OANnnwilZkLsVW7BP1MSlIVianlB61nu
kVaoBc75MrTv8G3urF8C6Bxjj50FfiH51IIetUyiLx34YciiaMXnbt7KrMgacite
IeDutelx3yVljYWRpCXu1FyYSj8i5T+H61nc4qTiDUyDguoFi3pCL3bZPeWXNmdU
FFauYUwH3LvfgcICfwYvvezGOBBws7PnC3WeeTXn4nNr0/J1SPS1iZGfVYuks/e5
bRUJEFKIDxgdsr32AUG3VzS2YO9mKrlqQ1wNhb/KmoSavgiHqFQzhluvFXShYjeX
NmFK9vK3G5IgrasQiLn7vs1b4qra/mn/mLWI66S3Kgs49ZcJ+ulZXhi7bQzaaxYI
J9fvvwarGCXyDZCA5vz/BlNm453uyafgJ8AOtt1OlE6VDPelgE2LZ91QcgBqoRZU
2NkxUAcCBigvgCazPDkVBuZG5EvSWQ3rTTvRUYuCuBCADT5oMkzwqp2u/Kt5VSyg
KMyMNU+Vw4XiYS2ylpmsQ0doODudcu6CO7HtwoX67t5aRnaSq/aMmY1rvQ+qRLGE
II5cwoD1vRE7kG9ihmIrpRu/ee97Zk+4mxQ0Qx/2zjOVlVfCgNTClSp7C0ZQCAmD
wK5UCYfajaulWxfinKsAe4Usvzn1v2mJDnZe89cxIedAoVDQzSBMWye8uqZ/Ye0Z
12V6ssl2y192RtGCh5IBLWWlQxBKD6t+NttEdovhfcCVmc1Xc9IzT8bRPEylbXE5
Ykndi4wLarEo539RBAQ2F0xF0uUMa8tn1oQOYGZ3poZGEonCG/0D7ylT+gKWW9F5
m1EFmTmmZk4ixJUYyjHo9z8TzbK74qVFkRTPNQau8Jy3d0k4FWlbJTm2/gOUHb9y
IH4FoikZnXedbQLPdFSF/rT+B7doLbi3nWXYTO2r24lm5rYyOHxjOCOjQ6eOcBnk
cwuoF3X8QrVgpIxR1+r/RuB2NB+LdustVE2jbsNwRaZyCxa9+SBXkHxbwNcUZhMZ
LcAil+r3dfFqKy08e9AZFrMFS22TO5DwBeRsW0BXQp9l0ZqmyUvgVhbwy0E1x8J4
Il3Irta8S7lqTVGIV4DeXa2gmhScVEltwzdc7jeyzZr/qhKON3YUoGEFp6fSxu/4
N0/3LnZle0gZyurN6fW2Vt0hdt/Xg/dSaXE6RVfXJC9bmkBy7GVqmtNggzQUOtuI
qIDTWwNZPmD77RXrCPOA/H9s4NgEbaXi39NwQv3gqxXiBD6WoDxwDz/M1NFPyJqt
jrJZp00ZPv5WnmBZN9/r2JEYtf+xhfBzCuNW4zmoyBjxduTRBp6P3NPeG8wVzS4D
bPbmDYc9isCM8h1ujw3JGNCKQVTtWRnh8N6i3i+Tq0Tl0yMPgQ+siKIRu1LX4YcM
vTUvpPoLOML7bAQ9qVg91E5OlBHOWYICQ0dgipU7LEaQh7EDJalYihs/JMcwpebi
TmQ7yTd5feKji41cWUkItdzebVybiNiUjcgLZcuQxCAbjfUmkQfxbu+QErMS9TBH
IULtjo5d8EoucphBvdyujwoXnRbE3DbTlJ/hSA4UtR/r+ziJMRs+MbSxXoelvSPU
o3K/zRWUOfOYzaeaeE69UKsDTNsqWTn4S6KUoNSwF9RuMR9W3EeWd6CgRQJUKt7y
960pSA24ZGDzheBRS2ABpXOdW2rSplkH+tiwrLn/sjijXNL+raFBzSSxYB0KfHZx
s516WT04kqvEmcC8Q/iEiUKW8MmhGJXtXTvA4p4lgZ4PT7zR5qHL82+gkwFfDciD
ua5lUqFtzWXJ/uSfl7WUa7HK0So2Ex4t+Cw/ODCej0NSB6YkcR9CE/r2HVJAzdBT
5KvQhY9GfUBCiRKAjxHcTPlVuaGMsZKSkeubbP0OGvhB6sF0DPRY9SiDr3mpSowy
OEqhdg4Jq7S06D7KzN900C1/XNkriG5f9L07075K0+pY2x6PAZgfEtvoG73Icbtv
VGGr1ys2Qs87KP1hwfOQ+FzWGMFop3oHdnzsW+9x0UybPX/iYbi7LGQFO37x7Fac
qGPTwi3hMZGO5r+2dA2UWUjdhFHDkD0PZPabYW/o3ePPBnqmQ/8uFpx//FdCrkyR
b/VqMwCorvQX0JPcZ/7mIeIIexKpdH/DAl3wO/OB4DhkSM7nSzw+Wpi5MgiuThHs
Uzu1EJ+vRwA65no0ex1FOE8+wZxsbqrq8/I1BWfRkywCYs6LGhF+TSOrpHtROnx8
JTL7Y6BX1l+yOaK0SXaVY8LKnqf2873HzWxHLbQsyWdSk7WifAcI+jNEqliWtxxa
U+S9/x8IxyvIzqqJFabNxTfD8vQiz9Upuq5jp1RpLqltLsEnz+LQfzaNidJ6X5Pa
Xg+lA/CJ2/ffggyeiVuPCN9NOTZD7rXeW/odaQvrODB7smsz3a1e5OG3tS+0DS5Z
xToL6d34IubX+TfTi70zx4vXx0V5oAzvRTn2sP3CD9NAgatENTVms4mSTgvFELrS
53GF+D8qzZsR/FFhsnvjV/CjBAlLHznkQVXtCrWYGzSQ7xG8SVakUKvD/kT7OZYg
+uguBBkJsVzHLTgT2Gmr0gDfJJIplGCA2kKH4ch4IltO14o/zB/9Bdn7GQu65nZb
uWaGHNZJNNoLbEvGWtziWPLdslJugXx4vKRMe3GVe0vErkyfocVkBh4fnsxVCpp8
Ga5j9N36/JTDpIm9mjl9ibmgH5C79OgQrCAeEyZ1VWfmqtOTHRd1L7CMCxV35TUA
82AA2RHtRkG4q/aOH25k6uo88CSna46TbLGdX5wZbO1IdZHvyQwMsHodGSMubwya
nb3KjJjxiX2kmw1qFz0RQK0Q1rFCAdgLBREQb2PHgEQXPLkGipaxKda+Uyukb31p
mzbC6yyyLBJ2O5lmWYYbrh4OiSr6ao9yoP+F+diBMLrfUfFb1IZRNG4D5OV1dLTl
4eYYo/ozS8AZqQPjX9s45cnp7nlsFfaSWy/Z4R7nRhnO43hqMpGUb4LjmSIgsJl1
sZUtfk0qGCVUmNw90u9YsJ9nvIIZ+aIYrf1DfzHIp8ev89g/pHQaT67VIRS8RqI5
tzTiCV+kj/AidHaNU57xzGlTSM5JrOsFhu7+0Wq3Y7FLNydP1KQItjy572Wni3RI
T/9x4i6Fnli8UE5BjWl9rV+v2e0/HzoDkAbJwn5RQyAdI8J2Yz8l0OKx6WJTyNi2
89ZayOeMS+R5aJlJZOoVFBT2tcBzvV0MUCb4Iw/2kV+rDzmoL2goAQT4XeOaezfr
Xz8i0TZq344o867BNfuzRzSheEbRXxernZgEQpqMHIfBwpfjF6GpjJzz2sQUyuCm
moO1SK7bzzP+ZhAAKe5Puu++gJqV0FMUkcpoHOXOuFgh6LEtrvTX7jb3kHHx0o8D
B9CmiY7xfLt9lvgyaeXziyQaTLfEJCLWyJ30pFvff0FlUTcSvs0UG3BusbYxGQdV
3d1N+J7YgMchDs1VMaeFs5quH21+jx13/mDuTgxivA7Ag0K4DbDqrfWr0rR4zITZ
AuamvTX6o2+kp1s5gY+BzgyTTAmDr9G6KGgV9lUnO7XwEgCqmy7qjArQ9A4BvIUC
1wAZO8CSTxqUWQS8yDZAbPifKlJauqGmN1CkH06gZZOlkH+21kwqCI4fR5Gu3qen
vUCzN2upPyze4NT8c6G7Y0f+2/CA2l9fOGwkjGhITo4gPD4Czjm7eEcpIkHjJHOB
5GR7nAodDMgeytTrHKZPiFkheeP30ambqBe3QpUHBtGQYSLKD6PmouV6YREff8h3
QR0qur/+qM9LOkPyd0FAgQXJVNNZjc559ZW/IYUkZVoOqhj6TcINqoyqUkS5ehU8
lh1w77TLbPH7kXEmZwj2W/HdFF2zVOHyxKwupKsItn7d1QmuiNAmaXYlkZJ4+YLr
AEEPBa6KWPro/P6OuxWhGqWWpH2iuKYL4qrS1E2jz0PuFEtuoFGcUmyFBDi1xrzM
p+tkq79bjanrqpZQ770dwTqISvtWS9AF7+niE86D2XLbWwuzuJVLHj2GwKJ8KRvm
XSC+wLa8skcWBecQ3CAE/jDQj79PL+hpjQKuJQr5A+6dVCXy2rBopITnNqNIxe5S
mAQOTQA1yZYJusPGOZq8HOXNuhEEoRW+mMeZOCmk4RxtBmKSO9x7eMnsmHS6WFnw
hQbpeCyDEXFYglhreNVL6TCMJbkKMWaSRR9gnERGBA3aOOB56lp74xwB+iHKLLyk
9BDXlKe5VlKA+VYCOBRdezNqjML7/kMDtD/tqY8YK9GwHQbBh8Lx2WC3z6kFfhMy
Dfrzpqm3AOXrUz1Nu0XP68wF1OjAE7E8oC3Sel/nvpOuuQwnFZscEFLYJq8dmeVh
Tl2CpMfewVBHNCzJbta3YdTeXLlHrbClWyNX8yvonpvEDhMAcDr0vj9loTIFVSq7
EkBg7jpMsyj/kWOcL+pQz07fOLy2BR3KU4kqQLGNiD9KoLCdIghjHOw0tzWQ4lOI
UVmyJq2MSungERw1RsuS8PNzdjcrh2Yh8BK1BT3zodSWE5YhcO+bqiDEtAfrXBrx
W3R6wavLFjWZHRxKo1sgKtmylIhhtibMkxEoGEWA6DbP3wpiyppvxa/8J+9BxcDs
kIVJVeSe1CoVdssJnswnGoEK3qdO6GePpNCaiTbEnN1ATj/t/EAIhXqt827i6Na8
9pCRaN488sM92OLicW3VqhpkTDnslCqIaT4S3jbWxCkYccwvqNezDz8D/FW+AA+J
d3OHfeBZoTvyPs6bZHLIzg1DWxmNY4yQH6AAZwWzDTFu96k25/fJHUVLOYnVbhP0
fGRaWi0pV/BSnOjt5MnNhnbK4RbvSsCPf5TzWUxkyHZSR0rrRWpzpFQllX1RhuGO
MknvEj16j8HA1GDfAV3+d7TzU8URQlGoUkH5RNTxRedNKIxKfHZnNnoyvNn1Pkbr
lf2WFh6fJ5hN+PO6yjUmxjZ9YTgIRG37vkWQL4t5v6Q66mW7Jxh8jkmpe5l40qYm
jk3C8d4rpf6DfAL/3Xc3dXLilUS6d+8b7w8hDfhCYLwXEHCf6PCFA+BDa8IJBDkQ
HT+qxeLpTvYjNL64m9wdAYWzkPBE6MvBfDhFC+iyaU4tY6CPY8mg5OWnoGb8mCjb
arGMlSd+YjmSqJpWrWwMh+IOmi7oU08D9DXf+uKuBr4fvW5fSwTo0uARlIza2T7t
`pragma protect end_protected
