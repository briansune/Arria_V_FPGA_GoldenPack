// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:22 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s3sE+WTNkbjHXvws4OhUqH5NMqeLidC/t3fNZQLLhRwQhVoGxMe7NBPXIfqm1gtk
9HfISYS/B69EKOwKJV6wDkcUP/7MADWmOc/WYHKO/wE5YCVxmw//HFyxR/BFvZce
5GcCMzxbdgCpmXksMHa1zEp2KUxbR8o4rMND3fWiixg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
6vv94+IVo/YLC+nIs/SLucSrHbnul7rFtLAlO2AMkDgFwY8hPXi6CPpVU+U41Pdr
8/mibkBXOL1LHgG2/xoZrPUuDyBOOore4xm2z9LMSuSP6PnbAnt3dmcikvDUacaU
8OtblQlTZrLjQGektesVKSFp4jMMEgtZiMxi5YyIiQkQuZepE4l0HCQ3VSMzMtk8
N3pToQSYJJa5SXUba8FFT6fyD+JzWNEMmhr8lUZ4geQNh53QI6R2K8DUpAn/Pivk
L3Fy0zU9qWcX9q5AQBJQKYGVEMEe0c30KnOJH6KFDuMtkwgSoKUTliy3nM6mxi19
IvOKnCn0rCtrujPFiaRmz8poFC+eJzM0ocfyuK8LjGLY2lAmUIvy5CRghVk9K/uo
phVPRN8SqGS4M7eyuWcxDWU7TIDGiIRRKt1JnCZmAqCWNumrsw0z4XOyG82iwvCe
CxzdpNbZ/LlfMpp6ljlX4l43sPnO9Tkak/kxbRRQqS2GXqOLt1vakxAgZmuRlFLB
x3b5S80FVWVaesBGmpnGpT/kqyZE1Yi7ftVzb7I9EKrFnZq0JBEwJMh61wKFj6Fa
EJ5hiLm7w1JadroDKYskGahcjG+IQNbck9pZamLLxjJjRtlbtQ32Vvp+4gxJdb14
DnxIA2dZ2037npuC01FWPiuxbDsUV4q0fov7zhyp+1tVktn74YWg08R3jySZhuqg
Vw7tynoUAvT8JpQNJgz5dmOIYK5/oVXgE+hoTnbT8QcMiJUhrEE+Rf4nzLHXVnMg
eohOXBGO1YYva3Y2n/WiF54ptPmmte5dRaRSio9HloPUGEOd4Z0NTBztYEvmhpi7
Hkj0N4JahynpPVP8hXkH+uCX7M2Wytd/VRMteLtQit/mZYsyEqLD6NGKfFSlV9Ge
06FRB9MJTiwxDmlvSVB3huGr8NftHLyMeofbgtceQ6BeRxbp0IM9i0QgFSivouN5
zjw6SwaPdPJfFkOWjshPk/RTJl3Pj4sBp2nfRRSXDEMUhl4Cdq4qRbrVkaca8HtB
tIun+8GLWreiLqbHvHhZOfir6w577RC7X3ehlyUNRoJCCK/OrPMPpaRFAknlCVox
ZoLAKgHDp3F0JeOFhrcNF8NM1H8IpF5QtDN1YBZoMNboKoEw5CLJ/kXjZFOLrzCn
DGsAFkoNXMRBnpQQ57ZHZHVUW/Yd77P4SfzlBdqse79x9cfFavaWNTyk8TvD7KPc
yvCaM1/jna17TCijdzjwvj/sIKJVczkCRigwLGtDSH135PR0M+Y3Vkw3xNdWa9rg
/XXJ9lc7O4O9vm+4G056lXYfzRyt0cR8wDkEzyYnxCM82Gx1QTwi2cgyE+QU3z3e
kURhVIBqKTkmde2irRK/T/2Jobq9LJ6jUcVRoA+D85JnVCsoNB2X8GkOSwwMHSzu
nHviVfPTpchTE6qJ/HncTBzSM/UTOMKPCsv9QzrTUqBBglO1o2H4D9R8wyMQbiI/
+uZfaasYng5Y4MlDaj+dfnnv5jzBSGmBspKqTBTKMjClgsJw378kmdBP5ME3MnV4
2u0pHsyRrzZuWHrszypffMPVjWTuF0K5Bv7kwhrm6rVIVcVoQ7iZPOHmm54PxD3T
LCF08Q0y4pVD/IzPm2gn187YXmRsR5wt/JCQottFFtdLI12Mh5Jn7bVLkR20Mnw7
ndXHXIbj36nEk7N3DwJbKREThem8gyMyR8nu94Bm2pQy/RZUlJ2nDj/bYjiBsQfF
VOS1v/za/yqGCMwSd3+EUtvzaoKFU8E9Mj6H5H1qLIIwRRGLKjUy2iLajOxgDsAT
8yY7zSxCrUqZbGi/XD1dMLyaBjrwwWOlg1Z/fBDwU2KFlcDkj/CWlBtlvMpt6t/6
TscvEjBymUD+Fje1imMBIbklV2I724/bMVRQ8PXPIl5IPVLzQarxgDL2tV9dx/xK
D3MXDE1NkJPTnmMa+yHbvp1H6CA/ti7M0DUh4lILMxliKIRkc1SwKHMGqnKRtJ0R
t9x24QTOWzK67hrRhTszrkijlFr56RUsp27ao9Aqr6UOwsKfafQZoCbt1uOmOh3Q
2LpCfz7Hb/dOqmIf6MEm1LwL1BH7VuGo6ORlPr9ML+0Is4Nr3wI1E4SLq7JIoYaf
1J14VjAhPsRKKDE8EJJlnMIO3WUtepf2uMvGjkvpXeXadMC9SBITuCzegUT6eC/G
+8oH483lxhUrXIgVT5BmJ4ISMCkcLlX7zhlTmt1wPhNsh7AWIeL8wHwp7JsGq2Tt
BkHPKaIWDS2lyy/G1ItNTIovYkr05akEKL26NMQa+I3ps5CYGsUcyhZN8yc5JBSK
59hRuKB2RkrNI8SBB17VSHUfhz+nwDGe9UQQe1xSXJcqrr3pOIoJwPRNaJLDEKGa
uv/wCjH8DVBNrw4blPK2NF5se5Novv2G0of1LdUq0YtvLcGzMBlF4G0896ifSjYk
/6HVLX/nC6KlXeXFlyRXGjkzKDg8HTFPWWz0hXx+mtQ0RnGYCcm/eFe+8Rqaq5kN
ARCN18d2gRf3TSlhrIPi0uMQJIMrLbMykhqvw4MIGYhFIdiMoBY6oIqmHJGjoKh2
iaRoOzSIasP2BcXK/NmZexWdyo2FqfatEQEQlgAkMyoIA+tlck9loehc+mwsAaBX
0rSgAdhQnHrMeMdsiSZeMnTWds+oWVSUX+PfDkAM4Qe8E6dKobEvvOQqqirN13pu
iR7pzGkOP1kF4fVvIeRgFAgnw1k+2rXv5rwfUnxrnsm513YmHhYtu42zDxSQsszo
Y8mHeounrT5PUPwEJtRO5ribBDzZBaNejxpCk1IooeSs1A8HxILd0ZN2jDhCvexq
mlFQ5QNMo/H3DbNloN6NkOmfWdAzrSNs9jJ394M+MpCptFlewZqXK55prziPEoy2
974HvtkFfI3EiAgei6E3InUszLlFgaWnokptB945XPxRzVZOfqG+uK4/DwomjORA
t4NPNu9OEiT5oTyIv06arvPcxetXM6QnuDOzJqegCkOqip4nvTYCxnSQKxjC+9sh
vkppUgaAbPOKk4cIAqNnY95O0H+SbVuahyA9C63UoBwMBi9fDsVbMeQjEDACnpMi
9HhGvn1pxNsu2oxAMv6BWcyI5hBkBufwahg8CKdvyh0fRdUF/7aNcjaYWHfJIi45
KFZnj2Fi6toVPcKVYzbc+6YA6UBZh0A0jTP9kD5Ks37NeSefYJtnjTUBQyLV83oe
7Q9S9wDgrnUHp7CCw0ZQonaEZ6up1X0thsTGg/zdUsXnXRmBrYb7gJecrmZAUJq0
c4VWlKj90SpyasR288T9qpUM35iDGKGVlKgqZu/2AftCtbONuHThg7G999cBDdcX
XunVyZRIxt4//7HboMIIWCir65QlMNoEV0etRjtu8KhlXskUQ71SZhKB+urH2FDT
/iQ2eWpIiiDhZPiqsmktXq5SteccSAqPPBlbk1cXh3DoVtn2/wQPrs3seFDYdCY+
7/SHiBITl20xQ6rwajO55Y3aAvvST3p7DwfED0mA9fRaZWQk0uY2M1agok9tPN3P
igsPPKdiHzuhy7mx+4w3dH2PxtLJP7JBtG4wcAoUse2XUKUCwQ8haGo1YX6wiYD9
B99trUbvrAthjnJpoqGzXN6rMxhXF20wFgj66PGb3E03gTaebbCF1SdU2ZgCX0pp
PgEWshNqFDtqQKY59yCkFEdgkV80SPwC0O62b31JbFRLQZ/jktp1Y3hHUFAFNwpg
eC3tWgsdZHy2DSecELUU6ogNDgMMoATT/4BbfEfLbptObgg592ESebitz4lYzt/u
Qo8ow5SxnMWM2zZXgaHa31Npi0s8h/aXUYA5Me4i+QnR9rodF6/K9HQqdGutrd69
KE7n7DCPHJfSxmJNJ9cpjohjPdKB/et3GW7p0RGOOYOBvff+HrfCJoYiFKMl2pGb
aP6MtVH+jBckzkq+70LznkllzD6p6RE6I74y9A9sD7K5bQjpZySLd38LSoVZQQUY
g7AQXv3iDzWoftmASD/tkGrK6DWNzfmq5aiHuzIj5gX5XRkRNoNoIlQbeHqbR/Bg
JfzJrSJsgAmXvLqyTNpL+rwiCRJBHczZIkM8XNJIUAm0zBkv9BujGCoGD1HvC4q7
/qbDE/pZvwrNsRNK4ZwdVHfrClrTm+s1fCFtO7g+4mTvcJSifGU0gEV74ezZdPSS
1nVM/o6ghuKPZME4mlqST7LvFRYaWvChbh+7J8mJN7yWVE+xM91wCjERlhfMEExr
2uz5lBKmSLmKP7SNUi0D6M90R851QRTHZ6kdXLnjpHP6qL5QpuDWqxaqGrYiO7Ph
b7UAtgl7WAhdVp4ePrcDZ3eRdiPwJM7oJpRqXxLShhHGjMTOlTa2OPS8tLfExtpf
yRlj2NKinCQTqKdHmTREXmdjUq/KzaSs9mtcOeZ4M0EqKcpX9m7AsMbXtn0iimVE
6pb8Vl2udU2olOrl8VHvp2L+jDiAhkmYFv2hAuuozcRSZi5fY/qIYZS8tjxBchY9
PAvB5yIqhPddR4qSa3T8lXZShH/0Qkzl+m5K0qkIMvyAwp9XLbybpdi/2U8G550E
MyC8MCptOfMN+DRST18ymfh+LymRyx2fxMFSb9LBOY1wjiUCQ1XSGQ29XIqscRdV
7MLWsh8kFVU6f9I79BtbVgc7CtZndhH6JLV799peCYR0ejg1QoazF2jc6dPwkVcm
kC2Kc4TZvMt4O8Q3R8oYoHJfT/4I/rq1qW+KnV0384sWRgKccTcurHUtix77KJ/a
1yRtVEp6vkBXecx5yPYO81Z6llwn4mCUvg7BdmmoA2Ytse26wfZum+J1KcPpjaBm
rxAvvr7/x0g0X03oVuegRiABV+YakYSbGaF5yTl2f+NchQJjS4vYY9FCNh3fQIgI
2ndQKU8Xyhq23taISdwzayzkG2wvfdsrJNj0Qy4LsYIW7g1c8bRqjhExpGCJFHjj
dnRilLg7/Wd/TH10zqKhWxeQDcyOOyyyEV4iyt1N6y4NCCNwC9bkDUSTMNfjiOej
L3RN5vducXqwX974ie9pS3WIx/NJi+mWImcXZ7eVPIKD52E2DCm+ta7teMz/1xqT
vEWD44QsR4Md1yCPFISx8lb+fgUm05/VDcLv+p+0Ie4HScrUXtkqr8CWcBv6SXeF
Kj3wTLhiPmy7/7fa8HIZEn7pG1KaBqw+im/Sin+aIf9IYIyC+AIEFaarOW/0Cv4h
AfHkCcTwVx6x5VoQ0sjdLw/bqwTMzJynuAxj+djl416181lqvHL7m/SPwMSSwSjK
SQFC2mwWbg8fFXxp0ElVe6H9xOh2ifUeBeWSIc2o+ldvqxm+4bc7cvEoxky/c5i0
eG/Lutx/p7I4CNLjeAxhF6YJcn9ZIPFGF2AJw3RsFSTuCfH7B/zsXOmi4jT5i55V
XyHafUP5vcMInaOG2LOXtIOr4bULy8Ll1oWHoKoUvaQ6x/158/RBpD3QBKreTjf0
uUjhn76OP7RNU0fKT61ghJOFSc/QJFY9RjpdEIRB9mt4o3lX3uFvVYJBRx7NWebA
3iCZYxWS4bYBbudVnOIGR0vWy5Ypl3YCVcpJx5l/H6hLc2T7110EppPuJ+/EmguM
7Q5ncSwye+ZtmxHwOVfaUeo4NRxhI3kFsq41a+KCqYqauhuYvir6Q7h8x76B5rU6
7doMqAJu5fgdsbylve0UJdxT/RbpFXahCKEHPAszzYmF0YA014fba4XPxiBS6gi+
Q875CDM9vYwd6XUrUZe4khqnDWdm2FZg5zpDdQ7Gq/oXv1WmGdpeYNsBgZZs7lZd
kWDOASIC7Go4W/tCvoZK8x/51Iot/dV4TFRNF9QK5zImhZkqgtI8RbD7TCEzfkSk
lPtTA2r9vTh3OsUeHXXYi0wNzI9fgz/IMrlrLl8gYHIxGxmZcnM03iUG3meAdO8M
IP7N3kncTmhaTSqF72FSfSHWLaO1L0j1iVdIaPetJVjBTwVy02kaeHocjQNmeVkY
nP+TW2kDwtUEaYYKhUvYzDxp9+CoX9jh0DIde1+LCXBwMlPf8BvdmN7ibUArPEQm
jcemRcfTGZibeeEj3pMWs7Xfx6MI/TUrw/ikLrCrHyaDJ+TX2XA/6lEhC3Phm5o0
SjJTC7Lu8GXursZ/toqOM1Y/ypzoxZ/lqCdgsbDSX0u0SqmA3azNFZVLcJPhDe4E
mRvy5eqR2zv8qORhJo2yhwZdvTWXl90X9ligS6+0U3NL51Uck9PByTR3uyhn9dYF
fctEliIINkG2u9+Oj2Jop9bASvOuTzZBUAD8aQmd2BTMj/KBYSr9wj9nI419slqo
uvJXPZX4p4u9GMxvweKrZs3+JJbvjF7lNCMJzYr+HM3GdVf+1aj+QxKzIXwFh4Om
ppr/Sh+hKp88lPSw06RmSBN67fUdqvXPxjVKMQFeFO+xvhsv1W3vhrrG9azMbCMJ
ZVsfVyPjlbRVVAG6AlWKlPR+hNb9JNAxAlg48HJANlARv+bzSSJlX3eH91/Kupcj
c/yQtHCzdV45cBtye6TFln5hKYDbMlODpFUbQmn5I3SCid7zIVdCBgFu0+JsKunD
4VGRhlKSPdun6wYVsOYGm16g+nagGp0DJ7sprFVKfTe/Btwep275b71XN/cSZAvd
ht1dm9Cvl4zE9MypKmg+bE4YIYoX32N9iWFEnAojM+Mw3VKwApqbKEEPRSxhEWQq
2i2F4JeCczNQ3mHP6L6JjV4qfzyqw3hHES5Q+9elwiOoxcRWQKiSe1tMYRbV8hb3
tlls72J5TfY6wLrsy1K7W1YpJ2MwxvbjfWMDCXZH4YpFehDfYzyXi/IB/PtKRZbG
i4/V/EhN/8pUBQeO3yzke3i3sS+btinHCH8kXNSf6p0DG38GBx0lS9YHFpo/JO3O
pyHB8GJJCQrT2gMbnEMycm+YyzGlQnsQnDRpUS2NDdcMFYcGyUDvkz2p2Tfm0W3u
hCuwVUa/+j7yFByWxPQnlui79clDsP7HItCz13XeUrR5APWtoJibfkDOiyE26RFn
fXNiaHxEI30Q4sXOsVu/JM8pC7xEeZ4HyYocaFZBqRbiNj13x8H0Ro5ee8ll3jsv
f55JctHXVZR88Omuly3inMAi2RBx4upIFO53fEBD7QQyzg7Bni6LVGPI8vpVIgWN
M1MFFZ2+PLUiZWcYQ9MrFPwzodNma1nzG7GmU3p7BgllDIM3a+j2ioo9E41SGs4q
xOk3w53bMEqeansB5DNATm5Inu8mMfDc8g1pIgoZhDKmVyNN3H4BTQ/HvgnKXMei
bo67a2VZ6/TcYNsSF50OBauUSiXO499iS9zQV+dB2l3aT4ABRWVIfUyx68v/Sady
6C5Lac3O9J3S66UinMvZoUTvE771Zet2D5YHw/vOvGOqO9Hra1TNUiMx22AVh29A
sDZMFfcguNiYWnOPEi+abrha/c4J+/00wawmrtdoPKiDP5gWtMPzRK+V0nrwCFZD
bks/tEpbq7zhopc0tjheIcEnD9zz01BFY0CHGZyC+9jqRIa+PcGltbpZUrs+Nijz
4t0h44bamv01YxTLyKyhEB5fzJYrJcIzPV/ZnGEJifUGOYU2CdBSAmkWM4TIQ5Y0
RlXfkh7KAqfDsFLrToC2exhVR5hb7te+4tx+d2oQ6/DApvTEdykosHrKjXU9N0Cv
AJMiaaxBMi5Slyt3x67SaaUQ0bj2YBelCH5iMupx5R/pCM8FX+Qnuz0OQLPGCCJx
MhXWWReJR2IMn6xiapP4l2EQFLIMWFeVNoGGkj6Vm/ohO/ojAHTXQAaL13lmGHjD
jFe8bVn66rUsDFn0Cxu/rAYrl2EqRQhYvmoArskhLt+SfPrFXFRwoPr6ZDpxbjZL
YYT/3wjSW16OZS2ud8F5oYcsQad171QlNZRLUtbHJrQ9ivq70FaafobjHXdyKh+6
ZOQCLVtNs3UhvUp5AHYZGLYzLh5rwyOEybUawPTGQkbvs8ZnxnURACjEP+GygTWJ
jBNj8UtRu58JRWXkF9svRCDOQdsU2wtdNofXI9K77VZNGv5ovjOSaqFR1LvTPt8g
etAQWO2PqoLzpgksVzIcIhgFhzOvMuu1TiOkIAWfgNaijOzrmh6msqzcqqtPhpD6
gQdLxFakCjlX4mT7ra6CP9UfcoIQPqFEreZaz0MykOx/oWvInkK0OgC9mYRBn6K/
afsW0D49pph0wepRa/AElyeXnqtpum/YibkLkDev8OvQgfSFCrgLG/D0jftPpTUG
lSw51pQ4b+Avr7UbL4KQjLM18FTOpxAAUkINsmYRtNlW7DkOVgZBSIlx824hgtdv
BBuZim21dDJGzcR2hB8G36OxiE9B9Z4CrfNSA6L0Lxm1MEF+1zQcce+4JpX0+w5Q
daU8E27RPT5XvxWxLqOA7RezwcXkxQlc8F0rH3G1owt7dMAm3pVlbkftKEKGwnVm
7cgGstguikKub+G5ZvWrqflwvtvwe1D8jw5FWvH5dIrJb996kqD2sl9ZISoTpwb0
pRUG511hpAvgqF3xiuqoNj0TiaO1lVRId9Fhp9JDiZAjyYP29SWFQ80MUjvsoC9M
hvaWnr/PnbENeAcY2U0oQY13wssWoqOijg7wH4Glb7y4NwuUE72nqbuqunfoRhid
7OdvEBsSGF9isMbQc2kceJbe3gL9eejXFw2V478X0aSnbkjuxgSCvpcJ3ccoEX4J
kCVk136Qe1KIE/UKICd0fA4ztn9kJl9jRTi2OvEIg0RvMFiP2tLwm8u8lSvtvkBq
UxZNIVy3r//e/dvahtOSDPuQw5fMgkpryOAInTvzB9CfGsZT74Z7eQQyvE6DbLdo
dB1fBlhoDOXKNIEWr1vk8luLtfCCcymJ+I0CFcjEo51wOGUAQ8H359LLJ3TC93gS
dU1rvaApM8Kj3xcoZZUZJxdxqUfj7SiL4dEzFzhs0YDAdodRAJGUEz8ZqlHH9U5l
+8D4FyOYeTl9yInIL/UInLfoQIKvwU6MjrSN4Frsq7DnQejpmPc+IqeaKY30k1cs
wj3VNwAlehd++giKqXg4fynhuy8JkUNmNngxHLKnDRWzq7ocAUyXGvNuPC5e0F7J
IedmCR4YI51kTqQ/kQhf4wbhxzSGk2UOJrCKIXEppTTS2AzRx/Xunl2ChL90PFi1
Y1b5ZRg7HAXpE7/NkPyVv/D4/JsjsLRexsmdGsdia3bk4acjwJ941uy+yB4RzIxH
ml5GpTYDiuAZBmy1mkdkWWxB26EScF21aTrwKBzRFqcdd+L19gDwguWnEyFWHC37
xU9LZn2ZvghVgpWkkJuE60j9KFosxF/sDgEO3+slGii+S/i281zYS14SaRhii1oE
CdMhoZTB0N1CVBn3uzYn5rqyVaEGhwwwD1QntZfz8QoGxP36O7U6lBlnHaBoPm8b
tivbeF/yL8HkdWdjoFnOmlOcKLRSGZOkcb3rSXgoEmhPp/qpbmykayBhkF8Ofz/P
C1K5rLGJRPrOdfg/8c3ry0uMHm6rKW0Ph9oNreHcgSVFb0lWziVyYPBL8+5rBF2Q
395S2H3+Orxk1FdU1e1vBLW7VgGGiV0hSMoTmVc5359GE60BK7zqOjNQ/kbuxzvx
6aYFWVjjHd2MIlA7th15ko3TEJekuGepIH6gUP7XdROG9E1YKDFkJqan7KaPYGd1
rWsFLK7XoeZGeTa3TIVIaRNRLH05aDRAQSTOOTwEOVeaoubFhhM8AqEs3/609AtJ
V7HcTZKhjS6XVsEL40DvwVSHmVWzNwYYtT8aA8Gkn3V+kclt67bYyX4lXSGbN75Q
nn09M8tA2VJ5oGa8DW8XA6DLGku+bYOg6fqHXQfD++R5acI2g1JVlDSEBiC/mRA2
2auZ3r2KxZh+KO/FMsXcGWPuA5nv16LvZmuTgq/ZaotlPHxYtvrOWBCuhj1IiN+8
UTNi7FOQz+liqexZOdKPYqH2pBi8K3X19AKay9t3WPKEx6Thf0sVlJTRgNzCH5ek
nh0Rhpg960ct7KdyR15gbT9ejuFQPh42Ak11eEInBDTxwITaqKsJiwvwR9IWCURF
Aa0avNtjEgTdjkZRbuGMfGVQcJ13l9K+42pjdQeYCzHWwtsfTkILWQKQAAEL5UNf
RFHI/GHlY5UJeMaBvfQZ1klfo8Gsq8hrWyny/x7Xvn0OpRXK+krvodhM3YxAdcRG
MOXlyJwyNxz08DeNUtFzTUOP4ogb0yi72pkTNFH5DAjzy+jMC2BXD3H2FR3jmziA
vnKyLYs6gyXBLVsuClD+NsCZENRz0m6AgSx18WcRawyyQwV4M32djO49FVfJ5AQ4
/whiyqM/gWgR5k4PCjxSqCobbHd2by67eiQ6W5TPG1hpiQYJ4a24z5swyJoaSJSw
hpAll1QHc+6b1ukRgv+6aCwfyWrbjowJH6XU8/GDjTa5lzd46fnOFtmlQwSoFBCU
SzVrYvYIanT5pDgv8qp17rtxk5T5CQlF7I8ZLDF0qh1lHLusuuj8MWkYRtsoeo8/
xC0IxlF6qAWhcJCIv19xVJd9QD65WjIyLeDOAJ0wCRUK5n0oSMahcqaw5MPVUz/d
FlBH+TY+qhgqSHbz4v0sCpgKC4VBU6xTWsKjtDSKAAuQsG5UQH2zRcMrWVNqELwM
2Dp/6Z4FhhCfjarr2PS4oFD/WqtBPLHsD2zuCw8yW23ENTzN3xQtwu6HGsUk3niM
4l8KCoWx6Aqv8WLhPDv/Pv1n3zCXm7YW99BPb7q00I6AS9JNxAvBwsAY2u1QbGtX
A2CY1Vpa6RcVEH5o8rxcM6eI3p/T0wXmlxwi3a4aE4yLDWndagwDPIcOdaM0K2we
04cxw9LtoHu1csHzHU9fjQSZOWnGY/P4k4JVwVoIyTGgEu1S0LtdZftNh8dJwC6H
zgzlQLDb+gX53bQISghltURNxl+fmuifOQEhlFDUVak=
`pragma protect end_protected
