// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:25:41 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qh/8hdPE7EBEud/zxsp33K9upK99DIGh/ufR6IZIcf1x9lSE7SpnxFwRkzKdrvWS
B4V/TZDXiLUKka5g+j38anTs9XmEu1PMJE/N5eOyFXbz4BPLL9Cq4ol1FXi55xH+
PHpwg8Y2Xrrh5C6Qn1aYR4lDr1sGqXktZBEHU4rrO/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9136)
NPOIAq6/qdTytJC65OXF9UGTbc8ckmj7e9EzF81KCZJ0F+YKDQirtAaDz7mZUU1E
inQwN8SYRLv1OQX7wiVjipHxZIQAdBbNCabpHKqvoENDhHSxw0V/i7o/RjyjJGf1
jXVypeIijgcIx2V0kwar7+Ane+oC19OVbMuajG/YheHBdxOdo5mw0VeivuAWHKZT
Dth4TScwCnYsgM0rIVhagfYZQW8d6ZOcqupRVeAmV1KTTUfGvHE3Mbhm+fxJfu14
SsUwDdPHrVOBm7nJnPdc/3XmzqoKDs7VFziceb+N2nt+A4yE3KIBrdcGO30lGvWV
VurKuAQR+Y7p6rfKVibzKUNFpCAtB1sINuc/PnRMSmDnZYHfkxFQFF8F3k/Gfa4Z
3YFsmkD//J/LXI33JizRKoRYegZuaDzAHYV5XjZuMB1+cNbkXNlXRXpLCKgYPBeY
DErilW9gxRvUracFy11l2mDjJD4AhLk67mh3UxGlnBbsMLi03LU9P8tT6yFQCd4J
2oYKKPUKzp6riYpwmbaagAUwcp4VswgHQ50liHPhq8QEFBFrDF10oE1azVGj2TbP
+cthfJoGhhIIsHXP+6F72CQtdXgDXu/LJF17pJnI4kSocPmhRvm24U2IhktjwSWE
Ree50zOJbWRqpZPyZOmCkg3NnsuYXZmnXmdWa2qeFXc9ncPX1ypKkPuV4BqkR+ix
LUcjspu5Rzn2HhF2JUXznEo87yprI009chBXsPU6UNENKR1I4lHitr2gb6qU3IDE
IvG4QbWVtCjc1lxCwB3hFQzkT3gQiwZo7/nNLRIEEPkSFdKm/QStsMaqwUwqw2qC
k4HlpkAmg4BI4i5DqW+6eO+X7AgN/I73q8vKg4hBJE6rHIiOOvzy7RT5zcTUA8ww
/49794mnrCtctH4qpWTomvOPI1pZ7v1+ZF0kiqJEiMBatB6OYqXgmw+oSsQnwuZb
TKd+zJiLu+srGoetOLxqrKEKwcTiWhwP3lWfVA7oML/AftnIpEk/h4VKHZW3o8Eo
L9D8nHgNA/bW3MZMNxxtCgovpkbRe7uNOOTt1ayB2c81ZHlRmgVqVHFy/34JIlWJ
DWbih5uKIzTeqI4NBiAKN2jeyytfS2OFr6/7q/qhQvXhqqIIA3B6yPjppRSepZzD
5B0V17x8ka4EDsqsoL2u/6wCIZYq67uDGxrnkZLU0NX7TY8+gdVlDsMy7fH2p5AY
ARXopdkgA9IhA3vyq5agO2wT41oLIEqk/DbyakKTu+AyZ/pSpUJ4kuCKxAE9cbAt
FeLijXMZOTiJRTDRB7PQ+iWAuKocZ6VKgsK5snqIGPU6Ap4eTyCbPPpWC/07xqgu
APs6l2BaFIUvQ1ybSvRsa3DOMc0QyZm1u/gIOWmVEbm8woUNevuEKhthunUUvcVW
8qom51OQSbsqs8OMLhJHuH3u+J3DEpCoWNloIgmIDUnlW2aiv0YiOoBFqjvRAA3h
NoP2Ta/i6KG93LYtwiDqzTpmUvx9SKE4uB12hF7NVSFDqH46JU89wrGqIzK34L6g
J3P6/WQbrlSp9ADATLn39KtBJrUbbJAq5b5aeq25Ieht2GDFMjGAW0IbeWNnduSg
pNRjQUxxVfGofUCk5hWwBY+tntLZpc/mwmRCA0K7cU8InVViphWW6UBwcqEsB2xd
c/UIvOJYFmVZzmx5kFUo/TdXzmjyZycsQdnuwRJLPvp+hZ6MCkL4LAAAcCa03RLg
SiMZQ4dxFRuKf0Hu1DsZzKZHM7asyWlxO72NpIIAqkHL1pXQl4oni1j2QvbFf2Ed
E8kw7KpB7/Txo3ms1/cSnRZzysF6Wgo9xAj/oqbY0gy7Uu64pxycPy90n2vqk7Jq
2jZivervcvxlIifYGDGtREdnojQDiU4cGzOQ/iQelV8Lpk3hrh6abE9cKa/oNmfa
zYUJxxSaD7wZsvtgtCG7Sj5HRQtQzNA4yC/L2OyBqwLfHflQcR5gA8J0FE23z0S8
foTTjt5Pe7KITDsjmX4qx47a+TWh3R3LSfJMpWQpTAdVJD6uNPzIHU/f2V9zpqPb
f+ljEC/06EJOOZQILaVXNUzIlWcD8lVYkPMHbpCndlujlQhi2IhXZfkvqTS3zcvu
Fqs8sOmfPo70VBNxMQ0ZN569xO6mQk/gzNNds+VP0ixXpKVAdLQccRKhVVKSLT9P
ykHBNZof5PlaJQ05cugpDD3LFchi0NgJ8gsqLGQm+EGeFWDGYVX38v/iCGlADOkF
QUZdpgcE5d/B9bo+ZuM3P8nyfcpgyf/PoL1qxsgyLuE/vjQdjoHbKuVKyNnFdSB4
sKLXmsReBhQuimQvzou2bijCT4rLXunNMbJlE+djxiUriKsEEfVsG1HgcnQtGMrl
a4Apek2KWze8q2OTQaAwWHvgann1gQAirsw/SZ09xX3y8v+nh5MGzgJ7yHGDqolS
/C9UHrGaUv8RK18kFJ1mvC7IAP69Zl2FiWSMjAg1/rj+LXkUGh+b3JPkqOIb0Qcl
K+cbP5lFSCIcgUigxcEtG0HPzHwqLJrsBavZZyfuzDo43hzfLupIljIMxhM7X5LM
f9iY83aY0UWBjS5iR06eRuOlB85VQCTcqDmsQp4RiEMTslF1DEVIrwGee9mS0Pej
dJpguuJiR9ldNjfDVrwHSfteFfw1Tb1kB4bjFiNrszzb3pZtNPO4z7M77G2ltrGt
f9LipBfnKc5IsP7ljQaYwZPZSpknj0bc+yccVrWu567rekXEsrNus+yFZbjqU4iD
vXGgSz+EdtoFPzov4eaRMLPDyHZfYlLJvwLGtWhrXLpZnJfm8g+whQXqtKbeqX2K
JuAeio2hE6zrV00r9wSO7UWYiUYDxi54YIMjUXc5ARXVKBQaUrlZUDUm+O6Bcay8
Fi+ZggPQHU8acn1ZYjhaNXYUcapFc2B+8DXjVIc/bESbGwnRZf5SvZR1s52YR0Kw
7TSFaNoO5jL6rO06tfCRItV/SKW2GiIyDPlC1+rYKArxsNaJbXH0dQIDr3yXYPFf
bT06wb1LboCkg6BoXQff5+6A41Ca5bFFiub8GqsZZfUIUqfoTVdIPNmsyG1E4MdJ
/Rkt1Q4TX0d6BfEv2PU6kwJ8R8rB51HEZO8fUBbfuQS7KaPdRzBMjJ84AzTvGG0N
/rKv0s0BzXK6lONh9CsPVFg6/1vWMNTAg8tCX2YdoBB6guclpRymL8pXCR4uApIw
+BMhddH+/Iwg+A77fKdo4fcQPUs0aORRv5+G9MpVp8pEg1wMfNZTUaRxXvH5ygpT
RNBfGfzlIVQk+dDmGuGqHri5Tg00w49Vt9esvS7nUSRdrhntjKeueCph6UMCYGuu
2AAcN25q04ee5CHAS+VxLXgjybqbK7J+a530ZlwjzTTBfJZpYqjjACn4ProEMIDw
mmD56V067nmdm+Inhy/cGJQIbLDdz4HiO28JLR3s5/YyymVIV4SY4Yr9Jlxh5Vep
Wjy2mi0WpxDG9VBQSPwPdnt8JxQMD6xIDfsSNklR/2ikILS10v+P+H1N60eB9wgd
oY78XfLHHr4D37ObhZY7XuieW9lwqPvz/1CWqSQjnWArRpS6X/Qe3EAq4P6S6MBV
JLjPYgK0U9lvjg/cPms/5Jm9hCO7H2n+Zu73c1u5AFh2e2JOuOE6h1FUP8NOeH2W
Po9LqMpZnQSKdxHLuiYIiy+Gh50ecAYxBwI+2PF5/pVwr8G7lXwf1eaRMpGvoBMI
joc3orim6b9GsbfZgQGs2LvgFAB6MWux5jyAu8OjiovHSWmcytk85b9uN2e2uM4h
dQMq6B53h+AbojfWviQqi4UicDn9yNX7v4mUXPJ9XBUl8Eeb8teQ09If5PADxoHN
OZt1x9QMvWjhcw/OSBvQZRq6iAAMJ7bs4g1/+dhuiE6HM2psomkjZKRbAIbCookv
PTXQJ6gdtLPHwHAfqrFzIpdZ3NiPTkousPokhPIbU2QYh4OLJi9newlh9/sio34E
PL95r7fHSc2Ih28DPU8FIDkT1sGvyYnaZx91pgOuHSNTSp9ZfjWKJOisSIwllygN
OrakJdvy/3PXUdhrD4TowzN7CMyBI3AdXnTVaZHKmLVW6tjrt9uqTO4YchGvCGhz
paCJkxRYwvaImtQmU6U3BA5q/Nk2WJX6NankEn+HWIcqdhnl4MFesnpPfwAmPvxj
SNjL1Ex+E7iZuXfup+3gNhi7zZFBHzNcJhCz6tQkYeHPe0YQMtWQME8aG+LXGTOn
UxfkTgDMpmwj7i13h9HHLGPi7UDuckzZzL3ypcEi2+dDC5IUwifCbx3msZQm7SiM
dumQnelWpMvLD9WfST3UW8//RwR7j5C5VmGfV0gF1JtxaXsE9nPskHVI0QcW5Qy8
6RG0LjBo2V63Z/K6cIpLbtA/LGnLrQkVM4CZ+oOEDLQgzY5LgJo2NcTrpizJWIAq
NVjv2J32BqmYNArWcnAlSIHNsUER1NM58tZh69zdayASNRDzJf1gc0ZAUDYgdTvj
lU0P4Z5iDTFw21NOzFt1mgVGjSRKodyj7bF1z8GZkvZiJCV5saKTfecd2eOTjOmR
OOOqToNz20lz+3KakwLzfLKZeQQQFXzxibgJdfjOj+yuFLWRuAZOwTg1QnnjIGI8
7MqsgB6ku/5V64qv+u4PPdF+aKaBgExssTs6ad4xsjDzTy0jHGO7dMEpdSqis6q6
l+uHXffUuYEhtLlsujvj35b8xPWq1oSGVOtKWkejvVovGYF1e+kqPudK54DndS/r
ZEDAR4JeYAOxL9LfKmhvHGUundGjUOWzvHpx6z+FF/ET1q+NhYyCJhb4qpDkc3Gt
wW4UsSH3AhEqt7cSDaDwLoaxBVB147U3/f9UOE2JxMFjAthbHYFGmMxueIXRG6Cj
cApiYrEjxDa9xZItQdggLk9fM3laaoDQBJHfoB8+L5jlvDVeSfq2E5qG9lohx+iP
UQr5KyKaMbgs5TXp0BFiB7yp7i5EvdX+Rb1vL1sjl55hRgcW0GACci0VJys7X+Xj
slUV5FgKT8xKv4X79qaufnobYB7/ssCtxPV/BQr6ss9sa6wPCkkTl66j/mfV8oT4
KdYP7/2gAlomKMSRAFKoJDW7Q/KDm3gsE8I5C1oVA/7C9dJdTraxHB8+qLhHTQZF
mQ7OTDmIG4ZykJhA7K6JZnXLiEaYcUp9hPbF2WbbOQMUOJAwEGjQ8XPwtH/zRBBF
Kk5A1tgJ+lveFjmki12NmzcGBdqFcfeVTI5KQlBQ4hbGg2C8Z3j2jLVKw7fLBYEy
GspQdsCthpnquy20zZeLzUC0/J9ZhcVPO5O4FH/7u4N1AdTMPBGjS/3tf24mt2UK
H2+v/7oN1Ph2H6B4q0k/DzG+SIIPE+/ISShucJwWwJqLnXC42gxOeMoBSWYodfc2
CnERv3e+hYo/pk1WH05N8FKrkegIvAr7dRScS9aJrYtPUUoNlW2h1tipNSacNQ9G
qQLrgcO0iiKu8vDrcqdL0q2idHBbGd5A/9ens/ySztiLW8uZz8+lzaOTqWCIEVZG
pHwIXA0joTB7lbR0llEpLK3h2NqQlPfZr3HKBeC+YKJEHXuE9fpPMwUFWBFFgbqt
YZYvPCzUVl+HMOfiI00EZp2saOKyNiaKraIn2rYrNystnCIcPv+Wo60mgpi2aEYO
CAd+3EsZUpGdacl8lv7I4290ul+YL7wkDXPvUgQBZzQO7Qn9iCQQm93aRRq4rt+k
X/IIAM4ahWdG7aoa7yaSH0+dLumJRf7+hO0/AQ5PWqItzSYKp/Lk80tiC8LXLYz9
xlf+8sBs6hJ6EzEsryoLaRhvMK7tMKYWHPwrCRG6eT76zpsfhl0hQF6cLS+zAWQ2
hPk3SmtamkdPt9ex//9fc4Nv7cCH2AogfDMp9CmW1c8jHwJi014zFhkoH5NHBA8e
7Hx7BkMiMRvb7HOiq+bHVzLcZrSTNPd7CHsfnHVfxl1B4FCe0sv2Hfio7ztwnSEM
dkJMCJNLzpPndTs9IHaST9Qmet8RV7+1iwBQxwWYtX2ybJp+pK/MCYAjvHJ+TFuu
08Xoc/ZWloxUOAJTfyqietsDpSh6HDrXDta3ql1OcaqkMs4tkK0zHIyq0wUkOvjV
TmhSixbbjh5eATJomi6JwkOOeaWuRYlnTu70kVoGHJeoQJZbx8nLz89okVP7Flrm
+ZBTw6pGIXfMuvBETq1NsJGBsWS7HcyH9CT8OPuvqqT/f0ngAw3Zkx/jc54t0Nsy
ARNwDwbL9fXpnyFVCAedL7yJE6VEfcEydhlfueKCjbKOt5ImNXlzUhbhxdgXO/2N
lmSvzUNfDLzXyqR9G1jHNIxG8KFrvTfqWJpLOFO6RJmNQeAO4s2Y/rkgvTdgWyCY
604JnA8W2iGG5QPZsBKl0YewLIhNI0uVUGJV/qcJ1Li8o8I2Hc90fPNd0WCeyq9u
d1t/xeiObIe4YkjvbIcK8BUYgPCYgd1dSGOb+bdYipPxsf+QpyK6q99mwBYEN0DV
iOacgDxBqlGUqTgYgYB7o44QTUPqgxsWNWRLx7FqEei62Dvv5gOSHojGfh5kuRZi
Rz7+i27uV8JOSjoPnEXcHCouJZBS621BYJSFCfby4lBZb2wVbBqAyxRAA7qHFfXt
vImLcJp2PZZ9G3MK3UoFKPywdekABe9j4iziOrsATnY3IWiRwbRYXVaCZ2SpLcRC
A3gTFwwH9gK7YhQyyUCE9GtmQFbxL5wsyPwfboAuT2oBU63RwF2V3dypepO+CQvq
O516qPFSRaxMyEl5o0/mLLD3RePaOnqiMlSY/6T489vv/uFzhNQZ0XErf3SkydX/
YDwYY6OxZE6LhDOpUU/aQ6rPtC6QlL51veLKzSWs3sE5z0/NhYErS5vWld2DqjfL
3os+YIVHKwmVq0ncPfL19ldGYbicOGqu+kXYDDbaBWoW1SGwqGx2IklbzHG5am2+
0ZNgbIjlpurNkvdo0qyiSa0PtVvmEu5up7SQrq43WCqJhA8KFq08Bsivmm3SjQYo
gI9x4OazQCY1yAS12uoul3rrDJmS9hnzZBbXEQ5GaHzSfftR2VNPfC7umslb8lZy
ZP0AifX+yt26vhPfgCcVQ6qERWCAtHI5MxOIVKmqBx73S4/H0a8bdkZFh6AiAF/E
FxOlycC86AoFpNj5fkoO35pV96N/AFyKzvcjew7P35cnoiYSs7EufvzM9v0eW1xf
6X0LTF0fNILF76PzbLPSMlFWxSCp2umLtKcpDezFnmkBIelYw9Q8VKCImQa72kPM
PvgQ+WAbyNG0fxnmX5oZuuQoGSGtSg1TQInPvN3a9ttWaZ23FYZTHNEr+6ZvT19X
6oWH1m6FAOZF/8JVpCoU/l7MxU03F6X6VefQ7sA+uW0H2lKUsXz3J3u3fOyyhcVU
wDIay4hXUOdCSS2CWcIQFfYJYjIh2SpdNn4ult3Y4CrwHMeCE7JlxSk7VfwuWT9z
hgXf+EZ09vI9KSzry0b7onI6ZQo/r6jQFWs8sc09nDVPW+Yj9ftCqEwiFNvpPrT3
NH3kixAPEhGR9omSvYHU7ZGp9SFvO1qFLYQjw4SGc2v6ZXIzpeftKOQLwbSfRFNi
81jVUpZ6bSsrMcrbUji7+KB6acUhgofKBIWSlhkQEj6K6HOThM2UDUUM8gtVF7K6
nGUzCZVIbUpnH/1P10c5QJNjeOKBdWdLuCjEGruJtzGCqjjtvD5x1mR7ICQsrQWW
18+5zZqmTpWdp2xW2BxHmlf2EugAlG+dXmO+Pd7oB+IY0Xcpe76cPs62qYtGcuAC
zbY1il68rEY8s/AK8wy3GeMkg6FQxzOMoCDhCnlG/2LfVwOdY2K7qFFjkb1bEnzG
Lp+uSp/IELPlDlvShEKmiQOXd4aq/2b6JwF01qK+63G5A+ltTe9SLXRLcsW9jjzd
22A0VDEU5SPl/qNAI2bxPFPCyx7GFX9hjgUXq/PKWKnYQj0c/x86yCmqt4NNt9u3
q/JeuBFKP/bLME4rVkS857Q3qe57hF9AHlCWN2RKDtvbwW8zqdw+KI4wQ1OBtEFA
P3I4tQ8a2XTjPkrxS+ONdRF8CnPjeTcAxQIgJ0v/ub8jhfru0Dubg/yIqhNBePJ6
NpF1zYnSZum3kxlqGqQiqK9cLh9GZTIYrfHVvaYscbZiTW7A1LbYOO+JRnylxxh+
KoEn3qQKosR3t7u1pERmRYt+JH2jh3YfzzkxuyuUY1CCd8MVPS60I5Xcp7bL55z8
jCPBfHU6V2Nq81bs/MK3pXDn4546oUKzJfrf/hz3IdXDQuBWCtPksKLLvXOKrIuq
aC3D3MKVXMC8EbH6MQqr1POnE1MTyk/qcDxL51CqMAqzmfier2h5q31S2KaUnjzX
SMEKBiOPfgw38gFHCn7dWXeJrlgQK6kDFeByrJjAy+kYP0T/0IlV53THSPvL18B/
GRi05tYJJCnHjomVayhOfGyIfJlmTtwcJp20d1L008ohGzS/zh1BNCycPl8tUKe4
6NDx8fPYOE/KSVeRqhWHDkqc3IZsrIgNmXTEdyKapgQod6Ht/YW9+boa10bi7mR5
TbSvqPyob4UHi4Anh5CUWYF/ffmnWoklo+8HqPVLbCfHq1uCxQ7rCBYBnQKYE74v
KY2pMohfbbw/L1viJis4uCI54/UmzWFXsE8KKxT/+lkcJD2LjY5jI1rTl6Bsq2a5
oCdvNN/3ktvOQNeZN1EaAxjtEHtA75eTP+DMOP9aw3hYQL4juQ/pbcrvijVVu/Vw
5rsFFZjJglXhQJVqlWjWdLGwj0txueuS8w9hEmbNAMTpu7sDQGI7eyjO7wUj58eI
a2eT0TrmqMOyKy6nPB6LEt5tScJf2LBdLZ2Oxz3Hji4hlZuYfLukZfWPC2yXIa1P
1UIUIPBe3nE1GPqFuwn0NDnJHaKr2WPmqBevBhCmLnQWyf9bFeSHijMMWLBlYRIL
0czGsM1MROF91Qk8kZBHsQdA72HIWnB6Tc4szv8qdMHm93dE4q1wktT1U+fXEUTw
eq8SMUVV2gv+Rg/L8mf4yMPjyIvujsBqn28PBi46Pp8dNSDKGww0LSUs++lKafMX
SZtVZoEGMDz2GjZI8x27GyqNYuvUBrNfxQliTx5cS0zawLkyrTKEwK2zPqaHbp8V
jZ5B2iu04x/TWovA8XPep0r8Mkg+kBTEmr6tT0dS+HwhDRQeQkF7loLs5/AnuUpC
CfM3KrgBtVJJD8LgHXMkvVK4fAepTBPfiD1e8pnIANI/bfAtEztcovjLGXIyfgAZ
3aOxzvTg5WNdAhxh35dRMiMYmOyaSkwB4GOa3qCa/ZHnuRh7DsYUL5cOiGyDRLNA
u6tyH6VWDJXTZkKnlwWMD/oaZ/c7otrW3Kb5GGFNY27pCcX+Oir1z/y8Mknp3Wtb
nQxONDVY0fTY5Us4cGb2hfmj3ZQcboBB82IeBtSg0IENWYdDJZYTJZsc+edJtioA
xxGsnx5W31WNGJ15QkXcg5N95ZhVRlhDXV0UlIojoFToEYCjElhulzDKxVzeP3mC
c8cAgl5wrOb3uKz+N+ehP+0dj2GTKHrQG/oLBaXDPpYwkrynkcu11aVjQlLs7CYC
CK0fc4Cr7i0hyoU571YHZ09cGtLmKTyDmTsR0XGdli/gseN+6j9QadfbS/dVQwT9
b7ku0IYus8kMcdEZiMuTsOQ2Ce6fRY5QIojrhLMQs5FQwRyLwk8xRPWr0OmMjAM7
a/wJrNuMw+hPi5nWvL/FAFbcskTgUA0vKEj1KeXOesbb3vJbtaYl0WYkf1tU6UwX
bpNFrf4yYjXY5hSYgTUBy8nCu48zjSGPRUC1A95BiKNEA6trG1xPLdzVxpJ2yJCh
yyoWRK8qXOLPzJzkM6kFL5Tb9Icpm0VgwJtbswYVH9SqdZUHONfbdj7tLuI2D3Fp
gg+f0w2+XyqfjzAfH4spXgLQu3TddLerlxdw70ZmjZNgT+F80iYjdv5oYMsGhb26
YzZGWUj8M+MuAtqMkD2eXmbcoNz4uQmUHJCvUunpKHF7S64t+tISS+qy2b372NoD
XOhShm6VjD47fyptCjo/LEXhm8ld8s/sRTXvDkuPSq3k7UOPUymRVzTzNZmdkgMm
3awqET4n2b3UJaOPAuTljBWQKN0Vj7mLOeR1Lppu3N1BzsDMVUq4n492i0wq6Rt1
1jyulWccNtMWRf5JvlI0szmlc8rfoCmUGxwx8HuqbJqZrg8GmK43uVuqwZK7lQNe
BS4GgmgpiGWChzArhyBds7wdyP1aZqHFp3R4kdLzsYex7X1LMbfiLnhGUV+w+itt
8Z423psZnEqHpKLl0rZbH+a+2pXpb1npqbZ7eJOEywFfMqS38wl+tmY6NY8z9heZ
LcZdJd8BO7IrLQvDtVaSKFqp2l4nXtZocbDUAyCi0whSloTgvQf3OLsroSx3thwd
wxwkrn8vxQAIJ1r7zhRPDBMvxgwZv/RgLF0s3WAIrtZGs2h28GFK33NNlkzy2egM
B6QahwveyI00T8szPGeG6EqFP+IAk6foFbYde//GE7fJSV5Z+67+dlVhRXk78Hxq
y+QT1anOHIVXkqVgnaeOWMa0HdG4bK2Lkrj2G+d8Xze9jRIeHn5UD1MNovH/vdCe
+oL2Mfv5fJImcRWVkz9jzg5oCalC10CxFS+KlR9FmtEEmYoDec+N95uLAeqaphIX
5I6oOAo3JZH70ItP2yBtXjGF6ukQ/4b8F9arZwDyunb+rIlpnarZj0uv5s/WSon8
QEEYZacC2otW6I23rfRC69IIEyfhCtU2ziBs48dHQBMUJIxvIeG74aFNR1dF/aPU
gLpxv9CnKwdaPuec9Mi7X7eBYDVxzkruiaVwayfU2fshKTt8a7Z9RIhEye5iHfAO
HjMFw0qwd3SbRA3Emb3GY8JUOeA5Kf2oi2TKwNd32oBjn4iYetTVpF8/M4PpJQoU
A7xxUBHgbSClsok9qdaOuBb23xTyetIVu104C3XiqdrQMcU3i6KimaaPInW5T2ZL
IGGH5l6Ion1/ClsUX2856gL0Qx1FHzzy8A4o4ZdJwEfoBZ2EPauUg90tWmdWjR/3
jKEe2GXV1AN03KKIQNURyEg6t/vDfi557hcXkcevy7ormgm6Pv4Ffyr0e1t5bzJo
paoEl+3WthZdFOsHXQmI0/kLYyLeMv/GuAbWmlMKsF0E5YpJfzswLgEBqG1MEJz5
Z8qlPPV1PVuaU9ppmrWj56z/aVx5zzL35s+VbKGb8jQBbY//cPnxsCY4AgO37Bci
dp3j0szIJfmzPmWSoCR6Q0VJdhC7/aLs/soTN9fYyDo6C/+/I7W/KgmhI0vkuymn
cT5YCNkyeZE9fIirQHjJlPHW1Lg+ZCwv07voEWi5oZK5qE3dae4sS64pqw3BOs6Z
zZZNGH2LmW7QPNMwectE2Ii+wQAaOASTM+fv27/9QjJ05dvUW/45w3GwsKOJrz9E
JBh4r8iAy/0sZHy7jM3gA67YBfyHwmm9WHfkR8FsoN3LZKy7PCOEoL+iH40DROkd
eKVZm5Ts2TF8Q+sHd0HkWwEulZhjNOSazjhqTRut/eNeXWxfFXS4AFuSivrXSLdl
3bbkSmJ9R3G30hlUTanY/pmFEXw2a9lxA19c5MR+kmdRMSFckL7iCEpmOWGLKe2k
dr1PD8YvISFil/YWm3k7Q2edB3IPq1/5hY2uKzVIdlMAHmNji3jhIRNL0MWm2X2i
6v+Ydk3JKXhJWtkgWQ3m2BHp0HYjUfrZUVX9p/5b36Q91OWMAo0T5tYqfD1UkQXm
rdy/mFNCRXosXmsvEThKt5r+4scebC54qQ4+l9bqWJwpdLluSUSR+g0v9lIOCDiE
b09lyRD+ReygwzRQpnHbhHLJ6j4j25mWQmz1JAODen5jyXU9yIuMcC0kyktK9d8m
q0QbKZUVHCQU4s+2NSzA5ylltkJ938D5hkceX7ynEFKRslnaX9Ao0WUpCAHag/br
0iSMN8DqHBp57Gt4kw0qtaIYA9GZqwHTlkad1N0UttEEmXL5GPgF+iEFencwlxj0
VetbhZ8h4lYd0V9O7oa0/riMTSl7OVB1VTGjyM0SK4fc79z24tjSLhGgrXxCn7nN
PajymPJG1DH5PeLoybpok9botQloXS2GKOLBFcKh68e+QZK3yjx8c38eVTyJwKNz
OaqTTiCXTY6bcIiUwhOyjNjQ1MVm1X1h5+NRq2hxdOALohcsoko238foxjRz+Je0
6RQu1tZZepBFwn0bxfBaJw==
`pragma protect end_protected
