// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:26 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kMBZ9qhssYg0Ko9drT74XjxxJzFfT40/7eiTjucDz/C+qhYuOSTWj6+tHP8wOfXr
Q59ZzAqqDrTp2IDjBBTjifh3kJNtH07FT+w7N/GuuRqjD0gSBjif4otlbd+89OIS
t3a98QRlyvkDEExEg8P9dZAfSaE+/2w1khkUBlV8BIs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57744)
8Fzn/yUjWrujO2w7PwJGtNfVFPju6CT8sLJIGwrGXYXuaidDS2lBaxZzVmwFrXjc
BrTipfbaGrPt9mXyXuGmNIrVuKBfj54o46nqSkY433NxNYbIO6PYM0ZEV1kykv1r
RTSYEowgnEzZ0oYTUM0I724cPygeUiPd0cMCrHW8M0DaG0YZOyOJidCCriLLaBc+
3guKXOcdABmYgFWxrTAn/wSPOSc0cgxh2u2YPdFeGaUHxDKKGUQlggYrzMbBs3NY
xmsaLWl/d5ekIsy9if5G/TyXp/g17WnwX3zjiQRWu8Z5mYKvhrKQ0r81q34J55yk
m+9of1/ma+jjHJZUwYPqqvhnE+Gof254yt5ZvswqEGhSvFsCaUv1ZAmN23Fl2P4b
jCUDzVYJwtkKllxAXkfmQ6WKR6q6dtmi2d2avL2PdTO/qx4M+IHshHEj+wow9XE1
kW1K2r5yidazfyNJfx8pwGnTvEaAjx1SwzusmSK18lIJAKRkDsmD3KxgG0xIBLmP
VuH8fwWFuGbtXA8GzA+cy3pLulYVNx3ouFZyKbQFTBYPBZZiK+Zic/D6Hte91DM5
Rsyy5h20SEDrxtk7KpRP5VL0KEk0iTiiG5Ixt9ym3XN4NV1hcVO+edYVzKq8IL6X
lX2IWRKe7R2hwT5xa1kb2BXIFF2QloX3KHNpLhtJPTcl/EoVvhYeARoBsgpn+yL+
HiLBxRcUw5IMEmgmRB5ZD96HdJU+HMLBjxCJwCUUOWGiOsaE3tw9Y+hrKfR7wL+W
H0ygNtf0R0taJNs1vPpsbnOjnpSco77OnpCsZTQ9f3ZU8JYCdY1agz0agoWy5A1S
+i+s3cyrRQTwEHAyEvN5DGZeAzkusQZ28/Zr1gPBHu31Syk4fugq95kMRx4iZJem
6sWtuRma37jNNeM2eBvtyYuDhCSN/mTRItfRnENiRSe+jYWSLmvJpR4H9gSJec4S
phV5Y/StmTRSLQtjyOZgBlBM9GS9vg4JBnyfqrACVpFdij90SBmaVX/fb2HK+vHt
ofOA4+m/LLgfDZ+CLcprswp/o5IrUw9VtVDznQ8RMwt7fu5QH+CNDvNocj0FxqeU
CVG2JJQoFNyIyS0iGYKKjTfSztZH7Q3Avqg3ztiXV+fCG5yljXRn0zrvmfxGq0cO
zZOyxGt9zXFp/8TvLVnTLox5CtbOXsEE1YwiDZlSxVzW+HbcVS7yGmy0zb7UEdbb
YbP30Pu16Ay1PXWdMr6OBAbVQjmOjGEgDvCh+5XF2MFjPTvKqiXo49aYxGOizUAm
hVfiaUyQDZSPBCY4LP3+USmpZKRru8Xs32iqzHa+PnRnoDZIYPJbeb8uv04aJU5d
YtW5mIgbX2QMyDc1m7nZ+/Q3xLShqLPU8+edHqQFT4yWNIt1abrFsMh3GK/rElGY
Y3NJw3sYudlA5q6MQ8qgj19NTH9MEy87hTqCRwZ8UUyra7Zy+LVoKcDdNG0e9jdD
m+A+D1ckZlWKMrey83q5iHLD7Mg33oyOiffTq7aOVJzr85w9hCgwYuRXx8GseBuj
cC4IfcPPWOpJyvT/IAIP3qvPeF14jig+LWIFdU4oQsz5SUE9ULp2ZuqA+/EJPSb0
xyGCfCTOn2w9T+9JOX6628kRe7Qk0oH0Kcr0og/X84UQG39JBtYKQ3skK0fiiL8r
V9d4NNNr7xRtgdBMnMKVXBaUUzWzebBWeBX6FLcOgAAIJB/eCJ7HXofHJisdZGIS
1sdwptPW0uHExFvh1QDLUShh/hEwd8dJGOHtynicP3HX4W34EQOaG6X1UzXQbW98
L1LsTybkn4eyL24X0zL5svJSMrp8iFvFyE68b/PVcPtVbFohwABfNAjmqWzUt5Gq
vzMfuW1v/KokxqpSTRtFZSgh0NQfxzwki3/2EZAAxyo3HQqcFSh0TwcT0m2v14L8
hVzg4f534c1XoyBgUIbEopUm6TQyfM7z3EowcnbGsBLaprlTYkGgATsj9tXM/WPL
J4tRrnaCdUC0G8coGAbrPDguzBrDmex5YhXR8TE1gT5WedvX45p86ReSCJM0vFpi
oNf237F7KbJI27LfxHr81VWwLfkq4sVd8mYijUTsHjwjrtzYeZaIHurg37un+o9o
0P+UA4Fb4nRXPixijSEx2DH8lTe1KLIZbDhnVN4XvjNFda4SksYCOzhVYoWnhLRO
xhXW2rT1ZriOh4cjZjB3WzbOZZmTbaeLGBEgZWsMcZ8hspeWuxahxsfOwdRjTAjU
/o28JQRRACc8v7T2cR1A4mjNd/9+r8Q8S/V1YFnHksEKDh628VutYSB6SafteTdx
OhEbhtbQSDf8u7ZVPDUheNlnzCteuig15itw72hU6kdSies2ZW1+ligljUy4PfTD
lF0zVx80rbcrVhYCAUqFcArOy8KExZoZPtrYr85HdzpDXhqP9t6zxT9oJ3e8bCml
PfVKufN9mx6tPbFw09yoCz6RSDsBr/qKBP0EoDM6meUrwT/xKuPSAgnt5mxoFiIO
2sB18jvMttAY1lp7PfaHhzmtO0SrQ/AzhLwx8KHAE8WqI3hKFOygwxF7PsIxRteE
RxNqI64Gh/1VZ01UmujdEuET9MUMJVkxbg0nvATpRs+sinusCDqN4SHrM6TfE5YJ
W4OBmirAaKym/afmHsqkfFjX1DqqsZ8eJksbHrqQNmANkRJJExx1A8P0KpXAM1To
0OAHo7aWT/GUtsGGUwSvPkd7q1TtWtJSICdtyyniN86ma7Xy5gAv4SqLASqNMt/s
BoWt1AJH2OZ7yzfjiacLJBn67SPZOBtMYjkOZwwMA8kOh2inO/gwgKYQmYcqxvKY
9mtgAgFAbMH0PpmAbwukTzZhlLWHhxylZ2sqmn0PzCmoIxbnSTRlxnjNfg624+RW
lc7P3UZGKk8c2WLFUbLmWcCLRfohqJxx2yHdzt4obxftvi/Ii5HKLg/dmXNipNL+
kvjHmiAYFA3vdo9NYhv48rtYGNTlCgF91h60uEd6xlatmtiUR+7eSYDosQdqLp6i
YR19/wpLNLwHohDeIZi9O4BjLRKqcvaKZp2sMYCRBdHYLokbJ9R6kodo2P2QT4k4
kDWo1LpwyVub+RuH8yNZuQMyFvaUAaWz1jGmmFOZY90qehvgSAOT247OyhqFpVHW
MxzUMoXYQaLgrFYsm8fCx4iseHyROULlk7eIHiXnNfD6m/3AnpLbdtUKiGzsJU4e
3XhrdpPEG/JyUPsbc4TjCAmFVki/pwFxYI9OsURsgAZEnHQa+BHxWs3IrlH0X/V3
KZLq7vEG8zkyusILwvNP53nUEr4Cfb6kN4UF3He0RFSYr9b9XSJ4nF3XIuIqPXwy
kJ7x42BFnSysMSJhdu2hoR8dsFdD38hNgFcPuIP8/Vr3RoifRLcMMK/7PHwjNeuo
42s4yHWU8mCIP494aNdsVx7Xs5PHZImELTjpBrogr1Sx4ialQax+mbIlANeCdoKw
wfTDcrMuag3BuhTcDmWKYC1YZgOc/Cl7wvQtcbwgRgIVVMQRiDLQbjjdAeQ2KAwS
7RV1XsDvcCbHf63S9lovy4AnBW735jcvsTvOVtuBAWtOXdAzvDf/qMKbxHj61l8B
6Vv54Ae1LOvf8x9YOv4Sad53cJAI7KFjgEO4qmtdkUeZv0BOg0D8/EZGgn51aAFJ
BbfhYxAbz7LjULOltwpJQpT2xtyBY5rni7k1IMNh+gshUlhl8Me5Tx7zyDmnlYuZ
qe1E+n17+o9mCEM4Om1QQZEDtjcIprhlPRIvE6fKEO7vmykoQb/r0hoq3xXfMc/Q
9iQ3lrfwb8ckUfnNDZOs0rXgvO+2IO/MflwFYf+CTyRSUkSBqqso9497KKdY0Xth
8dLeZCKL2YKdr1mGgDWKiaH0wdVNZFA0h7B1KwPh8tiB18xpI3Zu7dNdJCsjCr1V
g/pBq6Y08NkZRD8ffSWtpkUaysqFWUkWGP7G124j4wdhC51K+UpTnDL8LhI+W2lT
9a96P8QYeSB1k8TMiF0j5Yt/uZ/Epcw5+KcqwIS3SCGCL+07q5Uk4o8U8bClHMBB
4wOKslWwPLuVtNaBRdmUaAi3yRZMwKYQXf+Yo2LrDo1ieE1qgCaJIlbjVk8gRuDw
Q2d8ePDm2UmovxVSBp22XoSLyVjpUGGlFrTa7Uo8Aef9mXD58gKm9NQHGh1p8KgH
QSKQSp2/ZoDAGfS/KotEsn+ITAbUsOyJmGm4Gb0CkcmvgfrTAumoQ0eUXGx9I887
5agTFRplkyfVSplp25fJqIhqzQ/VbQzaPfeCq8A8/vWumtBvhooHE+OXMMjX1oAB
fCHkHzpNHM0A/2xVA/gYVtBKyY7NAfwQmulX5Jttt0FO4QZ+3Y6fNZypYezSRYNG
GQk33e9A4QO4liuOlvaNX6TvCSTStAdNfZ1PoW5ZMl4uVNObb6dqDdtThnufluP0
l9IJ/M9c80E42ORD4DUhswy2bCwr/RuDi8cHKtCiy0DiP64c4L1Fqpf7jT4kBnoI
6b3GhLkhzDhwW6UR5PZ03Cbiahz4FjxPwy85vzVZk+aXGh6njGSEnEXAYj2rr8AB
20bV7DZNC65DBeqEjoVaG/+yljT4UkepjcD4eWkShkC6H0WRQ8IDLE4jcnDJN+ba
4MFn2M3BxGX6I6HrFyJyr69EkEQNozNP0hV3u0F8VFvCj+QUUYZQT2M179TtZTco
0R/svcqTMYco4DwsZ6SfRWOxKUrm4RFYa/0ZWREtzEdcFdqc1z5gvH8uDDVfA/QQ
c3Ty5cR/pIbC16hgmB4yaO451SxMgM2NpibomRUPJ5PazBBSGHjemJbeXRSQGYTf
/juNJ/uxSmTmUPxmqR0CTsaXy6gJkgDuhLlLtSHViFkJpXkfgWQlD/udDWxFIzij
JeQaaiPuCfRP3yWxWxhKJlTgV/z9qFkxPguiGaFN5a6QolDfOj6oNLNoTnUP9PcM
w+mGrtKxL90hjRD9SALUvxYRZgRpuWTjrfg8WAWIgn2SHWXtjjsSwmsGpNP3vwnJ
pcwhYjBqIYdem3Wkv2odokyK8aOqTwQol4ykF3xBls4oF7DSvNyf9ZCZyB22QuUt
KTQT+hajAAnJNYaDvII2Cz0oUeeFhM1Kgs19S1x0l3GhJEuT12kRTYbKJ9ASZYLR
IvMnrXuOy2W5a2t6Q8AtQ5ZAMKNb8dkXLvReCvXgcBR6LboqsG5g/gxnGaVvKatx
jHujjacAOJ4higrppnI1KNxBIn7Nq1i37BjOBgr2ADzd8PBdUCRd0B6If/NPrBv0
9vst4EdNlI8lEjvNxfyxqR6TzqrhaJA0IHXpJRmgSnsGVKPTb2pbRdjT3WkyGd9F
I3A7l/qguBqvUcLzWugYNw+z3Fhx/7OiHv44+V/r1ErqVImuqCLemA6UwA+qYUyD
lz/2NGmnuYYLRddmexf+DW3fqXlD5SCDbKIEo+WENmBDvXbpbUiUl3SO+gdTfwap
AHk3MsObh1irr6ydERd3U0L1GA3QqrGI4bWZPfjv5JfFaDyGs6+OEzNA8yXim1SH
xBIN6pQ52kGRhnhN7Urpu0Q/6d6MX+5IpAk1SPPpopVqQIOuKXB5QsdireRiji/c
rLta2wi+83QtMWFFo5eC1mAwkDJXqblOx2Qv6J81hj/E9gLyMYd87lTk1oIygYhY
jMpQY4J8AJ0MrndvwvXffi3inogKARar95ewBcw5hvrwh6xTxm5JZScYWQo1kVxJ
XCBF9iE1s45ibIN/wu+lxGg124uu9Ne/mk8NImpl2Wutuq7MbZOdj729yTfpo3KQ
vWhgQTj4TDTNg3skn0KES4Y09PQCytYBwF3ZcK/9lCcXobPLNhbS5QNj7VH/M9Yy
JmUAE/qOKJrhgIiX0UA4Buzvj8zIREJaoh7AOVFR9L2uJ+2N4Afczckbhm6bKSKx
h6MKUU46DQdAGi691z7vcgbefJW1HznatKlTbvAqKBY/1uoqzy8NyjZEnBOcDMJo
3tEVs7W7ajMqWLrCrdpa6h47z8FHjlGyv+yF8mkoWYNSRzk/6wAfb87Vdy3xBFRZ
feky8K4SBRBVnKljdEd1YrDNZJo/ItITIkC0Z/aN728TLbVmftRCK9j3i4xnusBV
XobUxU0Ea1/W1NO+P7obkNQdldjxFV2/pFypTn91phNrYup5tIKFuln5NnWsWX6d
BocHziNqOdxPgW6Dejzd/Zj6DXKPe9Xp43dSN+4k/sF7FsPADUmmy+Gp3kgH07X5
3Zq0BDcKSgjx5OilDuRS4KuralPtynxiI0OAZJx0BqwsuW61yhhOvUXpxSDpgqsb
/HkmyQ5CMy6qI0GGYIKuFsfpLCGzHIu+WQUKOfG67OAyrcJqA+ir8lGmM1M+VBjq
CDlF5Io80hTBlBaEGZbVe/1VJri1+tfjGNFuc28e+UVyU2czYkMFCSXD0aXRU2aw
wgg5768uzlkRPqLNOappnBZRdy0itEbHoAieDCfEilid9xoMecD+vlxgAhIFKN+R
a/jtDO57PrQeO+aUwZ7Y/oSH+/L9jvV/207kJSt8wEghethArZtt2YG2wqP7kOT2
AUoV1q97lZtPvWtOgrVhBCh6LXI+ZtVaQwoQsJHVmdqlpUPFoJRCMl79Nt0vtQzF
H4QA4ml40F+ZmscN2LboTugx9t57HuxUgrsZKgDP5o3ldvW0Rbf3yUzN5nwH0gik
Nkxzqy7oLgMiyHWqhVGlHK4SycM26/3FKl8JH+N3zwgd6DVxjhHaC0BWONBgriIG
lf9K/fYHEKAO8q+1NiDLbgBcdsY6xvGX2SM4YOt0Z4cgo+epdl4xv7gj2YBPNn+P
5lbdiswIP4Ozr27NJx79UOujT9edlpzSs6d/kSFU3AX/7tpdvKkJwukXTPrP7HGh
MIOxONnK/OX0CQ7Q12NBTlVNQg6doQ+jRQFMiTr3OKk0M2gIf6pdPuCBMXCfav8I
M8YjDeZho5YZ4o3G168bFr22Sv6+AVrZTHH96yRxz3vVP08p9WiObkMqKETmzba/
5Qmd9ge4fuTDH1NPf39KMRlXw8YzCUcpn4oA4Sius+addKgMqRW/Te0FhE1iP+LD
RqmaMDe248ck43sPEdqYsWWA46HQOczCOHttF4i6YLC6PXfmEBSCcTNy/5k9Wm4U
xFh4/dgsDTWMWEnpaegnM2ZE+ZehYc+grhZO4XKYW7tVIBPH+v+QnQOS9LAj65FJ
DjAADIz2/EG6B4/FEipyYreST7XFgSiChQAFZ+y1bSR+ND8aIbnmL1spUBW/pxKQ
GK0x7NiWnPit3pqORj9HFhw8W0U0GeHR6hOHueO78PVP4638d7Zceu+tC/fqG/CN
DGHGiSpAQDf+cwqbM+MMXiYBCOW6WucwkXylKrB8dYmXLMZ1Mp/9HgCVr6OgIlti
8m2TjQpBGAN3W+S0qvtnjxLrbhXTobwLROPGdyBx8AI4liQ1rAjLlwPmhliq69ck
acsX5PIOACoyNmbPunu0f9bQr11TjD2pSLLPTSOg20Cmv91ji2fggJVcJkLGjjvP
8/iFim9SbNWqStN1FEylpYURg+2dHQDgMEs0la4Kbkgc7irgdqtTKA6RDF44eTHh
A6nlRWMbUB63L+zcs5KWzqHO1C/y8iUfuS1Gfhhg1nkyfyqjrIr2tbGOIwFQOgxy
rkBJzbDwD45mG9/mGcJrm+euXGbedw2gGizlTDhVxCp1URWycLlhbtgZyHZ3VIyF
h1eCIymhi7gCBjeeKBtyW3fP/0tkq8YIq5H3PghG1HB1YNnYQA+VJnvSKGOP1ukn
aVXLnW2xYiLJl5ISv8J62hI7WfBbbeVFJI2aTBipaqUb49g+m7VfDmRmAIEsj3DE
KD3Mbudf7xk07Inbm7wp4E/oLqCw4p4+nFtMMKVKQ/hUk+dprwuo1Sbx8n9f5x4E
Pdltitljq5VgHbRK4mF+Q0+1PiUQCTj0NJ7jgiwJ+Cry+RDdjMsadS7jB6ucBu18
tngmlk3lCoaSeKY1MnfDWvVr5BbYIM63ZDYhtboOe3gdbuhST5DYhU3YxNIhTiaa
xUVSxsJLlxI9iNDCVx9jEC4Z8TTeomENfwbg6osR1K1nd77W3e3xPJ37Yu/9+TGV
OUntLzoTLAXTlVLWEvc6z+axXXqsauRf6H7H/CJeFrPdntIMorAA1xOprrSMkSAd
iO9e+Ol4CqRaEojqmPEHYmNmNB3KpPbG80j+B/eZqYu3beEdBNNkkL9sGhHnpmcq
1K/NBihsf2E0ZW/dnJeQ327yJ54CtbWK7c4b/k0M3dACU3ZIESBRoRm8HLJi1OTk
wQE2UK++SgTE2q8Kw9Rq04IhB9vm6tIhSP+84jJJYYlHboJpJUXKL2zy0vsuwKJ6
RQWFKkRIblsBVZGEChZ8jRbul2W553YYAnJ1F/pb2mE23/hh9N1cjq34R0dINpXX
J3a7MdwgsHvdgQKx7hUAV81ZGjuMqd/HtSJcWLQSNIacCi3oDWI7lK2Sod5H+0Dn
ce+FV4D5T8sRdXV0xcZZ3KRXu4DSu4D67BCym8pNhbgaob0vMRH5L9lIKZsehb9o
lNrXCcxdoWW8ET/ngcM66ym47bQ6gAn30UibnAGC5fqHpEIqXohK7TgUxFI8amhc
JuUzh/BKLVRhwtKznC//p2cHd7HE0Q+Q7X0VQhNjANM282O0Dvu+pXhyXJvN6AUb
7W+rjw1ySsQT9GIMdDfLmvYWgmHH1WsuMirvpG1S556DuW+863bqIJjFr/NnUe/K
EJ4f4v59bl2R9tpBhPjQeuuBGjt1CxxvZltqSx0GvieP8NhBsGEPI6edDlvIBwI6
5DD3xt6B++iUVZGx1KVgsEooKRyvKDoFqSOj3/M8vvGxIU7z14sNlSpTBcsTa27T
ITbZZ3rGNp54XKarFi+LnoQ4yJheMpehAm8Y515B8JebU72NhGcJfAXeRzmkUPfg
3LHO465ylIZu6ETw2sTZljNDxbU5yFL9joV1/xQWNO3noWH+SF2i5mdXorak4d5J
E1/UMuP6Axt1JksJy9X7pz3hL6cR/Mg/pbXQXjLW5kAoxD8qejf4oH+RAWBqbfSp
ccyEKnQg16Fc7kHruhJRszbxGcujMLzvlaRgvbOuIIcNTrzuJi2I5UCmD987jMa7
UmvmNNiryUrGr0xyfnD0VRCyYAfmZnVxTTbkBd8plYNkYj+Fx8fm+eM7Kk5Jnpol
Fm9bgd/Q22dAV1lC6FfTLnT0oen/qz0yBBMPEw9jZiPU8TEFpGbA69+h73tnNrI0
CPCy6CWBR9QF+KWUzMIYsk/VV1qumazCeKdpSdJk7cACwMxMTX8UPsgjK8szy8+X
/MvW8O380AtagnssWaCA7CUe16uMt6J20oLVgZ1oN/mejG9BpoXsE8d7KGtRNBlM
A3bOTX62LgQnuXkEAo7lo4mFNBqPTzK8etQWoM6gFpY7Am3vVQe6ym0pZuQVDBUa
fMCa0tWuUULoEsRAhnnoirEHwdHPqMvP4nIRkZTV7rzaqqGlBxiQW40giuo9wSW9
nhxVd5P6COzt70l0YEk9MWLVRDx8R5CG8GibnBXBovaWvidC1r7Td5r0RWcTV67O
+sKkvu3l/BI+j8sZz8B8z1d1se0m/ri4gl7IfWDtOANf8PuMT7fBQAO1lMfgU2V1
3rcqZMCBRi+OEApChQ5JF+tQ/x1wvJgnYsXY2QNxv+YBAiWmWkOZGpJkK2JWqy4A
7779IiNlyzoqcDw3qcDMfYAC9nCS2qdGsKLZDuQVmznq8dcOD+f+qrFuSUPHa0rI
sQFsVg9kbl49IZPljrYKwBDXLDMIhbjMNnWczIYbnyh6h2ww/BSx+goyhKwUeYsE
0FkphMfbVt1+sbhDqGGogwngy5XWXprZbLCJzDzsCFcgPD38/zF82GI9XGVdNISP
EySgYl2JHGxkswOflCieAOzCqhjRgHvpmvQvixEVlfyGYIxVKo9146h+k4BDrwBc
lrJg//num3clpdkt32yVgvDhkQJ7KTZGucKv8pBDRd2wpjjy/r0Bo8KSB+HbAuKn
xoLWdRpFTRtGDrQPuYYXeWqvCkgdgeNlWpzsohq+knn1en8cp1Qq+zcMm/gaprFh
E4mkFhMrl6a5ow8AnLkAO8CD4BTzT8AU7qP354xDChX+6rD3gyI2ppx4l3mhm59x
as1CyAj2R4GefzTaj1nZKJjd5p1CdTNRZxYT1FtjM3v/T/Vvls4kn/2PeuuvE6EE
X2T2Kj8pH02zvgPE0Z/r60x8TsA5s5rNehaijwu3BP9kXjmkVsJ6NdwwTD3aHL/s
qKBIXCPFYuwhGBCn2S+0mACD6ju0hGso8nHxZkYonhn0iIyPnow4rTdhoNFx2mI5
1mHL/aYaBOGRuNzKMbbwbcWyOjA9RDK1lP7xjQKkOewiaCMXZrqCL9iGZzour4LA
tlD8OB1R2DURI46q0xS7QcuiBJ2lg1tpPlxOnHNMjpz/HY24Zz+e3wEiQhpFPlU3
e8iEhra+/obn7O/cz+eiC+7c+nnAPzFW9iInmf8/+VbBXglYNI049JbcxBikIh+u
XerKDr+p9MIlqQWV4a75YaWvEHpmBu1twR2XgbLHFG/MO6wlTLr++YQHI+xVmhPs
TLoUzxPL6NSNEKbVyLTQR8CJEG4dk9H224+ygYKhQ9pkVKxQ5qshWzhNQr2Io6Jc
+2yllpg63l96dnhAgXlOmsu1IOGYutT2XR3L6TTWp534whzDR984bZzAMQo7Xlva
9FZW5Tdmd4O4B9kc7DHw5LnL1CMpLNY4yqjAnDiEfkUXVhKyCbgkBXqRuMlQ/fyO
PHJam/s4/05JtELBAhQoFzzW47y7F1wXtPngsOBi8eIEHysWLhklLD3+WHDiBtct
2Ez2XbDN4uxOHvNLA43TSFmNiPvn5yLHpEBgKxeg3mR1dv21C2myEEIAt7B0UrKT
604Y4U3ie5Z3mHL78OA801IIQus4s/uIr5xu/bjpRzklRL9Gqvd+uylz+qGW0D3x
C+ye4TnTkFq8kJUkdE1EqjrGfHM67iw8qpgnSJzgURhIrvOUxQD09BSsqCAI4Efg
WEQIrxNMZi8Piy0rVucLhtZu56O7Md7g6PWLJeostADqraH9Us1YFt0WaATcMRR6
tcsT3GZG9xDoetzouD0dEBnoxQunVB8FHqlj/PUC/q7M/10v2c7Sq0bLIa9+TdSy
jgXVqMzcseYmcQ9yNvTZ+D9rTiggeisTpBvjczpp5WmC/PLfhpeKPB9a2CUUtRxI
D8x3YJk1Wt61LFYzQ/i2vvpX1NB7ApfO9Y0vmBRIYgHyaRio04sG7E7dXoJomXI4
/PYd8dXTO+oCCmDB9sHfVfd2Z/zMiaXJ0vWPgWxGVlS4PcbiPZLtYyrVCD794m8z
IHnUv3rEnRR6AcHOvG+JRooakfDaERuqmy1MC2LCmC5lGLXBpUq1YKdxPVpwr7a5
YlrcsSlTaEZJsYF+4kQM6AUdIPoLGQqQ3XZqNQ+hAydjA2beS1GnkFyKdfrcv5A+
SQ/d1KRMRsLr0CvFK6K0lHQcMo6TMKuwFLcz9d4snbYWdLLI8xxrjoZ5ZEpyprI6
vcohrKdbgc+QUjvbD+RfxlPt2iI/IJ+BkzbTGJCMhmCzlijakpb2v1+gbA0Szgqm
kAb9QsW+WYefu0hwjB8zARk2rIV7RKqQ6JhdENaTPrZfrUi5N8DoAztSYfSHJoLg
xqCN6B3jBhO+JXuby03tzMvVgYQCmjPM9JdTFqPf+8xJFcbKUav92wUZlFN8EE0K
gbSJWjZq4VwR/pRf11unt+WPnOoc2AopuszQNry7LunuBvh/x8YBQ/zJFL/qETSn
TZ0Diz9jDg/tDoeQN0lBMOreM4gYLGFaUYEoTxsOtFaXlmI99ylfQauS1TJM2Mqw
BWpLdpGeP2n2G7xjtRmuPeHyvV3Pe3ByPDuBkGrOzfSOwX3b2rVh8hdASa+FxXkc
ZhwHZ+nLNP8usI70udCpth7AWqa7boGjOhj3mCiDSxqJL/xvMBT4o0l/mKvfd3L6
vdpzOnHooBaDAgPDxy9ri54XE5aBUOWr+DRdE7vQhBZauvOH/Rzwb8tACflJz3oa
SiK1phxzyAeakumFUMrQTToTkesz9kjtmakEheTRuWrl/3ls3Oby6/fRdAbPOy/H
etfR4DKCfKXSLIhg/Ish88zxeg2kxejGGkA0XhNMWhI+GV8JXSofxlBR1UcMkYNA
sc+YUz7bKFSnP3IdUZa/g39rm7DfSTB5ow0OFH39KZP6RAETm0BAfPCKCjK/XfEH
X7nYDdAdW49lIdKVV+EgiIj9FiYxrkyMPaj0c//MxYPANS/SGINcuPSPrZNYnh8j
dWANV+3AiaEUS00j3ZHQ1gfHnUvaXTaWt7GrKV/l6peWknOGmW7rG1yb7oiuDovE
wABZLfkEbVDFMdYVAJgEwULC4Snj6ONfwsRlDXfqDPBkyThOjusCXvPTygHdCg5D
AxNVOc7qlXE3LIHTIVMMdndjppgVWIYortYDTvETq8WgAVyAnBdXX7Oduj3I6Xdj
wijXTsdH3OyTyhJrD5cBxH0qRKanXgdgJxMLZ6m7Skq7i7VjluR16eikax8n9gXu
6PCaOVaY+E/2fuhpOCQOxJq63sZf8Vtm/lhr8MF2/yXqdSaS0RJd6uSmUJKu7lop
Mtljzc0lZP9d99xt9SnUnERx2EccyXM5xkZjbMWnZ7xnK+UajKSJ6+pAqx7pm07x
U9SlC0uAsq+0aJaiftkzvknAMzXQv9fAqYQj3wKWoTQatQeYIm+etx3Ew5T2lln3
AaLjHIPOwniUk3PWnKkzCfiyjH5c9BpTeiKTKKYPnZQjb8YEooijy+1GxvATBqLq
mEEGXKPJYRpMTgumZwDu5vFZ4pOnC25XGq6ylzOyofbikeN95BDDKib9pA6wZBrK
45u36mCaenL2tsAYosDBVOPLhr2zUd8111A8Iraf22vMJheoQOl1o/dLLeOQMjdy
PE+YHv1ghIwo5Mr9dRYx1p6KBlwWUjXpfVUQWhpI9uiOGS02v+BWDWxi3PeF0COO
qTaWK6ZL/+Q9g+2GW6iPOn6Gj75K0lE4DEb0y+Qw5MRmQOkbSUv88kajFKPoDtiT
ht9N0CN1+y3F1EsBSToQOebvYx0RM2Nk+WpOU1Rqc/RY2pMc7oCXnLPo+VPYsgym
qlMVf/Zmk8/UHBQ4O4abxvHEJcwO58+8Az9DlftqNuipe3TSTYuhrpYi1hsZ6niu
ByUJJXRrXbF5qjADD0mGZY6PLMRNYI0Xz0b7hAXsTi+Vp1Qlx+RAZWV7uM3I3eiI
SqbdnNPpXpcY9uQ7Yp4kYQZqcBORfQIOrE/diY+IUokf8YQNHOQo7oDJJZbZoXst
B08yLK+C0EmN+JiDoM0o/wPqkXiVbBSpffx9bNSTJdUNDypWzSAuAOcjgEmnlPtj
f3cK5s9OKNv/FGnCRha9ZT8EZ5lxNrjQu5/a96wgOBWz2FiO1DM8Sf5o2/AKnDWo
fwCpxLK+Mqse6plNPSfTq119ibnuHrszF+oAudZwYFJVuNg7Da9VApDKQslLFP8M
hhEssn01kwait3eWgvEuC4SL9dzucB3YxX8eXz8prkYQ/7BrK9oOjfk06lbxH1uK
Tm6phcbKU0XjekDlDHvTRXQ1jaLsLN4qH5kwMo2iL4ARy5mqm3L+BL1ZlokOooV0
CKoOm+AkYWa2xJBcWN0dCkd+BMwH0Ifi2O7swFFmfWKWw76EdBDUMCz/35CxOB/G
qoBjAI9JvmLODVgDWTv3O6qkSfUILbl1rvXrymn05nZo2Zxlx6DS7TYsY+DF1D/q
y0MHoHhO32tg8HsiQ1uTwLX61VKREK2QYhfz+tNNK2KDwEqG4eH4XkwG6PEOClsY
f1g6HXT+ZfjibAPcTzTbZK0o0lwLEHy85O553zjLGdNrfNZEkfjiDEIoLrSUWdIY
xfeDMoOKhZpzUPgbdhjYVEiov6D5voKpt0MYp7m2dKnNVGtvteXnfjjT/v9giuDF
As+3WCTM325FfGi3JneBfFgeasPN+UOR2lTuVjeJmwCFocHOHvT5WYou+2Xq+HLS
3XZCBkaoCK4NavUSSMGwOxec/znyFzFUoPtDiy2u69KWPicTBhb+ZCCRFcC5P7zz
OZlqQMWjYzmN0aqPVqzeK69YUAmeHA96rkv/scznW0fQR8cBeulrUX86L0/K82hM
m0ufeDrjoBb4L1G2wOklbHskEfQQ68oZudea4V+ONK7CISk6UKyApcVRZoH+RENg
jGF3k+1JwkiQAz9P1C2r6NAzDyFIzYW+Sd6BrbbL8CxH0ovpRnsELh8uYgoQq9WW
IQAeAl+4PetxvANKza9msS5ZqfzSaZc6cO3s0apfo44SVEHl1Npq4wS858ewRpBD
HKC7UvGMyQ0p5SQPUdk/IZYWtapkrB3vCVrXvtnbehPGUBKHyD0LgL75DYa0FY8I
EEa2acl/oPkJZJqcVfLOup4+3FexoK6C7oqU79sXhA5PFsLGrjmc9G64MmK3ggn8
dQpmwfxcczYBIA5KrOnZNTbG7rAMZh5Y4sm30o4bQ9I4sC+cw13zlJs1FCMvRiiM
DWYgmdDBk+kYgupCXOmqB+U3K30E6Gtw6sfPJPlNLOII0nF2m/eu3YCgwWMAsW6o
SEurELa0ZVnAYVa8QiUvCKq2b21R7r0E6CC4aQGAmEc7ijb1LgYvKEQgJLD1dbQ4
sMHcGcXBbneAu9loz8ltMWPUO6ruYDgWeyon1+GqylNmtg4sFYLtRZLDFx7cAd1z
yY0ZF42SJI7DJkZpPjwZ0jNe2lfCsmz5erT8CkTjLxCY9L6+aPkuCiPyBPjBXdcM
XscEOG25pCsZtFPUXwW0s0c/9oqjCNo8pJS33NpGQ4oOfhUgNIQUbjhlKVWbkzJD
uBZ7I14b9rgMaQcp1+uLfB9uSIInMvSBIYEZii846ZRAzhk6VnuRy1Ph7ZtSJSGK
lENoccmZEAAvA85KwYXkiISpS2EUHzu0ImcojT+97mf0GBdGj0H+AxTCqNXVDQ0/
+DZ/2Eeeitnh40xLL6ENmB5B27J+swLQkQgug62Tu7EAE+Xm+In7n2pMzNCGIOd5
o+/M92nClflVm0kJg0mPp44VscL2kjqSa3ubRIvJWt5JjfSaL7nioBtSE3IdF4Cb
9wpMf/BqVc9qSQ8hjyFaE9ix679ynnbEPmiREuLoBNrNpfKOjNq+8+kOaV02j59N
PAXTFmcNA5TaGP6IfDK2sqH8nt5CJJbJGr1pMGVtCrs6nfaxN/2LJZAT1rAsL8B/
rFbRdN6EQH9mn+fTnKN5NrwNabMhyCvQH0FEimP8RKfvWk+/gYI/IxxeCcAPc5Vm
Gci0nF3TQw9nNLZYLCj0MqX2gGQSRSuu0mROkgk4UkhHZ2o2emkD9vAXbuIlzEKi
VWb78stP08vQq17OLhMgpcbdxBhZmhVpVfuPsapIv7eGr2BW+2bB06RNiWlzvPsa
LEDtMEcmqsknEAy+ctfFOCdULa5b9vSbo770Cxyjm/COrJZAK3UF9OwFfYPChRR/
bl09nMsy749EoSCiy2kiWR79LWVqGHGqRZ9yEHRmWGW9N0bdxlvunlv8+hyRrxnV
Ip1r/WTBwJ0rwhZYNZW2IFZVXo2PS9EMhxCZ+9aRYmjzCDtCwkPFFgA0m16WHFag
itroyq3nBpnx03LO46c/1LZ14s7fsir9ADqnTUh1cnkZpf2fz9+K8nRcLK4fuN4g
7S7vG1YN3UqWnfIHZp8xYL2rJqCTLAT2AX/ytAD5lHZ+3ox7a2tH4L8KW2DcuGcN
FCdCjuc/OZs75mfNNdbBVnziCXOzej+fB/VRzqeN/zmGipfShOgT0aVBx5BVqzrb
R3Z3+LXcagDQTdx9ndCGXYio1bB84hp4dI4/wZlHe5iI9N/P89ue5FD+HQpy0itG
z/meZEs4v68OXGFDsEKmpxUrcwm2oMNM1ksdqKtZY/UhFD1ihfVKb1wYAIZXlEIm
07S8aN9KLqZrWBA5nwMpoZ2Rx8VY+dY5TCqoqvCLQp78ER/oTD6T3bjxteaIGW2P
vDpcad2trgZ1UI7EuSZ40lSau2/ZjcO28iZ4ZMd3/AkbZ/reYfjaAsEUgvPvo5lz
yvc8S6xbcfa0kqmUBwHF5rmER4VFGESahnUy/wqAcovnR6NPCE//T+rtb7TgIEtJ
5FeUXmB87ikJ8fl6Kcz6dJBdibRo8+NEYk6TyXeT6cjpEsXnIxip1OOGPYCsnEIB
QDblSNh9CpdYktY23qWglT7F2O3FU9aJH0jhMXNLl2EZMIAiEnunB+ZW0PxJNvlD
262/O808Wc5TsdZyP1I25ym3XdQJ/czMFC9jQq3xD6+8OOtJb+NtfhKeUQK73Mb0
lKBH4xuaxt4bZP8f9aHgaMgRRzB8MleWtSibU3ZoIdKQH3PZriQ4i77MU32pVb4W
ZE3rgANOGKqxlqeKvInVi7LQ+9Yr2TjnDX8ZzXUaJJY7cJ7wU1aaJYX8zHm4AS3L
hSvwX3qUnLtF3eB/mVKrgnPksdZxoqr/27TPDjyAjdYG7t9XwECl6mJhWYY0aOex
/wWfvXtKAqBK+FMTZ495NqiGrkIIn918NgH2o4ZUawVZn9rpSoApTosuub3YWMnP
wS3ZJwTDRiCvUYocTvmQ75DE0+XGANL6TZ8AxQUoHVV8e21KcaEJ4yNDrC+nPitr
z4JeNt301rpIHwyAvyBULaG7RHTfCNR72sGoBmAW6uOD/APu6RmP8hC36i9nDonQ
9mD7yUSlgOd6zJr7uWCkGFYxj/WfIBiJM2vjqTxdNEUk1eCr6ZkdzzbW568FIFqn
Z8EhgPMCj0KDr9tpYeKK7GfahJyOh3K++6ihiUkeCrHnT+P6Fx4TubsNirX0epE/
842OQf1g1k5bzIZi2ETMpG0xfAzKhRESI/zC/ENFQiaquF4FG4/20EsfZlDzqnMJ
VPHTLhnIN+oBl8g3meThYI4jNu1qOTQ4Cj4wk2TFrZvz1lkixUX76j9WtqtxXczb
Cywd/N8iK1zkpyecq4NzSmuAAmnGRmsp2+YkpTyBrTs/1wmPV8lyJIMTBMVLTmxO
+P2RZZXc6NjCKF8wIoHdELjR21G3qYtKWwTGtWZEM0VXTlmzj/Qup070QvkfGcDP
SxHu4OTDBzydpi2xVGB7pupXxee6kM3/OB7qdoNE3aktAE02CRGqqufsI61ruhrk
gF7nEbrL4Zr10pyFmmRmG6b5CDjw18Kq8aRtRucJtwGlF3c5qxJVu7djHj85mzUX
EpNp5LhoHWx2p+YRpYqIXU3ViZR5opMVnOiGlxwt9camn/4OkugHPD1TBuOiTd0s
t97frXRmcWr07WFjj9g14Ew0QmzZK1hXgmfUXel01dkoblXkmddnxv1E19veqfgT
YnROoOFRkuvbWq6yjQgdHyAwEh1eF4mZabattJM+uj8R+JorF3i3//xif3F0E13o
F8d4ALQs3LkkJ+CeVpaPHx/S6c3d8qGF2HkX/oXpihWNUPPI4DR/QyS9JHgb9Gza
w9ubGbyPJ1h+DwNY0iPnXyw7/BYW/MvqbKkoGAcxLbsNurJYc9nM/l9z7RWpxOii
y59I+gaAhuRoA3xDgEDa5Q3cC93gSb3JVvm2W7BrnsMNrBMS0oCOP5ZnutfMjckq
/7orXk1I6glAC1UHdijzdL/NXan5DhPAWmznDuxCPnoF255vrHuwiKxlbATY9kln
HUwvi5TN3WkFMLu29E1u1Dm+rwl6UcJaC6zOgMXF7ZTrrTPrVedIOnfU+ERsJEaN
VlbZRl7MQd5iPzc0XnKfzkvmk8VaDD7OezbBDxhBU+kAPpHulFfKQ0ZaTzdp9yoh
eifMaB4ZaVKHgizCAGrMClxPnMsD0Jvd6iMfP6h/NfTqN+QE+TLlEQPkb3ikaRTe
qBLaujh+nD66B5HGN73zSrNto+RPsgWXFKR/IfdSN8DMA6V9Z+YFVeyRz4WpshUg
K5R7xHCqP5apHYTR+/NYBe7xspQSkbFfnOrm3pPxgv8ORR8i0WoZzAXwzoIbnWD+
oAAE0KpFP2DuKRAr5MaIJk4uLCJoH0aOAGPq+7MLWCk2zn8vvluxvjfNSd5BoOES
Kg6tsNBt3OVvOAbVz/zyBu1R95Jq2if507ipdXmvHSNDzQKHOrN475L6zoO7nwab
XXtMgihpPaBiTLQ5ysfUmlBLVPWTZIMjusI/eIu+8Wqq0Q+WoFovN3z1FJ80ggfa
gTZxqdR5ZmY2EBiMVJ+xVh2Dz6Bl6TM+wWEzFpWAubPPVLzsi1TGfoSNyFcnHG6A
oR7rc2avQIFVhQJBGb1vP+T6XzHbkjy7NOqeCRqpUYPBxSi1mIBBysU8ORZF7f+3
4kg0MsdgPTGwnxhQenRAh1WmLwvNaYF4ebl/KweZeIQLA4RBI+g2ht8lQo4PYdrs
rQkS+P9Tgj4jZXUup/rx9hzcVjP8YYSmwrcH0PkOghEniC0XutLVUpd5GYAiYZvj
RKfTFZu0G8zcuxTVk9mZvmG9O9DepUF+bKtt+lx/jwd/wjjl5UCECFz2apsQl4mF
kiIyjyjWLliSwF0kRn9unD0fa6e21RBFdKvdQlxDpdxxnLMTm3B1Hh+JBdVrHn/9
KvIFwzbe17Y5yYMA0cQ6DbkBXd6kXx2eCKFYra7ISPm3lfbIU/YBLIhPqMjx4rPE
rGs5EFTE1vJ25pebCmcdM+t3U7c3EoQFM9gQJx3RN2KicwhQY3zVn5gdqEHeghm5
e3aZyI/2KWam5/kZHS5jfCRpiLG8QV9tAuGqjr/LaKaoVqb/QiDyLZApx5gxAteH
rIwpspRtRK2IjT3oIn6/3LBaQLrv9r2WO341Fwi0iguWF9wzrQHoOK6pYpaFV7SD
DyoazIvZTe4MS3E8hGO+Aq2YwKW5Wct/a/OhmIaQMtqZE2JC/3TPUbRc+hGapplv
+B2egQmPn2rdMFHx897AyQg5bciVMM2vEF+Ccdp8oUZ8V5vergN8xd8Na4GXMDgC
wJyl65eRipq7UwR32sxrKoGHT8SisJOo8Qfk7HIyyMUK3ZRuWXb0GdJGB0Ntr9Wi
JuORjQuH/GdfSe1a3nCJS99kD1aP1VysDdOcZHH62viLeRgRE6tdEF81kuE9iws/
gMxke71e5EfNByXvkXKIUPiAKG88whGTAL4I5TjuAdcy3aSbAq0aaH4xxSqQJDw2
DOC9znY0h1xYEDbAcHLgFvLrztQl/OlQcsMFwQ6GgNFFsWEKQZEoM+LSo867AbBf
Lwmg4XWI3hgdsGGURVEFEY/Oa/hMRE+lh6bM7UZTWy0teJ3riSvxMtq/b0NagMaI
Qc3Qodrbpc8l2zAEsxhrT8EpY4jCI9TMg7HvWJSfqtdCYofA5WNuMoKJq+WMdSFj
jTihhI1FBqmgX6YAmMAcu/VB25SOe1Hn+19ytrsvFLA6wrdPxIh1y0HGvjx2htOP
X/MP+urargB7Q7LV6KfJicTq5NR5VuMLAq1w0mDTYpuGlgDz/tuxcr/dQ7RKBpng
c7HAMwT2KyhQ6+PtnPE0VZ71FyPsM6iCHHpCTm45Dsre/TLU2B1p7kCtQs1UO/BM
82Ej2rY69c7XJdW9ZHU/VreRMhabrAb1E2Adu2xG6Qw7dhxisbp/5mh+APzf/4q1
Yr7s2ik2jyVy6v02LV6OcPSBA4Dw8L4hbLNWBCGe2L4OGLEkP8grR05eOiHtfBd+
36FIB3lfkuRm4+TSyG4eRvhOVUUlEAJadK4k1eh7JWa4uGLZQ2NA0SNG02ghyqgl
1ETyRmx8AH1qXLKFmI8m2NOkvgb1Z3kTxcILtlNOLmW8noZ4F15TP2UXGiKOzoYQ
uU5DIKsw/lFUAU6ilfXFlrAkWDMgBXAEZLXh5k6qOKXZ5myB16I1CDjhkvLcysV8
8Dm+4zHF8g+87qSVYMSLW76SyyhSYgjau5VHVatC36mlqQvovZVdBtWrHac5+rYS
y7+tloLD7y6MPqFQI3XlPnkcaOkkBSG5+PYq0uEw6KYrd6yG36OYn0cETsKdqUZK
GfKXY1YaI1pQFNta+eBVfBgiVBgo1xhMEHIz1lxp/NsyoEo8lwYuBPTNsau8L7n8
rdnmWdURJKfRzSw/zSJ4dJLBCmC+m/gjQxlgnE7hpdl5r5wpp1oP3uobSd5hnpUt
XMyjmeglPrrycuX3HnFK6gEdTCb6NpSLEvwj5hbaRHe86sP3QVqeAmEmrTm3IO2Y
i0fjPp3+trpmpHzGaVtW2p36O5dIAUdsHiQhLBL6AoE2K8Rtv1LVwy/jSzvB0qgU
5SfL0g/E9W+tNj/8UWTiUNhqeNMIKc2jQzj0ZvZjrH0X3EubHo3txBZRrnQKZ1dG
4CQVijQNHPA0EiQLgGK7SZKymF54AU4CVDz+dP9GWd3e0qAXVMu/RZw2ySkx1wB3
cGyB04qkjyH1go5Y5OFVahsEAJ9rRUbe9u9noE8ZjhVRNGVUyyaNV1fQE2aVk0Bv
SVbtnZ3+zH/ZFUodRp0+P/jpIotN71vHw58iHSGMUsRHW0ZVfEt9TxtxiodxlTVA
ENGXqVN9LgnM0fL50wyzSK+wCZvDzaSBgJapbwTJc7tISbqISrCQPDm93FTEcZQl
Jrf2gMfaVC4tVRS+rPx88QStlzy6PGpD5aH9iIYePlnTCWXfGGdVV4NsKIue6KIU
szmdYvj/okacL+3kbCGnUlw63Si8yZpR0Fa8sTVtkISh9XVaIhBe1aA0N/M9nHFS
GI5nwEMyQNhlK2nS1xXNKCvGlYBMsKAAB5HL4MTMExbg2Nu1Fg9FyJVLUZv7rquy
TUxHCVc4cXClRVxyxDCyMd9uUDLkt46t+vh9k/tnXc0kfKP8C3g5bBn20m7hG5wr
qjZbyJvz2l5WI6b0brGLNnaYv/p5Ey+mY3iTHJ1BeHAa5c+vn488WCPlx/A4Onx/
zHvEX5W4q3KwNNYV4RmE1YPZdsot7rg6iTRaSrFlVtsGlN/l8DP+6E6ybNznA49b
klInRFQmCjg2jf9NCdR0nnhvPTQk/e1HaWP7mDufYBrb78rFWPYTGolidYeZlbq1
D3el/wDB+ISv4pFpydS2i1zmIZqMvF0Ggr9stGfgeSMsDq9VFE0K2fPdqDP084ax
3P3VlBLQpnS1XY17sB6TmmA0UqndtEMPdQlJRnQj2GEfvwJNuc3l8/fiz+D+K7fS
STVMOxjnSAxOxwEoBZ8EFNm2ahXiOI+RloMWV9aEVJP1eqxHW/kYY3fA/oUyWoXL
AXWTxGa8IK/mb5ieCrdP94LXFPHELFTj8jZVM+kO2U2gIJ7+Q8whSv5J3w+Y/T1Y
peB7xQ3dGTvxO4+XWqsqckUM83K0VPgdPSE1bn8MVZVRWk/hkLCqYlPLx/TPj1mO
jgfa0puxZZyfUwnw1eCGy+QIlKzb7coqpjaF5O0haRoJexR+13KKB8mqAU8o2l8+
IycEqYvjxkdqdUcGQCj7i3Et8fANRihcD8llVV+7EnYqOUtYcKtcE/xv4UwAx0UB
qWR2GMlPbmAim0AQ2vlB8b4sUrGvyIcup5x5FApCYFIPVWdFXPmne5GBZZyil6yi
9NQbesnRMsnlRxb31bX5O0x7oKpcsxDN/I0bybSWhJJ202uCSeKwY7RHpqbzyoV4
jlUK3aR8lwsomLX0e+bXIJks1qE+esO7lVP1mv8J7T/n8CJ32qWbjuSGcEmWyS+M
lypHjo9OaeeHgQju7gBtV+r5Q1kE26XhM+A8qIMCDzbmRJaOG9Bz1GNc4rCmOvBV
SspvNGa/HUpK6iG+Zq6mDNa1A/g3say0wsuYh+BxbwYA1LfrTSr/KtE6RzwNUfsd
JflkH/t7U6GH96Ua3nKmPyDAfEoPwrmbwy7gvm/OneozSeazFBuITze50kDahjex
3CR0uIg/K6X9c8GLwDLy9uG40GsVEIFPSjSy8+e2Gs7nkt8+oxaFc1eWkpeSMK4O
6porRb7WGkJa6ZLKfVOLuT/gHhpkRF77RTUS7VnhwE16TfIE2TmKRos6PbRImuLT
frxmNV9WoU1vQMYsXawx9xLSIlEq6pV9uPgaDIxXtqhPVt608jkbuEO0yXA8V10a
oQidexT7IwQZsR/RNTjXfJRzSaFF+TED7vNz7OkqYg1txoN+e3tdFQKzEjvuIdNB
inOOpihz7YrEt0Na4DElguP8QpwmyjcKMY0T50Ew6jGGcVKU0WsNMjhiKZzxrtFU
J8QZVR8GImO+ihO3/5v1koevUp9ELlMxW8aJf43v0dIF204N6/Fy+toKCYvX8vZA
fRQnYfopMZagOkY88S7qZihiUSTWvFt9fRhjtsgzF/z850vI2NXX97lf8IqsDFeP
NnEqJimKKN7ibVbI8uJLqg/Yn+doISGG4ZWcW0tC8afuJhEG+OLtVIC9q6Thxp/0
Zo1Qg4mEj5YgpG6O7YPQOeqhNiFn7wliF9xbE16oLOX8qaskV1aaAgFy1P9K4DX3
5XcHp+2Emy+eB1r1VT06jDlmAWEeU0CxlrLJ7LJUQlzplaOy2UGpiYXKQHdym8gT
v36xiq8fv2gOCknZ+kGnxEP+wJZ9Q/iYm5GU1AsrT5SIlz4sz0FWNzeOujq+IxpS
bdrDzJhQefJzOJSGeIAeh2tQC5O+KZSehXFWoEYmdhC7m4mkfjsv2JXh/0Mi6bk7
0U416nPEq7/1Ecl/5iaifJDJtCnbqdPlVEPfXZx9hac6CqXtBMCNg2roTACm1jJk
2gymmTUTH+dQaFzWP7ZuNxNRMdCGFcn1in1OlY8qDBaeu3nfJXKGPRKPLO1olR1Z
K1jiSPefXviI7j74c7Sk4kswilLAg+ejbgaYiKFk8hketzpzvfWH00H0OkMBvgqT
epSbGZktpHP30cwnMptAWmnvrsKDuEfLODcRiy0x11seg2Ksg2Tzojm9CUit8lqx
uwU7z0YvEOQN+1GViUE79Tui2l5UcXZImuJEdbXv6Z+lyNUBPNswxhpqpLV//WG5
Hio2WFMie1PQsVLtGRKbuFZ2ZgQZOEHUcbj4Puyd+QCWx0qn83UEsDlDy2o4Vo8u
VkHqCmkT8x6mlOUucYDbllThbRpW5UIHch+EQZ2cZ9Vg+oh6RWYBNdWD6ZIGuLIx
OKsEGXf0rB6SU6bMjnf1Gx9PiSkj0UcOsU7jsjCqXKjdEnU8JgD6J16j5lbgfTuE
vFKtbh73ipsNbyWuA1r6Y9cTDDrCks8Z1ssLsy0DTsOlsdeZHchRMEY5yFNT/XJb
clXrwxvFN12JrNER4fjJiErMImjZhaPAansFAUSYWoZ54GttoPAHoUwgAEsptPwc
XUQtHl3sR8MO9R33Va/S/svJ0bsD/aufSyTuxPsKch5Ns0lyttSg7vZyoryxgokF
kVZMfVSDLB6fB0zsiJu07qwARSxj06KwQOfTnDZSVfQ7DToTuvAatybTt/CiyvDK
868JjnQOX1OC6oWVxyLGjXp2Ar3KoqJCysi2cGUB0docYILnm6mFnWf8METfw0Ci
+Ij5R8iRJEHmfRsk+6cl1a7BB751WY5Gp+gDfiBwZKI3ytYl+eh61yf/5/Ko5ATP
xQ28MB4hFEpfbzlwJsYUYPRWoKq0h79V/IcQy/i8NMrTnPuk2F/ggI4EyJpcYgCS
gmAeueqI0YpCIhlwsNkW3SVvxTe+b5YhCZCbdETb8eGWZkUKuZu/ieOfRW7dCZsW
wp9glBeVVIBlsoe6G6zHkgq4/3tmXDGIvKWEiZvlG7rXh+tLnGWUuWzDxsuBZszb
hLV5DRiw3iV8MSg5cFjZgZA6CH251wGzISGC2Djfy6Q9AhRoH/VoK96iQVSvfF58
DpuU+VdnAXnDEP56mwcj0mQDNdsJqxKrg4LSbOBGOoWtPisBEXojjJxfQtxjpzc3
tiv6tHZM+g7R5MUgeNM3mlFgFZfGr8tV/coIlpQY+BQxgOffVUxyGrdGuD+X3mT2
RY0pRGflP83X6RVo0kOHrwWoVIIJIDQ7wl53FXCNzTnloDv/auhiSAIinhcxyzuk
QYJaYYy0K2EotIMNJXOWkOA6KjochEK6wBfOhjkf9Ktm40rOuuvrShjznW4/GsN1
KhQlBDUFZy9TSyxsVm5O10UJtpOABxbWMW1/oYM0DlnOtbf+o+/sSpx1OI9i+TP7
KMcGYJP3bDhI3TCR7eZBffJ5Cmty5M07uFTLboAD9Bz+kAy2mSTAo8db7kHVXj31
op7OM96xQfcLQjDFzC7Wbnp7bsGnhgk2W8EX8dFbTbMSiVF8xtbyz4uqakd/hsVk
DmUoHCAsCmr1TDs1cx0b1mTc+9l6IipS3/fvDAc+MB87N7Bi29cp3vxDsSk/Ef2r
xRRg0g/kf3PP471R8d+u21j5fFvsjMOW4sWq1TuyGz4HDF/Sx/BPh21NJtrvdD45
TCtHUjrKor+/nWWpsXLTLeOt2jjjsOeuSBkvtwsffSzoEX7mHedhtab5WJKsffkZ
vMRxRVGePZVjiOLczepJtQztZk/tcpo9lo6ycnh0FjTXlxdCmD8Ke/FWDCJxfclS
VyRdJaLSZiexfh5Xo6EqvpAGqxm9cXesfBFuM207MGJNa9qU0FpKIUwdjfntsxud
+XPieJlft27LzagJJ5SAaDfEQs2B2ECsBSKWSF0XLxC/+Ue1yNRDzu4fTsqdygmG
evn/zeO7boR0v0/opzUIjJiuOE9tpEgMkXk+AH4aBgikdAV3vlx9qtAlss7R//Jd
Mn6e0vQQ3ai1A6j5Ky4FImEHZRudQRMP0Vq2jDa1FTAIngR6xdGvNoLMwkW3y+ac
XtJ1oEIZnOqFpX84eiakZdc8JFazfnQqWgCV/Jt8gPL/7s2CnyS/hMizHys6Oxv/
ltiiTSjYbwof8evLYkrAkVfzY2HXpkeJu2eWhJGzMWibP6lr6lqgAGSgJES20qAN
WdJ5acvgilNIrS/S3666LempOBLFOuqm9PHnrIZ/t6kaV+fkLPcV7bsL+4nj6gSd
ejYfgTeHozEY5QcHqrPvK26DDMUPyO/UC+hdQvHDi1tWZx1z447t+S7Yu79V2Btb
B3fIGMoM++IPW6Ob9k9Y68BFXhKoMB4235vJPhgqv2OD2Vs5ace02rjqBN8nEc61
3d6Q/zRBaRvJG6AAx9922dia73pIs8SYEgcvhHL+1FaA1yaa/BtufJ8F3327ZnKn
/Zt0y4a8Zi59h2SW/6LDypQu31uxxVndAvDQHNdSCsNIrC4W6cXeOTkEwmEJopvj
jE4+oXmd/+hl17ZwzkSzQbuIDztge98jJ3b/8sze1/nEX7w5pegWU/+tziQtLMOg
XnxHL0s+SVRAB+0luBZxIQkFdAIMmRa6wEMIVSFrecvXUyq1XZ7X1qsk4ef4MAEe
3egPaIpLx4cAxSfpvDdY1//EHFRTzpP9MODxVsaiA5dY4rxwqX4Gx5bZ7MW5HP8Z
YgTAdIGzhmn9btTX3N+QmSmq4rNoXFXI8XGoTTUtKH9aB9czL6BJbDXaDlQL/SVn
/0Pg3holmtondiHG5DmHc5tnQmk4cuYKTGNXknsCyoUq3jiVQWh6u9IGA5ML1Ipl
zVUb10/942m88ddLeKxpwCCyqDaCtougl/68ljGvZxj+fZ9QbBZEN4PYqp8nnMhg
hMKOcvj6e7EykTf9e02P+ck+tWM/6kny01lpS5xMmHtDnK6wsZzLF7guvM9oyWmy
EJ87KZ5RkuRXS7EjFgjXUL64/u1zJXKee1iLbSXK2edHHViBIrWXMWeO/Lkabtps
1+maPQQfljMRF+0hESCzUf7Ga0meEo2oBvX3iYyequEmoeqagzdQgi9pf3dXw6rc
5JHE3VAhfdxQ9+00n9ZlOzxTLeixmTPZUGH5f0cEm9AG1NqGCRUBKU09mYc21Cn0
L2xlrSdiSih0dkDhVxa+OEb+1ITTFuAJi3gfTYcb1nAYyEi/i0J8L4DK6PSfcdps
MsHfi1vQ0Wba0/kH/q22NZL+nPePEcmGVnot7gQqX862n//ouvNrMlPm9A/9TpHX
6wyt2yKTG7yZ4MkY2AxtmWmVdKeOCx0bLBuECR+tjwbdlAXqMlFvjGs64PIw6t+q
aHb2niAweom1MF4R1dyVX/JEBF4sXCyROMSLvzXjAdT044YdiH+ucrQhbddVMfmU
fPlZ0JPJyqmHb13ytshxRVXc/afo3H3fsCftp2f35qmv952sCI+WDAk2Ly/49Rl4
wdvOKvPmVLPJkNWdU3d5RKqExSZksOwuI5XLeECJJM0E8ZtUrZ0sXOHRIF5uF5oF
fXLAF+htzvs9Sf1w5fysFkgHtSUQ3zDYSY+9pN7GjInU7Rm/F3dC467nVwbvrCRm
5Zbs4URli43cHdp/iBRx7Yr6ehcB0JeR0IKeOv0Kd9Rdex3L8+/Q8AshpnWaD4l7
/llcV5wxrjRLR4ygUVLb/11DUPuu5TgNWX4gvIZfueesiLWD6EXiXdMqnlrjYZb3
maKwrRYYcabRl/xh9HZDzuAi8zuEnvIWxZrdyOnop16S0v0n4WID5FAP+V56hfK3
y0/SlG2n+lcG1/wPhymUsuqM4N+2gDgkXVCiKY6LIUSDAFOUgYBeiQcHxb4kLiN7
HqJtyFBFRYlMShXPtKUTXbcd3l+vGyshyP6fpwEiOdlVLjMSsj+RFSqBbB6BS+Ka
CIoqQpzSgNl40YX/5YjZZ8PAuhg55xA+DaafP95jZ7A4Vz3p9R+CSUSylpzOKw8x
nX7IMvP5QnXNmqO3koLHN2Zd3I1hT5bUydQzsO1t4tlaTFnWbYXzlgMqxYT79w9h
TsDTsCvRTLkR1kqYaAMSRzrwEws9ruHX1ZqpmlckQEljp4fVtuNVLQN/fZS5TSIr
2FRlt4x6IC9MlT5H7bEN8VEcNriqS3aEbTCCFH660x6rXTxedsDtt/cXlhf4AMIy
7kN6UPeqOZQfrXjB39HUIANdHJ/60n/DLSZw28/ToZcPnBSeLhzUO3gkh1UsDQ7+
APMxBs0bXvpOg36Kh2PgrySxl7tByit6bwGihih6tuIgPt6n40NwA+o2CSjvHGWa
rHZiMNsu0rhsjPTAug2EOpYJbmtUPoROiH++5DrzDFNfG+VzmM1azZzHW++BDYG8
tQ+as63sVngFSwElrWqjAtRm5GTgtsLa4+62ZbNVhpwR4GHFzEJTWdfbBpldL7Xr
/k2U8xhr/g2cvwefO9t+gDL+ac1lBlPt+4TIeBGc98CKt+Wd7gPVIfKU4dyuE1YK
cBNuaAJKtsfAI2uY0IH1tCTlwe4CfdFUd+BJL7r2QEn8tImNzdJ9KJqQEwTEprhs
yGCDl/RSzhl8VYbKE81h9FiVOjmISqQR4VSIVkA7ePxApu3gQXfi9/nWVkd8Dc2z
8vcdJdwAN8Dv4wVqtKtVyZ9r4vVIT+3JX+zVO+tNvPhRBs12SzZXTuc/nI+VSG1i
emllFSAOY/viA0RbNJ5N6nKzxlEUHld7jxKMMovHZo8dGJ1gIMmAA4Q70lTjBzrK
6bg0+czhyTkLteXsGilQgFdqheWv2IL7xIzYnmwzeRA2CpbMmQ2ujPnf/SeJ92Wm
qt5NGiyxY76tBZ6Mx6aNT4O/vL69OX+YXyvtsGi/VsoBe0h50aKK6qCqkLwsuGzF
4WFKY6M3sK4WzhPWWoH/yh41jyS5X7Zpe/KkpUd3UU/N4YAxfq4tmM63bzv1OVCe
YwdhuyugkTfc1g8YGD0Urg0Oek83ELn8GqRXJmH+kSMQcw+LmAziQOTihhLvRN6v
wNao4nUywiQ3h+LwpR5uhIa2Qkwu/PvqM+W97t4Eee/NN6j/Fcj392h3vNGiGE1O
2wriMJkk6qJnJBTsG+jExd/pGBtHjholGdhirDiAZIMPCCPKe4M1h74APUiaGl7c
pu810PSttX/xCLvQ8XiBB0W0W57BsXi+7cTJql6lQBtcpQYo4ZQKXugLC94liFkp
YsgxefE0XqlvOU4tXmZmLhnwl4x9GOuaaQcsn1YBtmeI31Ra/bZufPzTG1GPnwhJ
mdoG1KeT0f4Vglw8SQHuW5PWU5quf1LRJiNl7fb5PcB+x0wHiKbRJ6pmOVKnWI0l
iWkq17gpkyjkXrHJqKbCtWpn+ZLQy4S4EPUgaj6RmoQZ81AGQionwR2ojuj2kn3n
xW+Dbo7sShsZ0GSbNfrfbcxlwIIFLbbqhrRgAPXlSnRHDgpZS3kuwntZSNdYh0Jf
aWWyMfipX/5oM12Mukw0u+uYwokRGOvL4GzNJs6KBY+fhKDhMkJ8Q37MC3nGEqKg
VQwZAqNdzinnM0CBqDOm47ozVqDTSI++H71VkPirwnq0ZtqsnUY0Z6NEDrpmcElY
qJDhIvLtCQjLY9fmaUSYv4kRD08QTVdZxvsIT8kdbiqfqMaQqpc554/aXA5mJqm4
VM9iB32gW44aMVwp1oryhJS60JOVhVFKZpMGYH/dwVoPCLI+JoR1h7hUcqvFjUIl
GYc3+r6w0YmigTbMKOVfz7/K7bUSpf2zm5q1Ue0P0AN0J9vVV7SgJOqu6x86G92E
YcoHNItjO3YsF4mHI4+7j54HtaxS7tQObEEcyzVoiFi/nUhP4HmX43I6Ot2tJruo
b9PS5IhK+YO2m8vs63rTGoxMLY3SM9cRSCHc0iVdAU8H9SlDv+3XhgBFX9VwKhvQ
AKgSwyXUzREW6tO5nABxNIENVCgaDbUtMlbo0q0xf12TcqI1Jl4HeJhPcCiWv+H9
YIjwckJxIGPzN11s79okOf1FQjGEZZZipKbY/XHD96TRWesFdsrSfdem+ztDN6pW
zIjG2pp3jcKgGnWNrWzdYtO+HteVwc5PmIilUtNRTfSq/7MtAMEBd83PNFaTw2i/
MjPfCRChbEy7065LwVjXPaJHhleD20Mr/wIocaqD6JNPUtRtlmzDWVie6ZX1aBPA
pXxOnWQQvyZPRq9nLMpMDJ8Tf1DUEm7HLrFQMoet65qCB68M2ZyExOB2xTxcE8TX
Eo6KnaM36Ca8FHoA7DTw9r9BLppGobEDty73kgBvbXR6JO+Z9ScmW/3O+8C79dOm
HFrVd722marP5mT0Og1gQEOA5KZ5wuC20Mu2odkXDCLKfQ+677J0GbAoUCv5dKnp
uog4YKAhuawER36JjMawwP67ucyP5dgBPigDDZPfBgPT1Ibu7c6it/rkJATbAaBt
JeH4GGZ0SWWvn2QfPwI/Rujq5S6mH/JHEFhgWM6TcLZYOziBFo7Df5rOBjHtaBK0
orIUfR/c48ur3qH1U9VKvZRKiU5O0ohgrhLFF/aHG6h5E0Wd/gPSYjFmSakloOqk
7pSJgMmY9r13BGFkRH+HspbWHS5vf2BeZw8KlbkBnG0coVzrbaVwWc0e16W5uR6V
djibPpgCOEfyvRZLbr5lWbRGOVG4WBq8T37Tw9wVmPeWV2fTBXl7VN4/6F0jsUfn
OFvFwEO1v8YoWgOYiVh8OQoJL17xfwuK69W/mzFPTbYkf7maJwIe2yyHYif6bBb6
pBRSyQhUBn8zZQI6e1R8IDAUsM7OKM8RjOTT6euPqVIp5D+LHJiKELsfy4VXW3e4
SluopjfKHwju4RF+wmtGR/aEtVxD5Ob21NK5m5K2MYLpgsn+6FET7QnwwKN959eB
1LF2zSq0DI8gESoP8P7WCpVsT36SlDdShVqURIUqi9U6GjkS60NipCO3RaKnFfD/
2b0Y0HhAnLQCvxuhB3XQuxzCH1VNGxfHiiGRwEvsQL01ry+RoXnAooxG09pPtMEA
AePlJzW7q30XFtOzufYIsk1AFUSwmIl6wDo1x2qAWDlqujXBYKNiB46PUx+0XzV3
0EfVcl4g3mMFnGi+XT48BZzZ0+6R/b7ncBvHaADxcVXKifvx55PzB9M1ZfSR4H9O
jreGj0Q4XRZmAfjiIihP5nLnz8N4WeGTZNQWh6SNTohZCHQdx2ERBZD0hbunwKlo
77R5Fm8w99FS9lw9E4vBkoraT65j6t6niBNSzzFUQnz3tFxyfyIZO+n/H+R95zpN
ZMWPz1c7HXxOjBC8fDfY1Kf8JTWlTYoJYwYCG4XzAxz26K5n2fqIcSo3XE5RGTJS
HUQk+x7Hqj4eOWEm9+px/X5D7PQLgrFC2+arbPqFuPSUZwT893GvyB6F402FTTY0
ZJzHjUR6v0EFfNtoOhoAVly5m1gWb/7x1ly4gCxbvupfa/+72WmuaP10rLcjHwbP
YOHONc6cnK2o/9y+JHzueNvhvHeotfDd3ZPAvlRPF+hfokFIjd+lVeOzqlTDCfH7
sAmnXVnOuzcymKwrQ8vSQc+L6r6WrbOgJF8rPqGpXZNiMCul9U7b0yQBM1QoSwGv
ZtMWg1q+BDBWzFoCTyLt1t74vFFxZoAE2D+y4EU+jDcMPNPchqvsZXD+viMFbvA3
Hjd0dcs39hxejU7fYy2zCTGsI+RQrfJKfLIxQT0iH/1UqBlxyc7W1ZfY25jXxAQI
aW89Q2rKYUuE3ALJva89wC/MKPxY1ajRkDW8RO9TVk8n5AjxIw4DppfeohK09V27
p3396slkkyHWTA3vSXxZTESOMkShmwDM6N5xn3VsWieKIBNwLE+Ek2x6CikbZb87
Du3UGOfq4VSBFfRbf0+oy6Ww9YOsUR2+ncEWzRxfpiHrDqpFVRpaYeta/yobbh30
WO1MjYBhMJxieClcUNqw9wQWzIzKv546nl8/4CaUuo8Jbp75NlGtQ2KRRHqpGlfr
gux/g+w1GfKk1UwXHFblpMO5yGLrRwUDd2cT3oOuUPon89Gr63rL78uyofcwlt4W
JouDnlGsOk/TC5aw3XQwgWf+RSGJtqLoC8bSq1uxv2SrSG7FqP0NMfSqeqgKuJPS
TeBE7VTRX9SL4NcpknX+z5wo2IdG+eYQXm33Ez+9Ku1iH1XgKLQmNBpXI5/GZW43
Q4AfXym1Awf5ufRfQK01nUPbMNZ/WtyCwkTnUlDYGxUM/R6465NQEc6ArSfug6GL
iaDbaDJ22j48rhz2dOR+zOEw2Vqv5mk7UlY16FgX9GTEo8pCYXEcwqNFdd1NtfZO
Be+oIeMLX+MpVWV2g91VIr1oYDkTtEalGiYPZiuvXiJbJ/Ji/P/hWuCgROdv1y3K
A7vMvwQ9ZDeZ5ZgAwED9qW039kHQBcdmXcEsgGBPo0HwlS53NsSm2s6ia+L9K04V
XynL70Oo6rcv0EReQIoVQ7tc36iR2mk57/B45Rm2BV00ikcGwskrqVSVGi5QIwOo
PciMlg2fPO80xO3xd+j9EQnZNKgmx4qhvfH6UzFHpQab1Vj8aVEzXbu0LFTMVD73
69iwZeNWvj3VArC5q9azk26CE7STuckpHQ5fe1Nb9zxvomsFGiY+eFdw2syxCzx3
U+DK1t2r5b7wRT9kdlOgby+3IcG7tdfjVhiqu6wsZ2lhcOuAqit1PFwc1di9bwxq
5y7ycKkaiIrE7eTTKQsT2+zKL+5rCT4+j2lTGCgDmao86fKSkRT3X8AgOYIQOk0W
NxWlWnc7SGkC7E3vlSkfUC5OzewlXuzSZubVoCe9BBFAKc2xbLQRl3ShXXZvGQcV
whSywLq4TrXU37hLId6kAK4OXssANhTVH969B7bqinxiBRx74QVvl6UCABygs7X2
DZw23GPNWo0QHIwm+ctR6xhak9R3XXnFyMfX9a2BLD5S25mS4Tkpk3cOx3LoyeKb
Ul75Otj6i987pBZmzY7MvqX/mUrxkuOrret64v2NBAnMRV8dLfeRXEw7RqtPnSzm
pYJsT1g3zLm/Jxi7YY0zb2nI+TtIvjdR7kBlpa4hV0vz1utBqXnGdNN1/o6XrMmz
JX+HzeW/3YOi4hEdF9ceXnO1tXZHvZpY73wYyZuQY0FqIho8kkNlEZY9XjRVFg0Q
F0sJ1jMbAuEkUvDdqOWkSvlBg6eg0WxIbTzxbXtQOcxnaNLYac2jluo1wRKuSABY
QR7tst8BEVfRj0j+o1WRcwsebK0eXKJSxnerLWgIpdIcLVLyyrpOrx6PzdyzP6yT
nHCb7OlRMNU4aIqPBNnAa6khEbZgWkUwwO1FK9mOWDl91ltSB7MEbV++/yfiTDiO
9QnqAQ1jhskv+wlDJv4YGpn6MD9iO4wl2QjRPZLnyt8ywEvY5VescAFbO4l/mu0T
dPiiiUjgPVi3WTCNwsxx5r5eYFGOSkUzG8Eqv82R4ES7bX4J7ZhAnW+Hba2MX6wZ
KK8Pn5ED5tHRP+sz8v12LBDBGcOKcyVZp4ucW/XMAA8ok7yr1gE+UoaG/24dB6VR
i6Cp1EHx81VnYj65A1uCXbXbuTemAuksLMAuWpGXHRY3Dm7xBOXy7wtBClZCziE4
T5R0WuEGmcygf01atAdul69bR4zQXjS6NIAVuhBkcApzCUM1dpwNymZxr7CpnZLi
us4yV27xgMv1QsUQWbViGIUbTHJGW9T2D8Fvjqjuc+ic3RELeucDc1xbz0No2fK8
mwr5bRPJwyTOdMiIfJGcaGkV59/GcWrvXr9HybA9KnSVVcIeWT2OPs8WHw5iTpne
kIg31uFfPYp5EzJ+UopZL/q1dKTv8UYAaaKO9u+s8+09dCEw8Ahr4WdB4GRfWi1L
19qC6y94buTZX6ScrXUTneXUKNnJMxPzqSOIGgVSc/1R3P8tcS5t7on5gQDsTM/t
mTNllgjDlpD2gGgjbsnjAFY94o3T2P8O8il6GinFo8948lHbwBdhco3Z0TvyaCfq
wB7oZXUitGGiXAkJCd33YyKDYNN6otAgGc7IlSxKzBHN4wz3Eb5AUlMr/49m4Zgp
i7pGKZwU044KHNsUXaF0ukyg3ieIscbHRYE8tr+MyhySoYgLqXJZQk/96UEpaa3U
WaQli9ZBX+nB/1bPobYFqMyPFEdiBEQC1ZsM8IoQ1kHDlSM8PY7KN8Mo5ajdPbss
gYWeXKaUamfL1P79BUDcoEPBm1uCjFQ0/J2MYXAMj0bQsJEmTf7Fl5iZOuplVoNX
uakQAPb7o144q2gwky4buqqfnmrMeaDrudfNvHjAf/5QN64FZN4/mirCzSkYbN3Q
6NKGbPtbqCyJTi8MPZfmNJDn2DFnJW6hOmbjKwSB8cDmffz27ClBmKNcKl690NjU
1wKBhmPmjX8WICaG99P42LQ80dBOBM8O6oL9nLVHpNrY28Hhxq/N5JaW94F8hjgz
lsvssTybejG90U1UVMRzv9hHZv5MfZhH1qYbOPZmivCJlEfKBFtrECV64J3U7Ips
a8ew0TQMPEc17nshC1djSX+i9CCsQj9f9Mlo7o2VNgdUKjrqiz0yDHjzSNMNtxy3
/UcVmMoPwYldWc6YqT+Mk/vj3EgWNEF+QGhMcRq656EPKToAMH5o5OWV6MUcQ29k
XxxFp5YV1p56ftUnnh0gCnon+Xlqkjzulg4ZwNYWRvj7Lwu5TdzGdwaTCJ1sVrYl
IfFg4R+kDNlBWZQgw1vwi203rTRMtcKfkb4JF2HNx95CYx1b465hJv8Z4iMr3MNV
RLjzfIzks3UIo03fwb985OxmELk7emdBdH6bXCwx4NhNq5fK4UNZyBSFRtBKRawK
glUBV9VSFN9VZ8Rxyp0Zz5ajOUSl6eClMLYOrXUeHAoEpY+8wNf+1PfoPlpRpedA
DjGlbml7MDVGthSKxafTJE5lPuJgTCmMv/z5dCTm6WUvOIqc5trT4I2crqkIqdyW
DSbaQrd/sRGmYqZaRFIdZPTQoI1oK/zubaWDUOwnGDJ2gLOqF2NxWQtdV+WgHBWm
mJb8tAHxiJoIeAXOJ2nnQ1CJbngrRdnl34D5k+n+GZfeT52JQhFrqf3U7DhlR+uP
2PjaXXZZ2VF+Zhbz5CbLNS/2Rw6VDBav5fQJySLhV3C8XVzBOxSUdcvSIFME9G9b
h2TfDXOFlY7Brlhu7S7zeJ0q+vObgOhiaETrogq2DY7zZNYAXh/Lu7qKI7TZm1v7
4qzx/4UFeXr8ovQ8+qpQOaITE3LQ8ZhtKuS7vOtNgvb2dHGeAoCrrQvLSGpkO4We
o8d9mkzlYcrgecqZt8bgKWmLy9y+uhaQYzDukrx8KZBXXk0MuC0vBVI/t4rWKpZD
IfLyU66GUCWQZMSkFSdSnnTE9xObOdGJswOlRAWHoZmdKeWVVpqjo87Hs+vHihRC
rvQAEbOuzaUGrknOAIhnOkQEScjzEmriP1oObI+mOKM+4AVDT/Au9htLZkAS7OGc
1LjwglDLYP+XdHuQ3xb6JLASDhWfS4dA7Gwsd5Fghd3AB8eXMM+W1Ocu5kAFfIsA
/ubGE5Tht97DWk9T7O90j3yu8m08AsYUCX44jLB1e/fnXHEGXFx9+g+PasA2WSCy
xno2Z4mZtbDT/7tjETULDBRGtXIWc65XTz+v5mbQD0Tau1tR5JjhwSlk52WWDG2U
qjfpPh5Go4HwrZlB3hHctsZ6MkWP8uqomWuAoBfHHWrJEAVywzziJ2Ka5UtKthJ7
FKmfsUHPeDGWg5yM5JOsHKAbu9Z3x/6UvsjD6HMD5GKetphZDINP4nBxhgJvk110
lzPwGW0D9UvFREZ55SQ0pyrLqMrTkLUTJjKegtc4RJF+QmAbCFz7ktSleqBngh+A
pfKJp3v16fln2qnmOFHYrqKVPwZY4Ck1/PGFQT8jOqMEOnThkVr25Bis3Z9kQ0h6
31j9UnTMqslLgkNcucdHsypgXXu8AOmxu8QOEKPRv2jYIrc9H8qDZh2+1XW7jNM4
BZVdGd/y4JD3lxVVEbB/erjAKMG8lOJ+jzlb6PJ7TfRMzmnHg+Q6pD6m/gf6J/Jf
P3LRee1m98MuKh4N+cWK2IA/2HkajvbpXoJCZfAGZbXP83Syv2FSvCT2m64bCVWt
OFasEEgsH/DIJtllLw+t09ftqCHFTrz+jm49Vd5X1vJfv6cZJvD4I2aXTeCBoVO4
veRA10rZXmvf6EB/au5X7QmIMWHUPPO94XTVgIdc5MoO6Neh9Bzje6FIhROwWp5e
B2J/ZXBLXBwTp8JrIGVt7lpVMQx1BXznFJvWKBgorX7biQcCoWL5YMbtlOUQTHT2
fWyBeuwJFXlk7xsx9XIlMN17TJmM+7HjtGdxMJvHIfxqswP7GOBxbkdZEt9/a2Rd
3G+59doeH/COtootz449+d4COUJFztBniJFZSHjomlm/lV5AS6TNHBHScXYFl9AM
CW4hTgULISodnYF8JzwGwFtYP3QbXGw3aasIx4RyHgM4n9z5iz82XfioehYRHSXn
9TsEirC2NgU70NZo9xj0GvItD0/MemRPmxYSM/AcqIcJFpAzbLonSQiy/Sg8vBoa
GkGnh8pmj6WEu+yjybCd0B318dS2yIgSqCFreDuuhWOFjU7J1T1Qj0/1GxLO1P8E
fFl/yiXj74weH6t7lJkvYWnexqVr9ZB1w3miOjfw95Jc0OL5SnsZfl+y2wpqwxlt
DsujeDzrPvQQtOhHBuAhUoWxHv+xLKhzkEcOLqOaLKZXNBTYeqeBH9O1cRmyiNB1
tjmEZ97cAaC/y0krRjXPIBozGGEk8cf39/ewCu2jTBFzGCLYGmARBThWEcHcUeug
V8B3O/5uSqQYLf9l0hOrVFE2UVypJBe6DetbFOUJsuON7jo0q2UbFcM87oZIpMGG
IgkFok07rrwX/9xV1InFe0IUPV5BQJbu172ryc3BkfFZMRqFX0ZEwQajb22qgYQp
rBuoMYcF738xtuWDBhoKwQMUCE0tK5HMnMKFKoy/rF1nTDwXXTLLItcyHwL7pbSv
NWGM5/Gxhs0+INIuL5lOWgdjEajCBC13aOoXdJBftso+WL/lLmfLF15DVwRpaEyo
fGmETN/4/JbR+SgtPU710PdJos7uUVfB+LBybGT1/TnNTa86PlZGonQodeRZNrHZ
wwxgBYLAC733KhtVnX3RkQ51jXJ86al2P2yJSVGsCTWU5TflmmgnxH13Agp45NKr
1t95fQfwfiie9BwrwgtNtPrUWiHZ4gNVzjROHEbumOkTqWJMwzBV9bS2VRIzYnm6
84y0+8Ntd+xLbeB9PfgTDry4jRVZhoNWmFwSSRDdcQEKiBn6eFbY1bZaniUvdA7z
jA7adUS1CdElaax3u2/NWMIu+MV7i0dde+SZByk9ouObAeWId2liSJJ/32mhxPS4
0oAJnPh82SalyJHoLzgeNatD9SjfdEzU0svP+R/b7Ff8b9dw/84uTxAaDxSr99j2
kyGrMvWFt0tifSonxyChUE+rMTuRxY3a31cc7vzu17uKX0XDrctvyOp+Hwx0jS7J
GxAphX6YCsa6iK6tnog77ebXKn/iTqFfCAj2DrFfxJpcJuOmuOpjuKCVyWNTn+ef
y5SqN6ybIdX1wbGVBfHFhUhVzzZyP9g94NC+FbNf64P8a9Z1kz0td9PPWGdljGNt
n30JBUeWI0cFgWZ81Ws/ydMgub3CjLH9J0PFT7dbYeGIIVblpixhcF4g2MQ7OKPy
hWmo6lYoByWLYNhgIWQuYcXuoStGTNgLBFoYH5z+6sGgo6W60cbbHFU84ybLBBQH
Gt7uk2ZV3CZv4oPiMT8w9fQM249qJBxHFDS36O0SYM2utoKKrR2qLvSjzVAVAtvD
gtXJnWiO1YY538XD6EW4Rfq+OvjXl3EITMp/Wz/LGyZ0kzI35wFhaTgtDHbVlhJ2
A1rmcTqM+0H+IO07duGCre0cyW4Pfqkbpv1MRrxKs2BHzJkTc6MvOpw3dqnpXW7K
BsmA8lhCcd7u3lYCs2mFvJ+YFOGq9OVz8jCUUeZurwkHXGkv2fst1G3sBppcxmbk
C6iTfAGW8jzbHHDRqX5NV8w1Fqc9cRBa4Irg4al2rHH+mG+O4ru/0sOPQUsakxYg
dNYCYFFqjqg5RU1LFpiQi4wYT83ccdEbPeHSiDwU8WJeoCgFKdMth7WZsvB0cLTd
teuKoGICO5QMCoUZI4f24o+G1SjU2Dypai93qRlKHBUEHMOkp9MeBL4XT7FBbY13
RR64d2i+tXSDHaLSITywYgjPFz2rqLUWhsW2Icn9Utsp8lV3/GYT4HIvjGTFnrau
xHKugfje8aUWy7Y/OMp15YzFZ4mIrwYAZpeidrdTp5sMlgQKLaSnP7tteI+l6rlW
/9Usl0vcjhDyrb0nx8XlPBunmk3Yo1L/DNXghWTDXawlw2W6/O1FNcgoF5VsPYiL
Kv5fpW4hL3JVjpDMvnsp1l/++eD8g+Ps7WmSRcXJ+6Ul1ZcO84iVjsRvhWDtPdO1
a0EJeKP1eoZnPncb0fK+WbYTMd7d9eX+z+nyU7rcEOPK5R4pAdMuHKYwiqE+LIwE
zBHkVAMxqUg+HXkM0L7Nvz5MsDUQga5ppfDMUyFCp5N8fhvHdkRGFdGdOmKxaV+W
bvelsiiG9FQ2YoUL5cO0M2AdyRZpnYGm2UH0bzDz25kthdC5eU3J9rGKB+h83So9
nJwA10ZStSyZrE2eMmwFmDTvWrL+zlFX++evkkAwsZsd/1wB4uB6Kpc8yOcwQ+qO
W+Nxry9SXm8AyBI0BPdd2TzQZIoG1/Jxc7G+6HmIewDi16psccpiqpAXDyYjklZ2
U50U8dInNnmUQwGsbk5euknXGkUGP/oRsV8L1PaKQzna+/YpnUYdRooTsaaSzDjy
B1V6f+zvj6GgfquYqPU8eDCs0nezDDUesesxKYOWXtw8Z2j9JdpbfT/NuS1LV4G4
zMVAiCVQ+qAQ50+JXkoGWR+zT2hPnmkf1wwHQZKWzE0gUQjDwh8i1RRxSEU5UCxG
PISFWz2eGaH9yB1Gl1qfoFbnjVym0ObKNxEfFlLOtI/n5oWhCw1IwBzomq+ZPaHs
S5PIAVSaB5KC9Xz4NMToAtBwQrzhbXLhUXAQ3Z40A2jet3AFkEI0AOle26+9LeL6
IuNJVS0bqLRIiNHxxfFah8mF3Sholu76X/O6TwYn75OUF2R7H5UhltXfpQeChXll
/KU3L31YdX0CBwJvsvDZekQ51NtDCFSBTc4pZGoWL4c3I1HTj75iI7Z2d8X5ODXn
4Uqs4JVCHHurvrVnhJZ9QD6cKEAUfjUa7xSQFwQaQDXnoVAu5dyWYADH9K5FxD8t
mmyQFY9AgOLKifZ/o6Myy6htILPIckimeQapyBgQJ5Y/Xn8/fbusMbpo8iLZuVtn
Jld7JYULePm/RguLRu6dO9PhUHCgkRMMs4dEFSI3kwIGdMfYLrh10oyDw0hpUW2C
+RzJ0Pom/k/iMApEX9fJhGMEv10Mp6DAihj4RjA00RTAcFbR38/vHJWlnAGCa/8+
OVD6fPv02wWYkn8X7Kzwqp3XILF/JcEUNE/YSNHtHPVSffntzwrfY4tpPJyRfoVd
rSYcHQNOBo0DBG2986VDMRiGhNr1pkvxf1DyvGRjF7Xm8FguR/PmD4+q78tfDZGu
QXdvl8uOz1rL8TE/yzhoUqUXHMcYjq5bZdFLScBoM0bU33F/g8kYnRD1v2Vmwf+h
OE6mztoUQh+n5lFkEh1m0nV3zBCaKLfPgfqBYhaJo5ZWADpY/BRkKiPsBGy/XJMP
4RIXpBZTeIETxz4zXwGrVYciZmu2iygtu8sl+JhEwtEsgIdeIu1D0mjQA2QNJxW4
NnxYBQ6aaLw4lyPSRrFjndVK7v5pNV/6pLAtxah47lxUz4G4X2n8y+gkPRMNxGvP
HV9vjcyDfVSl3zBew+E+mBy2OJIeuLggDJrgpPfYDMCMpJ5e6iEpXCsp72ofIleR
nktsvvyoYJ42wLUU0/hG+Pzek5Oc2S3DxH/mr+IZvH5GRRcVC3gCaxzQn//Z18nZ
PX3wiIJ/ZtLs21OnzhC9hVRTtLT2JVKDnIwdpZY7F+/RwRvsWGlLa4VCutzGZifn
GITqHNlXqeAyFaSFQzF2+2VDHeCgvlbvhbx+yVwBQ9wfypD/crkHd87q4bXlKGDd
zozSMt5NqboIGuSWXqVVGE/9GkX7VDvbJZYEtlWK4YyVm9Dfd4BjBkiiAOA+AyyS
cZxmn9ycUGD5s4KXwo9JcxBvTq/OmA05fdXgJEVhyMcz/gYLTTPZ3R4LtIltPkwd
/YmgtEHeOHmWaNx7ctTcg3eBMnwe3didyj3fwIn13qyi0umEmVbKThRcpB2leSJG
5LHP2tp/7mdNS3O6XxR/4yJv+F0xZxXcWCzB6tNkW03XlDIkx+im6RMYhtZBu22j
Y6bjVPJap/PNwZ2rfrzorxZAvgi3hiMIASEF+r5Ox6I1yQLK2v1n6hBGb/Hlmkrg
H3oaJh43L0gkmSMgOlZuBGCsMiyIDVA2qBc9UiKWKP9XRhWr4EbbYgAX4wsciOwq
W3MedK/tJ5LztFpnpwmcwuzemmO+JZ4881tbPkOxv2i6hPXF7shs8sndhpnxDkEH
vCzmH+Ufz0/QFvzGmUimCt25dRrhU2H2Wc6Q7Sx8FmCmWHQkC61AN8wU912HZoGV
lPEEhreIiZ394rRBYDmiX0ebGdRxzARQFnyJQZuBsyb43/K1rlkok8tgshLe3vCb
RDd5fHOSDYYg8n18vateaCklDKj3uf7YEX73BXdllHA6nqRBHqKOIWl07PWWKcia
E6I/yYf97sb3kSm1j2CAT9Jj0xbx9ua/IKY0yjIqAB0Yq3V/LJkD86nUS93A0sSk
V2twlRF/zYCTqks98gL+IUD3JbFvKTA0Ivlw/ae2megKZzqc/pcFJU8YWoyQ0Pkb
nV+DjFBPvMcKYZMJwH1ulmAJyaSBiv9+T72a1vnvxRU+oeWiMchShqUSMb+rAiRK
sXN6pAuObekKaWsocqdTWvpHshBWYcXNiLZ4aVoqYjUvsVCcLrwcAaXT/jgvAZus
Yu/6jW7fyGuhI/Hs7zK4pmDV5iSRHpWopXtg7Ir8P7Hcw2Y+roVnyKD0VfeJ1D8U
6bf6lTB7oQFI2FBIfydjqOe7vIEoBnZJgQjWuq+725w2moYaAh3/LZ2hOZM+R8Mg
0UOY7kDUjR0ktn/LmkB4vyjPhBRdXs8ohflLI31vgoEtX55UF9L+IMJug9TCRRdd
2C8k9NK/IVIcCcmI9drdaN72EIe9EvWhTGIj7RVYsAdWPn+rppz08X35KGda7rto
6KD+a/JZinT7RTMc11xMbkgGHT01/65uSZvT1xUDOyxLF12o83mChBzAyZCkJmoE
sIQAgUT9CBLA75SXOMWpUuHRKCHdIi0/Q3WxpM9LsDSKL3HM98m2ta5VindK8VhA
aOqSAJYcNFj3OfTbpjcIcSz6E49RUVqOFNN/r6a7EQzETI//7I96bQXgTpIxDAN3
nArzJpXdCxZpH+zxPBNVrWszuz2e3vXHh1ibdHyAZmGWxbXbCpRuAeAW7FBdzlFy
xcqFHjbhIwZUuHe9nTvGs9mfLkvCXUVkXX5Qn1MwBB8rjMqPhkDN4bf3NaLTPJhs
5ZVT3n5nfJlMzchm/2JuMUaAT0HUZ2dqZvbse3qGLhRyS+2qw7PiFdYfH1ceXHq3
IZYlD7vi2J2JyNMAaA0d+ruf4H/myHBUFdB4CzVdkC85qR09GJ7bQjvPALRGD7H5
9ADIcfDtoMYI3BNkKgCePa//h/QgDvB8Rx00j5i5PGYGk9+0QdmTFeOrQ4fba1Cg
nu8fGCp16PExm+izcAoLxOgdj0yRDu++Wj0NXc3EsdkIPne0PZXjb4hhdK0Dt+bT
wiKrIf+SOUMSJRisjtDjlslURfDF28PP6FMZ7xkLsgSk8bjDyR9CNfDCRt8HDnoC
ex/cQqdjj+iIbDic5B15FUHmw6RffRwiYVBV2ht0fMcPkU/rv+wEVY2BFEvslfcE
CDQiCcRcMAthYm8FWtzDjzHERwIpk/DjFU55dszFKTOrloj6x01D8MdRjbqyG2Mf
7homAYjN+ZSpkUX4OnBWjW6l/zV/JJdMGLrRpH/EeTQ/KKgCZgTFsVNmCIkKd27F
apuR9NmBS19MgqbI0wvwWsBfg7/xA+EniWSxX7cTo+UXPgCeMtL6v9mC+3qKaUOj
c3YEY47ksAgEwBWYhmpzJ8KZs0QrYpXKa3J7lZKsDpzsOYSobW2F8ZwLDRl5nM25
olDuAwYZMHnoa85+TGz5WN8bI0OxnCOBXOsMQX9WTV16ls1VUv3DnKP02WOqgM7I
ET+ougicbanAL3YF0oM1YCgkxHti6jXmP8Srr9uHmzD1hlaAaIoSZnYWesxMq8c6
4pNNbqYM/bKLL2P9cawyCxVKOTgEMrLZp/nVIxTSCkerQe5MIjFmYN2+lYQf3s/D
Hc196skUALu5CIGf1lO2+ZnURKxu6EUM5/pwIAfSXWYKUWO9+epYAtjUgMeK6+0B
kQEWpUSu02q/FBIy1Z7AJC1WrNYJmhoRzTJOIvMAA8iDCESh2xl/heVLP1UmDMNN
0uXKAa0Ovhl0p+/Jabkk+8uMB1+YnBtSORkPkdPSJap6BNlq3Cti2o4Hzj8R+CN7
riQCufI1OvLQkseyYW0DEnwaMm8QfhwDc5MMbo0EbhuRH9nozKikN/u72S8o467m
jX7wyx5qAyMhDIORar8VBEsgn5HY3/Jetly+GGKjXpSRahzbgO2UmqvGxSw0klLJ
IoGBeWbTSpmjDcX0qSxZk8CTcoYCB8MuB+zlgN481CL78+scZLWRS0u8RF5OVShO
k3OP0TSPqIcgMouGo02pS9ZVRmdVhdadp1AlPZ/AOn7ML6Vx18OXPUNeMdxsURXX
rJS3tffDXq6oi/XP4Qe8/6nKkoXaBUoTJmrpQ8nZvIeoXffkHIic+6bM7fJ8pazZ
SQL4BNbYhfV71SMBzW50q53G1H9PDiS9icw7JSl4SPSx0hMl7jReW+JeravKRfKH
0lPYja9BKfRMcMdvfoE5zNC9wIxVUShWg97HkYjhhLuW/M7KeCN3beoAIxHFJZMT
krZA8sLWqeWjKPYzKMhefdSIH2Oy5o0tui8FmLCZ9NQ77iFG/KzcHHw+1QOxA8G+
E30hiMFB+oQDAonDIIoQm7Ks4RDK2Vw4nT/ZMb8Z9TIHmesyzOaXu/GELusiEmDr
CqCox4jqojOy3DnuHOPGTBelCLFAMNzSQ8uLbrb0h6GloaF59x4ltMaw7fSmO7uN
ge2GUXaEciFFm6tVb5a/dIEJN7yZWbp0n4YglizS6vVkfVMiK5rzFfzEvtE9lstj
diyoD6SIcu5+YLNckIxuKNL5mwAYmr3RVKdVU4UCluMRs4jLqKfDpSOZGAZhfCn1
SzIFfeHTyiOZ8kumCdRfuXLYr7ICUPyBt0AbIXnHo2s+YnNTUlWfsIFHVyt7CTyh
lPlQgG0HYxkwE2nODD/koJ2XLvbMOYI7OEK/xR6RLyCxUABB6KB0hurlmZIJIbrl
yEZStFSSqlBEhxpvOjmvfPUjCUnnlMur1IvXpaVqjX/wPRDotOvDnjpWOQ5gaouq
DJIUWBy9DmTw5L57DnNAVWklt5r+fKC9VVYakkK+Mq9IyVCjX+bgkBThb+EWO14A
aACerW2TWTey0SyQ5f109Vk40GdD5popEe8VCke+F13xz1H0K22Xv3sHT32TcWP9
FZo13z3ongHS3qv4QwVaWeS1wEJLwPoJNqoEAxxirxVJjrQOJ8bmN4Hc9IBZ7a2w
kyB5ICaQJkxVwiXlxqfgM5I2OakfXC3UiM4gseZwb7oNyqXfhvENpVkVrIB9ddhI
NUxGs0BA5LZ8rwoIjX4xvQxk9Vq1gfZUu4WcqUWmHPZBarzBNDTR7kD5qbCMQ5sj
YE8n6jcpnO7tUHMjLFKCXdZtaI189oSqKO1fYlvT5itG1eS6go26ifpaSsG4zqzM
ZW817rC5dxTTuRVNLnP0CG3m3xnTnYW8+Fjml81hbfh4eJtuBPOSV4/kjJEZQcZi
AbDJY3vb3kQivhOCkCfVPFpJpZ9fiOfaOs56E+8jjOWnTvpZPcYZq1XfYZ7NSdwX
bzzyZi/7IKPdKgBIM4lmdrGXWDPKLYgrnGO8y54l90fQpbyeQPXbwwymLuFmMfZH
qLUdfHX7xj7xXVcpPeGPqHPCBFa6cOZ50GdAiMPZBsMCiUQeYiSpRLfK7RqCTfIQ
lM+S9cGxU1JCRODQyG+Rxm/T1MdVppFJOUPO7wCnFnZB+VMEgnVmw4g8mv1fKQZY
XmRQcFqEXmZsRyqvXCnpVoKsKSOaGJNxiGpVCSIsel00+yPVlYp3yPyILrdz8hds
lATqvID3mPmNQ4/OBn4Ax/sTLaPZrJuampa065Wzw8aAa+R+q0hc1QDMG7No69yl
ZuWfsRDM54X6kY94tuEFJWNrnU+//x28ibdO05FWxdTry+742pmfpBv4uPJ0nTAY
ouAKCu04zzTWu1RaEsjJySCR/JpEkPQBZ5hWxFmAYrfpiExMFcCWyDIgqEqAKFsz
tG8e1mNMklCRFJkvw6p80ZukcTnQxWvn3YoS+fdYlPeaDZlXx7JZW0fvko7Hg8G0
xEVnseiMCMXKCUNQ2LEXuNfHX5bKy+1nBRvXiYDWkoLJ66Evpe2B92dSC0oVyVav
IKz7EkVc8u8lU9lFFcrRwS/SlVHEmlcJ3I2QfgO7BFos5blkWGnszjph+D/2dWik
QUqqQo3IxPaK0hcugmTizEnWLKYIWgDzJaytxmfWU9SDFzpoLm+Z5n4ZReqtbQfo
TRnkuxA8jWbdT8PVOX5+FgqMBnAWsUTa3Q047eFq896T9tVqGs2frv6eA9PTordh
IV1Tymk32aAc0SlmsE3WqHn0zP7ISCrO0i8Uuge4G5/atCIRlJ9w89ie/hZgPAKK
0CWUdgA329rmadOOG/OWS/eMxbXg4efXd7cOAYh2Se2mWq3PAFnSW++I4scycU4s
E05z6WhEKq0hJvDZMaw0PrBFu7VRXUVYxWkjNdMFzY4jwgv5q0FG0vnlen67/DJ6
B8kGY7kdXyyJFpgHHAnT2H3AneTfNHQehmtDdQwOPW0mdDHP0XL3trdKxzMkbXXU
76QobuwqHli3GUadykMyGPN+eugtA1vF6lIoqwwrt3dIKAHod5/zjVwTScegde+7
7eo6vmfJpbMejQwbb+FlrT+Y9N8dnFeMFP03eA0pucPJzXvv1sMkH0UqqNJUuZaF
Mq3x7SBs5gn82DXR8/455JhYqy1wWhU8hE2sYavukGJEmX3yHI2GaIz04Jv5pE+v
YNugYahb9/7YljqIAvQAZrRCnIOjfCXwVkakDb3jTOpcwtcgU6CDNJsXHyk0/Rup
n7CLTEUXd25bqDpQzOLkyQczJOwixCfNaByBX2afAa1+RvtV4T06rSBNrmw4eL8J
ru08mvR8PkKUaXkda/x0MVhrWucr5zSz20ZynQIb0hEPeWZLhBotDaetcQTgf4+A
HtfMHuegRnr5oDLi/Zxs17meju3h9wJ8cpkLirBHbS3oE8qqWlfOBFuAD6cbf3wS
3q7/wHOFs9FPOozbdRZD4i3BfKfBYBY45ooZqloft8Neuj+ThY7neCxuKlrjkD0E
9+Y7KOQDSX9M7pfeWwizW672xPBrMCt9uduW3UTXWlNTGVJ3vb+QqbN3NX8fuYUQ
o+5FzEYlQPreU/AUQ665ly3uW4/xbEfdurvZYc8MoSkHovCwxTWA7s1dbUlcobY/
hNnmbrg19VU6EHPeh1Lk2kgKpvZ65MoQKoUawadLsC++TdKi0atBFtEr9f5pNrkw
g4/xMbEOaNl8V5sqC/3MEVxC+qhGYgLgDEXmMT5iRQixwTYTX4sO4nQUeRcAc6oN
I7Fjc+hRkdIPnceq8cZSnHpxlxiTra6batGJxbqiL+uBsKp/ra19O8ARqwRi/Ltx
fmY5B2Qu4NIkBt6c+/NFF3I0HtBMgQghe3W1OU/F8SsqCTzFuLSR2t/uSX5sVxNw
2oqHmlL4uKn6uqa+tO2c8bUc93QU3zNQaRRV74ZWN6zdArIOrUMa+Pqhpy15xGnl
ZAF6hRB8FSJgOUhz1TBUGRaojhEaUJ55gF5TKNiAMbaKyswqbJ/oosaBNupzbcyO
h08IiYsd5aLhqVU6Fq/e5zsXLNiWIC7H2ImPxDTN3RGmC5NqEMDd82vZlCwYBvom
dT75cbIbfF3bmLbgN2bbM6LZHU530cQjVZIs78kI6mRos5JcYuAvqcawvzaEE1AY
WLOnJ6LEn4fSJKoSEbaylsp3jGIUsh6lZcgP9yylJ4rRMcOfqxbkqkeunaLmYQz9
p5Mo3nIesz7OF5asGe9x8js+Ejc0sfRM5Pb3vyBRxFtb4qgHitogRF/8lycrpq+N
rt6WDkwVbQx7lzcfu9cqg0U8G1VQEPqxZk4nf5dOiXyDF2zZnv+gMi/QNezFuP7O
olGoxHi3U+l6sv/ZG4rD27A3elP2V1OjdgoNCvVbcIFZOyLIKJmjD39vNFHwFzFh
iP1M9YJJb707X1azVjS8hi1RHcCv2WcqlmplrqiD8YzO2qnrXf9Z8tFGhl54ipiw
V6GpQdaYB3FYaupnI5fTh2HeolCee3kofWOlIaE0JI1TJsCMzUDNjI3XgM1ZkuvB
FvpRXUToP97a+IXnYLc7LSmkc3YXbHTdeZJ9zSSMjw0Ja0Uz5LkzDbbguQbns41I
fyvOrpA00wiWGwb7HGUOp/JphTT+t+PgFKROsvDJr7gyJxQSzDHhRNYTtshSf7Z/
XkFdWSMiucPcm/W3DmmoBGZdDENZTCHoSYn90hpId12fQzstgL7VK6PX7dxt52wd
yrsE/ni8jHkegG6BVD44/A9e9jkxd4LbRasv4kqdlITefLtd/ewSnuROpDJJ1CkV
StBzoT0bj97Kp9cEuaTiH08//jtQNEnaKBVoDSN4Z7TYnDF5xJ7bCXYKR05nAvj4
7LG8Cxs24xIydvvcIIBaswHtaGHNMVuAx4avOEo6DLTzOTdUk/lBNsNIpJq76QfE
2OR08bAZu3DW9n1V9hYDPnZjRk55rC2T4/fImJJ6aWAwVNOONgzNkovIN2M6C6oc
cSayr92fe2fERaxCZwSRocD3EGAtaMNKU3xpIKMLHaxxrdPDLZVpkKXCzxlAwhMs
aO5d7REQkc367dfvRDlMS5+Wu6cUoZDPlhco4CEom8NcvwK9bQ6Kp/JLPCXYTR8H
iw8ZmZGzssQDevJ7C1Gh5oO8H76OLS2vrk2cgI7qIqLMyMnVDERz+OgmJds0Oi3i
cuOs/6FU90RRh6kqFQM1nHc2Qwvc8b+oWbmo8z47BLgfS4Xpz1EHXbfUfYLv+Zop
+N6HHUzyAkOXTMOXhVPTZ7W0w6aE8lGkf8t/FM+6YLk6Ml0cT1jCpKgdwB1yGvH1
ZFysGBJ1kKOpIm7jDQG55o6p5l9jYtX+lgqspx22WXfq2PZxEtLHXUJDD5KQR70C
I4jO9ljC3stRTzAce2dFy4wUejqno2cwuxc0B9mhgbJLB77JHbsGNkdG50ChWUhU
RGAwCWrwXiCPNk5+/1TZJmJvIoehhJi3lce3jfyHloFp8HtoBP1VK6BE6NQ6DLdo
9vKWggsszPUomMbCF1EilzFAJi/QiQALpUdlNzVEOxodN3eLlhmDpUy65lPbm357
L/GS2EqmLyiSus7DOw7R4iZ4ZNNS+jq8o3F59O/s9wUrbMGqNnpIzPW5mRVSp+Qe
ZelMDumV69riWHv1XbO1jmYGWCMJVu6+93p7gQbR17IKYXWUz1WayudC2i+25fvE
L1SrApIyOuHaSMfnaqHs7WafWDzdSi2O0f/tPSRAyueV7YBSAoIYQT/dHiqfF3QB
9w3DEeEgfgOb5e4aUPOAnBA+gWebgbhabnDWyrYWaAqdej6ov1+OnIKZmceqHe1X
UrsepffpBnUTWWDUMfJC3RnYJxDBNmKfiEXKZdawEbU6hlXnmXSfFKhgs2Kabe59
7zQWEwfXTpoV6amYJqFgKoZ06A8A0+32A2bsIyzcfHDhIoSv3583MgGk5/FgAPl4
gXYf1EV9M1JYcyJXHXIrwxowUXmi+N+TdGKMJPCcKoFvz4BrMrvtrfjji3XtQaHf
9EYphUF+uTjPk1DFW+1yHSkzcyrlGFor6XHOwiKWWj1jVbQKj0gn296vr7bBWDKL
ZI8ZF6Yy7aTggXfrR9k7pR8ROaDW3byUUIOXUcmOPOShkO7INZ+cqSi9J90oytDm
5M8vi0EFBL/oRXU3kiyzxEn8tN+P9scEhL9OzqOfY4zKGTKtcCmYx9Hl84Uww6b6
qXE8YY3TlE5rZKgVFtvgqda4Nx4R7lnlmq21vnAldNWwBXc5gR/Z9YnXjCXIZXos
XU2VIYSG3KaFnd+H22CWQ2wfot2Pv100UxAZAGL5yUmUzRG6TLLMZoBPcdVhysyi
y9iVVFpg19eKbHUgUGojcEncd6USra3OhGXBrMM3qFzHwdZin0Y+tPD7IAteBp9g
SiWj0fTabo216riv77nKsy7SZmUTJRNZ7EG1yVrQ3zUbsIOlJRXVjofV5vZjZ5kn
9VF5pF2iQyB4EQwNDwBIDUY9zohKEzWs+tpA4Cr5o0swac0HGr1CgcNUH7h4DAXX
RyeOCIALqnl5OUnOPmSdvvT0VbeqQsNbYVi3uypwIE3V1HpwekEnNfCyHWNCEEhn
y7JtDHbxtxLzv07vdkmHwItAEC44WWLYe9bF06QTWOk2/dMxdhc+Ss32rNFgzfU0
iy3BVtihXKfcgsLkISErh5FL1sPNpY9OHPnCbwzbwxTo4rI8Nxe3oqCOCCkN2CyX
NgXtgmv4NhOqDZij7sWa+FZVTSGa7mB7elw9UwL2vKmHePvgHFWfzYGreQ/LfVK8
AJCeQj8T/pzsNjb2GzCfeoZ2P8sXOcvfV0sddXlFR4pvaMQN25y+yg1oNm9YVcvK
eoBGu6JiNSHGeRMcSkC251fGQx3jgaX/WkpP3S7QPO27vQJocvba8cc68jF0zFFO
GVRrJrqwZqUvJelch+PKEo06UwaAdvUgoqcRVIjgzTuBnCzCPN+ovoseMLbR/XZ/
sZvuO08vqSMD9jkRu93mqCmW62cwaabX6Uc/Kkp+L0U0uxK1cq32LfeUlTl3rAsB
JaUC2cEPJnqAmWPlnvg9DLOCNd1OvgyBf5xICxB3KnE9kENp3La6QJZCT/CQHrIP
xBZ2Q73Ni51+A5TFEerARAe/XoV898pvkEvcY0TJH3WCRzc/wGmhC1rgv2jF64FD
B6tGM3a/RDOw3QX9ILJmJLTodGx0Ebkq6ifIv4sG/SyS8xE1pbAsYRXaElAJLE8H
RZdsjEA9Ql8n+HgLIJrQ6UHHbTeSploE7igdI09BwSbbVasjKmtPRv+P6sT5uXZW
+ZIPcSYcTYSdjy89J4pltA2YUs3/gTdbFnCGIZBJ9fZO38JnojuPF+kwgOQX8Dq7
LGfTpNiDv+pMteoxXaJdB+dkDfUa6YmdtdjZPl7z3IvXDLEM+8H7FN7jIVIj5tqW
3vvS+yFJq7EP5PYj1c8cGJiBeo3gtIdszGKbjU1f/J+Htfug4mMIWV/+/11cmCW5
HW4cwQ4uzHs0zKOOAc2el+cnusOh64K37YlH0den2Ws0T3JTWvsl4UI5XYPFLne1
fuk5o0zF1Ftsv4C79fbrZSrD90AAC1WGuhIHaN9evUiCj/nlQUv7PVIurQEdwIis
Ry+zchmB1Q6hhy1oJO3K3TNChYYrr6cP7hnkUtd0thxNKxwfJGEWM9gAHm4SSKRF
gqgmA2luu1cpfnyjxq86AXQMYuo7YdrmP14+Mto4VSPnMzfjq4pZhZKhgLFuQWiR
uKNf38bFpr9SDfLj0cag4cocQqV4Q9pzPVCj9gkntOFOhGGqo1rQHXBl8NZoeFFO
PCX3oc2qI4LKkXMM51wjDzN83b/niJZdzoVgp/aLiCo7xfCVqxzmkCPGSHADcxoR
bjNyzypA5d2+xgamkBXo+tyqvPart/wpVGOEP6mmWgQWv1frGTaxqMOHokmNPxrU
CLBjisuBpqln2DuPmlo5hsRsCRfh3L2esVrKVM1UmLapo+Ue8O6vAEZfZBjKR040
tAqrb17fjthZ1k+keRVeVzv4+uccEPrjT4EUPa7eyyHxiHFg/IoofhB8R+Rg0K7Y
ICxxDtYlLLFcGr3DSfPN4MKWBkutUdQRKuOy8c/GkXFpyRcG82Mf9PfUJtADI9GC
wQqOtk/vGtjZp/pFXV9pnrbc4yOvRZzbFo1GIZEAbI3e2cGD0xrSgirSuWsmg/yS
fRa3stVFM8LS2qPuZugeUaCiJKlJVbzlghC+rOZ5A+HZA03jYxMxY/Z2dJTV3jCt
wDmWlSFzRJLS0qZI/9PYQp3CEZPk0bQHtGqyznFn0lOVJ1p22vSNkfhs3K4rLkF2
ThiYACrc00ailRvccxQnN1GHk7U0GD+XsKl3nIM66EwBYFmkuDiqypj1wbwreMcH
rpkiFwG6lUw14qspZixgkw/JNQd1RRPpo525doNiGRMw7V7LX1UCNsJ6LylYG7oa
DhAp6LuZHrTjQchshKI+MHPtyhSlfRHS+132tTUEAXsSvZ5Zkarujj51r5dZvUW7
yIqQukCxdaKs3Gf5xKeV2S7UNXimCtsui1AUWi7kktnnYzEd91mHDFoWomkPCQze
riUlRVtggxg6z1yiSk8omxwjZ4meGNneu0ECh0ycYaNNyPYboI7TfOoESQvs2NId
3mIFR2MsyZ2H3TFCfnQxAkwJ2Lin3QVXiVGZPoF6QjPVWBYdsvVC2QKoSBa63/w7
2/CTEXSUBs8jlZJCfT2E7oO0sZu+R5iapwCQBfbGxTRPWALT73dBr9YxJ1iGbrLo
jPPdt+VDFvVhtwVmewY1KUyk7SKTVsSa2IMa17EtCSe03nBTjJkCVZOZKilhRddZ
V8pviMF6LTai/OL9ZZQVf3+BZUDH2iq8bP9so7mRwxEyWYwtdQo353P/W3h/K2WJ
BK1Oac5HpLQgJW7ao5ckuxMeI0/AmrMVmTboyMlRviGNwsk041GzihE2fajb9eQ+
iwz+S+ovAiQcBHg23/oSHAx+s3TvQ105v1JlpncYd6gbHCXQ5Sy9WtSJUsuEYdnA
KFc9aaLXdCVw/qxwCPlfWiXhI3TinVyGXTnzRYfgrTk7q+EOwJRjtfji5ycqydG0
6kX0XPpl8ohmdH73ZHMmjN4oa4/kii+e0LGTrQEas6TSo+QpGCjKMIBiTvoLozSO
FnwDg0Rh5ujL4Opr2/EqlGB4WehHxVLn4lsHgqHgKTDCQkKIx/WlFHRypTuk7n03
uP2jQuCqiDt2tVvEGQHJpz3Qtr8qvJKLa7+cAm8js3IBEKd+5BkY+LD6E0AKQqpg
Za7SACpZJaJVB3FtoGeYDj5EfHrEx6CqPFjLsUKDCgsdQAf9pOSv62Mj/SmXIBdm
Lmn6CQoll3J5PA+U+vzLyCfW2OL38zLdPmW5QXNiM5xhkj7ptwrxdv2LqPp6QY3a
e2iMUXRizfMkdp3lyCF7EoNhckP5ROgtw2ABLjrQICd4tNPaNGs+nAbNryGQh+rd
IaYjPgRLqHc7u2AVizlPAo6xSTKHvfzFhp8RRIJEZMfe3VH1F+3XWb6+O/16vT4L
65ndhFNtX63BBEENnn2v61pVh4ThwddxFOMZ77F7YD1tsOAbvZ2JLaTCDm5IA0BS
19Z4syaXEuiWiBQHCjeIx9SErM5qSiTy6bqKkMrshC9CKoTZKug/dS1UqgZYs1PK
v4N8X6v/Ky5hLolh78ATW0RpHuMXrho2hy40DSTLfdWAHy3ivRJDfyVxw6OiSfLH
ogYg3665Hruy5japQ+1l/J333dONXDchpjIEDtD8nKR8y5NHfY103vuHoXC+XP7t
HKiE/mWXNeKlP7Ptoi21PQYM5bdQrrBKO4yeF16GVOLoJoXDGV8Dk0vWpxi98u/t
0CnnpXC3RynqBYg+0etqYUOeTKJp3IzdFVltbNnlNtHfcCdQxxtgJf9rCZzF3yO8
6gW7X43+GXjFEtjQ/8pn30ClbSqi4tLB42JTRL1ggMSi3vDUHBv5Hxu74dP5L4QV
bQP44ujMuvSKRYVQVsucMDC4pJNqh12o8eWXy9Pct0g7dZft+c5OK4IBzFPTcZ/k
vJzynYnrfX34j9quJePeAY1bvUyXNOOq/zOY4Dlfx0/8Vm9ytB+AUNYTnerY/TMV
Kl2tfv/9p+LyMU8/3AKrxlVSyz1boL/EKN51LAgqg7q1adj/9I9Lk3qYcE3d4sxA
nzNfoF7TAtTj2ywpuUodso67IE5z+aGbi7uk0/Cb6Aabj38mJSVAUrnGOTM1WicT
XDNnO9LouWdh7y9ZaCLWxL7YPGuxdI1vb628euK4vp6GuldVrd6SPNp0mahUC+wm
QzAkEiQRhmgCicnfB7gPta+4wMoFMS09VFORnkSXUX/hsEtHECg5mS+oWWsWrbWq
3iXgSL4mXfNYqW96DN6L7DfYv1ws/q6S2AKGtHFeOgK48VOQ/pQHaqep4MB2aTZF
ipoX4Yen424Lp26os3Dc55mhDqRmF5S8vHSHaG90c/cK8bwvllKkroyqZF/eJQCo
eaWpbP1L5lS9bRsJPShxzZPDKji+Ab3HFfTevA2jqGu3vY4ktIcogeqVUjEyDcQA
RX7AsYC+y+dpHVlKSCh1XO2OT0Npzz4gMiagd85wRtl2Z7jJTd8H4Y0E4hqyUWCq
PDl3U7OYiCHhvlS9oTY7iVMY4lvK8dgXW3Dx9kQHX5s2sbTyOA2/du5wJwDg/U5M
/tH6RP7nOlvTYfd+ZWoVnhNG28wESiN7mYbtbt/GRwHXnvLHlkVu4lwDRC/p5xAQ
k/6yHXaX1XQvBcRC6CGsO1WBgKabmuuZELSHi7JibcwwQBJD/3R/aDSD6I/hdI8a
eN1AVoK+a+AxiPm1hHvtiU12iXhRWSLBVKaYmwyWwt21v8728O8PizD6iFQXrso5
ytrNfNF/fEUs90/C+zQkhobUVTFFq2hhBHcVvlbyzUap0XJ6X73JA0Pyy6z5wbLM
DXW5YGCQ9WarUgYRSKqFUgZJrvE8Ioeljn4nxSVC4cRlrHmcRs4qX9p0spLhuhsG
3ybBIyz3HrxmGNVyRfOMyEi3RdjyQ7tq/T1Qvg/+XKryMmqIh+jZdIXbC9fWubmt
9Zl0BaKtxzTwvwDAmzbi9wSft03AdtEzV2/WA9y+6HLGmyfwxpYSbft3PITWKrb7
H3UUWX6YBSbhvfUowxbD4BDLtGDrZowKImb8e0dH3lEy5RqdjggdVjfPLQUO+xBT
O+ZoVaHSa+wyJ+Nl9n5LUGcRgiwA3qWg2kdEOhBflU+tDnWQE0ecYSNM3Ie4NDIt
x2mwhLJmugv70eZlGKu1aPTfz1NVaGPAKGQQPO0GfL3WA32yCiTnuts9aoxgjTq2
tXm/ud2wdv1jifZGd4UgKQRTqW5JzwUCFswqay2e+GMqbvq71iC06sOXieW+F9qw
CMXkOqeYjMxoIEmBKS/Mbr22PXM+zbRQ6vvBxknc20oav3UDxdoVmrV0RV7zu+SM
WNDNVYCZ4Y/eAIIsDjORLyoceLHOhdOIZINYxH+L6UAV0Nyc9E0RNgwE8KPFgWRa
rmJitEjoEq8Xk+wcywksMtUmPsdSuXv2cCXpyWCBL5WmxeR+ZDqyMkv5j3tjeoAY
44eZA6Xx8H/Mva1uuBInxjVPobrvHTJ5N1ytBCq32Bth2IVjbxloJwtLlWO3W/GM
2CQ3KpGmL+8aQWClpHrj+D+EC026B1umBEfF077toFhBxscJHSAmyCZLo7hZZk/F
Bi6c52e+uLzLGb/ryTB7rLFLyymB7KYOyAjhikZGFREPiY6fCit6fFfwLvqU8Fuj
cQEGojvtjDk2EM1VcuauAMVcYbxJNd5UbluUnFqUdlIaZAGMUNHOdq9hkLuUhrEI
+1gjECr3RVKKT3c706mDj+qG/fontCLwxAPi0RNCU3D/08Og1ixry9P9DZ7XBNgK
ef0WVCm1qGLGdmsDT7PNrpTuA3lh9rYw9Sdlw9cWoDu9M1OQ7CaC8RXhdfJCifXt
fTavNAVV70z8n95+RAIb3QkZwtZgFihkObKsMVzWOaarWUGuwaDycxjaqnUriboy
bu4A3OzAU/C+5cjT9Feleh0gB6pGxfy0KC20LlXQT+P5xINZlqCTjpJvPoY/9Fxk
vmxcus0tD0qZJZL9Ltth+GqgKNdralQALFSUyfpCjVbPriynvrW8EPVIBYvrzRbj
jDI/BkMlIt2aKPEltUkwm5HKiVNrSQlY26xYJ9pPZtaC4h3YvQHnBrH561sQGKQO
Vvidkk6snXxYnB6+xPGkGbEXtykiC6ITaElqogpqs68AAWo/JLmkOo2YqSJ7XOcV
WRJUFAyEFP9tpUVbiaFeSuIyFhjcesydAUTvDz1asclp6Ivfztk5ze3SzyB7QFw3
bKqoCTdHll5WQvnJtkwjvtYOmPuchm+B1Lblbc/f4r4bVTxTXnTMDnt5LFTFZFiq
naq/8rZH7JnzJdUWOFCOVMgZXtzWFPbyIt9wQBju9eGIt470wtgXFSlyAtYWp0O+
1QdXCa/vwarE59MtBGcKMtsf2W4B3UyK+MbulWlg0PuRWJMLL3LntLRvQIJBojo2
zamR6dgfayA1cdcL8biAIKR0FY59ZKiPJ9BjaRxajDO2EjNPRNAIhamW6qp9TZUz
Aq1h86sWGjquJBh0BM1LDBpPFFnbaJ6ejtWzDVWoHDNtKVPQ53npONg0k6jdcKwJ
zCsPS5ss4grEemQr/dKgt0MM7vDZgN7UHkNa2Fde4NZaImdFoSL/QJatPVeqVROg
7ye9EjHQbrex+8juOG+3WcED93/l7Pgd+mJUGruHW/fPrgQo2k7EPQzCn2deaYtO
zeSklJW4Qzx/lwVfzoWHaju+4hqzd/zJEv9egexbABXr6iUS0LYwLmUOsUa0XOwo
ffzWGvmB+whu06ifPZxEhl31YZ+Ywhxb+wLNc+zd2mHii3d5iuhZsNwaiozIUzRs
lryLpZ2MN84dLgizZWN5juoskY7YPFtlryO6lpH78kggl43QDcZIVo/AUHBLBbmg
Rj+FrTg92ASGsfk6TZ3VEAf782s63j/uq8hQhZgwqutYfILyroIkXN+lABANxZAJ
s/OKK9I2T/iZCScpjv+bfqMCTbZWU7iAACVukHgsoYRjMT/odCXXZtvV/qZcfPIS
+7HdS12Y1sqDIAcDKbS6zHmtmY+PjFSAKOreLbsqscvVp8X4zhCNvsEo0mt/jNfU
5IJe6WM+cXYNrXeseCCbZ29ovhAHa9wp5+gvAs/GXGg2RKaU4d6p+7SV7zYYo+t3
It32H0xACIEURykYL0k0kTXYC1Xg1sPtVrOMAvemVHTyxwDlEztrQoPBeVDF1dA4
gYtL3zvf9rvlB6P0paMxhVb5dEZqf+eFupmII3v8rbJ7x9yXPGjASqoo06pvi3bq
wVdSrZr1GskTghizoqn6asjCb+3vPjstugZOdQ510wpljh0SEsmR6PBplkNvMozh
CeG+cl2dS6U/3rW6682oIMC9IRQGvz7LQchldyBHod+WyrCp9YaNHYt7hpAdT7ql
t0dQDSGN61/UiM6sfn0kvW6yozItPFonugFwBgHl1F3pvzjCR7gr1loKOjJ/fomE
oI7sRrGWACWHalSK06wd1V9ErgYwAe4K/aNCsTcuNjOnWdnNcnhDryYqp7uFhlq0
70hkIL9Agwzyfkuha6Kn7x6CAppto9lG3K0JhzLZsynBlfCdvM4QtZ+yZHIGfLpf
ityJjmThz6ibaMPrKJmg8T5YfU18RViwfS9wZZ87ej/LNUyRDDSRXmUk28KlxTn4
Sic7tqr1TooWfk2bbx8pvRlQGRYT+jdc/a4gV5LtAJ3a4PAuXbZQ1MxM2ro3U0Pl
JivL4QHYj5z9+DWbYvZFY/O8TBWK+LO5Pf2vQYAeySTSKxNqsov+Jsjnjn+/93Pz
1Enmdtp+MIB4+ccfDtcG7IaCZJwYLwIl0cqk7oPcbrE80mQp0mmTjg9z+wBGqQQj
gj0HRrqGh0T0/3vz0e2iu3RhjgnA41hvqCcIKqRZVh+S6QI2id49AOa2QnCPTmOp
v7upHBLDcARKS6eIut7TSDV9WWVstIBQW2wwxKZJfvWcTuJjmh/hA9bqSs4/f+JZ
oblGb8A+OqqKvrextxK1NDSO0r852NStWJZ5OAv7s/I9mx0H2uFAwDRVvTL85vYX
85+KRC1SRkpfLfY6FQihWoRygmar+Btt7kG1DfWGYy+igx2O9z+0cZQckF2GayNX
PGZ4x8jJsMOFFFytfc5y4bFCZzRxELtiYrVV9RaNjWR1PZO6lUqEKEb0ivXuaphf
LSVwFeAt9zk52zDnUlKaTYizE1G/jyi4lbhIrmueAt03m4rCTI0A1fepjxSToR6+
MIN5qh5H6IXxSYrIwSgLkM8cqGvKmWr00b+tnQrf9ENCwllVF9RHFBFvXqimRPJA
vwkmIwbrZeiAUAl/ChrlTOn9RiB58sIVNgGXAvLbuM7UADWf9+gonLaQjjZUnTzo
+m9FP2BjTVaYCXN0LJ6BXg9uUpnjojnn1AfzZEiLgqUjJgtv/HKCpdpV6n0zkVZE
sDS6DDVht5+GowB/LgS5Vgo2rahSFlBKSapcDluPGQDwdIlmyxJYGwmrJU7y7zSy
obJEmaglDP++j5Sy1P8ULzBGiUHb0yinmO4hpRPhhTPznyP1FERWu9+wmwzVxXKW
GVxkFp9BP2lvH0+kVUCaobU4Br3LSaLjJqfIaBPPuSY+ZN0lPFyj6Vac/kGviYyB
nnKQ9H5G1ZFDBWlhoJy0e3NNUwoZZ02ME55jA60m5GNKBxK4CaayExYG7WCflUo2
QZIAEdX8nnFMaIRZmBfO3TzeRUn+Vh7qzpH4//inlQXMGNUGQZ43XJanXcTkN7ut
PlN9JbF23LjfIqJBQowo3BZo1z7aIxZPqas5AtsS1H+dP1N1JzERdIgVO0kjc3P0
h3ksIA5+Sz5qyUEzYljWf3jHDWiwOBD+Rel4RfqZprMYpwj6zzSQcFIrcJ5WdhMa
dj310wjChn2e2AULFs3i6suinzHmAq8nbUX0gY9WCgS0oSTcA2ltyeW1Uu5Nrne1
MTzc921kalzGhFTaeBKXmy6j9e9NWx10BZjuX0T8Cy5u7pF5NVzQEpYoFRMr4C8m
6VEK4BhlbQwaplfNQv0OddtT4zTLkN27kpTLoHbLxWkkgUePP7BPnHasBIQKbeJ3
EAbiRi+1d8nwtbeKSG6C8XAN5hyBbhOvgyaPabd5d8MB0gU1ZYvQdnKFaFTq0h5t
CwG6CimcDVqlMTmO74HeSCdLZcyFXra0PQDnxRc/akE9B75JtMduhNILxCiuVknU
+3bsnwYQd8JTDEMYrbo/XUSduHEraJAwZtTOhkNktFY2hXD1AlmtauYLq4fw2OmL
Ki0MXYx1LBRlsraoovrVuCW7GU0Fa2wzEiMz41WzVHxe44l6d35sdEEGoAuRwrdv
Cbnr4NX8vcRundEZUJxezkkcyNMbj9/azL1VlEmVFFMTgEFiyirxJkJLV8zFv1hZ
X2av8ViyH/0Gro0rI1ANkUtpU+IJPJOt84W0t2scigvJh4nziCnbmbkXrBvwCBF8
WW48kg0CEVXPSAndq3zVjxsO9H90f3WlUP2C5BYjdUDQiLK2CJArQn3wbl4zqO66
bsqIWO1jwn6NtQISG6fs5bbwkUg5pAmd4PvYgsh/5SYNkNFjWsubePq/PpSP/euD
wFDiA1N4Y86fzhCOGSYE5eyUbvEWHCwNCU4leioTuUiq6L0yINAs3zh6YNBAKM0f
Ba6ZlFZaF9PLw5MhcDP7lbIt5cUt5V0TvNGcW962WbSBCDba6BGjj/SIuIsxM8/E
8+nxcqWGaZpLpGwfQ5c/pPLqhElsWcenyQ1KYnYQ9BpOpozvCk5AkaGnkl5oXDAT
TksG072NnJGXzKt8GO/TI02hHtz+f2yseOiAqs9+tGuUf8KXoP3pe9zqF9mRtKOb
gj0RWp+Cz3lAN0CwmYIF+nFPRNI2s/Dbbu8853jl1L3YmX0AUsH26J7V6/+kZ3mM
qnwOJuocRMygguK79v6LOrzKJAHc/xHpwSipiRAyG69l4P5zRQuB9aaOTytveOUb
btsdUEFYXFL4O1zbKGN4ARwMxjHqH1DebkG6pRKVOA4r1TzJpM9hu698S1j4jk+0
ccVcombiIqXw04KYr2BM8YjM6CU+yGSX40ov98unImFtA/G/FekXe3UMmdlQMSf3
ERFn0OkjIsDSxphj3Fmuw5Iv72AsEY8cgKoFx6Z6ln8DazB8j310C7Hmr5Mabt/z
Kf1h+CLMh0vcbAKmQaT25/96XzFz7Eb5WpTXwRkZvfs0XCOIG447ESOoN3mkrDcs
CuZSUaZSohTisFMLXUfcWSXGv6U/MXKqKuYyNsKdXlVL9BHqA44DaTWo1mVJds3j
I3gCUa9uXK6zcssJoS8j3v0JKdFeLR5ZXNkm4cHmRaNnBgEAZReRgWhr3ahLbfkV
4ziB8+uJ8ZGdOi7aIplNnazxW98FAz4weOx4hfAPy89/QRC/mzbMH519HuXnDgBx
hkzZg09XetnjVGz4bvcBPAYQTUrVfhwNix1D6sAxWbTvW9He8Wsgugn2ZNwI2Ekw
6CpVqrU6vC93+4+fQd/7/jV8eLuZ1cZ21HR/4v0uabDnrlEeJaFTAgyxHJySFh54
E+daT8gGkciVh6waFADUkjopMsxfYd8lbP9G6pDfd0gZJ+Zn1ta85L3v//ASlVoE
0eYhz3AvbmrlzAnPIFa4nSw9jqsxkUNeSFjRacTugwg2yM1oDVNAAvkZzbtQHj5T
q9ySERfbNAyfsUuyN3lIVPuKoi5rJ2FvixCwxycycZGm3rHYlvMYA4tF8lZyfT8w
fXGNuUcfoiAHibPHyCiwNWCQl2SXhKA/MqdsLDAYI3byVcSA006H3YyOb5yNx3P2
SzMgtIoGOCKFojmWfjB7aewxCcHDlR7TLaZllG0pibR0Z4PREwR/tQ7ZNTBfgkEd
Skj/sh1lrU3S5AvzN1YS8Bva7Tks68lsVpm2D/y3QQVIuIDqBSNBmSV3j68WWWvE
WrlQAc37BKzif0Wsl9j9uAoC8eVm5J3mZOkPfjg8RkW0s2EvdpNX+gn+IfVKCEUF
ndsct+ju0/4KdZAuxfVfWyiI3MDkbY18mTTnKX1DFGnpQcTjUUB98VolBCN4rPam
lpvxJgZWrJwldme8w+yHr+jw/Ms8c9u4jLtsZx/vEj9GeH+8d6gtYv6QyXtk0+L8
J84cHfRfxz9QhEklTpIFFdwZJ8hzZUxQUxhQVqc6ePE2Hhsy2ekozX+aMHsR1K/p
RMFVYS1pyGMZLrHfHm0fUgicH4MaiL5agi2+Yw+15PAbMYUuLkCf6riFa+cvXexE
GYKxKq+Jfr9Umk7ONHiHSQMob8lYMKt6Nm14q/2uxtjiRjRaCBBjXw3ZwpoHFlDM
hA4es+VfKLY2PyewXCqSLw7Meth7KGwyjFRxm/6+qA+zNCx1g6B/D/PiiBHfWiTX
tyCMEuwmCWrxm9tPadaQtv7rncyj9MqBpFOgJuYSg8V+SbUH9Gy8ZTIwhaXBdkJ3
Id/jJ6QW9tqP7gAJLYwCORanC7cWL1Jh20iffTKU9k1YH+gNibhnIsXiMPC1OQj8
OJqTzvATxciAmUADb+BUcjH3IRrQyBp5AXFRUxDqRxONGNWgazmFXjSkZoAzugJg
6/Q6TKuPEEuQbP5JdByFq70Y27zMW812gKOxhEUR7nta1iNW0LxW7K7Q+/Idtltn
PR1JQIYj0u+xv6QG69IZ/Gr+yn0rIgE4BYUsCqcPW1EsFjRmHfRdEJZ5hpIvAQqN
FpEpQWwA89aejEnXijZ+gK1fC1Ua0pB8mfEli5Wq+plGEuvSt+r2A1gClrsWgozl
AFobPaBagUkr9z3HVETeBQPAM7Sq3yFbfrVFjQfIS7C6BE+JW5gEGJIefpt7uXvq
zogHGR1IjhPlWfgf3VfrlrdX+7dxV2pCkYbkYMVOxfML/H1TVXSSb+9hlOLIVtXT
uCmRnLz2KCL9yr/G0fBP6vvRzZogqTMmmdlMr0jar2vVF+Q5QClru85UpT20Ey7G
h2iFHtcyvPeT3toU3u4uAG8wf4YqKWNic0RlmRc+1NR/O1UKunpoFy4sbPfWWdrp
oXjWDcICVK3Lz7xu8Z48biu5mckkoHhyx59k7hnsPDpOL+eyGazI0aaSG72ThEAa
JNAMspK+ehtT0ElQYtYRXJD2zlBqs18elDoWZyEt5QZ+KEduPqdyzg19FPQRYMiS
dlY0zsSz6T8fdQWAL05AQ/blYR7GYWcmccsqxms93f9mvPisSm7cyBwU691dVs2r
a252UF7Kn9kJWNwHxbfqLsxf79OegnX8v3A4hj7Y+ThRE27P0Vdc1gUn5oSHL0lQ
yhATmWUo28chaLBiS3KRWxp1ANYkkbAAQtfMAHq4PSxQsvvb24q+JNWvkib0fjuu
YCCM0A9P191gVQPcdULuP9pJWVSkTLXIpSl1zCNgM/3GnqqY3ergchj1lNXNdSVp
8slQUOylfnXOkLCgTHir+qpzD9RmoWl1di1td8X/3TQyezY3sBeOoWLxGhHJxnw6
GsipfaMfLqipfiDKui3DPygwwJl+262IsWlPJ1QMZOq4EDaIul0rLCRzbMtF9DuV
igVW78Xkg6pjL5a15NYJx2kf1L2sn4FrC4HHqE5QjoSGUB+VYwcfSpo7X1Z85r6y
FSFacgAuGnfc/5NngCOx08jRtP9lo1kkYVooczQUDyjZqgKpnQrHfHs11WOynr8K
aDvqhJdWTCxmTEved6OA+M/A2SkgIjh5yYgoi2PZ35Lb+gszlc6duz5ERiGVz4Ds
qhA2tanBYttJ8FZEiv+uSmFxFzNQ42vDSUZ4+/o4Idh8JfZmz4s36IoDOM2EI97h
2S8iu9HuNFgRFU0B0AtwFRkBs+acn/Sry1+Xzl79LGtzX+e/Hw/ztCAqVsYKmsUE
kZyq1FAMEOa7xMZo276pZwlThcZDtZDXDxvhZpUwH2urCGm31AyIa9JVKa2xGVJn
scuNQekVJvBfYJfx8+7YdUSD7ua5UO9Qk4Hp+6qedaXfRBJpcEKWJgiqYgIglM2u
meY/8OOrebu5KwoTZanxrGk5It0+XjT0aYsScPEaVsOPLZeCx4xKfLUa3mBQ3nbP
0EawbPu5FU0ZP+l0YpK3B7fE5PZm28hBa/W32dHb/EXuySb4yjjsBudM2BZ+40X8
aNta2YtL6y2stDIf+mOMBlTVMqfgvUtc1P/FNFhwZuttQD9gN+881Mq8ddnRuGtK
/KNQuPkS8b4gxMGa5kdbzM/tpVGgiO8Wso6Aqa7+ZZ9JzA3Ydr4ty8qP3di4fdM/
XMUmExA745UqWzHGmwTaqdVzRIo34NV0kVMzgSxoPyoHoRw51AL8WVL4Td1nGILs
pkUHXZ3OJd4fZAsK9EzgqDQFGiWKvs+ilJ6tPWwNA5gs9VQAIhKNSBAhPEKnRWhS
8NEjXHWTHMm8HE6Bb5WppeS2kCL4FNZ3NsjnYTmKGMmjLcpTJsd4ak/WWxUSjXRl
OZ8no/mkfWUBRBVZHqpDoA6xZwiJSpRgoOkEocd79/qDS+nbc2i048neYi9cI1hd
WRcWDXMd8EhqbsJ0YbTp857tBt09PMrkBpN0xwG/tBuVkDBb04/jQuu/z48dyuiB
2gJRx9lh0XdLoKLk2tfXqL6WE4UvQBLP2S55bXVfLi8NXq+KoJ80TDaWr1zrUzmw
C1ft2JY4PYh9dVbJgGD2vUZbzU2FeNe1rjNnhivfZnINNr1oGDRArwsh4k3oCXmo
VZ4Fh6fa39d9QqiMp50mA+kxOMiZueLLyVJpsX/KRUg5ES+zafuBhQ8gaPsQr6nL
yTEWbxqt++MvwIgQD+H0MqMwdCpM2WfPq1/tXcOv/vSRriUfTRdQh28ab+efk0HK
4q+laP3iQue/xrmTeclUi37EVj4FCh7i0TqDF/Zd4i+YWXQrSsplpLF1RiXt2Ra8
PBHRhPXmO5D3JkfAjat/zWhDBaX2lOpDNqidcElYjr6BX3WRObJJ2KRoPRibT2DC
1Fsj1IMqWJkiE5OLjbinEZML2HtNdSJWod61BULGxFkOjGcwQ9Fq9hvmDOy7DAvO
X0U2DILoG/KPBnavFsVCYljIYHjzretBT08S4KbFgBdJaBb7lZ/EFucBEz1BbH+9
IDp5FE8pO7l52jllecHTwONWtd2D+ENuoKxSIWE9+AVsWcfbKJfLacesaPVt130b
NJiKpXwTIFG+ll+BNdA4dttrPUXd61V+THO2ubrl7Aby8Nu12x5oBx0pciIkky2N
q6DcMbq61o6vexpV83ZEw+Z+zqFa0RvgCVFDC5IvvCgKAVqtfUTNXLpWM2oDu7aS
QBg0kvc+SHUWZU9tJDe9lYamCSw9YHnw334Wu+pdM3iKUxoOF0Ni5O1pVKgRuugC
Jdh3WnFKtpVzMBn81W4fnXgop6KRrM5knbWnlIrSGgGF3P0ZJ8bKbzpi6xAYC3qm
WAJiKJkRJ0dlwK+SZqTSylrmblHwQbwpUq+u3koFP/TcBJMCeBZBVxgF3d3SQoRq
aE94WHB/cc64q8aVanoUv1UELji1xi6nMDoMc9A8WySac2C/hnS7nAm6ug4aYBvx
0CTvJIUW9hce5gO4pdZrlXXeZSm7+jODY64U/YJqd0tGwZAYTbFh8K561r+eK9IP
+eZ+Vd0boJSl0RQXoxvn4r1uUCtm1lbdRG2Cdm5kZk+8VAwuDKRjQ+n4RxZJ8hlh
Bh8/k0uSPtEvtfZJc9SWvfY8fuQHFuWAgHaqTIfihGbEBy6A25GsB579lgHGJzBC
ZejFiF82jS0giPtj6uDneNanm3WHhflXPAyx6SArhReZ3VISW91vmFDcaP3pqf8W
bAFSVBhPrO/AMFFlKIWZjtjHqMy8uKvAYDtu0p2ZHJgkTT1zFWQoZbERi+1YqOun
eedt6NkElESO7Iic3VJAmbVDh/6Zc0oPuTQqorvpA1WKBQAYSbMiZEGnHw//GMdM
ndEOcKH6bqyYFWpXLS95o+5ZpWeKbyCGMI/NzbDYiIzrANW6f5JXN4mz20QC4pKf
/kzS5SjSE/u/RMiSSBsiX6Tx5qGJLjHwVa1HbbrXiT7NBU0W0ZDMOmfxzgLmCHs+
+RsgZ6j6ZU6qdMGOVcnAknbQMXhfbdksuipXnrQ5NgCQvrYblXEOym/OljQpzMqv
xUUH7UfI+UDDQCts8CzfYYVSprtYXWpJjNmzUSQivcrusocQsMGIR1REgx5Dha/x
B+qw2id366c6zoek6iTFDoA02P/mYPW4zkyOr+nCIDkDLIXK13Sh0U+Ap1Hiz6Jg
MyLL0tRoRdbACpqTB1tsLKI1FszosTvRK1HDtEoM48JcFvsgR3fuDaW+JBiUbguf
CKMKYW+VFntxLKg5dEk/Y8HFBLppXEVqBkUugD01m/q6eumBSJielrUN1fnm+3zs
ImotI7Iegj5jsnZLFIBh4c340Y6Ntxu5z40AHU+a1GJUnxLOLGfIFyuh4G8JbzI2
qkO9tacbc/g3jg9p9tkOyzAfpsR49Lrb3tR6/k7t1emrRBMA9oxwozmmuh9jZgmb
N9rybc/hyXP4I++ClHz2oEi++J3UzIS1U5boVfdXARsIey43rAtiToqZAf4KCQ6V
yi+VnBL3VGKqrsH2sjz1t1FpzbUa+XsqEfyRj6r/uT7Ow5oLkImD3RSo/BrWzqaQ
gLCYFN7V67Gsj1178HM8dvgOJxxfNRbgQXgRzcv8a6cQ9kS4a0EoLMsqW1TgW+42
crKZjLLnA70sZdLmqlw7AHARLrIGPKojHpwnET6Jh6bFAwiL3yXy7h0j18J70xCZ
SbSH/UEUP0NHrjqpkSKhx0/SbhB4TRlHNgZ4ojjVR3HEj11y5Hcx6Gs8clWuMT4a
t/Sm/OxcR4uW18Rs24TgWbx6EK2t81UMLGQJfhGZcbT7gyzWMeZZDlHF+2P/exrU
X48NO5R6OHJLM7LfdbjG8LDO6DkYw6nknMM3r4KDtWQmkxjeOeC5l28VbWCTD2P4
x5HuhLg1Gc40ef3Eo/SELPuYvWmGTkdFWQ2WRbsdr8Au7wQqwp+YxYgdP/w4dvsK
fgf3TsDIUj+k5OrmLWt5z9qiLFB/IUcDwOLIH6ODuZ+mWO+LxfSs3eEMzqbP02PL
eJstGHe0OjUNZP3tN0lxkHoPhSnM/ncG07iyRc1ki/AHCwTa/MovnTcdj7Fab/2t
17oibXkKbqKWTTE0k+R3/SMc4t3XiX2b6faUOKMi/bu2/O4A9sV7fht7mMl3To2K
1/a3egEpKRr6Gm/6CASzw9lSanSf9uhSOTjRM7gElBD25ZEUy6ZbIsaZXRgdCD91
+wORIjYiSTeOOEGQNSXgbR7fcH+j4o1CM2u13OPcYVTp4ttZ4NAkI8lecms9PeT6
u81KSRtKMzrrV1OXqK7LOYSTrmANqcMRcPunNIBDkigQkAyRclwgxls6FODqOIVj
KgDEEkDqKCudplXltDY93xECnzV05SXE0hMB1O3FAnjeP+RIouPZbR6/ZAWsvWkk
U71GK6i6n6V/lT+tfFDXCiwLafbQ5hqJDdLzMq0677Knr8ddXZ2aujPHu3Ug9cOW
mO00z1C6AqB4NI3cU4OorOF0SdP8HaUYLenZJ/cv8RUcz+RKEuUjGTf7Oxi1w2Ea
vHgK5lGXABzNWtM+jU92Psr84m1iOX/y1ShJWq9T3un3vHO2IcOtmgb5aM1Bgi53
FH77Wd6RUDMAEdF4MaUDl03e/L4ZXbGrv931jXbxewc64Cpls8bfgKiUy7kaON6o
uZ1Ffl7eX0iNpVMwzSsXx0RR7+r8HHjJz19ZFrnwJ7QqawCgxcAxZXcowlVPZjkl
IEfCM9wP840vLxj7AtwP6BxRDELOwSjb8PEAD7mnovb5SaMxrExqnSkUXvIcymYl
uaQKv27sj6/ZzXiyyCYiboLVM0VLHvzMtwnKtQDm8EkEcg2P8PMVCBlbFvIZ4Ho0
JRn6MKkQsLk88qpvce+/ezBc6oGVZocB+a6PC+bWLAzmKVs9dBep/grdfTD6wwqu
EcwQHX4SasPeyEwy4Pp9PzDq5TSyH+p54aeqbIj6+BIvewT3xy5r7DZGvSo/Wp4i
/Wjkawfm64GyUD4IeJNSENzNFrGbxU9o6gongZ7Oxq4CIOW0ekuDJ5FCeCqvOoho
O7AKDy89ojQtf3HBH9dORZGCC9SpTtQqMDt7e0duzu9V+umCt/yEOfAPDlpXnviS
sAKcYgKmKcRjYWrlds4Ulrqs/URqPjI4ALWp8KlZMU5yR4eUpe0dQrl/6qwi1G7L
oKWuX2mR/JOwergvCSViaC2fRsJi1xHzgXkEByL4H1b7V9EJ1vjEMm4wBQ8XYCq7
E0//OigiNZ127zXGHI5JNTSz82/kQRK/w/rbUpm4SrPZqQxhcjasSn2zJL6WjteL
1zSW8Ca/KXA5bHKhkKiyKGABHQxTa8boYF2JPL+n01qcKEAX2YWFmaaoxgNQc3oN
i2ymkroJCWSQff7GsGmH/fz2ISnTG46UCqjMXESw059SsyEoVTJ21oixctvlUqVz
6Hw9oIAyfqUs3cUYSJVI9cHkwj47OWxyWrQbzcUwGgHHG29r02DGB/JRvvdBO8O+
M64AzdV7QAWOK3oTtYFkPY8vGTfbwEgZaD3RTVknzvLd5xfXAj2qLMkaEt+8VHrT
KwOq6xyvk7b45fcrGiPZtmfY+tUdRQTeDPYxVM3c0xCYb18zOAatrp2etCj9lumK
C65XsO8Ptq5JUWvJTSTOT8sHTGqBBprMuqm1+ovgO59vW2KoUHDQHCQUeWSQ6Ayo
WwdOT8tF9a0EOUd0mXtI9sQMBfCOTGp4OpZQMH0Bfv2eKxtaOVi6I/JyYxT71rLe
wLbc7AFnQkSypjgBdEE7XYBvsSxxfg5Y1wws+g+/ItupCIrJrOcCvNz8A7zo5x2z
/01e22Gl2EpvWDJoGAERylg3OPLev15hCyE9xi2x31ZKdMjoxcqby8HtvpCbKR8D
oUEInOnbbBUtUY5e4Jg8h5YDVjB4rs5lSfhsGrH+IRiXyXMreY83IThMS8ritCkd
T5U37dQvKL631i/qnxpuXjTCTr4MCTTcrwlA5PgQpxcEdCry1cXHoq27jry65JQl
Rp67GUzJzkzAjxvrW2c4wPf05jljSLqaHrfhHfFaoDEyzCXD1hTEUKsk2DObwqI5
XKVmc5zUYBq2QRnb+1XeY0foee0Np1zOHiixAaxY8My3rksy43okOlu7twzCP7Tv
zRT/5ajJGg2q2b9Nqrb0tdEyqxeJPhHxN7AHerrz9SzkbAODlMNr+oIcbZACYfnZ
3yJjg4gMOjNV1Co01tQ+3Ihoy34qNJLkQN9zIWFNLuMdp0Cb/YS336SSCDk8EcXP
oHLT3FW6Y0JxFE1EZBA63gagmwSRRD+MXKQ0aCTjIcWhjdzxfG29LecObNxzy2wg
DVLab/yCx+KjZGxxH3PcqaLylOWCrj+587C25+pmEe+Axt4LETWU2NzQu9Cg8B0i
9EgTHJvmghYKNmkQqiKo1vpdJHhcA1TN5BCOBEu1N/51cfyrtAdAwofEsZG9eLwD
vN0YARpQ4jz/u6pvIZrjiU7sFpHOOCMjyxmWHlJHqTtMWwC0gw9a4Bb0yRAtwgN0
J58wEvMvyh5B1MMd7O4CLqIk5jYIbDcOIaOPxas+c3mjO5dk+yb7T+Mo3ViAvcwH
5CIskfDZ/Ao0gxawHZbrxcWSBL4Tfs5aZaSrbPEHljcDbl6ULTHR+GEwbzmacDdh
/8yRa0bJVSFnldj7puDzv6JEb4GPD3yQRc0J425X5XRbaJMVIeo1Pjb2aE+QFnlx
asrIYaGPuWxGnZlCMW7fS3lr+2DhML2QnpYboCydpjtNoZvYgXz2ofaPIQ8fchdZ
b5Qp2/k8XECZvaFvM5c1IBwWLIBjDv38LCyLLr0dNB7uVMSxXFXCNfQgerAzl6mF
YXw2bZj7YdUsuLwLXQs5efhPdW9vC9XJ9OjtpPQ7Vb7l/HyhAw8O3p//pmMCMScW
FA+An02oBRWVcLWtXnlS11yiXv1cGMsK2Z1gN9iBDZIv9pUOOeaHdSxiYMhh5uzo
VJjuGiGrcbd9vrA7rEB0O+x78MUFaNlh6ZjjQywlCNmlJglfcUN60sjIsb+zvz0I
f2y45VcF83Ari4UfvlpewcokEBTPDl/Q+Cqa3YUobTHG+eT5lBy603y/BLAqhWfc
FSNx/SBoiyezcg8bpJYko12C3d+hmVAXqG32kOSFE/KJIYGHlswrC3aO4TR3y2oz
Cqx0HtiyFWWg4GAEhSfn94r3bQVLmuwok1b7647oT1YYfZAeX8SKDt4JLrO+Kyjq
tRmt4go46Qs+sIp/JB1ujaMJA6Zn+eyDdFRrNovUubn2lZS0iV1Wd8TaOLtHjCLs
smLM+WDmZvsygsCe2xRWYGJJ36yL3rsCMV0P88LVyh1mbyg1qJKZ1hgFF+Kdf0zQ
Cj/hKDA6uDX793Rz4KbBvxQyQHA5EaxxaUme98mD9mJpq6FNIYdrJE6m3mGrgdSy
KYa4E6TMUBnuRZ+MUDcMFUWfRoyw+zAdTgKQfbNvWTH4LF1lkzcqxGOZLVm7w/ms
mLhOHrAQY8uQ8KM19SDnkOGWzE7wOALsnt6LSPAx9kbrNwIYFWQ4F/TobIgMxr0l
Z5a+Da5T1LLr63SuuGD3oT1+/nP3ZRG/LR/QGuy5TnyglHEjLi+vI9EghzqNMI4m
Jub6bqez+LbPkLkgcI+1m498QDlnfcctTHCNT/b/kZwz4XkdEvaLnV7Xj1fi7weD
hqiW7PMWyTg5ghqXvn37AG3+fHU2j743W4YLfLbH146LaWEcaLYSpt8GiLnmxskQ
xX2eN7HnpiMWg0NWCBImNH+ImsZMyf9FQw+T1CModgehFPHloApaZHCQ2orM/nQC
k6zpVmczSm5ScuQYbtIDZlaE5lOKrAkbjmAI9Y0EqgjKn6Kp00mXqQqrn8+WrPC1
vMg0xaeywsv62/lfBU3uAP8q3GWgWyqj6NmASJa/uvwFFn+OxoW/VC+Du735Pft3
omoPYyk3AagVWGR2ZV6iSrauPHUHs5z/bXW5aMdjCHnNTg0K1buqBJFVUwhs0EwX
9UhSMPyN4bAyLdxxNfDkj/A8wlNcfvIezCuXGfpyPnUKeWOX6+pprq7QdLeCit76
c4vOi1qTIAmafM3j9r9dRvmFZpL+KDnVtjmDrRfGL0UVef7o3wLdLqJ3VuF7KaK8
o1TeGV+ZcqHH+tmTt/EQQX8deTXDWJF9Cno0dhqYhb8BfaZnn2+R4MmHkYLvr1YL
YUeLQBpVAbSsIdzRso8nDc2ejzC18lFHh+Kg6cAJlURjVvE8RWqjhmerQRlsJIlU
OuHKeIqAFFt3P5ZonQ9ErirzRDaKU4c8Cg5zgou8ny5RfGWwjW7BNXRuc/BTAdxU
RVAQ5JlB5iHJJpUb8LRFlDx8/5YJkVi8PtKWQGpcpEhbXvoRbzTt4F1SrGWHrlzc
L+02XMdzzO1hm6gQYZx4agwALnfTgstJWedHkpie8GdG9F49qfa6hBiP4TeJqApF
vrrlwJ2f3/vNofnmqLCi5rxFHX4ug0PiVsJ512rsVkWQwUlX/SKuIW515eupZvcO
tLMeqGOSd8RO+edAmAOVIYdPr58aFaf0q2yY1dOJCXUrKupXU1nBsNzrokTMMvus
XquUp+J0LVj1qnloxZ9yavSW28my1fwdNoQfyJYjN0WRsqL85ERfMkdL2AHnaop0
TZxrXm2lXXbwLQDI+97RjGrxu/aYY+JWukDOjksyGEYxhhdnXrEwcqomlnzvepPp
qpJfHfywj4VRyuLWFtEWVxMGNymlu0847LL25AUyKNb2nmkXkP3FHY/MliT9/56r
X4DrmlDpWSfJwnt8HtT6mtt3EPSSSD0CD7EdCNiSpc6Ld7ZplHtUZTwjMzhpthNt
Qj66Z5WQNWJxjWEfi2ZJjlM9WFX+FBukw3EbCX4sIQ8BVQrWGk1CY/a6x0KlGLxR
QxePZCo4qqQNdihfEPqzxWdrk/FJ2ndY0OfeCwo3J3Kj8WlkN6yQL4EdTS82UG4G
hAFX/Tu7oi9epyN2y1jQdTX57D7zf96nvczbMfRS38nZp42jUY7BoIH3r04UMfCz
C3pNsM9heH4lu7j5FwjSE+MxB48noaLnunZlX195JZxf3NU6XCSblrth0gs9cdI6
4Ec8RwQNB80fXDk2GXidTncKkmQD0+a+T4Oyetal7mK2JTVbO2GTmm1CvIt+phce
ZGxVmyy4Q4rWvWnxJoDeuyCGzFL4s16hX+2mB7LJ80+qFX9WAySOi1TLlgX5Mly2
Lzan/GEC4QEhDRNftwC7xDZbZASDuCDxS2iPrcij914LxfFBP3OuDKAfOTyOKkWD
OnNJbnszEzdIHQgCsh/geDZEvDamM+XDFsBwpX1JcdgrAWvJVRsE0IQXQpIyzwyY
UvLyA/3t1eu1yuonx7ZUMKZgeuRa1c1j3H7L0In34ryO93x0pQ1hXc6j1kzqu6tV
OCp+3jQ+Uy4oS5GHLH4IthCMric4UhBymM7a7xLsVkjQH0XPh67B81QvViAGQRAw
PPJ1Qjp1Nhe7cKFTEVm0mJPvNb4hgWLDAGv4Ny2+M5u5fvwAybM9kR1qyKDbS9zx
zK1XbFOXhTytr9i/l1qJ9c7Z1A243xSxHyUbY87o5/2TaqfpMBgl1kiX54zSV8n3
kmu21nm18xq7zzpN5zlSczYBxnav9kJr8kdXFb6iLptF+RquLAAE66V46Dgb58ua
recHE41ttq053HcnegsZLAozYYagLHTaGJr1Gj5RBvCjsFZ65uVifxiPHbkV0jZJ
S6z7iFglPqHWeuYcbrGXidKLURSIU+Z6pr0UUi9/IWb/choXeTkC0nG8gX2CFRA9
kOTkalOniBMWZbcbXaS4vwjDasaXTUBp8RCoFCnlapNGCwP6UcsnFsebR1/blCsj
jp3st4tB5gcjMB4ajGqNakrybVp+1Mn77wsAxaqhQ3Odpp2OHd572Kf+hoIz6y0Q
zocufSVm7tH42r30qjWKvsTTK0P+eLNrnWZoh8AtCuw8lypgYe9QG8z23sKuFO6G
Y8VpFSjvuSw783RTZ2CeGtIm1q+Xi4eJhEQ5MTaRCfGNu10Ht3f4DCRBPT5UbVX8
D0r7TNPIWgrmj45FlISdqO1Mq4JXABcwCuWyzz8gn5tOvm+rEH9qn5zRR3pXQy37
j/AwU6cfLqyPwpDDZBuLiDTQJqREzY+JtlHpjJkemPnjCrh37etUct6Hw5nw1TJq
N733y0Yr4NlLhK9fAU9J+m/NurfrZzaKwL5wmr/1owA4JcXXOnslgLj0pL+ClvXK
qh8lGGWW3uM7/PDcGgiLmhkLaZU3qCMP76ptJgmxfeoXDeDYku08TzIkDGlcXIzj
nhn9HFo3r3+ByT2i/3Gw4/Wsq7Q2f3k27HfRUbuKgYKnmP0tLR0tNeYE2I+JrSEU
4xj0fGcy4rxEhIOvHIFOltU+KjBCzzoX4HGbjfGv1FV04THtN+0F943eCW6Wgr5Y
8EIRgyWVLja3puRG9HZwZV9dm5WYBAV9h0imXI9FUzxIAvr6edA/mt5sMUJvmWyZ
JRJs4tEwIQaGacv1pd2+ejmq8522SDWqgPHt/xWfRz1q5u1aGAHlft4UUkxRYsRC
gih/Vt9C7Cenh73Gw6ENwMi99ZVixOQs7CMkTYD2Zo0wLQ7CofsYJ4WJP97C9KhF
VmohELYhGrJ6EqEhcQGmSRaxbhVxqH4S4tAoRMYgAfQkNqKiAXimZiOLElS76ai6
lFr5VUKEFZr5IL+H9mqNwrz98jlNLGM7otftDo3vinZmTd9ytUDUDyggTnyRB7Op
HqwgR8WAhHu45EmG1neJ6VOeVUUU0EcAlNnB+gOHB0yvQFgWZCrsWoZLQYz0Dztm
x3e71QKaSW65hXD6j0JbsMb4ZCSkODK0UPAr3DonlmQt+rHPZ2uyx3xcyMaQ+6Ck
Ts035Cc5WP8jJ6u0aNSmy9ua/ZZLHP/vA1BgN1qzSsaM3gMEHQTAUIq57QIXoBbe
e5hoKZiKjcLNNz4cop5Q/Rlucrlv9C4JjAtWLFE/PaOb8VwojhIEbXXUF66qZ8w2
ennqzexjrf9yRVcBX7EiuMxykDx8W0v2pJw8C/BZEOK11I0uGYnyIIgcNwaOMnT5
vg+x9Bax02uSdzpQbvVyKBaqYKUFNf+a5ccebNnbPyovzgBO/oi34hyPMjqs5Ers
NWWVZBW7ET6AOSspE9CN82qYXBJKHH/qx1Wy88dKej/rjOUzcUlX6ukGL35U2eUf
IdUlhhXaW3iFPdKlPIC9B9V23Pf/CXsOeMVhiBE+T9W4O+r6azWuWppUDntmC6cb
AJOpWiH/AMkbs0RA9yWm2eP5mnh2lwmP+CsxFvkoOu/kAAw56yhQwHF2yvEdIl8x
X2Z4MPcir3Wtxa5tC20Vi+ppCeTY+zReXl/QFsGKXosVaVLvDWrkpxwb7JpNzwHR
K0BLy3YJoq5gjR4WvEkLVPLIpVedXw1PnZEDXeGLzQlqqvoeycOG6iR+PafHXrtv
8SFfCx6jl9Ap4RWJyJ0XJwhVuJvJnCWwXit0qcHo5rY9AJ+GMuRsx0KPoFQ+ZbGY
pcuDHUiOeVOuIv3vXLfG8pZqflpjIdyKg/upILRBnNNt5eBD8eE7WrTJXQriaiF5
1ayaRz+iur6HGwY2v1vZvndmf1jW8GSt7WwaratXRAVHuTrsR+k6OAqap66/IMkh
1KtkBbsipqNcgp+D6bF7g0+zS3lWCkSrgZVNDCbHDkwJ7+Oti7V0PW+Goa9T2u7h
gfUN7DgmMLtHJZXsX3YO39e6YE/yyo1uMjXVleYL9A8KGqcDl/v7taBFRSnjjm9D
xZ/FbIKOsNFo3OSLPKOvypBSVhHBaRVii8NwFaa0fpTS1lcbsaXX2+cPJibk//1N
ncQkqg9FiCXRWsZUYP0nOOVBqVLzpbhhzKdHGVUO1yHkyMBAbbX5pL+RguAJzkR0
yKyeW0dEX0SUtKV02NPfO/lLfdOwU0bZnZv6BUdL4GcuqLpZEwT+zxdPx+uYe54S
HtBzwIfbKDfa6DHfec7w2loGnugWub/tS5aZzcJGJlsIdONhMC2R3Medjdv9PSPu
LldQlunbJcw6JLRx5umgx/pdAWCS2mQ9cdxzV9QYn1ZyT90v8Q4HtOVpOZ8LpzUY
paUOsXwt2x8lRXkK2r7mmZrVw7yEBXd6SblIIeixbbJdKPY/xRb504FN5RFdKPI+
MMb+XluEK+msne7PJfxxdZ/UeNzAlm07yryZL5AbmMu07Z9G41a60Rwr/Jiz+iY+
xGlSQ/plWNL9+HJoDGOT8ALPdn6We7p/F9eBS5052fDWTQqMUpQYxYU5UYq3768s
2ooH0g53Em2AeMWMOLXdKrXytvlHbWqni7dMSwvDAOZ0XtsvsgCuKvxxp7Jpa9a0
Xr1Og6P2ax/YeXYkg/QAptF/XMKTEJQpmRZCTV1q//SaPSMxmEOidUT4Qho13A/Z
Juz/67ekFK4x8b0eJBnxpnNS4KMUAmtkPCnFq8285UNo9y00zAyh3p6f3M6oWymn
ID5//xRONwEI4P3pCHANFaJd/7RthZLi6hKhANIH8RAG3Pl7JYlJvUKJ+R9Jy2Wm
/rdROYYOxrVddYGW7OugqurdYYJZDmhOXCa6JmnUUn3fskIyKvgyHSsqmdjJFseo
Re2Xqo8FZIn9YPHqcZGnSDk1+1jKBJpXLuytrUrPOgYjrcal3USlkJAC2bIr4328
X1bYxo8zwrYOIT3QMHZz3LBaNYig1qkGE7MAH3rxKC/YozwK3S2OYQUsjl0lQ0mX
6JgXW5TrRLfp4UEKaEdI1WIl2KgXol0yN0KnXgyB1AlcOJn/io8hlRv/vgygmFEa
LG7mRf7ztmXav24F6Uo7K7hZRQMyImSozWAmmYJT0FK2b+mY4XPQd14TI6WsVJcg
sjHvILP+Sye4FhhqUDiPx4b/LWqXMTi0kluFFdX55WUs7Lgc2/Fwyad1WYlwtJv+
6PwFns72HnLxQjTZGpmidK+AyTtzEgCj6BSTZS/T+g2JEuoHJcDopb5rowSfWTPB
0uD/eaB+t/J7ysgCciCdMH6QrJnt6LIIoJu7U09FqoW0RUTAr/kM6p6O8XVEiJSO
djlhCo9/wtHifNkDTnktpp+2mn/48fwc31sxyvQEXEZwWTJEPdP1o15rwWBXMUsU
RhurqcTTgttMqQMXX5FS3h57KjWK9L/FO1Ga3rU/jWMDuJTRfN8Rkw8XIzvCdTYl
crGmnpZJR8Fu1DrlW3DRpQuNy/oU7yCK+/n9f2GDD18HC/REqIY+0spCbhj45Ph9
iDEVQpPixBZ+BEncZenPDuJhrpkgDJarZv4yE8mZ4XuVQqDupdXlFVi8M+UlqfSP
Gs+WN3rM8K7W+hzOySVAQLpbC91POJf0ZvXx+sUl60reP+XYx//qM2EE6Zu3AE3K
b069bjn+4FtLPoDKYgD82/jNOar4A3YotKQIoRmg+TsZhheag3XBpIlcux7kFjD2
e0V8W7PKeAHr0Itv6zX+TPHw3yKCf2WSbaKkZXWQmvGn/lviVX2g9fTrk+5DFNtk
gPVL5bGoFI7fTgt8BHL6bXyFIQoYMwzzjl4htTh5ao+qz/C17oOmHTQvbwMSHG8o
mlHrVROIO2099MPmmADGvaKdMJAbN2FG6Sw+jlKMrFrg1hf3AMvGsKFTShb7czEC
8JLS8R4UHJw81PviUqXyd5kFbjTOxzCgj366FhOYyUZazVmEedm7bTmXY/dDJOhD
lEIGHlusY/s0CjclciCDrtMJAj8QpNlBl7wj+2DxeiEnSzKYJNz1rjqwESZoSJKt
1bLsHZX8VP9IhBFeC9sVD5Ftkrp8SGVm4LsBirzUgAIi1mdOt8bXf8LAqDyFZR0j
V21SeC/nmJ20jmw2E8Akot7cERz9pS3ysG5XBOC7N8XZaOdfQnGhvg/2FinuSkrp
Q4zFF2031Ha36KZZ6ypq4HS5owvp5zodDqWzf0zPhfJMeCn0cPKD7IHZ5OoGL5oi
16Y0NxiYzFEDCfee0VwHhY7Sg/kAZmXjQzRFF7KBHoQFmiqaG2g+M7lNVlwjrjBE
g+CIwbNDxxxzK2rN7Thd6EtL8aqBOejMPWsNvf2mvakTPXHmDDWoIFiQsd1Nc/L3
TtnWfT2vg4QaoSgxrqjT+0cKnE8ZdLMRCg+8BYAKwzOwGjIUyf+iZPYyGYIIM2yL
qr1pc9j7SIRPQOCyEcQCp78OIjxMgXVEKrP0j8NS+mW6RHdMkXHNuMeND09DLNbc
f8pPcZcsjCiWn8ZauMYB1UlfInl61MKEf4bPbLVxFyc/1eedUOPPN6HSNFLEHm3+
vUfdh837n8k3XgyGgL5ctIa3c3pHZMyG/lEBLg/5ZRaJ3lnqJPG/L4ASmDgAW5Jn
gDlP2AWGp2lCOp1U+zHCHot8KsH9fel3gViX9MSsDglVypWRHz8kFgZrTccYWwKN
slJLLQycpw2ng7t4OZVxYj4GznBsbdECfP0A9HX3oqsbtpzw0fYII+suKCn0E+0k
1ynsJ10lLwc5sms+A/E3W3/ggpbmDO8BSyDdXM7VSWo8OaxoUGwgzp36FNeyVgSK
AjTMMSbai3Uz+5wM7oRlfxYVdofXtKsy6jNspPehOarttA8M8DCQ+VmmyAr7A0B9
ye8aNbNoHWE7LjBGdDn/exsUYXhQRll1PW9jh2c3tfUU2Alh2yaAT1IODtXN2kEq
25sJOfW8E8xHIsK2FsRMlc4VaamLvCjMvAkjj+Z8VRDcjjvfXPXr7xBdx6QWEFCc
epbCvjNvDGpUAYLfTqxM2Sv98eqTRxEtvwD7TzjseLrXJHOOiapgw+W0SXEV0BYT
NKBqH5TZUNvNPkMej3MnC1UVSx/EbiG9xymaAmGKbT0ELKd5IA4iR0O1kK0MvkxS
lsHos3HOnJqpsKkasoWKvsr4G9D6pfJj14SFDdNJJ4HZTcGHqzJds6nK2OtFglug
l+WmJd+80F6quYFtuk/MCnKBbL7OndQVssQ+sdD4aWJCRa4uoXfKbukCqKC6bplb
p7QhlQm0dQVB0atihoKKQKLTxBxQZUilK3JMEOw8hD4Qsy/9+jcZZZPTTHLSTILL
gsn7E3ooQJ6MXlFjb+uyzaneJFfX3Iw/6i0fLe8tP23kC/oQJAnAssgwkiJ+Rx10
+a9bdqF3RvWnm72j8x9DYAl528CeBeB3RN+RprESEiImTFtOycmS+JzdV7DUsvCD
Kh1EerpcB5Kgx5dWscSioIemRyDUAKlxy84BptfHt29wnJ42rxoNDf3jnUhtLYPR
IWhEygWjlecP3O/4FGBVS/RtMyXXVzVtEU+9bZtYIbjSrevSYFxOmODXEnx7J0Yx
oj/GPFUrr1dEuA33GV8sEs8t6aaEnI+S/1ghNQrZizY0VXE0RaspH8cGmD4m0FoW
KBun54rVRuOE8JaPNk65PKguw4d4xDfiFnAe7n4mVOT6Ig7ettTYb+IySc+Sizq+
cOjgHkLUT68KtN1bJlQrJbYvaiuQgCZFk7Rzd2IhdSPyfcYqs0FMCVVeDKdALZei
jKa/njqNPn2svbHU17vTV7KOnjfKo5GJovV/UJEYQcksVqCWW8byRJ53CX4FDldq
mMA7v4fl2nWhpwYsnx+BFC8a7Bvn6rfvQM0EKIWbCwD8hPvWHP3D+4BWKc7xKsca
4bkaxE/ivLIGtK51zanQBev7X1mBvBStdeVhE4hDJQSq1Bmj+SbolzDE+YTJfsKS
X24MpO/bY1NphCP50HiU1ddy64Ns1SGBlJ2lPHgITTogSyRfQXgEjJItw5vGaplL
tV4GEFzCrdy0pNjol2ciOXsc7APcSu32OKVNQQxt5OPlYK8wsBEZ2Cy3OMbNb9LC
17t5Mt94QqCg981gruJ219BgutqWoShypDJ4H2k0y64O9KeynwGHEHjbZf7h62Ik
ieSOey2/NkM53/XBbIpgQX+XLDmjLdn2jJqNXSMJ+T4RaZC9jyb8zGl2TmrIvybs
y0Ydx2t90PbE01i8fvFwMQYGpQhJwOO9a1dP8RoZb9SK90qc91XIhZkKotu2kEai
vq8BXC5sw5SphVAH4xAwOGXPwgX66Pth3XONB4P24izaVwab6UQtyh+K10STVwMj
OzcjWdzBcWdMnsa/SPm94ThG4Ds8fhUKvwxTIiPn0vjvswTA5rhDuXCwpGw4Nigq
i8lWj+Tkuz2RYl35mnNuRHbA+Jnde33XahtfHmvwLOW/vf0c/r3gDLxExfObcAc5
6j6y2jH6kQhthMEt3G1dFP0tlZUPNW4Oe8hTTsmY7SaMuhOakLHVngCyyWAXdvdx
Ozr5Vkh+kcDv7MAZQYhVGyX4iO1Bzxj29Cz3OcMBOYdjqRMi4EScc4Lhj/c06k7l
Ra9hrmGG1dg9u3dRuADeF3XEeMFq4aq8gSuGKQngPeIzn6GmzD1KP8Ohfq2q2AaP
huILcJNy5I65Ab5PKKJBSmJ9zqAqZ7bhsMdjybcOJo7Pt590WNFAEd0H3+5MDAzf
9QcBTC8j/Ipy519pjkS8enTeCzD+Z6Pq6NFacZFD3dooGF/PKBSKAbLeMCk+ZH3K
Xs0MGpDHZZTyWnu9uRGnOe1MEs4qlAWjFcCEpCSWRH/Ac8phZa6ymUwONVAn12U8
+K9nIaMUooUOQFVitNnT7A1s7MdiuSWhH5SraebrOq0I1sTfiJbZOeJQ3j/shiQf
os+gbUKvizQjtTpugvgKCqzq8mZjSQ9M3NdaqwQed42NAHnICylFpU9uZbwQUBYK
ORIXemKVdPUQI7zhoIumXC8ZgyJpbqcGJk/cz+K8CMfaYqKgP01u2ucpdMT1AeUK
AbI5BGEF+Wq0C68dBVKDNcedrY7+1xxQX2DIhkyxoQLxANjRsktZczWIVn/jMIKd
XTapZO3NAJfayGmYbF4HmnympKGTKcYIGg7sFtGPaAM+NY3nZ4y4mssi8b/o/R2B
i3kLL5uY4FggR8/0fjM1xuJ/L0jzOVF2r95+YS5DG0RW86bhZLVdO+VhSdXpjsoH
JOyDBO2XZztdagosyVBmStsmNpR5cZcx0Fz0y6Nv4gn9VPFl3MTLO+81ie0WpXsx
hTEvjYbSBmiFNtgP3a4v+xNiA/2NTLImp97K1HsNYzMCFa3G4dZOlMLPvKWoYqit
fFyev3f0a76rsCZmYdLJHkctNQNms+2fIv7d2TS5zpjcylQws5ckCNZ+C5yIkZes
0ed945YgRyug/8RuXE5l4aYeMsqjyXBplw5oTnxsxtzL3RhzoHV1Tc8qdTnfWsmb
uGGbtveaZPAVXkgdp8iJmbd16QYTdaQPM1GYKt9/Z1WuBscl4qxlaJjh+4rx2PR3
0OiOO1r/7SWFtdY6Jcv+PpFFxXJSnnvS37TXqvjdDrTtUNoYUXZNBGLVgNrIoW8W
jbH1/VGTBCdDHE06natnyAZr4Py79P39auOqlIFdYMeUvYeUP930EWRwyK2obduQ
SRssTVYsBdA0LXJute/H65fm82/AvKI99Y8/px6/5P2lH/DOiamuqZgdVVhGTnvK
YMvUy7CWJ6gSzuSi3Cy9RK2OB7it9z0l2cxiNfcyghWkTp2w+qlqzVTAmu7nDS2f
k0OGARx5RLVDvtDezZ+j0tfrexQpjMYDHw57I3KYAgJmct3jzj/gi09GBt/TZpGB
e5Re+ru+hLAzpcZ98t53nslZUGXz9eRS64Nc3YGHdWW2noLtSN4kkWvsnnf9oFwz
4d0egqUE7oCeFAUeBt06S0NaitmiPODdS8iOSmHlCT1+lCXGaI8c66N+qXP6aLUD
/PHEXjp7vtSILDaBj/SGb3tDEcPCwwmhXRpiBlIPTFMQB//+C0qyY72R/VA9Uv5i
wBrsIwCtlw0nEEuBn0y0LO1OytRjNk88Kytywj7XUX+T8zcWf5glZhgT9aGwYuTc
U6hAXGKa/x3H50v557fB0HZHzDI51u5UE12fwoSvY910kitSmNcLJb6UuheYguv3
5ytnuQwZtkTC3mDKhXhs0IebpSKQ88++WmGRJ2bW28WJ+nSlvnC7kJ1ANAclzEra
UbUCziXw0V3rYlPlMYLmssv6OJwFDzkpUJiwtlQxtUfXGUOJAfaswwHVEQd8lkPR
CcPgvYMEl71d286Syz6rY/epGYUMN/7DSTdfJz+2lksx9YsYd2+MBIegHqsrMiRU
aBnq9Gn3hxZ3ixWyj37OSNmpH6iFuADwvHt7EtMTvd4TphLtv6dzw2y+UF9Zt2C8
`pragma protect end_protected
