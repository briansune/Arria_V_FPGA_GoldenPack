// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:27 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pNA95sAV9LfG3VqtK592TUefAj+77v+VhzwEijKVoHQjmZWMkXnk+GPSHRcFlaam
z2BFZpMK+sPLbzXzpYUX/DEXRso9NTV7CHxVX2QVHoGuMXRngHq4RkbDVDrvOJgC
snlqgUEPWOLb8EAXir5u/a1bbWENO57DwiiqkxZd8fE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
q/ssyPVjVsUrlNzxTQexZ54Bp2NMAd6XsVOkABicLMMdhaW/EDPXEk2pou29cgdw
MdpE966CP00oeCvkxWFaib3VbRMZxBMFySFD0rDYQ601Ps2id7/obfQSM9tO/abc
CaKOAq4S2GgtD0C8FdsYlnCdchxChwy/IKc6CeECAUMo6n/s9GbX/T/yCC/NH6VG
KXGlt9vD/5017fAa46Br7LfXhL94vW3nHgR1RIyQZTth+xl+6x+AU/450/WGd7bJ
gihLr56vJs/8AfTiafJx1N0xGp3fj+oU8ccwG560D6Rnw7ytJlL7mVysNib3i0tQ
dv1fOIFZUUa0Osq6cSm2DyQv4ZIQUKNl5TFEakKhALEOUuGtE0MdhbgY/5E2p8kx
RkiB9bvN1PXbnsNS1GkolRmNHhhCujuVIfpCmUvo7zqI6/PEfVgH1+GZI93VG+Os
lz7QwUkXUnrUhC7nw7q4joiLBVaAD6W9nZ95jBhX+pqHqdvQ88vZxVFx9YrPE9sp
aBrAmeCbi3Mya0An5zs4PWnoKDqLjWqEztl5ZoueAeBp7jpS/LLsiHJ5HtuisKMe
iz0v9qNNN7rkwJMO1Gl+FNtDgz2nQLbxgU8V7h6HesiT74l1ZkKJVrX3qWOBuCfC
+LFmjoHFh7r5envpEggevswaFO3XGb2aPv/OhzrCHVoz90HDrqkn7PZ33eDFxllz
0oVKCy3LopeBR7KdP5JU7f1qTxXuNj5xkpqIy4Y6cJQiVjtbV6uW0M0nRwtIJLzR
1e8cKUTlP8SdztjvJ5SFrZxbCdEd/ma3DHNiGycRVHTj5Wa1D292R9JqFNOQ+t8D
jLkom1FKgedzUzyJRpj2VK6tluy6XXgObrFQAINqETlMhnNg4xRq728ClwCUyb1r
8Kg4M6FaICugr90zgUSdL6z/2qN3mIYrCrzkoizBhGrSXH/w4Vvx1ZmoA4CqmGez
Jb+t/i/D+OtbgDKLfJ/SFqBmuBMPtcLz8mNDzzFPJ7oIcpjwUrC2rSiAn97Jc8N3
ipQHupBe7HaUKRQ4vZxd0oJhIeOdIt42NaoaqNUUo3K+GMWrT147MjY8KsQ7gfPd
typViBLDtgnJ6SO38VivmwZxwsgTNdnDi5HLco1dsaPswZgsSTtcgDVB9KcLv8my
xYtZJ0qc+SlzbUG/g34uJEFZ8NxtWUaVBto9vj8JLQ7AeiAy5eqtk4r4aplOiyLA
QoBCDu/bO2W8Fdr4ZU6SHUqlejGkKY6yEGtzhIJ6Nv3Q/F/BLhynBdOxeqd2eaNq
ZOyzDK0NAVZu+K6ZStJBQPG+PVUJdhPo2aCQnagk8ADTT+to7TX0ZiPPUxmISVgm
kASZPt2wN3YL8z5PbVDjPYpa2sPYynaNCzGl8qQ1Pgmb7c6/tNMr3VnFK0XRvUtS
1yea8MuSg8m6LcGFU634HWcHOa7n95nEeGCMxW1DBlGef1AWnIOjiK1mbYdYkMuJ
SbaT1qZp5Qe+eHADfQ9Otjr+h7QNTuE6iOg9qhLn95ifime9pcf9Svtrf19uugll
Tks0U8klg8EaEANt0tM0/FjnUjq92ZrCIGiUqinfE3bwVz6ybtrBWUgIkbQLDykw
V5+nc7sBrSIM1BPghvpqN/2rbi7154aBN4JMx1qmwweYrgyj+a3oplfpi+Pvzy4N
bUtP3gbplpvRyppDuoCvsRtJBNl5gRG6ROxLr07pP7J/ZTrvy8uEiaLA/NNLlQqb
QLLq2umPttfcxSN97fQiqtPxzUYKUJxihjjtDslJ/TkQhph9PV5UrPdFYgBjxtE5
MLZCetaFWmyOeFiu6WN8zwX9ddlINDZXOnnfcn00z4ucnvsQKrfExX9kPfATlga5
DkRvKehzJqpfoYX/DW0Ty8Ex9zY2awrDu9MZCl8r96eUruU2xB09NIRVntjVDabR
g3GwjEnFaioBoSe3z64x0Czsz/96ACUjZkDdDTeP4QIWm5AtLdsFmNT53EZ6xPcf
d3LZtgQkapx2hWzrePUOK7ChVxCZeg8aNAn0MJG5B3G9s2hToCqggtC7PC3+WbyZ
nLCGWWG++91/aaFH98npkJGwjl0XtyVqRgWo3i0l4O+3DALiFAeLoJjTOFgpWHJF
a8p6SG1tu/NmxLVO5RmVLKA2E38o4adCAjyA+i14Td8Xd/XoW89atOQSsTbN86CX
nd9Pvze0AvPpJTQQO5JRSkcrZu/v4RAAhcUg5acqv4S73eA0Evc8B5t1MzX0aCwn
4yepEEZxsxMaw/2FvxImR3QNLaXBaBMfUDjdFjuhS+jvr/bK0qGF+VTIyCOZQWtC
dYLNhn+jMLzBc++3dY0EeBA/3H/zghme+ni4VUmdt5zH58eaOBB0wdojYuElblbj
ILW4bnOgoxOjtamdcB2wLKODi6yiQ6PNKTI9jIBbjk532prxp3Ao+8NkbKfQJGG4
i6l6VnpdfQrgBltO3vFRQ+txR5SFidfv/VPc0iBiuDdL77HfD2m95y7SblXP4Zsk
/mmEq/k4OHutBoPqsVJ+PEAgTC84MeEpwZFkW1dNatdKnRFfjgod9v7sjKMuD/IL
PbKzQK5wYYUO8AOVtpNCNAW6K24lLVt1nKRbQUFCZ5dOZjrS7v+hhagL9V1RWcXW
pmej62wDyoPAwxspvjyBnEiqQneiub4gKN3tJVl3zBCybONU3x9wcIaM37Wscwo8
AsqtRcLsX7MJcM69EhpQLIgCXavQ3BaxL6rBFiGhk5iH0TnJvnZ94DE1Q9Fuop27
GMw28OTemBQdL8OKZLQz2Scxqon5q3vU19voVB0IFCs0/U8IQLe+NPjdty/8PR5o
zosH838EqQiyS4ZcKfeLVkHyABAdiDVeJC9+Q1JPhvtCrWsS1YvI6k8fajFnMTal
QiWOssIapixFqBjTEU9zqekizEZUBjugsHbNHlfBhSbkG69cvshqUGW6i9Nk4VJy
vHQ0W35HxeBaAgtx7bqnoodetC4Jp+keZkdx0WwakvqfB1A9ktWBMd5Vk2AQ2Quv
BLnsRitFARnM+YGINr6BzTyvIGFgddcRmzNWdSBReKK81NR4n/gbAq4QnoPPuH2z
YFHNA2d0mhuoZyLDuKpJNlCzokLhHWsrvB2nRaDQfBhasT/UQnXL1sGe9rnoLSSV
i2Xh01C0c653J3zZRd+ERzhhXhZhlVzyRQHAK01b8Zi7qYIsjJorpoMsA9qpg9TP
b5ADDmcWx5is3ixm6BzUwetZFWR9PhInRPOzCpV4vpM+kocgaXg0iCQaI3o0JA6g
I3dwUBrp89AQkL6hDx0JQJ2c81mBbbwBsc8YD2JhHRGU0JACVzRgnCPAfeEW1wJJ
IKCkPZjYvy3AvaFyeRTN8vTSAWMXA56xBp0qt79/J6gCIGXmmQ5PE/0P9Gxcq/lS
V1MSZq58q59LtkPUOCvrXy9DIEfWWikQct6RUrkYIX10QN15EgmyS4zkeNyjv+Xv
iuJm6raPh20hd7aL2ULIjFculLgl7dt/rkqICu2UPEOyjd+Bv2AmdKRBwk5+hiKz
LrGA4NV730xKANBUf6OEL6cROVQOlbnFP5ErMrHbGIMPefBpq2IFsPlhJrkWbnIH
0foPM5WTClJgJhuSfz32DxMJsrAQkdvAeVpF9W4fC2qfTmumeVIgL3U44Z0O4bUQ
ow1M9iuNHanwIcb5a9y8X5/z8JAZZwM3+1K8oDAeb2iohSr+ZjRO41Xl5xXuHebc
cozHzlthuR+GODja2U0G3a1ZTEwMdju3uSCmnMF6JGjQOyVsgpAwQAv7fBM7tEzF
EWG9AePOy0mFowoctv5KYXRkGfFTNvuD3vktub9T7OujhoAAKtIo7mpAXwh5QTvH
PMbf/0jGwda9DGuzSXuOZ2IYT4P85SBcnIIB1+gDVVoH9O3i/hezCfRcO6Wu45sq
/DONXr6g9zlGJv6bAvP7nq0FxvbK3ctV+uDq+BJiKBDT4r0jnPc1XBFOnKLr2AVy
guVwUrKUAZXQv0056veCQLAYgQoPtFoYoSbaf5rSVl/ACIV3mRGRSPiP5MJQ9qfg
uWApTrpAous/3Ch7Fb4hojYBmkw2UB4hbjhEUqteLsNT/m9TwB8uNTKXwbtLrso1
n+eKAIipFJoK0iumHqWYoPdX5G+rBxKneZT3FHJZz864tM/jYvSoTaXj6C17C664
PYssLh3lIQqUENgI5cZG+XTllLj9xdbVdYmvGRGPLb9wLd3rpgluORv4T2PBX84o
BLFKgvJ7yhT3ZykdrvgVcTJZYKqNxboUXwbcJcSAmAbgDIu6tBkYpcoI43TQd0Lv
yjdXjf1LXkHlQVH5qYkRtiBgJcfC7J4/9O/i8ARUfMabEY+JReYpaoAoH+sSyKfP
alceejF7YGa0rh4qF7+jHLGW4HcbNdrCWh3LRlTXyVFEq8agrBVHwp0JWHYaYf+t
qPNxavfvmwRHSlf6t9H3Ws+vsWYTjEzjQW22sv+vjM0DsfrbhwvlhiMfxT6zLZEg
CADszDq3JHER6vM8sE/bVI2p53s3/y4rjxoZlPqaZ6wORqOn3lnCztTeXNocpum+
JhG6zflyTzlAUsAEioBEIbTtSHyXtqtm7p2cGxzJ0+VqCor1+snjTmE8szCM8VqB
MIBjFs8R9rUNUbMVZYZN9q8v28SD9ViVr32yb1JejA851ReSGW31a7e7JNFsgFQk
9+Nvpw90ktg4CIR5qwNlZ2cC+Q+C7A1/MHHb1+mxZe8TvMn4twNRUzMO5GOF8uCI
SuVW8i4kGOXG4oRClVP8chC+kZ3zFgZMPW0JDm6rTx6P3IJDIBpFwUNbrn9WdsBH
PSssd1k5UAaVU7RyPb/CsllArRm6GX157uAdjc7TEqW2KLX3ylqp3AH1100jhHMT
cGZVO0CRj+y2FJcXdguTRmXbj3ZcJfs1QeX8R7bwxJu0qXBmyo0rW/KCaKGGPNXO
/cSaBL+VUBHajgbWmIT/wdVoi+yeHeA+afevu/EaBpydyGyUMXXOfpozUUaLs2D5
0LEDTgFHrnBg6Ygy2f1xIAImh7H3KNlOSA+rF7DO2OqEuK1OGsC8OeBJk7kVKswP
+2fg72biw24i5hq6/3dWXTy9uYMhqCyZ7vrZF0dSLtSoaDcqfuCgfwAkjCGT6+pR
Hv4z1Sa419l0MY4qgogaPMUP7zsYYfbUu0/8cqRwTk3JcGz4hn1U2RAqZq9IAxKS
dphHGCrUyLbUSTjLAQ4vM+jovCwHYKwDVLuMhGaYWXyQSmxhjDs7FORtMdkkJk+d
cMUMdTa49MWgawiiyc31sYfAFlMTWjnJ0WdLZGwJhWOtvrE6oTtjsSGX5MGRX/oW
Scnw7GsqQtEeN22pZDrhAjPsGVOeie50bCeNDR6YeHa0VB/otuUSJNMtcEHwxB55
ErhYBE6uqP+WPPdm9A0tnYDb/44h/o5jRYpXw4XFkyUqmLtMRrG37DdZrqG0dvgC
gt9vWKghunGC38Xw2lGUy7C26ah84Idy79vnMEaG6q9+55A0iH6fGIYQ0EW2V6fP
7fLNzIqb/lx7oRBQNuNKpke3ItPA+Bv6bZEjDgVaOGy20EvNLbyt5a+XGKnkWKUn
DoUQy9CisZbCmLRAuGZMe2/j5jSwgTt3X8zsF1NsaXswFxlBZ1ej9dUlok4SaQ2i
APC84VNqCaQYB5INJD18c+TDICkGcDeuXGSd4rYllzGTDcXvZJaUgZeS1hN/A1Qh
GGRh2nqfAgIKSYmNGMCHK4JANnAipyVAdS0+R2NrcBpSBD8+XKun6og/izHiuTIC
RTSh65VLLIDHL+wWcItCF7aGuyMad4IR56nRJiPR1LBP4XdJkWMGUvGbPjdYj1VY
l3+67AE0BsZTF7tQ/ikiaFcqS6NSQD7UXKoRwSWy7fbpiofNnauKgKunTVcI4fA9
uPaPrkh0oUyVCnGQ8vqUlY5gfxtJulS4RXbCPxXyCeykaUe1jmhzjs0XeG41H16T
ptGYV00dC13WYB2cQlqwItv/s3NMfBRKViofkMvqCJfFa3HyZQwMIFxdn6GCWZiA
E4KkXTcEjH4okfuCWIux19YQkaOnjRxOoARz7u/IrCvoMBVXXZIotV2JQEaqc2hS
fbBk2fjXnwP5u6iwq1tJBtL64jV6C0qh34NCC6vF/6CiUUvBJ3IPuW405SPi3AsI
IAsyceVRBNkJbk0O3xpMIG4i4zLmqAXj1rnVr/l504y05NTNPi0dKIOJb4fGKhGx
JraQn/NkNcp5+VSU2B+ur15dH4p7HwqESrqvxLlDDFbEvD5+KoKXjmLc1rRYqNW/
q9boExwlE01q5hxF3S5NI3CuGCdO7dUUvAnnPQFG3drLrdmKV8huTPcjvLsw8q4t
EKaYDmD+L+RBYDIKTbGREGVw8Tt+YyGx5coRYEAHd67Z5BbaLP1Sd4PEqST7r0Zr
kuFcb/23ae5UTqIUA3TvL3+CTUQuSA8ZpTUEf+gDjCM/Vxsmw8ftImKObpzUWB0C
bKglaiy5y4uHICkEvAejZyMm/EOVxZ68OE6ENEhpTp1BHVabxQpPO0ZZlmpKttKF
tk9LR4Eev2iuo+NxnPI45L20CotT50XlGjJinMG60spn6N4vzOzmTRldynixtHPq
e4oAB4+9fbymCARx5jytRtmO6O4TTafcGeC7X7k4tA+wuAZbZd1CeUaPxGMEcShV
jifUNRDy6X+pVvEcFTvWUGpN+JakaoQdBT2PYGaU7lfBoP6rWtKo8ncIX3ETCqEp
CCaiI4KCLqIcX2o/6C2ZUYwgrnj/PISYVorxsVEiGByrm2z6cC1uc7IN39DFwAMk
2Ll+i8jSbVW4ElObm3FCTrEshKGTVWe0jfg3lUhZJCjD2Xn3LXxoG9+ToSE6LkhV
XBr1uCkCMtKunqv2GHYN2CQ1w9JvHmYFJ4KlkS7jr8bjIga6rxFgOI+0kTfvcIaj
zcbdbqVZGboXRaJggKO9KNrSmGnrSw8CPZDvAY6ckznVBHF37VgoTFxvy8jbi9bA
bVfGTtkAwzA6G6eyCtmkXrKG3aqXqrb8J/uRMKa/z29J3jzFUTOMUtEShRsDVOTY
1lN4kNzPyugjDycWOe8Qvyvqnpt+72Pr5+l61A16eyZFezf5J8c2zxY/9HVXXRkA
IEKhhTXLkN0atcwbxkHDE46seJzSJz1bk+F/YHr531dixc3hqwud44H8zpDdJ0ci
IgZ74AdJdFFNeYBgQ/mCyF9ROvgpRCTTBVKE62VDLv4oNO6g1xpDHX+RYLjTaXdq
WOaIAYAjwwDaSiOq5wkDGc5fJ4xqlUdytacitX2TVrc2p6ESGKmbByR+CtxikHPK
DGZd3fbGH2zWHLtiJwUjhHAiZH/WVy9sIeRnxyxAFo5Tit9K4TSGtMqhMB0tbJFA
EQROSyGRBahTaOz+63y2Y5L+6TyXXNUAsks2O0FkwUTmkFRcAf/JlHqfmrheOWMZ
Pl1TpIlyAOy/zpIxysLqvZL1ksvRWSxXEuW58x85w1EZjWh+/SA/gA8uncBpA2lN
h/UGsAISEix46091KHoBE6eGzpoigNKewBoB0rqbVzX+gECeIBlUrlDoSiZ9D4Xq
rpkL0jQPZiUhk7rs9YJ57ZMEIfLDFqkaZzesP0R5yO/X4i/E2ugAQ4fpVxtJd+oM
cWEnhq1pg0aXx5WNb3bIrSOx7t/3g8h9gcmk3si6O3ulJEkeoDB42HAlVICsMCzf
xkkKdp9+wPttrASQBt3mZi1GBt/2R8LGiCn8pYyCMY7i2dkbAGPkXmiBGP/yBNgS
4GDHDmu0p4x8TizpfopWKq99XoX7mBNWX+s987SP8OZeQoVH5qhL6ZfC1pk7avwh
b3YkVlzE/oIJd1HkUUVUdJ7qOzPD+qxuqgLtIxAjkcM90S2G0A0d58/iuokLqKCQ
dBbVB1t/oa6b70h+Z0Lk7awavnIBBGUW9ZsfIZQN3lETetN5bZ75LdF1hakNEhj3
CaGgEi5xZjx22AQnWzf8ZMGaYqw8p+6nQnueKRggbju6JEUcD7jFb2y4NrXaApTh
q3eyx5Cqy1GQPtKsVETRTv8xJ0+/6ANHKIGBZcTeA2qqagy1ec2ONuz/e6zf95Le
mxA6u1htH0whptw1No2RUaNFqFjjvL4oe4htdtOkBhxfpNlDLHpeWogQxlvNFvcW
U7pDMvVlVbGU+q6LCYXwSejf2TFaWyhLu8RtBDGmgamTW5P7BJAvmOtxHxg4rdDj
5ZQ/EGN0BzTjZfVCz7mOhl9CsTGUKfz7A/TkvlxnNvZJDzhYkxBEn+PxF9DGxEU+
JfLc54P9lTbB2exc3RPsYFQLhM+ro4MZ3O3Uazk9/lkl94EtBHR+JyNHdpFlV2v8
GYeLOoE3cJVNy5pETYhdVad8lXKVY0fLd4HgY8jf54PpymRGIY96laKOhNaziskb
T+qRs6mJoiAw99EtPqZ8OLmaLksjUEW8RRHJ4gwPEhOAN2u7fTzA8Dj86P6RsLDS
7Lsr6fGk5W2I130o7mYzCMpRLjz4ILCQZN0XDmR4ooqCRW9mxmgE7TnwgBgGrWkP
ncO31hXVItxws9SYg8l58FnaXz/FnCNvXTBUZGNaeyRuM5cBWDpTAOhdyoL/r4Zu
5GU1Q3W4yT2FCHGY1wmKvsZKVkApNxbf3eVX1OWyBNMWRfTpHkYEiOy4hgBnaQc6
lErImI9v8tqQJhMbF/htoh6s8R55hubilLNmCqmwO2X7i7ScGx3XMgPh/DKg+9aU
ahTm6wG2msRsN9zTEOWgsWL9a0loUXuctXuz16knmCYaFRrxt07/pC5Ip+15st7n
XF4FXJNMgP+MLLTKnbcwXau6QEY6ykYtYflxLjBiN9oU4J+dAszBUglxc+q01HQR
0hXfNTHhUJDEIrJcZEavdg1jhC03gIPgKn7TxF9/oHzCfNWH9tfSp4M2iS7nDZ9q
MhHKoemaaK6khYJvoEjoXBObdfoey4BoCd+faZYIQUpkQZHIcWti7Z5VPzZKgUsv
1dlz087/r7e7q3ASeJWQsUkoD312ht/hH3or03apgDmElUaO6v22poR9Z+ZAYpyg
Mtm372t86UIM8jBhHDIQgothzk4VFkdfNoDeHqvHOoKZ7PMEdkR7O+6799vdvcS3
cQuYHm54tcN9QKrkFTu91SlU0gY/nDA7e7lA78fd44RtkpeNpAm0Rx5i9pGkX/CU
xrSSiq/mKqmiyNfV3LvdaAdHhpNQubGHG7PCLG3KgwdfI6j8EzDCN+hSjxwniHDB
XiwGpTFh47gofekAubR+5RwtDEIu5wuKrKGTyal56k9Z52/x5M1e201tDf7CCqK1
u9A6zznVzBxUuoFh8SF2R+Vhv+u96xnsjNpJOkAtNmcBegDLQcQu+RijTzqHv213
XwrXrnejBFugL/lS8x2UolUVzit0bZxc16ma3vu3DAzg2P7Dwizc6rfy9zftJkIC
BXEz23SHi3CTIf0AtoSZH/wyV7ESmytUAz0kMyfppIWLEJDG6VtEUfnOfz+8ap59
GRqqOz7fvOJWVuOO6A639OCi3cZcsur5FimYPfGxQLp5wLPkkbJCygVsKpwizLzk
q6jScXHwsza6jxnw6r8nuwjpTxWyHo4nMUTK3jEfUBew03JOyvxW0k9zd7N5Rbw7
U+hF4rGxVZ3nR85xdbYyferAH+f99UEbmWJSbVnI0lRy8gGW4jwp6kqao5FpQE2R
eRXYu/2RQv4OIFDdbR+M6yRj27f7VCiVdNeRm9RAxsKYj5OtQ0LW8wfIy5PJz3rJ
6lBlXCspy1qpxMpHbZs63ZOR0RNyjDkpufOUE2lnPL6CmVGpXtN6XHE9xxWjRrzz
NckUNcuVg7o7Gk7z90UIdh+WhrYIHM/FmivvnGyKCfjFtJA0ffhf4Ue+hqu5qZb/
w6mzFN9fggxm/5OEfEzNmaXkUHbBhuY2K4Tvf8xNLiEjZlqY9kex9uws01PfyOs5
u0T1V9L+8nhNLi5PI3S53+1TUI4X4luPNO8Y8L73mZUM8dak2zjb2hIcbkHf+VB9
6Dlhk4wbdXbOi7oiqcBpsO/VdQU+1h3kx0BnyItSF5cwSQW4dQzW2duVRWAYZyvX
aWYpN+AgrSQFVYKlxtJC+htOwx3jdv67hEPKP0FV1Vg=
`pragma protect end_protected
