// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:54 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U9heCV+KE1QW+PGU6kwpL3NrRJF32vlsbgwhiIfOkPLIKuhEu3nYPxBS108Ir+li
yiiAGzYWKxUl/ZVILHoJDtDQXDByNa3kITUs8MWb2rq/IZ87JHboWpHwJjoUZaE2
Gg5Kju416GQ7VBgxpz4tekTs8B/wldxFP9e6hMzOnG8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
LhrUUCCTgPuhYe6CzRwH97aZw5/JBXsO4JExqC46yqNmf67Y2htjXgZPUf6w2krf
MUOjjz4Ct+Mq0bqRiF8SYQramsKCG4zchYImMOJqqLcRtlnr8TjBeycllOqT9lpk
bSltil5w5h32y1we+66csx24LwcjG0WIS4FKD9Rvw69n6hWHzHTe+MftUETxD0vV
brAO15Cv+3j3fkTucqu3tGoHSwzPhX2SKeTgJLAzKjxo7kn0zQ7HlqlAJ0/JMlyL
veKk8DtZgnAtEUPcuxbRswWIACbxSqidouLw/izB7RmiPpkRkJgGkXnjgH+DmeA3
frV06X9LEdDGXb+lXsIHncsOoA42IZ2b1eiqhJyFq6WPCX1mjkTLL6omESO0J9Hw
35Fm1iQgVYJaKIiZhpAxUDsb8T4JywsAMT9UbkwGY5GFcnqju7DsBA4R7l31HRWU
iamFTUh+uteBASKQsC10ldwp/TaV4WPn6L5e2cNVfNUuabtQCGFeMnO6RNz2AJrh
rJFTFJUg4LHt/VYxzB+u1jN2zyu6LsygEF79Yo2mjIi2AnKag9/r5WL40mVI7NlT
UfoXW8A16v7tHCsv6tZfgJ6f7bquiO/F8rTX58gsvzSUpnuFpZOj0taJZwYcFKGS
uvPn8LDScs3XEiPfqHbN9pmfTVbtaY2jWW40Y5bFw4E0xF/fOptcNmiRzYFijdne
oUn9X9/EKP+MEIcbv1eCkOLIFm19NE/eW4dgKNCDnXr6WWjm+ZHkj42kqb993spj
6RtmdL4+GY8aufoCZNkuqpCVHhz1yl6ujY69kBvNWuKxZgdvCRGsessmhZDJfw4k
Nlt+EyOJB4zYaK05UHJ2aRu8AFKACe734rUxxNy89VZc695m/CNKIur4s3tYmuYp
XLQud5Llnqoh/59/i9GqyEzwOTYuvT9qY45E/Mhg4OgfkfMCscOCvnQZjS/9cS/I
oQPUR+5SYuUMk7P/9Mh5a0B28SxDtgGBB4xxFhj9wUlyQmFPWaTRbob8XTpYaFBK
Iw3J1NcV9m2Iqn2IHVAkR/Wd+o7au18r+k5LSID0o+IS/BaMdyXXZ8pbzaGzshXL
xJSHnKnobZUPJMz7PMoZiRJvStSMVr637tdSq9JPuwWAZk9L48aq3y92y+qdcQF8
zU4aGCrBaysZhfxfB395QognSXwvmC6WHFnSm7L2jy8hK8KumGNkFgLoenZZ0cnL
ngt3H8ZAj2UhxJZI2P/g6Zizqe8BwXSfFI126apcE4aM3AME5lyYu/dueD8Lp0/w
ZVCcE8u58scmarNBNiyt3uqYbGY9hgwiQO+/ylie9Sclr8qrc+I+CawVBh5zCqw/
DXYY7o1h3qaEnNjZdVcUt9jVaWIpPJM3jLbgbJiyxKWUyy1urnT8i5d1aawFAcGy
0nwDtZnDLaV2U2U2whECoTMAhnBNuevReeJZCKRrnPHn2gmXzp06QHUiA8+eEXVT
tm1I8PK8eOECIoMnz8385Lbo8BsJhKNWchrMHC1TZblJGxsOpooV8hwElZ/g/4wo
dcEE+lKLCkklFTcnn6byssb4a9Y7jEyn6nElOSbsubJnp/VpLG4WZAcj3CzGQeqC
PJvobtjqqU3fty+80BqC9EhvRKPezNK6Q3aH2DCLZcyhLjBXBxcERrbSuOx118gS
bu5QJPiO92+1uvbuNnRd/XxUr0I3vcWnNYPBZFE8NHWKJnOo69YA1VpPgM13c9MY
fEIToGvjhcahT4l5vYMfiUhJzveCZ9OHkeZGF9d/B/nbQU0JciWwukDajaa/MHZk
o2VX603TL47Z7r0NM+KUMnMFqVAQmeb9lP+gKXWg+t+dN7t8SqaYsREPu1MSZBxX
wxxSeP7TbwohMsofK7Sqkpe5puvhHH4dnyI2xLTi2rBDzUCSgRi6wJ3YcQ5sIA9Y
+0QwrR78LFtvBzwV75LIJyFCtIGaCNdkonqFldxkO6Pr9v+XGUPF8PM9h1psDB+O
EfWpy8+RN42EDrH9oUwdv1kXnEIUTIL655M0oWGsfRGpp8/kfOTROCWUaMShl6yD
2wxohjKDaI8dg4crH/OYRu5ud1FiqjCO5RHd8vouzCVuh6Hi68PlS4kIC/Co1mlF
HcjfXCU2TZrIs91FMDM9ksaS2vX34Km3Cv9Ybn+4U5GezEN4Tz4ERgEObphBG47i
LktVh3zp1YfkVj/m+CBo4NP7WwcJuPgAITQwxHghWwhk7NouLL2YRFkwXyEGrvhE
S9h2G+Ab8AtQKNgNz3QhuFs75FMWEKfjS3ZneQdeIiO/bwa0UXs4zLunNSjwteLR
T7lgS9t0aKT1aktKKy8QUYsyTEXqjHTffZWzcrjt7W6z7UCkjloPWolu+7YR3yT+
TCI7fhoSAKFgASoGAhgRuoP/KmLAm8iCW+JEIViFxFy9IXtSVQZCdHszFVGYLBao
X6j+syOK3GRUmQvPrtetU9tpLIOxamwsk4iNIiX1fQIAlHa1ffn3EHg8tHpSk7D2
M3Tw8WOPVY/yz2FxsvIux6vvZoYc0ZZ2B1qUWYz3z8O+DtY7AmzpaQdB/KAFGvr0
DUloq+ec91shPy9cix/XUuq5x8CCGIRyoghuq9LyHQnTKuLENhqv7kgo3TDGmPFK
rzlhmZqDf3uGTl84f1S8vTULrZJkQiSw3K23hoVeqcv1mKmgs42quIgIu0sdJdV0
XTOJ00tT2hZzhApcukvokMx9CrZbyn90JTSyKcpWjul8h8t4hVy7iQW4xMmnNvFl
ec1WBeJZszxFK7GVXl/cAE68niEk0q6jEkoWY68ozpze1Hm2u/iyFa5y661aLpsJ
8RDmw6y7i724y7OrRHRm6QkvW+A/CHaWGJntKjTAc5naXHjoKbIaAdGjgnSUzyP8
cDEuxGF4a7GsqIkjTTkZYLMDSKcyLFky3t12mxh9HhCTKOuYTKgbWzCUO1DIDTWS
YNydLhsjBb7YyJj+OSEm9YmTbXJ6zRRhq1NpBzXzndbJlSF8BU9YTDnXWVgKBiYd
gtnm2P+zdRPD1PpiQzDIHWEdCGffMLjaYD8hwqntqC3w4UYLerCXM0dVg3Qv5Kb4
EjXiiVT6ZoOWmtLLFSXFTv+VFhdAuSmmo9tyAQXvU4JAqVcSdXEkCgOo2IE8+jLS
uWnRc9XNaCirzg5trHvmqxl1ed/MoQaPGowJ3P1tsDY5COzMYb8BSaW0nBlDeOKK
Vftp9eVClT/xpcJ1FCWP+exU3oCscyLyJSWDpvOC/hlXRu7Wa/BNczMY2s3VhJoH
DilFURemQCbMNjY2an+JiQINZ4XjllgD8rhxPkAI/We7dF5LjMNm6JTBQnrKhpPw
2TIfmp8EzZ7Y53P2XupqUHj3+eCMwAvsZ1jwnwQ+QDnXGBosfn3/SJJ7ZOvq+FMp
wc+Kle6Cb7HU93kaOi6VL/4jNm3O8tcTbhVGZgmTiZ/eshM2pluWpYiZPlUVoWsv
4QXvR7fc9aZZjq4F/NwIp2nu7lxdQRu7Cfy7V55wRqS4hAhRQ9YWxhUD1h0kQzNW
k553xVaaiE94M2zTdGnt4e+1XpESEzIKjHThNbwNPHnXfQyg8oLCgE81xHtXX76f
9/8VbMGl3YlB6eOdafhkL8iXkS0Psy+SCOSap3AlrDBaAqPa9W+gc7j35uXUMwYk
kI63zbIOKptKA22xQpyG7h82Mw4aiQsGPf023kYGvj1X4eysARj9+YL+p9oGK+SY
cskegw0EKCumsDog6bnOz8ThIQzIqGKYAAPP4J7xTI6Vtq4Q0SrIK7gmLcquwB19
o0hZ3mXj8SCpHIwJBoTu4oVQAYpT7priRuBjJkfIR9m1WTTx9lssvIDzi762n4uo
933nRddha2gf95EdTke9GDfSoXcslGhFMtJZsSaVuwMZbvi2A5oazQCvm/rTs8xX
uCcvmCo6TR3fFJEG2PW6YmUZ5KC6/ay3Eb2eOlpaC/bQ8/a+NdKWea+AoXPEHv2s
1g/c+0IhnO2A+13kFqpAoWBj6xWnKu7AoMUihqlMc9wEJPKRTIVAMINOWcz4QXjH
QL4xI2xNXx5gVPoYePMJ28Jll5Q3AG5NZKJNzac+eT6EdHe5YtoxNvSQCKi09ZL5
UChvfo5FLnunoU5gfW5NA0UJiydjsWwa7DQ/JfC+K3/Cfe6fZxcXdWZphEFYQQau
BQNFGPx+gcCLeE5uKWl6djoT/JKXbn97LBIHqNwEHW7tmauVnK+qyS4RmoIX7x52
1ATorue4coYnmihhKJ/ZZ1sL9RPp1D40ZakNjSTSxM8sUkuBCRvTYuxwOWh4FeWo
bM9Xiw/EaQKRwDpsFtYy0cP263ezgbL0yNNKf64xFilHxHgDRORYqIqWUjISmF3W
GjyL3SEjTERvw4Ykj16sC62bdygUDDRl6E+kr8XZAZhVAhHStd1wOV9tW7rlYpOq
D/CgOcSg6kwWxS3hpe8dBk1vn8z4XQawWbogkA2uENXB5K8MtcR7LNmKg/qjgkYH
YQDVnHECww0sMSVQ6wDMxtgnc+fl0H/6XmY96Y5VfABLbziXuGqq9t0wz3fnyQ6p
e0+Ssnxho+0HL8uk41/pSyw3NIDsc9RAUweACQArkQLTS9IllXNLCvSDspIXTyqz
nLt6JBRNWCXTZn02v/fA9cXpWqarc4hKuJ663L+W2xnZQpQDdSUBtduF4cyonQnf
IKrfXjs5YsXox72oHlRWUfYShkXC8oyrsDxCtbttUhoMxHv1Za/4oURDfzqrP1vf
oDJeAawoGkG/Z2vGSfoauJrT0FtLK+pRuplferEaYa7zrm7KqnrzFBdFHJ4cYL5z
NpXez7uf8yOLuzGgUsj50WQcTCTsJPzI503V4XhJzCfTND4szMxVkpNWZd4ArABR
kU91m353EXkKo7UI8hW9c/+4fV84ZqbA7T3LfyKdv0mi60H6En+z2hp+aCJFqLBg
3nMDcaqUiu339pstwg2CmRKhmanKvIv3jdtvLxc0MqWnFp1AjojGKOw47L1c/0+a
w0j/q5Sd824JhwPvgasakPieKOE3/Y5e5+mx3zkA74KJSyOjG+JED8K/X37Ahx9H
qBU0qRN/3tZWc5J7v6jIaEfZzHUCGJSpjJpaamHJbRedwU9JT1bCPMV7nmSfbC0v
uxcvPUSVkSQ4U/9pi/LqYbUKgnELE8jgWpkOl5dxrYImmBhIthHqcIjOd5iMAOK4
xSYydcT88ZH056OOl/KXVIqpBttcLUaf4owUIX4jpIyxXCxl7+v07R9UAgHLOVeb
F4ZmRuV37LSlmxwvAss/74P5blcgFRDA+91Um8e9rnE1qa60hPNIpro5VTNZo5Ff
k6yyc9OzUL8Zdi8UQ3mgppsTY29cV3ZJkUWYaMPLtivlnh0uW+gvA9b/I9WeJKP4
2c0sPjl4mDvEXE6fQLk7iWVUV7Qx2HEQBDKVEKhf4tqtIkW5EHucknWj5b19xEEF
Q0HBVWAJrS8w+69eZfxNrv2X6cAICCGz0WGmvGvSl8CSr6gdjqczXC3DkEmlsS5i
5ZEQgiuK5dbdyCfZ0Kgy92TrVkm/YWqaOiY9hf8iC0nrYuTD6gBquhNohJEqs3h7
0FeuZaiBctdwSblt3BaeRQy/OJXB8VEM4sLBDrN8MJPiRmZoZDGXxW+I5l/TL8ll
15pRLuDXoZZZQcZVZlr0mxgMlai+mxS/4+9t/wKltqIaDCyiYMlvWxrheHgp9O6r
Xs3mlm6aMTIpvFAf7jDiBlJEbWCIvSwNzNstV/w90o73TmsurvbzPQcaNMFslUBw
Fra2kny+jN6cZWBNmNMUyGSkaBqGoNGrTc5UcdxOiIWjFJKB96UgMFAScIBySQjP
1ia5mS5I25hpclUv2WnHj7v7A8OW4KAByZTckTzQ3+4WtwLG3LdmXdMa6DQ1rKcb
kQOTNnLORYztHhlKS5cg4jjcZSLIlAi5LMUC8wA9P1r7j75q5cWzjj+h/x4f+YFn
d/LM9Ch0Tg/no5UJUiP/z/lU9mRvj+88okpcbiOvgVNnGA0nSn9EH7aFn+5W/eBm
ZD2SJMPCsVz4RLG69FihuifudRoP9Uqm8NddS7q0/frdkqhvNkkNKADDGIxLIXCd
Tj29nZ+FwDnFLe8+GDeDy3ppdzc5C1c1Lccj1bhEHQ5fXS+mJ+WktMj3ledmxPUF
NmL1mKsiHVQ9vhNQ27S2pubk9UylOfRo6Fzwp9+L/IlOV9OARqU+Xop/Cy5oKdcN
kAYiA9owkVUKDIWVyIcrx+tPNfrRbPjb56XUXoRVDXO3WSFQx+D3klvs+cbwLCX+
aAzrFXgcT3xR4kFkPIK3trbq64avU+6eSttUphLNTEccwrrJX6C+WQegcLz8kqMb
4KLgcRvOzmDPDT0CjGVq62rCqyH7FBjLboEPR/DwUncqLptBFs/FvU+Ewk2F/rK1
isZ7EPEVKdf7rsHtHfydpYTOIYj5ImD4q3+G3SMBg2aQH6AyugnTodYa3/YRICgi
G7kkFZ30a8Rtll43xtRqDKUiGcIib6kccthwlQ8qvYM+1LEDuq9aRjcYvrVUSwAF
SlcrHF9YuSUqQtwQm9hiIPJRTXQROwd/1XNllTtYtWV0wEinXuFgw9DJXkihw17o
orjY0b4+1I32IQVtl9B/zDOtsEWww/6DcHSpwFQBqGbyfYQLDkLENu/4yftUnase
aHePn6GRH7BLU/wbq6SrzLyWGA2dqv6V5/mTu3Fmr0fvBj7mG+qDwr/ZIOkhdshm
EQEjCMS4O2bzF4MMz5BDNjjUeqwvrqrQeUDAoDp4OVE6VTpqeHxVUFnzyg0bvZhp
fRJx3Ridjjj1rurR5ZVr9I3RZUpm8GIPDCtFd4bmaqN2PUfNfeOjswjitYDYL036
fgVLGh2HhZoW0yVWPCBO6mGibCPEyw73A+UgWKyWpD5rUCQJl9gdEwaK8Oy6HNTl
1NUUOxqpwTkiNgmjhORxRLytr5YLDU80NxAvpw6pZe/I0aEGMCGsQnNdXuv9gyEs
LKLXDh2epnUZlSpHjvq81r6p8BsQ56TpjzSP7x8Id5ycvN/xk4wzn3rgO0ektLFj
p6H6HQ34/Fm/Ib/BbPqMLs999JrvAGCpxuQQzKc/ol8auMFMTYhzXWUY2FI8XCCI
jfL5jpwGngjUTVTD8n71PIVxDegokqa+eBTRiWZVbW4q1DU9aot/4/BpnT6U2AjI
IyH2Te1qrNoX2Y3hgEaipC7IidkwgL/0FKoxZRe5VYc=
`pragma protect end_protected
