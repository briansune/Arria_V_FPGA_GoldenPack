// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:21:15 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OJRXee5aXd6PN8ilTnuAo7jHsOrp3Py4RkrLJ4QITq6SmUAPn5ORzLMGswXice8B
zHirXKZqwNWKTqXAgeKYx+tr6rAatoIdc/YYYFUM9y5SXj0qgosCw2PWdR/F4b2Y
utRT93bedcjEg68g3UrJFeSM2YsbMm+Y6VVl+c86f5I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16496)
pr9gRW/etJFrfmPug5AyOlgRR38lhnbqEasfixzsmoKwdCsnMA+2tPKz1RVkIrp8
H6naC+FVDURpaevzp2GpVQOPvzotjDKiOGQVxOnXbMLMMOBppcK5mghLBVkv390a
46kkPzUvsASeJA5FLig/ZPp/onSfK6TdMqA0tjTYWOygfJo4rlFhOrKuP2yMLlr3
RpubFn1mCq/8ufpxK29JkS2DmpXuvoEjrvZhp7Rx2XrY1DtygkJFB0r9G44cdVPy
8V1fp3AnqaGIsRpNtgFNi/ToHspLk2FKP7eW1gH2+ARk0D0DBwYjzNQX/zhnniZF
AxxUBE6UeZVV+ZcdWpwEfGHS1kLDeTkX4P/cGVUxKfwE3HCwq55QHwuD6eTlLcsV
guKvuynWkM3LjAfdrX5fsK3lz2vZ8wfI1k7lxcelZlYJN45Vi3MSBQS0Yy7LIP8c
MNRpM3KEL0UW7GyEApwWRxzMY5cQVyFGrPpfzkH2dNsOT+CXkJm+IDS796skPG8D
84maSE80TOluGHwYriDgO4FOPwOf/BzAqPOdkMM7J4cByBMBcdt+67/0jkVvEKUv
ygbtE/A+yJljHmeIHQ7srAI+ZdekdFdiLebqJJwS4F6WHx0C4LlVoB/eJlxfh+d4
OM0w4PrRKbrhYQsejvhFiMEFv4XThyEs2tcssdPcY+Cw/OYzH5yLjlSCWfzR9ORV
Kpj6mYUcSTtYKd1S7k3BeoYxSGdRUg4rv+JPAGhVsrKUhDffBX/uuBBJkybQOGuZ
ncb1v65TFfaqgjGhj/4D4EbkdASzsxUpBWwzpI2qZK18Gzje6X1vGVl/l1YUgPaO
Na4yPXkCRfYKypnJHedXP6IAP9JOkt1kGjzlw/86NNwJ2KRDCpxRPnAZ7CfZoFg3
MnIRRz5QujQkq6E2hGYtavS4JfsrwSKlpGkDphPkG9c87/8oppysZp61mBXUx8wD
1qX/s8rp6q5dHT+1R9O4TxH3IMIFG4Z/3bqUbJPPP4li64YjpwRl9Wvma9GTmo3A
YlOP1DmQH4s+oqvHVPSoAKm6ZXB137vb+LQ7QJvrEGHc4RF0yvLWJSWhTllxa1W0
SVhUqz4JDwVgUF8UIIKGI0OQ0mHZk+X9Pc05bRXHaNEkOVDJ55jWAYtVkFPL0Jqw
rK7qLYnF19ETv17crH9lsvoGw1ZuNHxUfo2gO8nM7fhbxjyMGK31jss7/IPkHq1N
SjQEyMXYopOT6f+758uTSRa7pMEPpumTsFPmz+tJ+EZ6LuBBBEe6Jng0+xbY/cEJ
FG42k7Q1EnCcCVZ1sEqvlN0t6Oqe9X1cgCr60S2cGhGKq8P/NbQryOKHeN9SeKva
l2m6VKzZpjJRp4jU8FavLOMeEhQW1lon/iDzsFnP1JPrkCoRCk68RGyLJrRiebz7
dl63aem0w9V9EXvhwmo/6p5KAwMqKy7gA4Oex+O9njQwiGTyGyfkV7bGTlL0WqtZ
bsfPfb26vrL/bwnu9KFNGpfBbWhKlgaeVBe4arQKri92tjaB6EmsmgtbhmOC+T+b
H6S0AnBPRx18i0Gf/mVlxRhJkiauc/nUjbq/XIoN5czPzuCjQyFNqYLz3l8q62vS
TKVJn/GPyl1AOKjfyJrET24hghZq0SscGppSKXQto8hclxDWpQ5FUNHG+oceJokT
KQp4BQ8PNi+uLdVmA6STQTSuKt2ghR0NfU/D3cNAg+dv1thfVqh0kc2CzKalTyzl
G5EGtGon+WXaE8oken9pmFwYxIKNkIZxiFUZqaICM8CLpbQekhK7o1/bXl+smmVf
CwCHM6uSSp+nxT7AyN0j7Q0Mm5jOiqJeT7THjiO2ClyWdrXhUz5qXiSo8jntsXnS
awMEE0cTupV33KpKAnmCtzoQpoSStTqa08j5x3cEqsAwo5/iQy+GKNoLMd2dFzd5
uGx9XPIL3Kc86Os9Du0Bp87L/Hle7Zb5y5VIFN0MUGWWQ4CWJOhErSxTSuECk8gO
6E9p1AKhJ1W8nJqnHX1EnP6HXOgOqhmCtijpNH8jHYb3UfOPwD4OxXLu3r1J4+Bs
KLhyS32FNyKgERFX3DgOxA1euhorjkPAblqu5ZW7ywGqAOCzp6VyTG64rxwjd/g3
tXaNLEN/aooAMTwHkgVagLHzMWyQ3ZOvkRCCPUWPdDLmLzYosBVaIDTdPxnYkXNA
pNuhKiaoaitGzp/2LJ09Kqk3Is/smiho3CM8ss4A84M0cmuB1dgwzRauhoCX77LG
cGQZdJqHvAANXxPZW+xWghLtaHoNZilXXvIHzcCaT1QuVHKsfguI+vZLNwrfwz8I
b8DHc64EwukHl20bj58Kvsr51sXbfM870mFvaCoq7svH/mLQ0DzyKaMcjzUsOPmJ
HHfwNxIBFpnii80g2eJY433OdbvmtEk+j12QMp1ifQLKFizxg6unfm0wNJZ3kOSo
PQYAxDnyZK6I5pAl1sljjIKR1I72GVaDZVs9+fyQ128/4mAoDR6kYSBVNlwQTBd9
9GxxVH6/fU1U8eQ2N8E/GxGkguQ6AIHcpfZ4y6uMlu0NQyBnKza54YA76akRN014
aNC2zIwXFkk58hCQET0Tf9+3EZNOOD9OnvSINNkOCMvn16F1IvYHLd76xkE4dsf/
Op9Q3bbyhstyt0jIPMGYkYYG7fMnSohyQ/z+jh06B0x2VR/HOaJx7w2AGWsRSGyG
vIz8Z7VzFwrutmGwrm0d8dhrKhZgm2PpcVNiyEC+M4kopjriSHvP7UZuszUjva47
ik+Ky+KcMWx3VDOFLNZq3/AQV1E5JvaAyAU9QTjMsJx6WEIbaX1VqlLU8Lcvc7e7
R1rGZXNVXKaIlKeGfvxcd3aUbclZTxrafBFddL9bjaxGCssPs9xwH8MmzbBJkTZt
TNYjbS12RXO2SjwBOAtnI71XeYMEQ4W2u3f9XnTq+VfS5i7ira8JZGr6gpiB91eg
47XgpgXfJIgdFnXHGfvf6vNhRVv1FkuPFRtvUINPv+KLS+iigCdhT1Xv38JqvFiS
1TG+jHFW9kqfy4mDcfsr8/VgN3+BSeqst7Q0iGA3u/VSAfaghrhAaXaFpwqUPocw
PfwmPaijssytu2v/C1px/PNNAdGYL3+giHnsELtNdKRmL3GFiNanL0W0E9Ii30+T
42d9BJVsN9PXCSZ9MYbBu9WW4qWEPVMzTFIJ3Ep+E8w9khZkoNDajrWjN5Y1G4bj
9NJQC5DIigphco9typFPLSI7kkHRTswHJh/yDwq81TGEXClclY+BcBPDaMmZUNmY
i368qKSYjS++mOEmL6Vl0exbInzR3VybQE3/tYDz8nRO+B1HHzevZ/8LAz7l+bTA
jSQ+SYtMajBM8CYXqcaI9vsgC7zgmuSowW5F6Vl7mZq24FdZF6xNTumik0s6Wb+F
RxgJBCWhAJyJ4RANKhiNjnQHoYRvr8Tj7MwJ+UrxfZLtP1RppK4p2hnxwMCXV1By
nTuDFYx9EyytXysWPjdbg8c5xyYlHe2gz6mT17iE/iXUCcG/JrQYJI2sRKCeU1bR
l9WY3uQRqFHSw0momffTo4EzFLyCMwsyxWESGhRhEqc3IXAe5BzUubwBHpr7pA+c
tvb3rt4yBJsMrHHCFnpNUKsi+/2EDOtMREJJJ/NqT9Twpiy/plQnrf3MO5p1LSj/
NTV+i23BypZr/22eJ3pMlAt3EHDWphr8izTd6g7kLLxKkUFPzU46zk/uQ4AGJzOc
EVjJy8iOYfoZvS9A5ueZIZ3+hwsjDYTHN2f2/V3bJ2MQHNu3bSWLKqSuI2mdj+tc
gwLk2t2ReDKsl4ljuy71FRcFkJsjvy8KthX94HQOBC2L5Jq5uWKoUGnxMaxvJTmf
xpcSS5JsvDNzGLCPvHma06Aqe+gkYHEMdAKuWHHjXTMmhcB9LnXfJmUzllMlDAFv
uSoVbwwTi7L1OqocEG2W3fUTx3teGJk4eeaBiOOnEQ+AOCcaEblfk9rZvOmZK14S
vno4E9USLTLzO8xFDD1KmPy4MJWjaWa4WmYA4zUDbd3Q745Jx78eKghevzVVasTS
i6p2tCZlrzOykRcOH/vO+9Ux4ED/PRfaN45ql9RV1KPulCP2k0QDdIH9txJvzFVy
DyeDtrJIi35nSOg8nf7w8Qy12fBvCWWeb1Hxtdl6xRsEYjPAw83mGn17qovL2w44
jQM6KNNVQctAExMmKtEDtW0h0sX2mWzi72pMm4TBpUwxO+9tLUxr6ymWSM30xFAc
wHfFhW6e2i9+3X3GbGJn3j2naQ1y1L+mse0IB/VpspmuiEni0WAKtaxwes6NjAl9
MUCJsc/RIQk8G7m/aKyN9195cEy3rSTGb3Esmgn7XwPt99BZWNwcQZX1/svHcD6+
9XfKycJeegNZUp0edW7mVBVRX+ZA1WGtUqQnzXDyGhvZ06GNYrNreKQtcebJwRX0
j52DqddmQ8ZvRc9qhCk8MgzIMkoEjBFySeOud/U/n1GTuXbqOqYFqL0jufXCsUXO
PG18GBSjZmvdhdhfaeqteUVrS/PstlCUcODch3gZWfE9x2Fne4aXFXpGv5aZLzPm
tei2LEsb8PoW3jiQP38dhdc8EyozRXSkpSLXSG4HFXsYYDiR7Tne8QfblPi50ays
L/w24ZWc+2eooZtuI5HCI8Q1t21vA9L1KAfLwBMTVvpQ0cNLD2lbKAnhhZzaEdr8
b7icK480x75choZKjr0JxLviDOLFqc+Gz7D3r1Tld+aEjaSw+vYq4N67IuzTe5GV
Lhsg98SkARncS+vMetfltAXsMwKcv0TTMFWB4+N4iQr83h2QOLZ0/KrVBCheVZGY
qafEu/wnNc7uEyPf43vETtHdXRyCOmo0Bu5DcciM6NhoPA+voUDy16tHMQFAxKYr
AAPYOX3UQI7zgJUOLyHx6nq8AqHXNw3rUFFZktbjuws9xCl9O+EH4Cb/loo085BI
YkYbgLp7gkRbvNCxlBSthQu85I/IloQtKPFTpZJvth1HTTAgu4BcvgMogHqi9AiV
2AYfe2bUZRDNqRBXwhNSKvDJIcH+Z5t397f7NzJkoHlLHH3PEsuXS+zzBYzqVK16
+1A8tcv1b70cuOZPu5w61bQFO/cFpM0kaBV9nKSlB2l3MH1N2yZU5E1dzvHGbFOd
IcGeCafqTheH5OHtDppjEeO+TicI6PuaV+bhrH7Z9OrZvnZNdgxhdpXis7qtU5V+
Y86KY8HpVp1rUhoZSxAeQ8Cma1/O84P98hpXxrjv2tMw3Osb4vyB7iz8i9W7WGnE
i1ZInm5WSqCgrFZRI9KcLQENIcTVctXCP5iTktYa3GX0q3CZBDeeUbCStmWyzbFs
CXd+N87Yg9y+inIeV0EsiIpUQTFNgGyofVuWnSpk7Nzr42kWB2doicaBbUAvx1j2
wVMbsEC2HfH6Kr1/RkHAkP4FbdhOAkYoxqgpPgPABinemNp7Lnyqdlb6y0IHylvo
vwP1EtLMJRM/BWFnQOfC4Kooi0NuU0VX0KmBA4oxhX//1KTeS7PZhh2ROpLwXZzX
/2iTC3iso4UbFZO25Y/WWwn643BYuuLHzIfXdq0Lv6fHsWNSkDMyfA8GMkm8ml1k
2hdENi//p3kTjYvSpA9k994HK9bOxbdDQ7vrtJ7ChD4mtU1zW7c+00Ho6xYtNW5W
dg2oDIruiAhlalSZMK2wWUQrZe1K7pb2tVbosjvqKZogpO69B25tvN48MWR2pixV
v2FsY86RyuApOoBDFNwKy5peu9fG32zGBMmb2zo4kq53QIO+Noehi8K2UG/5Et4P
gOnRqDQ0tNhdn0dx7YBAYz+9zyFrLMY0AZB941UqHncrrmdWNit8vlZwnGau36AO
IqXj/k+YqfmPmx6PK6nCACa39UDFuEAuljKWv5yjmBm1Zdbf596vVLtYtEDXOcSu
DTIGMcC8mlae+NRmOEltQ8hvDg8OOpoZ0V4Ty24Xr51zGjxwkyerfAP5s+epqaHM
ZQoVZplzpOyh71viBc2i1kHBfYu/52e6x8xDNimfdBiODiv+zTxKEsOe6wJZcMe3
+JK/TqqDtgSb1DnVzmrM+lHw6Nes2fDVYkN1cyTOUfBGD5bS2EbR2YXph6lexYFm
WgR1QuypR2h6JFcOT/nPGcAIqtNDQZePox8vX3lUlz+MP38Y+tkgwWGQcK9QuITo
uTmlN2FtFzDqLgb118Jeq+kjOZxzCvcVYMDdNT887fY8QjgGjiumNBx5148gswDe
dYhusVtsVB9uDpzU/abJyez4q26BEi5Uuk/qblcgbX/Ay+xNP2JbX6HwyiwaF3z7
RE3nmQabZ+1oaXxZOG1Kbvafb4uWl+A/E4rnG9Fd0jaK1irqRJGoLmiAjicxK0ly
TJ+6jDRFAu8H5gdng0D9NAYTEFTyKn1XiKcmJsDA1HsF/Ro/addVGmGJxEh+ECzf
Fyw0zMx+51XtzDzJ+56lZwgthKXd3K9Xjoy73u3js6eXMp3sU+GwFCMQcAcxSL/G
YQ5LHRcHLkNPA1WNtuvOJjdqucVK4fUPJBXcTHApOrXzeKbivEoHZxX88yEZROIO
H1LPvisXJSjg3KHpEB9QOG5w9EW6yaAteaUjSaUrUU/m1Q7SeSpEvq4BPx41iQvz
E76ymY7l3t4XAraCWviqrq/g0n7IEVmCHpb3OBnpjuDrCbNx9YV8yAzSMRBppfOS
Bl5Sc15/N7lxQfO2zJbeDE3RNryw6Yn4CPX6DeM1cmK3gqEAgP+AmSjh9IATb6/r
SDzKgZt9Ggpc4yqFuPgGk85LttN9sDMmIwAKzspQQcj5h50i9kA77Oiz2THc64wh
xy5e+SHyyZ8wC6yAI3cSnJPQQKPdgmUmT3yFWRLHWGNF46wdQnlKKSTJU4YkJFo0
wg9bV9AKtKPIpV7eACQ9UTTiLEwFFJ7Bb/KFcQLyhbZR5j8O4azDL/enXfLGQJ85
OkxbUA7ymYohqdeyZXJJioYi1fNqQ/vqM0HhWpRd1mkub6ANJpnqkBSZPjc9UugZ
WNW7MDFew5Os34T5hxdKyI22Xt1qSxQz4WNzDG0Cq+NieNX0l3ickDvsadL0a4Vd
TozCI4ZUhY9wk9lcwJ+rq6+Q0FsP/+L4eqfGrICB9eJEHv7QLEj1U+XOhJoSXt0q
ZaleOGgZyLAjeEPDMipS+TJ4rogXcbI1Q3FRfiw7D8ZAiypTeHyOkSLc1CehkQYq
s3KMiUmyVFriKLYX66tDs+pERCTW7vlQGPV63bng2j4CyrRHfJ/M1fZ/QLXn0WaP
9zLm3uO2pa6BJlzU4hhnZYxkHTejUekeaqCykd6hqzL3TPm6DJAHEz73P1X/Y1qV
KjeBouqpZ0wxdTqTNJk9bkA8dGy1imz4gYpo+ic+cIZOnS6k20lWvMX7U2O6+dTg
wrmT7+vQIRPHqbRdS1nzKdP67SryVSyhQ5bRw0Rxydkh8EGpz1qpfnV7rpEtxcmO
+zC48c4SAnzzy6KxNTJvJUrM49qIGEY3pDPs5T0+OMMLPWpED8+KFfnbfCQaX0Cp
utUVEfZZGp9GGpZQlgRM0cEL2kAk44QG8MIM3WlQYSNfpd0vXbd0hzqkKVj46ER9
oW6qk4rmJW4akyKtt+SbgjN/Uopo0qk4itLyqBrYV7OLWh5uSvAOoJJebeOQmCuX
dJ1qERIjTuKUUj2DQzb3QFnOLpVD0hDaLoYKsk1ClBcXpxyPCVcOvIMzG+wxjjuG
N3aF2uJ4JRfUNMZAnNmo5pwHIyPKXtBDupmIY0k6V5ODZ4eMAXIpk8TBVD1Zyyo2
SX+KIIBZCqwER01VWWdy3znYyu9h8/FTAYYS5mlum79UA5WpKPSTPYXK0SUau141
g2cMoDlHotle3iG441TvcwwUrSm7BFtwqV+G7I3fUPhu6rJLx2O1mScpuW2+FFjl
P7iAtT/oof5yU5Q4aGrKODO3fpU2oZ8EPJ2TmFLEYDMS6HPFAJSCKiRiD6Bxl6NQ
85AiVWKvCm666tW0XYKi8Cy87gMdE4Z3ctaaBOwbjLZvs54PsYducIjg/C7IQyHG
kn7xYYkICme/vhzPgMZxgnVNvzqPBFpHTIKxLIML2q4yPfHifp8KlSL6hoXLuQ2f
Izms3TPJieFqIKFVSoYr9fxeGTK94vUpcD8phfHUmgeGJH7rBNCsVDbxXe6XVSza
Q+VnDreuty6E+HtWCu5IjSCT2OKH0ImGxSBCCnDM526wpkyPrsinPgO+i1G5sjXI
wyysD1cVrkkYxuvku0p7RrAV2GgmkWJIM/JLNLhIxIMGpFnofktjUNWhbyuNsQXN
peeBWVQzBSrCLMcwu7S1fhoGSjtqrA/ZUv7khM3+ApuL+jezyNhpuGXWPLnqci7i
U68CuDVvB8ZhzhHnwN4DvbyV2Wrd06XAu+mytsWpwh/K+whMOi84PozxiimALxeH
amhWkumAhOs7+O6E/Bp6Gn5TTT28/JlN0FSyKwIcQwjBL4duqfPEZ6MEobS/gmKD
g4nYmEGVqZk3Iu/WFiffyjEIVoIRPoU15eTRY8gKQi//nLCS3WMmy2YYccSkTJ+Z
Cr3lFkbWIgYGki/7z3mplIED3qOvuJLXpAnZVaU5xqMzko5MOjTig2Nm+dS0lDAK
QJgHXSnDwAnVA4WFHRp1Xh7hOvDNyzzEq+cYMw35N9m64524AZubHf7JTMV7r+vr
srFeR/gofDdBgPAvG2SX5aKKhkQpuygI7hnYrF4PMgbftbmjwEo5lrQonzB1Rr/X
iM0X5pii1xNJzJ7OOnrDQ9ZY6kdjHd/SSFepF7xGjjwVhGmrccXgTFZDJ1Q3skPc
HNAKfW+GltPXLcwk4FeXEaCzJz8eCnkPlRWuH5Ock/UnJBqqNHzhQYfRC4VF04u5
seQta7MrlrXMmrUhaDy4SDRZHHOaZa5oRwSvJ9c9FrklP2gedB+L1bezUAEYihcr
grdCuNumeNg7FF7I5PtL6EUq6OscacXoPQkK5zxF95GWHQBAUHP9PwpTWZE9U+DM
AZvo4faAViLGXo8BFs6jvhd0bIUsTVWml9+Bibkd+Qj3p7CC2ydkuvq1xkt+Ri6M
yL5oeg9rXiKz/xFr3P/i/A8awbicA14a0W+YkTqkRi/yoC9ZMnHGPQpsjMCRhfq+
gvppkuvLktA8KwYJsykVdBqaKO6JEWyg8aUhDUir8OTX0xMY5CKqfnQKZuWVKUX3
jFLYryv6J+65mdEsuSXwt7U7ljDNeEbYibMNevJMnC/Lisx/bjVOhPB+Ial2DOE4
qQ9rTsite1FPCAjzZMwCE5V4m9/X2YOeYq8g/yOJOS+NmJZ8HubAVRLLigGqlJSU
GBd4pfJDWFxibbPk3Zqh3dyAKYXTgaHWKVqDXbhNxC5dqw4i2K9epumt0z19r4FS
Fnz2wcMc7hl6/70t0jaK1A53IaxNj/aUFKTGP/4+DIlsRgGgynYeXcbmfnOfcki5
uA47VuxpvwurI6vz1qeLoUUolBK54Zry+1NYRfcbnLH9/vBy3tFtcpjyXYoVb3Zq
aU1ueQP6ClSDHvJf6h+vsBAH173WLhVZDz8dSIgCSdLbna/1oAcG9FX0eNgt1VO3
LJQT/UOgUJN4rYBff0CI1TyYKhQNB0qqdeG951xKa/33GUz+J9Ach9eB5herakau
Er0ORpBcubFMWqP/Snd4RbRoEL9BfBufv5OEDd5HIydGH1obOOOUO77iSsbUpLp3
4W8NMcDaJL9F5aipKNpfEXYYOfuHiyrNzKWDOtNH+Ld283Aw5O7v93tBRUCWvnCh
as0OIQI4+sm3sMhRzVoK+D0gm8vBpra0mh/wIb+E6Neoz5vMRCgbrWNi93naaUVh
YE/IhJX6Ory1GFTm9LG79LInD3z21EfW7KsE9DMzbGzTW7i0BBPsU2tL+SwYPzPS
bhSwN+lD3ri3yR8l+vyB65gaWYhOrAUSkbeb15ktf2689KGjMxTR3l/jst8w7PRJ
Swqr96jQl3K20toM0GfogGgSyuqMPexX4TvQ4qNwbSiAEtym7lC8uGks4hiLU7qd
THItw9wPjYSQpgq9d12jCB4/Wzjr1vUszNFpHUx0swx7OW1kS3tda1uWK+0iz1Gh
C/8qYKmVRmF7UBACrWcOFqEbMrc3KUmVEdnTPeHsqsr/CIYyutB5wOCt3oRYKwfr
9WAJfIsiyrCEfC6WUgvp5qV+Mo50LL94OWVWufQx5BGYW01roZj/pfXO0w247Zuk
RTx1WpmYH1xABAKEk9MXUkssWH242ifYe717dtgJZyaRmayfCTjxNKa9kqzB92Gc
vMVgfkDU62bCg7h6RmjddqNmt8t2KZ4TzFu0mEZAvNSHiIyu/juSNV8+IInCP8w/
mhU0BkkuAnHfqmmp5Uo554up/YLTlygkT/Tfwrc6vCspxRYM0J4avCKePIGr2MMh
iqUITA+Boz29DzGU52GhlPpu8jpj3GRPBYHG0Bumd8Ol65dRYpqN3qA5PUXnxxp1
cku1+yIm1wLlPY44DQgQNoZ6L8vQHmaXij+cxId+yJsH0hp6lHGglfvK/lFJ3txA
7qpsF1WNwQ/7DJf7F5hLoGu4GKLkuYOGqA2Z5U/S8vMclGwX5MZHofkFaKY2dz38
EKaj2Wm+yD82Z9KzWN/0xnuNAzkCKdye23F7flLHex8vjYHWXQx0/WNKYm84O2S4
0kq3Z+5glt/JW0tTl5OOuRDcKtc3rLvg6MEXZNfQMwgvS1HfzOilUYLvmupNQ4Xw
0VGuMYuuC6x0lVhvnJt000j2Eulqek7nF1e5kiCfinHYeOqnV5sgl8V0zvZz5T6h
WzIXOYmWZBGrLt2voXVPCFxp+sG1TVb6Ba7a3xdEgkizwdP3lNj8J35h4gK6BwlF
kaqDUz9eN7zvklU/w14jKd2+aNLhVZklp9oWNNtBcGd/wpC5e66dK4CFzdIDSOwt
SnF3+esRURh3jYgh6ubPWJcnrNwkNEQDhS2I4eu56qTDFRGavzcKPnkDbanV+I30
Uafr+KvtIrTIMs46DBLhZPcOCbFb+ADhYkoMhrlJhNG3+6UKRRWu8gQfVJI01utj
BJ1Puch4CnhiMgQM0GFAoDzArLADv+xg96Np8TTFv3iNAQeP1v9Ya80H4tFEXn+d
7zvzRViuRjLJu72OPmCCg6uH1YPDSblbuiGoO+XUpPXBpAmTd5kXi6+Y78LfG+dJ
itDms70ZBrCDz8KTLgTSKToEWnHIMSvTTPsB/tZJtu01Ii2RFBqrX7AOz+Vs8aPb
VHXo/41ZktIQzP1XLTHvilE4lq31V6terGbBdSiabDh+RU+GCEJ9ZaRlibkR+oRb
Zeik3daaXLV/lOcwpJHI2omkdTbfKdrc6R5EjpxY9YbTn9h1sTPMi25kpHp/FXRg
Ah4JJGQ9GYXWZRb6wGpJP0NWKddS3nG5bW+iw2S/NQrF8fnRhVD0teembmrsZ6Ot
Z/VdUIBzATWKOJfO4w235wYtHrO9BMh4KV5rZQdZtUFVruPpw6gZrgeIR0HA3PjS
aJ5YsZRF7gMzFc6TMCc/QVFcAyW1gBrZCyYOdOC0vjpX1UqJU7KD6Q+sbrT+ACV5
UTVao6daW1w7MTkBf6wmflafH9Emlll2NjfkLdKE3+/rKGXu0aH7bq5Jmzn+IvhV
pRIOm3ZlT7L1uakFsCdKlZCW4oOpuChUvaRSLHvuA0OTqXadv9iFl6PT0/HboBwU
xhnkRI2i9m+SzGJFCGbxWPygh6jOKnXdNFU/xaHe3M9z9V4NDqgC+884o5ovkZaS
XDU4UmLUAdWPxu7CffD4xR+HqA69ZeCuvxP3FK5IzvWjE1wZjgFrC4RRMM55y67B
sYV+bVK0yISIoLFlx7l5wFN7FWtZtcqzkdYc498hlfL8xdarnsCdV0Oa1VHCmuJK
c4pGEMRjS5fWyn0SQPyvZ3NVFZgyrxAps0PZv27CveuuKsd59KO+s40Oj0XVyEj4
OB1db9X+x7OW9OJ5Mo79hNgmUkgGyKPfdO8bP1F6AU6MfkQ/tOZdrg/gKnXuUNe0
gY/GpUr4FkpxXSqf2JX3N0Dc1KYyMJShxTQSkDO6HvE2Wo5AvGPFAFI5coBcfOhe
eqtFC24uo1mAMHGDze3O0yr3stc66F0BnCDTZ54as1CkaRnaFTgNI4E8fsSxLCcV
BBO4EGCVLY43Q/+0KXGVWpDNi2ExPjfMYcuDFVvUneNp6H6slKGPyNFIoIrtkc4C
dKLA3Kh9MIdzuMBo033e99N9UgrX6PPqxk3eNq8RnBk/KGm9FewaKCmHD0ozY/m2
u6nSXKISaNngGmN1gv0zN+aw4ddYzSP8ezIxLVLcUlHf84i1dhszZbEHwEcjJDU3
MiSXTPRwPt+s+Om/2BYKTx4fw/iqKwukMO991hBHUbD3daCDH4X5NRrihg503Bk0
e0Lz1TSxaxXPVou6jAGblbMyU9h+Tn2tGQGr3RwxjDkwN/qppugMz5Ew0ZqWXUW5
qFQqicBonESSTbvdKIVT6IdgAicwwnDMJn2fBBHLutY316lJQojkKwm/C4/ZOEbL
/PPpwKBsWb4BFksi0jgpsDe9cRDKte7RtKIEKyhTLt0p1++1Nd8Xo1XtHBoR94B3
e5svK9XMnQKPp4rmaZT02+j5wFmxVFk1TINA2ky9xa28FXMD9Dkfkf/m5pmsWSvg
H3yT2jZkl1IYmIxWdFWWCgNmTXr4RX/Nv6iPEFzCxJHSlQdS410pTTkajNZ5UdZH
CtYfhmQMpUN08s4NxPcVhD3H5H13JVSt58aeFWML23T6IA+IWwE4QAnGE19Wo4h/
EUt3MX7qMMND5v3jsMMlbgToMGvjCP1fVvI6qjEn9tLUKMswFRCpwsUQbD+mG0CS
3nJNfxqaj5XF4TaaJWvxM1vu0b1hDqku0k8kzy79BteIVDc2diAt73GLONtbFBzn
j2lMiMrW0agGO/E1GUHQOjTDiJom94PMd8PYYL0ZYCkYMTUF5X6xM69HNcuksYAP
NIiZQUkmmtncT6Gern5bLC4u2m8/LaCfD+MocnZoTdLg2cwSUL0omEhUCBnsOLfe
ZloHNiQ64xes9SrzdsTrF9WC/f4CRlwCdHH+gscSf0aMXvma4iFEJuxOnY2pps7g
j9BwHDGWaaSt1t8uupSlpY86IlsiYyb/CJsNQ7lb92fFSfg8oE8yOUAcm4A/07Nb
3hLBJU8yTq+yHyASarIFHTMMgS51QmTaNgEqL5wn/9hKO2dfPK4mQA9M1MSYoNUk
KUZ8fyk5Pnu05RgyOxRdkUbk7MT299RxRm3BYUDYaTyPsW1ySiHqmqcICr38gGEX
Mw2Kp4/6Az4nA2GOBkYTfZBefxLpugJ04PMF/rAYRjzUKTY8ExueYi0QxYub2UIE
44NeianSkQxMLJX0lhhKK9tgfyLJPSh93+cPtVG7nSVggLgBHruYQN4RvdmHB/nw
QH2m22lJ2ECUUpowtNyrmPPXqjbwkylii2QlyXI85xBiYkLjDLOElPV+zt7GhwLi
xy4t0ktymvYguNx3R9TThWwR22TpyZ6v9/f1MJwdA3ola2GefVH73JrlOtDd/uj7
yGAWF4j287X5omudFf6jnMgHWoGwYNUIS51d/hmDB9laT+pbCKfKHfVRKy1PNGgN
uEButiET5lugfbo3SMHWUHqegZ2Wa6wh8BpamGm0k4XYQ+wmnA86kVtdjsqlc1TX
cdCGNS5cI/9wfteN2zg4Lo1jZ4hNDjgGesLh4cDwtir4B6hFI3gQ/8OsYkiO1XBQ
qMerJ0AiE/yenJOI0AR/64mixk1cijqQzPTIPS1iOHRYc8AlRqiPg6Tgt7kJ2Mjx
nIdmFij0C2Xh+bi5qEssiZaY4Hjs9AUkEvgfZkwwKEpcgDoJmckTCH6h/SuD1y/H
UDAKfoeKlVrRXxylMqjiRMEdiBDzY3doZPDxwiqAN5T+zHgxNdjgFR09PH0A11bK
MNM5hh2eO5qBxxLvHwRAg8hUhNgoMeEMtXJwYdpejGKu4jvho+gfvxyZvZzstLly
5L0ptn0KoDwg6I8Z5vCqkBUO70dxvZt0x5o4CQMEJJ9nVYHaqSwb6ACxbdFuA/0m
8InmkVL1yZ3xyYHLNH0NZUOZieHooDMLi1BnoFalCL+w3Od6lxh1YmE3Ju9YcB/z
i7Cqo9ntM31fzq7SmMaHcWTMWWIvDSkxt1/RUJ/V96ciGtkgp/Aj8H7cfAC7AOgu
nXdlnz1p+/TcDVJQPeCU2bk3O7pP7yo0TgT/g8W7CX8q8YRqz9CBHYPn0KV9xhYf
DzgTC/sz7bp3ZfMDV0TOkgEmwMU8MPUYkUbgSQrd3q+aj13ouiUbclEFVRfQS2Hk
wepU0g2s5tuLRlqUotOgqmdD9b5guSScO+jLJ/32mBwKjcZzwpZrk3JdGbFxwKW+
CpwJ2gxLk3nRm6g6FqoY6LlLbvU0hA61FXksaullwR1EA4WBwrwvRqwV4XkMiIon
YbZYw+1oAi5jCQu/ZLkBD32lUoqcyqmB0Llh/MRqhPbEnoPSPN530VBptrvIjeen
IG1eCHWScnYiro4pl8muflpEULvfWz/7Be2Wg5YUlJliB9c68hzam8zg41iX041F
383Ez76PCR2cX7OMMxlW6GriAuCjJN4EyUlju92zS9eZxj92wQZEQokSfTzsGAzh
SttXid3rlXRaLn3bbSeB/dNMIf7MXLXaAPrJ6gp3E3x9Ew2nsPzKC90hqRXYEzKf
loP553Wu7RDEs7j+O6I/HzyU/F2UWw4sz2jdj8zfZpCtniwnJy3k7jeLdn4w1ZbJ
C8pomHfjHRVaNV6olJYABHgm5iLvdp3h0l1YUBy5fDRTfi8dE3F/zySfq6qdbIEX
d5L7X1A/ZYW+v+s3eAqxpCWOqRJrt+4RICawQQQxclrsv+HDV4eL7TeJUeVL1/BD
maLNVNFQA8/j9uPY1xPCpHXzG9rXz8dJtzibjC8hf8wsZW/aNb3DwbKElkLBXz9R
Uuk9x06byFLiNHelInD/o+sXFPX6edePzDVDueRgWQl//QYlBRVuSesySlzPT080
FDJ/59jyitU3+1ZulA1m674EP/AT8GxODwd/zc5U1tl6MfVASMUVxQcFNRbG/Th/
gZAWWWpUIe2giff7Vo4UL9Iu6OgzP8puP5NkgrD4copywMQvCO36Jvb201np36bt
5VXBnYl7SO5ce9lXDj9f+E3Cj9OYYhKSZ+YjK8mJyV8ZCsKVJcx58v9J45IeyiEA
sHL9UPQn7vzeTPJnEDuGbRpRtT1t3DKqDLsJCGbBIBxB1EIZGiuUcl4MOK3eFML1
FuJIy8rOTM8xGJz/KsTxJZkbKYV6L5XCZu8P3DGNROmYzwHzi+Fc2XW/w5rc8JkO
0vBKWqHZpos8cOJdFYBBPndg/LIyDbEvfZzw82mDUSK47ZYOAoLrmLpQYX3TGT3a
j1i+rTPNZIhv2RyttzJBe/MYs7ZdDW0ryfeHGtQG1oAc1dUeOg9vjBnOSZgH9LFV
UF8VsXQhVLPtY/PErl6FSNzBPJUGtZhl8nG1RTSLiYYKwrba/3uPdXWapVOgIx+E
aJu+vd10qRcCUJqvabZVuVldw5C2gMQRVi9o1JMNmqYEezYvrjuZ8rnCdgtvqsR4
IbrGpub4nbJyMV7K+L2YHVWkfujhl8mID9FImiptDfKVufFrjPNmF1fYymgHHspG
v5uzlvl//+JwPRhW0dzzMfLDTVULUFD+hlaHOhmVJelzlvV8e7daQZwIC90t4oSs
sU2y7Krr064W7C68In+bBKiph54ULxrRSEXVqoRPMmkR9xRcha7lgShE/xPBLdTF
T0othaoDBQ4eAm8ExNhJeJq1YSzSyc3ja9gdr+q6U0lucfoy7SI9ERW+lHiH1xvB
g4IGMIKY6oaO4/A8h8qdf2j9S8XBdjBtVFFm7yi/VqRRIdG2CPlQ9qs8fsfHsjCR
AEHqLg1FKSGTPGMljWF13/W+8EEnMT2j7Cu5eIVnn7a/SQ7T22iDv62He+8FMXgo
GdDdRJix6vd0xj7/FfZHw3BTpfWsvqSWzwh7FaiR64VL05mzOqlqbT933F+K+1ej
VYfT7DhNnacTNwSp940hewPp9o3Q1Fkz17nEeruAtDgTJrz9JXrVt+dBO2RJeAUl
aMhgL7RX8UxeBtmnMZjnQ25MyhfTNlsQ/6dAn7n6ms/mNMof2S5qbLct3xxv3RsO
zQWoMPXZxv5aMykgzND9yxj4R8h5wbLBJB9ibJT30i0EO1rbHNqrZJc/OpNIk3Gh
aE/BhTiWcVLFeDJ2ealke4wsEQvfePQvUrd/MzIQVMsv6PBB+39HcPdF0qgZTDMZ
2yY1KpO6npvsl2nA3rXF4ntQEN4DFMCGMLMz0Q1oO/UeESIpxa6gn0WtwsNrIdC6
3aa2Nw8wl07vv5oCjKDoAE6Q57l/yLGFRBwf92UUOnflOQKO+d6s0Zhu3mZN0Bnc
4WOFoy5Csrus59eINytASXKpskno/usEayqhYTEsBgebs69G0E71JbDV6UoC7FKM
361wOxGEUo1NsoTogZuDFa4L4UvP1+bCO6teZ2i7Sa5BAkfn+390R/h31gFb9KU7
ZpFWQ1M0oKb39MqAQzo+rr9hnzCEcFgPNtAyvIArJIGFoQGQwWIqOMJV1uy+WqmI
Lz7koYVbI2r/2vVLFteSx31F/gk1xQ+wff1T9kTYuR6mFMeSsxu/Y31/TXqqTaCZ
pdAVefh74zylh49Srq/hFK52y4ChZb3pp2qTWA4N9c8o4cuHg9xHzHhXR5/cvyFz
xGLr0M2CVledB3V0+beYbuTung/JZBHKPZSYI8GXs/G+ILm4YN0wsTvJ+3EZRFqw
dtA4TAGM7mQ00ke3uFVYYzZV8295Rde3TYYoypXmX7YFdLm4HmuUhVhTJfDaHYb4
dq1kxD4rmG6qarBat1/4K/myw4t9KIeThAhZwuyDuv31Xsr3w3MKBVVznJeMezII
XaLfudlv82N/m83fPsZ5aS5Ky0qOsJo99DlDEj9eM3xoDKTl5JUgUKIzZTothWZd
iUgO3geTkhVKO2EM+JB5MKE6Qmva258cFkhuwHx9l89rXdVfTCV9HCjZNioEpkvS
TYDa01zC9RIZrws1rBczWd6oSd9rWDkwVoTZpqT2MeA1MHK3CXK9AZO/9BsRh+sb
YycGjnGrW9s4nc1bPtGQpZrIlUopPckncphzw1E/t59J9UGpiIxKTpmm/tTKuL3s
8Mtbb7H1D8BC3gFA2SQ7v4d0zPqwzXo60mjNahEfAEz/VDO82lt/QgREgavQKuIo
xZYsKmoFQ1WLCyMtDU/sj4x31W+ulcDcpy6PEZkXChFnQXEmFYm0/nZBngNfGJJV
wWVeRRiEMfVmUxw6cxDfAA8HfaScdDdMo/5D8Tj1vFkc5tVWUTxENs0lLvIL21zL
DmgdYdoAqHYasX5okVAzq369c2gC0MxpOcspHCkucR4Wz3OBYuRRvEjtXnTslpmd
u90viyD5tvOd2IiBjc/VK6Ey5IUDROExxPQxO20dPfC46AEhiheOudccinuDCSoP
L3ZxtH+niPbEVLlOnovr8l/mfYfX60vThJuSAZbPl48gfZUZdL/47A8xxrdQ5BGO
M1fLd7IuwkczCN/NJVRNr62lPqfP6grGiadpv0nl1e+QQtY3OgBwinsl0ko9Hxpc
u3kvOUnMnw7uMUKLUoWlXcGuTjrRPNq+Fk1xw4/MN1qr6s8H/mccyCB9ggtyKy8r
aUf3U7ncunv5jvTeMY0Zy8pSi6ipKXJ+x+/1/p6n6DUAFuDm+5bWnAl0N2jgRrWM
0CsuhGdCziEBD6GVKHHjbuVwBUQ70aL6MdU+aRlH66JzB8dRWtSetCWCmLpOadxM
JGMf/3XjhEJ4GVbcmDYqSP4957A3Q3ueXD44zCX2Skp0EITMJqLhR5mqfi3C/sYv
dCELPvZdm7i7hJx2tDlOMxup8cjfh20QtDA7s+c4iGsadrGse/5AP14pJAdCb/La
YISJ2zyp4aMK85aIhF5wFKqt+lI8IGjYZ2SOatbbZQ4Mac48MGzHOkRJfgXD2q85
XFGQ405U9dsmBgTzD385b7f3gmmdPRW8fE08VeoSn4hoePZY3QeqbuipMS13dwlc
NTpiZwzW4O0TpqG/thSdSbdE2Hl7KwLF5425gmEyVbCr5ms+g8bQcJnSiyJWl50T
uyB4Ld7vMPQEDtiVNNxMA7roPdvmlHD78n2Ttr89CqUD/Ak8wHQuf8kVEGjrqz5A
UvReNUHrvc1pXvSBs3iuo0ZRuDOpxcjY7LlxhiePCvIaGmGDeQ1RrTpRf6ZRzKM4
24ESO0GSDvr1TDss2XuzP3nmdhoen9LSfmajkxe49q64vHCK11uzrPhRWO80aIgO
3SU93wkvvudEzUV0K0Ey2AQz2DkcWuAL/98yRUhK97ro3VZIYU+vPwymKKBWshNJ
B8wYTOpklzkPudJzClfUzbYEIkERxjCK7mgH8YpjrIyBdvr0TELbHkmeeGExYuTz
QUglwvtEqzg/idpcHrCU/28YxUBvxFNxGR9djHsCYYzWDtSnw0SzTG0IOBtg1jSA
HuQUs27FhF6TfJURQ7TbjVCsKtLGYfwfxVarISMgA700pbXb6++1Ae1KU+5RV7ca
NIpHYl4j/GLinnNVWkrLrKHQDMNXzEO7JgqgQhLafV8zDYYP/y2282OE8QSPsVuS
1L6LWva25kQWldxIcO1SPl0U+RcUdx8tMqG8torxsb7T1bAiaEJ55VDOSSW3o7pa
lKb4t72Y/GyEKIorqEtqUXbiQPbINSJLmGXLs9qVPXNvLvAgJEV3J9WQm9CD0Fkg
06HDIF3gzBXcoVawhlNXP02rz33pWzaC7TuFq17QTSZseCFQm1TPiRq8yID7U/jL
99D93eqQVo+dK+X6rOIn8mBPsXwxKAr7Qva5Hjytl33C8IWil/CKa1/ALxvjLQei
P6fNv8EwV562OXouIIaJG5Wl8zcdjB2blU2X0HjUSX4+MYiuv9Pg7zlwGJxuYbuq
xvDeAvz5d7nm3mF/rU1sG2J/lbWTEpl9xGhYIS1BKqSBSgydgDeVX53/utwJb4cM
PXoFeOxyz2VeULNoO5lJ1eWdjVFxhRjgRkk/vSshoaeqnHnZm2uO+22rp8icwqQt
T3SLnb0vVePdtlNjSopdv8hkL59dOkJYGgDH3VikoZpf9LvCj97f53RbOZI/EbUA
IZctIXlxklRafURDemauUUrUIL5rOA5WRuMT8Idptya4ZNzp1q/MHQNAS2bNytkr
MxQfSegKOGn60p9ALJDraajskHkWv6AcvfRxCDSt51brm/p7bY0mHZLgRoN6kiCx
3OKi81ErFyQ5uNOuTqXEbMzBwxTkqlwgB0JiCz9bIuiiMHiad+1wEZnmuvTmN4f7
vuYk8vd0ScW8et8Y3qL9X54EXR9NVVvjNTMekzu9Uf9Ji61dUv/W1eaAtBBowMX5
2+H7/iuOwQPW5Ab5kOF0O3X4xmpXXEscWYO85ZKVq1qTd9i8ccsEG/j6oaDKWOlt
mn8j3/gBjmq3Nr6gcWKx9VSpXk90F+zT4yQ9pb8U5QtsJ3MQ00gR7puK2g0Crmv0
MpLfgbOSFK6XfTiMxqqarxBdoKxw5thAcRD8TwbEyygQdJHrJghtgGaEF7osDRup
2InhA3alazRuu1PR7a+l/vpeP6/FJt90RwCKukkeHqBn9541JOAKZ2e7Ig7vI8T3
K2PDUXdTAadfR/QE6ivAk5Z5K+32eKa3xCfKvpHM8jkfLa7xNbZWeHfGL3i1r9O2
xhM972xyI60OCvJOnUa20JlROqTsxC2DmDK8GkZXsGwEQU6Wv6IbtyYD+hvQ9qK/
gX4nKVwNoUMmfY9LHg8mqeZdHALA/Tu4CbipWdyrzXbB38N96mZnUs4sjpiJgcIE
m7fUDGO1qHObI9xP7iRxkkFRtpWwyEREKw7AK9T/08NIaJHhwsxB9ERHid3wNW+B
AZCYK83Yb3URMXv3Za2soYaP12Tvcss84sKEg2vcgH3QmhGUg0C7rmsYeLvmXGh/
VphK1xwwUXFz0HuTOax0mXSzlb+Y2MxOls9+PfZYf6FaN9C/TNECs69Ez8MqhOSV
jUPpVHiAziqqs78g/zJxK1JJmjBMNYej/0mQlwA3t7RCZBEwryr8rZaT861b/7H+
NF3E+916ybcLLfR8kXw9aXzkVYXAQYSz99LpE80bJX5MOY+trPaNhQkp5FQx67mf
V6LITPEsh1eif+bmp8K9XWl1yF/lHJNHvUwZ6DW28az5K09QYRBK5VjvuO7sT5q5
oCoiOq5sV4UPHIz0IbTLIjyG0iIchpPGs8rLToe15H/eXKC6dStvJjLEkUNf/9Xd
hvqa/bWwbfWpkO0Joe4SJcf+g/NYJp6ICc6fz/aYi981jMMpw4u7WOOFubWMUFhO
iaXW8ZxlH3dzK3lMOLzZMT1XGjoJZevlsTbQ0/8ooQB4E5GnKB8Z8SloOGlKoi7R
rtZ8z4thSu78aPOeeNrTHuZjSKBUMv7pDC4AWRfDD8iYuC8X62W+Z1hHnTjqs/rA
5mfZhIC/ANtISkOgapLAGw0i5GYsaWnLs+kvVutXtzz8339PYmCBUAYDPrZhPtxb
W7EPLl1jhnZu6M9rFZcS/IqKbjWB0snUiLTDjtoiZAFRTqM1ikGZneOLqgXn9EL1
gz0zYaSwWRz1ACFc+WNSS8LuJWXv1DB1kcX+0mQpTYBw+bjOV0icMEuaLUPxP4wr
km9GwgKZ/yvnGze/13DLOeIe7kvrPgk66UZ/eCfvAYWeS9poLGx6i+TGyjB1mA4J
hA5rkc1H6tsMJ7v7KLAwTV3DAYg7IWvm6gtWpKQprXELYAR4iwWpIhhXVrEge2zs
0wecvOi8gs3FjZHgLx8yyMpYem4bhDvnJZENMj1uRyxTbXNWjeMeKcnpPlVaJpiW
MXRSjxuu0pEyIMt5P4Ats3GViVKsa5Oo0svuEtgNBsdX1fph3JfShsIKMI2F4g3o
AY5MyAX/GxH5ulsOU1slZIWwNdu5UeqDFhcsKYtrc/578fbjguaADnVMd7OSBulx
thHhA9X/LpGd+AYsD52/cAxmJBO9qqsj6pzxw9wZoDl0LSQnx6v0Q/50GeCfWMK1
GzXyZ64gqdNtaxfSvbhkt5jOW1JggoPTk5f8IElSQFezPcFxfpHpRZoll3TVM8q8
hP7rHh5rHpLtq91h4MjPbwaBxUbLRv8Y2o3a32GHUd9YO07gCd01OAT22TBl7vM3
Rs/NxAsdbBCo/H1w3HoIEOL7owoZz6baD7u9kCMppcRKzzrIg1/ZXboXl6zA40+v
0ws+ZHnVfZ6TTNs/gC0UCSuk5nJ+ll/DMFN7CkcvBlrNLP1mYtYejqzg3qUcdcLN
CSHR1Bz3fqBEFMV2mtODWjHyQe+u5xLU1rqnONLntl23W8yddCHlO/A5d4mAW3RT
3+AoXfXpYkPwCjfEFXSd+UeBtfzU+ogTtMBtin8WAihhE+YWP3mzB/kGrBbXGIEu
cCqS4dC1t53/C+NCjioEHiAFGc28+FEpNZlDc8c+m/XXdk6mXgnSagkiVjqPCWyk
6V7AdwYdwbU5Enh33MsHAHvzkguXvk1eJkMRld5ica18u8Iw3x1EPh4HlxCO9q9j
nkUr/YaF5HZVSlkZN5PgEK18Yms93L/fWHpNGDyoP5t0wVF0dbC40777vuXtFZyH
iuolYUaVLmWEoNwfvfKf9+dhcvgfNxdOFeHMFkEkKQUyCrZ/BmvF1P+eRCqCI7VM
XHJWSzBH2v+n53eA0i5XnGSKNXwdzMzdYYxdRpoRrVnMI5Zr+PCGUo5KNsQ4s6FM
9vGzl1uykZfOQ/wHnT4K79JVPIQJbMXFbpd09jD56UgXi1Uez5YNNaUDElvE86Qj
iYPgH6ICi4FOjklX47rPF9O39ZS/NrefTKu5qwOBwMs3B4rkznmDh6Zs5rZZj8a7
WcQfZSgCHojmfow77TJG7YX3q4nxO6ZPBelUODB0kXz6ug3mlv3TSHQgqeq+8eE5
FgctYOq6mnYkZwrZi9adFHyKm4BkLgjPiabXHVhU4pM=
`pragma protect end_protected
