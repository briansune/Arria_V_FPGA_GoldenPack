// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:21 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bl8tGy1WE3ykXvGgDSODDQYtxOHVwQhZ2yxp4P5+qlAfOrl1k8VlCHthGnZc957T
GC2+uzEwYq4NJ2XjT5/SbMaLxkHNcsvqBsIRU600L9yEZisqEqWrKXS4e4aMeprZ
VHVYjFrSG1f4uSPfWreuRhG3L/OQGuNrOPbmoCaGc24=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10960)
fJF0jSWgV20M+a2Fg42h49nn34eWJp5jPAp4qlC6EhNWwH1mMc/mIrYV3jM89MnQ
M/Kvc9YKhQzyQpTkRN8mtIPoSuPYmiTvToCLDYvVWdorzoc6wWC+hEoBLONVyyrL
1D6qDgn7QkCIfLbvZ2B6MvkaBI+MXgWOI8XfvV20Un3QlmbjmyKBY6wxFV242c83
vPqSWXtx9n+9gw2JVlA7e02lcdxcPSn1uZy/2m8H98oEwcv834dU0yNfT/zvjprD
NU2ocspyNZotcp4gAIX4QxHUJFoGsxkNb9b1/rVmEiQ2TFmZxmFcyN/J+oWy4Ch5
Ao1Nb71eaNGxKo6pMR8HQNCEbKaEVInPkdrFiuEjgW+b313tJvFAeoMSl9ss/jGB
//DOLi/8ZpKTu6abJG/tRPS3HCggqNffirM0YKzk81x4MoAWnGfxPtMTD0sfGr6J
ViO8smxcq0kOgGUcsKaMTySdsrdZqg26yOHXwLugH8ZtYYwAmdAVuDvS2RF/F8iJ
E6nofbvWarjPnXm8on+JebkMGdfUSJ1Kh8lJ3DV4rinPoPeDAEs4elFipC4X7zCr
wEfFnKosBqJXA1GKa3tXQ58GusbhUOsVHsAHSqVAZJRBAETA7vwhOKapPFUie6Tv
HWtAILLemWCm1i5E4H0S87ePI3ICdnaBUaXI3gS68V3va/LLRxKtntU4adUlghAu
ez/41dqpwTlArvPZ+58wr6B96FN4gR7CQD5NNaTtgpQWRjq1ATxYIt9GZVn9UHzf
vye88ZzQp7QKLfoXSW0oUENFsE3In3NP3a6A0AQ5V/wFTOlTn3/U8hwziH9sIgXp
mCqD6ggrc9pORJDXLLa6hJ7xiknGjrMJTxwPFq4xXF/DQ/kslX2UH6f+/kcL1dCr
kwI81+Y6z0WvjyDXPiHng0J/Gp6dku7nLNnSLn+96XKEhcbbmHFDIykj3YWO9mxn
TWtzqGS2AZb52f9IOdzhWt4MT1VkpagZG2quICSh3QzkprCWgVGLqp5f1NslL8Y3
QXDAP+xXalDN/67fHGXKdyLG5N3nJOAP6V1vLUpCJch3BBTQCdXd/krdnNxijtul
fSnINxisprsaTUrEcz4JVqpy37Pbxu6es6aMI3tll3DXMSdA2ROAlqEyo9hsi+B0
Qq040L3ohoGOFoDQcGBEWfgQoEw8snpNnVimLAHRViihAWgTQ6H3j7DGFHhXD+cu
kL2YPL0ilH+6DWbEiOBaOC6CQ72C2x4lI93BOpMI3RJwmUkY5DU0uGTOuf18Jui5
UlreoLdto8HlBK7bJg/VsZvpNNoeJB7mLuypn6lcBfj9eJXl/mJzt/fi4WjHFmNZ
NPMNRWFI9OPY76bSXIh5Mj8dbeRKxNMIyGDEClQPmrMnGdrk3BKMdRrJVElJUh95
Ily0JN95bX+0snQeViK2UoTMeNpqjaU6aBZ0ePUTtap9tvL0aNlHdGnoxmUNQaOP
ISA8rMgsWp/nwhZiVPzq5v3GJSL6w6sNU4mxWE9FXVrq49/D3195vJI6YNk/8BLX
U2/IzfN4r+VSD7908+ZNFXMIS2oAskb+z62MUJN9OQPdXuReFwBT7dAcK1/0pssv
LzBGccG5K/Zn9+Q3WXMYT8Q8kOpojEMyjxHhqVfOdArFf6SkP/WCcGiFN2wq8a94
fUVzzjbCVoSQjKfLrR9wyzOlHgK0GAWQsW103MhsPdjmKzFcKZxe7b1/qU/FSawH
d8zEhQByWKMnitHUmbjbaYmigsK0Ur9MhHyMiCGtbI7NnkyGUXXH+wgM03jxFVEo
X/p+a6DFbS9HhXGHY0GxNxSRA9BOn5H0QLtR3N8QdebC3qpnCUrqjEchZl0yukmI
dwlH4ZvxWG2cloY/vLmdM60zBFfp/qIrQUGFfcdaIkVtWnUeT9btWIUAcgpJP0Mu
Et/NsovMxZji8CvpSQAtQq47CNujOnA96r1FODef1c7Xtb2blDJVpzhjeFVU1jvW
TMk8ATLRraOywHIk7w72SgzX36sDvQWganFIh95Q2dvO0gsCiM/292H9Owo7BPIu
yOAcZjsDFnHptLy/ET2aO5zgsBVZvS+x4a/ls7tS8WGxy3axZPovNEIkhoubdU7Y
emOVPXD0mX7F3/kEjVPQ5QMvzu9iGntsM2b0NdSsuOcsFObItpZNeRFKBjv9uA12
5Jcr91kWjl1kUF0ZUstmrStlNIyvAH9VuDNpcR5SFmF6bc8Q1nVxFZtWeBmgphLn
hQW5AyfT+27lbVbLVQ/Mk/+NAebdtsQVpPKErsxFCBFjMRZ2Y8SGIn0+VkmVPgHP
lEhopjF6R6DA97rv33ReA2H7uaRr5jyFrhJHe09G7dbTfjNEa37MZBWSdUuZ9p4f
2t1cq6mNaXC4r4/4epkgXEuYopGqgSfKBFHR7agpeQRyBLzS9KYk1snh2eKx9Qib
5I4aIUsoLJvu4N8Av8XVzw7MHv8OB8wENsvI/F3fwierr4AduYQj9tTVHTFZnXga
DLC2jaRwJx/qWqGwV173EMyhWuHQBquEC9gTs0mnQEKie7Zw4M/h2Vog1mIhpoyb
lw1rDJJqyzU87ZPk7fB+8cp9unprI4kiNvN9BgQU6ciM60WKqzC6NzQ8R1wqmmkG
F1LdYsFiGpxSs9bG9+t3vcyk2QX140Jwet7h9q7QhiJ6WGiaiBeAtNOuEDt6kX0n
a9PAtYMI7IubBxI0R3u6Sbz19tZEt1DdvcSwJ+yYZGOaET3rLbxxNoyoFK1s/Q0y
Q+40Vap9ccER4pIQr94Bm+fW4e0cW3o+MHDJqpe4SsZAAEK16UPc+2Xus8UI+dRS
iORVYxt3qNH93uaUXp5cvxZqu/qJfQkTnCaoWXn3FUHRmBXx4mBfuMH4CtkYg/9F
tcRUlthUlg8qIiqUr3uXjrqKt9upRtYg18mHfU8bv9E3t8xUI+BJ6tusKI+0supI
kXY81ItQ1bO84O/Q1c/NKWTGeU7lFK8RkOD2aE22y9IewOWMJGZvGAqS5XDjZ9Us
B4cnp74l5II41RIbMmFuA9g7RQIpMmgbBf/OFhpC3XWctDb6vsnCdtRayOoGCIwa
mc/bWshINpNwc+Hz6ZfznmBgisp5lsXMKPUB2ejQ+Z/O3eV4n4b2+I2ZZuZihnYC
SMAiapkIYsI81ov3GksCJngM1fysSzVDWJ7nHRdXok3IRvDwOdBjMzO+2jNemVZh
g0Ezb7+kVtQOF+PZ4ATq/PY02sACVP/WzV2l4efAvqF7TK0iyKMqvgFTO6Wqojry
rQNi26LL827VKvGmmC0lWqo6y+pGw2TOCCNsxtdyRFJv6z9xOTjgwFk8AibNIIlN
BtBmqDVwzjJ9lhvesc1R0t/Vt2IE99/Qg7AKRUFuFMgkzLsdsw4UfZxWdEkUINdd
9xXmzYWxTCdnK/1AyXdlhMbVTNd/psUW5uOo+RYKaoMjNtqtZzu3AV4JmeuThSB3
fprR6syHI0xTwQPCj2DzU9UCRs4yUAoWDr0cJt5agYNdGcaOJBwSkb3vK1lQYZ/M
byO9DJPZRptZeeSNVrB+FXMMZzFeIPkS/y9lVGUmRKOR0k479miqlJVP5FMAw+bS
nV3ocoJoMCeljVf6w/B26rpEjUSHcfKytR5zsY0p99BhOkpM+q3U7R4KChQ+ZNj/
l1It3n5z2pAnObO9H8w0YETz3oVoqZj+10mjE/j5J91SB2id/21pKWKim6TvoXE2
3WSIwlqe6DQ8kCb1DKNdJ7p82epTtE/gNLAxwOTF+TgzAYk8RT4bNHJ9AutJfv75
AGnuxK+2cfujQEur+q7g3kXB/3NNQ6NBo5X3WllolM0TBIH1joAdwbatRgOp6yVV
Fnf+gPhrqjvpcrk40C/bY04Is0PI5AIHw3SFTVWyLI4iY3GAg6hR1KJtdzpyUqUO
U9N2opQCc+aI4FsIbpMRMAk5UB3i+PTHsa7vWcvAcKW2Kpj+0L+7FN4Vgba0TSr5
0zzbUk2YAHryeFelXA7LbsrwCov6Coh4sdFS5OOQUWbDfB6scsvQBvvgigtrR0pz
e50zxg5gp7jbJnij7+UBEwSmZN9sx6MJlAyKWhqGQ4HXC1EHz449v+EcqUSJ+sLY
w5Ar1QINud8Oyjw1OiF9JDOKeb3uVeHwzkQLiHOOf9ZnbA9XLqMrXPJ2TElLSF75
spRtmdD7O7LDSorlxIMh/xSKdL95D+bkjIHCKIGiRWaIWFMqw82QPIH7rccxRwAD
BssJ6nhab3cC/aYrwu/OQ6vE+ikWj/yM/UIqK0IZBfmi3Fg/HxOznyKzNdyDphpC
I/FiBk5xMl3zRTgNQSUt2RjjWFtNlM0b4dkCkG5brPkkNzjbttZZ58lWEu3yesed
8mDE104NBYA0tEwEDDUweZbb34bechhlZy+msQrKD4+epHMzyYxFHIeN9S44m4ZF
7D9XKonEgqHr2Jmo4s8zjtSdMZ2NXqtVu1PEOqFW0nlhZvjI2/NqJi6qLPT9xzem
TgTIY6/UCIYH8A2lEVB0mSsMjCHlcdVcJ7YdbRJFWtv464g2Jlf7z8qKeEJw6TbZ
WeCmYX4hinTxgDWOZoL7z8jJpnMfIkHb0EjSVeHL0MZDp2hr3kxYFxR7NydxopkL
pNEMmcnPKbd8zYhte1COjnlvyMKZcE5XfC/eJpj+cjE4/J0cEJeW+G3OsGGFTpxH
hVi4wyodMqEk/FYNP7nLxNkzVtNkGfJo3bqe9qiNAs1irvdZG10jNzixsp6EcUzh
LN+P7dAOKVMup7BxjvdLcIk30w3VMgOhXTzHfuLlsazOpdS8HSszY3urjm0PHGkH
F1AvGhOXeF2ZhbsEGeRaFPfsM7nv+VlhS8WnVn6otlcP60aHTpvSd+oBIDgygxir
k6ABzaBili4zp2nEJMqrgYpshYdjklV1oCj0m8+CHxOUJCG13LA1UJtDxFd1v6D3
gCTpl58TNcEKId2OKn/GG1lBlG6lpi42ewmy0Zm8H4W09rK7eBTDbBboFBq+xrOl
KEOnCw+Um1YdbvpTU0pJMnNWINwOFvvDKO7/XgnQ7lFOb9ZSAab5aWrdnSPmKSC5
A3x4bgX6+uktcaw6W1JlpbZlnp2WZUB+my/qOUyNLR1GcYG+yOTbxYb0m31K3gjE
Oj3yVLLP9IJjZILjgBJ23IW7UxnrBfH8JsxJ3YxruK3u+MyP3hwliUAoNxTykkUK
ajB7jiwJzS9mp75FZ+qS3lGc10yr6v4DfLH0Qz4t5+x10iLfWrO2hcv/JLuW9115
4LfrEr6fWxMfxfTVCqIGLvEaXkU6r1rjVgNEbT2geNDFeqqjser/St60ahu0FtKT
N9LtWzJgjDWWw8wPQhk/vb+SSFXHtTYPhPLAFGm51zTo4/8VnMsgM83tBIKJ1pvJ
aL3AlwjiCd32RCJSAA6vnJJgqAXDuCjgD+i6nyTN9xueqJ0IQt2Fwg84qM3BSLMh
Ty73iscLYLnK2VeJ5iR2VSL4GijfFvXqe4l6yFe35CRI26hd+un+95mpGtc6348d
TNM77zIIkFmGsoKuqBHPWEa/QvAD8yTfGx/GDllO12W6GMqlnxwC2nP/pIW/s5Dq
7di4PWIDTdAt5Z8tfU/p6FKfIeBCf0AHwz65mVcU9x9fdrichAEPhvAS+3YenO0o
7WBmoRnu8/75f5xNy8ffI4iVwsh7FAFaoI5szUyBATZp28UyjTepiZW9rFw2PL2e
+MTOM+pwgOTFiRvhf68ucxvaxnITVbSOvUWlf1Ts30xwiAoydS3gQfP3TWRAQHbN
ReY4HKnbocHWMzeTiej8QcjWRsGFkq5wehnCst2KGCkywQ4jI2kl+vatlb79elae
HEU4r8W2iFFKgy7DZFt4pxOWow2GFIREYy96hRYsX1rQfdHqF3Wmb/suGn0+zSoO
Ve+6FmLOolBFTlygO9Fsq/Sa4l916jq7rffDPWfcNZmnW196Uh9ZaJ5IO/liUXp/
JPjhmTMbIilDRlHvq2GQZ5/YjbgdHzbuRsQUbMJxaJjoIYYl304rtjSJ3aEpvJaK
o3P33KPBIx+bG3eBocF4frEfMZsUuW4tcSyV8DzOIBolIv39AJPZdNb94e9AAxZc
bmd+eaTGcBvnGJMGC+SNAt+mHs4u3laBiI01Q/x60g/b8CDJXCWIXnqeGdnxi6SJ
ieU4MnRDI0jYxNfrCgD4I5EX4HOjsioRwR1pnPSB+Tgd2913jBdGInphFsB/xVlX
cWhUWRj24ui+QVNQ7bpQnuveuyzqQfgo2oW7N9s2PTv6K6id2db6mK6h3ASqYbDk
RT7FMEiF5JdDnbzX9/N/u2e0wViT8HobyxphLQG/eAZTDIywr9ysgmfRW4f6hckV
duuH1P6qFOUiwGS+oqzXMnH+Jo+kl0C2Qa8X1TzLFpT02Us4klHzRe69KJ/iMNYV
rUy9rms5sopKnLuKddD+Kuwr5qRkVFbw24SddWXTwWA4DjqREj+85UG33D65REwO
zD6xWGN8NvwKDg3qCLBOXSzv3806dPzwqjIOXOM+wozELtDR3L9xq6pQF2UgzdZc
/cq6l3DwGAHxHEfYXnfq8FVhlrzRleu0zKU0WAxvC9bHykXJ+o9v2TExPldyZQ5X
ZOsNIBlcG5b8hHR3youjLvaLLRF8EQgyg99iAzZ1T5st2DDwghNWLoEQbg6xLy0z
JAOBBDZbYSkdDQxaWy2umm35ScWvJhwJCjhk3n+YFfKadGO76tUL0wrnSpjIXQA7
hpKFzrfig/iUcx6iox5/zcl3pdy9VvYOF7G6bA2Lst38Y1seAnnzX02+WTF7TSLg
6dELEpPguYhGzUzfVyHFhTwEzmstoPkuwzCS9cykb58Y/5hKZRAeXyQ0sJJnzohv
L7poqeLkdHcFID7e1VnB5iAF1J/bnQelqoXlvNe/c/DBmR6Yer/DaBQ/zzjuDSqr
95QIYB6OMIiS9L/YZwTnEzQFgY6L2gnKqWkoyJFe2zWOOvrVC4BMTEFuDE/CyjED
A/Lnu88gUtSlEq4qjTDer/m4GCrm2K3xrlFE6F0J/Nxrwdm9BIbnytzhpvUBmiN2
yqyG1+k3Inxuln9heQmsp5ft6pGwtqP2BQKs1EqClDCs2mTbod9SF4BRCyJWGGQQ
aggupPjLGP+Zu1dbtJxPHgvF+NnLPFxoiB0N9OPGe9tNNzjDb1kIm3gPlerGcwMS
ms7Mgbr2EMt+v8gNIsyJPvgqHFSEz+QtvBEZEiZ0NVFzpwlvei6qWRbObJ3ckLqL
gszPoXUMDCEMzQMh2bKu94bsXn7YzviBakdO5Z4mjt8ijm4BdarLK+Gb4Bf91PeC
zbN7jvykimAa0IH8i+BY0AwBTEz88mNAKlqiQWieF4vuSMxrYDCcjdjlN8DT2XwT
E3qawCROKgMzijim7oS9e8JEfhTtM0SdxKryL7zNzETZ9HbnqT3StiJ/cSfnBdnJ
NSv/7EWoTZIXoyhonAH9yp8Wrv+TjWx7EDYIeuJ/wmYrTtJ0qfmHBosLCKI5q1O4
EM9hJuc9P4vKINt5fntmntQo2bcd2Jv4WKQoFpNmVz4YnN7GxFHhDX6+Lnpwh4k/
9lpwNSW02scOy7hpKbye0bmEvsudg9fNU1+Q44IFTSJ6bUxuhltnrNXgIL+OCLE9
EFhemAdS+kREu2Q2QYQrnJwAB+NoUBE4+fQpzAIniYYNVa+uRYfwn84n9QRLK2mI
r0PpF87CSxt6pjd9l9Dlu8h98v5S2CXQRcHUwXN1JZYAyvVmguMKX0yfuwKx/WoZ
qTRemAA8y0yUsmPuedeKQUHhPYJRI5oBAXlg4ER/6dqWdmhdK3J0hcrThx9uUTLS
ZnFrYFyO4EBv/sNX7eOeLTHsO91/KQVrs9q5S7gNDa3kjetkiJuqpYw6V+jWOJb7
nakXjjzb7Ji14CF3oRrKyyNa4/g0tVY+sSJbcI5Be2F0hNbVZFwsd2DfIwy0o7JI
IMTlrebo1X/Lq39kOZdPFazXB6136/fDKNnnEND9Suw2GqsSbcVBYqhzRPlnCFZH
O2RVixYlk/RV2qPolhJ/Wq/7sEuTqgXyHoyLfut+JSeONiz8w5E4C/962c3uKMr0
ZKXtXL8ixOcYQntUxLwWG5wZ5FBGEhSR7M7LAJ37yTaeUWJGdHuwMpVahztYLvTb
il+h7BVjP3ENopnwK3SEl0nrlAl39JfcngLOW1cp/fJbdmO0ifodw3KSVASAh9Sq
9wiCjOpmzRumBVa6Qfv8LQsBj6jG843d2fmioQXWpxd4w1E1/rPfAzywdj2YcleC
DjiF8XICK3ghIEDBRW1M2xYyD0CzwOs2xyBOBzGDVBIzK4Yk5CMcUVn46vEr/78m
y/0dRxAyH0TQGdatxmeCVblIeNkPosu+7ajIVz3GHCWqKJmBbZVnAtRbxOhuMwgS
U2bsklxuyk11FRcl7ZYdjwnrZ7YN3DGolFWaLl3qMV5F3jH8E3+UQi97h+6cpxB0
2uUeoc7envRuH6Kc1MNADpzZH898QAz6H4v7pUS8i9Rbdml0LONLgUuLB48oGS2b
V5caw7VHvmY1S0vLU/yxGPGgdR2nXnUHrKw9G0UvVCQJYxhLeM3c3m0Wl+QwSAGb
wqYqXZgLoUDUxzMIy8LJ2eXgcwUq4pPmqZ8xFXmw4IiRUssE90rGzC4ApnqknzqQ
A2X0J0l7270Ij1FrPVzsHDoLNsJ+3YPwQPPswQe+stIiCG9wd4NqqnousljkUt0+
W+ITQuqsF82AugWEBWZWJDRVlKAWB/8a4QZJKChT1crGvhR+4Nd6CcvCZaCuqHw/
z6XJ3nk8S0IldHSJ19Jgv1kW8Fhf0yUsQEYmqJul6zxwEcnmA/5d1enKDGh4msvW
kkZUeeRrxFBEcyuggpOf+NCrniR6TVFJKryZQ6QJtSOujXKwu9KtUOqeL7GZ5SjC
VE74g8u0iXkVWTpxJLhWDMdY4O7MbOeGQRX/eNMr1vAEucsg9jY+tckh/q7bAXUb
HoKD6wxmbN0sjEJ0YdLtD0zkJ5OkIMot56nh0RTQJY1ZFJJBZe9+PedG6yvsdCmR
xlf8ZWX1gZLv4UpjUAmoqw9o7OZPVDe4IBYAkWPXPzHyPyabbbocWsFXjUK+0DHk
a2arz1FpyGgx+Zc0jZ4oxvuSU+u3Qfva4vP4Mi/M4A4D7OFZhhNYQvXIuozzqcZF
acPB3UZqkGKT2brT/bZg89hllylxsXsNxCsHy8ZE1fPWzQPpptCUBUlhaXzd7Bh9
0y5r+shU6jo84Nk2BRdo3cbSbz2kEtFn33E6ccBgTYov+NwknhqOUu9RNt/+Rx4o
WrMUQMkeI+ae54WUJaKHEnB4LRsywzfqDDI9Urmr0YZnn0vyzVsEFPN8vXEerLZM
Ynqe/U4cGHU0jw6lX1W0xrCpQoNnOP1ZntZKfccCO0C6/A4l57DXOp1W6kt16HGn
K+K9LZeCybLXyTsTiNzQw3PnrqNPeiuFyI3xj3nL5/c6FD4Z6XtJf5uyat5Cbobt
QuzydHq8yj/yYqjftOS7UU06/zgEiKW8RQOLeb1nDRDq6PL4MJbfQIyjeOBi7xth
CSzMTvaRK0NEQrYoVjM+HZOWdxIC6qcmIij386CYN7rs0Ur2cjq5ibopSjM42n/i
anWcxNXKdJLS7rZ4R4g7ZDn++bK5BwRin1E2aEc8eg1tEtF5B5vaiVKX+pqavB3Y
Rpi4f8o7X/D+6v2JpposqBtOBWTOuw1Lw9YXQ1K4aApy80xilG4W46H3xJIW0W2b
LuzcpEl02NDopgsXXfkavhQRu9QEBmywinjPYV6Am5XN5kDAtiUsYKUSMKNaw9cK
9bgLeenT8YVUFHGmOrUJ4jLe4PBsTUidDemQcxwBPqJASpd9NTBDDmBMQq3eMbZd
F3eEj8r19fAzr9Y42S4iCsX5bL9J21LFGH54Cz+GIGbJp3sJlSpwWjvVDhP+wRzJ
hf35Ir3Y2if6cgMhnedCSXEIVzxhPupl2fR9u/TOb2H6abE1a9pnITTW+CWHpoWO
eXoUaPSsut7B5Ox30Qf0ujaq4irQSqXnTywPtxEmTzhRcnwq3nmhGco48isyKEDn
ms4wIln5jVTvOWnOr1827jvdfpZyIQJ4IxghVJ5sWgtSCmugVjKDYaaC5OWdCXqh
7Nwj1+MjTMbtYkPkRUxvPU3l2g62VcvStLQqZfjyKdcd/5SvOlX0R/4BNZfCYLdn
BSthhMHRfgSkbeaFrLoP0mJDeyLkYC7fVLg3PgOYjknbTvIPqoQ6qWc4DxrdLUcs
tf/bgRg8ETGvTO0va9OGQ/n9WmwmxXdI3hOzZ5QB9a95PQF9tBvet7Z+HakAX/nO
EKHne+pS9WfDfPq90SHxti14OJ4umkAGnvLVKWfkWUTQxtAiAUM2RTYLv/Lk8EuX
s/WOOF2byWd1EttD3xOG6c1p+G00OjW0seEPDPjTV9ovxWWbokMqQwFhwshXDcWA
/epAFPhdiX/16GImmJuXt+AFIYEvPwWxjphD5C4uPwM7r/SIEKDgx+oXvWsI2ktl
wiIbEKLvPtFOTZECWGVzJBp07yDnCDNPVVXwZigwDigKvmD3KVegvGTNRnTYoMl4
B4V1V6eBZyU1Hfupni98gFuFnpDaJwMvcVTVyBwMZKYMR4vseyEyw8RjReqLmk/H
N9J9o928rdTPKO/OZK2rTm4dohiLPqCTMvJYpaGg0rAbGQxnPMfxhYeauJWRb2kF
uZdAjtY8iKqSWBYAIckMDvSr2SiBvflcV2bTSOoMKFtIlVDlR99oOj1mJQ6iLHrG
lfn2GTDP8Wph4cMJHMkykikA+ZTc8DSNxgVX9g0+CSIW7l8HEovG6a2zgKQNcuoO
ZZg0lv+bscBoeMl36b5Tvwumgp5b4rRNNzolNST0Oy4RGPSjpr84ravnC3lwZfpP
kQa64G0QTGuRrC4EYAQcTW9/22Fg/YzBP6imw20ZaSbec8PyP3xu74V1rNKdmdbC
cq3Df8hu/3cCR+29e+xdKglwGco3UoDkbtMVt2p0ZtVv8FeeFg+IjYzM/nhDtoza
oATBeTRuFcripeBgGkUSI2Hy2skzbgkMrNHX6yQ3NFsmZlAzqxUwJD7iDGagOT2A
YPD3KbljXVHrYKiiYkw+x4hLqIL0Zk2dymnxHEQlGKUKgjm9RJqNRQHI6pY54BLo
oH5dQT0QKrVz/+jRxNFbsaDVm7pv9kMYA3BB3mOlALMWxg/fVQdmTPUEL6WN0trW
OipYLPO16XQXjyK7coSKgZivg2HYdPsTd5xeBtCW9BJPzmJjW6Df/mltuo6A+WzG
rF3gQKc3KwQfftvM10peO1fmBNvVktqYVltaFo8oox9xdsxGiVDzucVKqGfBJ+VZ
o1ctnqx/jcNnscvHPRgm9oWTcURlM472eJaEnsSoaKmh95SFELbe0j47Pt74UPVy
aW3xDrl/BFbebAxPLZGA+rJrijZmM05QvNiE7mPUBiMEKwTNIC3NkcHxy5fpUq6Q
e3glnJRP21lKE1MbLz02027rbirzH612/Ykydj5J7zZgjQG+0C9uDHgaYsPAN48S
FAe0edJl/heYwXmPvN55HLMZ0VrpWVdp11EtrB0PwnD6bUzqjXNx2YyF2QnvsrqR
NdGHYDlM7vL1WMbJF54cq1wNpnU422N76nqqYmdgigb3tmCrYaUL8IsPZ9k9OG8z
6+9FApgKnrGKKFldKXP1HU8OtQvkzfD7Lq3I3NTfqWKXXckEjT8JZXqPzIc8YQC5
gFPZaluCTsjF6LUB0PDmD4g5Nqv5Ih1OcUpDVeVl8SONWx6RfFllQuKX+nRKpyWv
eOiabOWrDQ7SCWNTEJwNJ/ch+UrJYpUVTmhP1X04D6EhIHTZVrDLAUc/zs+Hf3Us
UIIpN//sGs5dYvNYGmdoYb+G19+F2IIye1TZqRIp/d/bvXUmPcBpjehW+vGgCcQm
IaKu5MYR8xEcxFgCRxYcvw2+gotFdY8yZ/KNs/QAhC0BsVB0vN8h5HDdxfM9XfYp
bEQRRAOaVOq8r7S0Xzd05g0I3X1qPWNK1J6eciSlH8kxlqkKCKRKYCJM/X8HhBXn
3MM1F4Ny2p4705q4H9qYbAykqFTJmmDlR+STIGHnymocabb5WUCDqI9sFG09kMxy
G6zA5qXynh2xHaCW6lSput0r6+Rz9V95rw+ITjzOmpgWq8R7WxqNjDNrvCzsj6GT
Vat8DRgpRBFs+hNOjfB8GGn3efP3iLCPC3kBgSEv2+scWG4S1CyYffxmea/HQXUi
As+UhKKR5fONXW9yfZNjdvnVoRJh9SRg5C9Eas2zzu7VJxXH+21Dm9iZlAUFiTvV
27DgpJ1ZXGo8gm5JXF7mZX8X2D+Xl5iFFtGQrn43P9LNyXTFV5+zrG0V8bVtzYRp
iTl6h60wZ8oSieMyzcc8gZSV0KA1CXeGyWgMV1zyQtYycW9iSeJgjjJBYlV/JJ1p
cXKYy2gKsT51a9SDLIPEkJ5TAgq3F+M6iBte8EUbvvdftEVzSaKwBEo/qKxhWN+o
2JYWV/nxfiR7LMLHo1AM2XM8tSmibvRcZRB09YPYASli0yAUs8x07B/3OtOb14+T
CUpNwYtIRnY+mOZNG8KZwPqDeTTK8vnCESHpWrWdo68Isb3zBjuEuzQEG3dNXXTm
oGqTceJFRkg5N25lN+siWMxQTke/DWC+f9Bk/lXiklOxGpyGVo5MwXi3hLOcDHF2
hwh5AikFqSQGkJ85qtcqKYM6LTqViXZNj+vERDLp2aCjhYPvhN4w9l1EE/YY9nvI
PfguSx4ViG12kkcoNyEYHDjkJu/a/Keo8CvqeKvwzFixqldAX7H27jKyEycn6TK7
jItacFxQtDYNBA0CHWaE0F5eMGbZirNOjQ42HRoLzljF6pZ4wDlG9ZhqqSs6xIL8
pwDoRbUAQqtJKKQS1kk+SOXkI7O6ye12V2dlEEp9eVGsLRrjbI7qR6wuhFGpDI0O
Ip/9kp5VeBxmj+12O9Lx4Xs7UNeHU9AXoHwaXkM24DUvgEAwXpyfrCmAwClyxjDR
ahgKqyzW0eQ3aXAWxrGmJytU3CnCyUtLNBjZ8lmvxBLFzH0FN+MzGYsve7I3lodH
GfepdBTrbjLPjP1Td4/8jMWIVanld/ZYHrohBiLdml63y2JxKLLh5FhkASqdoDRA
UtXLPxan868v9MSM8AKdr7Wk0tCGKDKzREZb8W+x7WGTsQGXXOQJBrhDT/eif5Zz
oRRygnsHWLDBBRxVkE/sM4ct72dQAMo0rBbRgIbI7uuW+8fBeHEc82DOwUPdgsAF
4581kdIbvuuSGq9L2wfenyCklt4ZiHWJ621LYdg6mwFDxu79Lob8PPyqfA+Uw3+b
8oaTisAD7YAomwKh2rhUomnC7Be9pza50UZQ55feppGr+dW26H5cZuWDscudN9l8
9U5WMsPMTN6Mf6fv2+A6p7gZprUSClAWIjsqJRRZ987AgDLspVv0/KaNTC3hI9Qf
4I0p7ZpqR9q8mXgdqaEerSJNsd22ybqdBPkybRiNiYQ0lfRmCgkt6O1B/RM/Gyob
OIcwVIeyj/HQEoMaNNTNOKsFn5ZIVGGCQfEgZOywsCgx60ImK6oJOL8RSxqCBaOu
LEx2LO8xB/zgxfc5Zdn+d9fiFoHvawfsfA1tSceOI3xG0Aiv4LKR/kjPEOnDltBA
9TVSTAljWaMS3jPkCx+BfN0DMCZMPbRkpZyfbq1aNt3JT7C1x2MLcGo+NP4L0daC
bmr6pWmtVyxfzMjj8t+t/4FgAh70DgxPidp1OEymeVibVy2DSHetdQLbKp0c5+Y7
0NGTMEY7Io8Meu+4iXKs5Bt6B59D+JSeI9QDR2nt84um8x1ZPMRKjNPkGJ22s176
hihH4yCKI+oU31H1G6IbOKT3IZ6CV5GxI5NPkGfb8TafMdcFgm+czBlwfVW6M6x1
8IbN1xs9kqlsiH3UkWUqkOAhkAo+NqdZGuwxhM4/o41gX8L/88Y/ChR+jUO0buZ9
wOKJskm2vgosvKepRghiIaStzC+F2y5oUNSDH2jloazKiEdtfmKbBv35kJgKcqaD
zIoNdyTiMiq2OpUM1wTbXsNJgcj/QEIQHFU6AhanTIVEfrA8B/0wuy7BfQuVEe6a
EnB6NbjEOO9Dvm3dFPQQT4hXW5eVKEQw4VZtW2rHCQELDYnnBu47wLfwJYJJjze9
R+67zyyeFOdHU3hW5uzDQb1jSFeGmbcw6Gs7EN744E2feRitAHnVU603KfcwZgFC
LhsExbLP6Ss0OG+RemJpBTttZkJnt5oFkzvUxZObEhjBJ+euduySdv/2ufyJlv1V
iqEsSHGLdbZ6SzditJSl+/d3iuFSt5PBUlZ/XcWu6Lidu/SutmHyiqVTiHonZxe6
jhCr2KZY2sQvltxNLUQm55xZMujoiunNGnLWbJj7yIDJWwbTHzmSKGXNbbigKVlb
g7UrcrsikJm85S4UZtzmhNiI15NlnHbOdNeXOmgVDX5gkkTJe+joQ4yjuhPZ7tXf
g+2unrP4llXvuGFNz13phOijioUozKZor4ZnDM6auoTycX2bqQYT9tCIzUAmtUxN
rj06iTmzgHXTtbvZ/8z7X+gHQxd2FY2AeSt6Ub0SE+V4/u2R9gCYoXQJweoJLRNv
IUy7794jyRbZXPF3pt0jNw==
`pragma protect end_protected
