// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CDKqk0e9h1NkwBgesiQ2amb4K2A75kdshc7S+l9z/pASSpAoQTV4sIKwJ3D/Ven/afPfzjYyBig3
+23aERLD+OS/WJGw8PXuLHXUzrCkYAPxzobqSJlA3gCmFIjhLvbU8l8uMwy4OiR1a2HjVrrh34zh
O+w1U8Vz5I6+dgeU7IrF6zXKDuEEVj0vjWFmoQ8bBQ6mspMUmH+AA3nuZ/MlmyuTOVIubHF+o435
NWn9axOaYLOxWdPfrvHgK44ztTocsS3d8vepubvoCfO/8FSjkdVTNNwwwsXtabqkHFIoWhCnGeq4
d5VKKrq2o6bd7Pdm9XXj/0gRQ55q9lL55FU/FQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 23744)
DCm8MS/DDkDSVJkEYqVL6RS0z2uBnNalXdqYHh7ISMZduvLXA44ALukOHjldmzKnAqqBWT6dUvXc
cM2Sz7+Wv235F5+KjOFHFhWHmw1TLZDDUXx05yoxmMQDo+SP5fId8pVOFI23q59xxAufDHWmUhzb
faHsnWDmhYqMcFuP+Q7LiyEzlR7mr4f2yjA4AMaoO/pShblgHEzlTklaevyxseig46t5Hn6nYFCA
EeggaC75tHqMKiRzTLfoE5JAZRDk5rPgDMilPwiw1OKnU6NW1t3KEPCpJbT9UGvPS0XaUUAH02RL
2Fb0h27Bbtq4rIyGR0MIGoIG9QRvUV7eyznVsh7Ay7zx1xF0Tjc9JqaftNW5P9qEdlYZe5D5VsPD
tQ01ZcAaVGPIk965rvqDZBTkPJKFY4l0peJ5b4PocvQJi46gdSEII8ardSaBXZfu3dMvVbHi80sa
iaNXIHPkZgSclL6cpnFOoBbr2awc6zFDQIOmtukaN07bwH+Ha2dvFhSYz1uWN03ldVefqC6BwheC
ks6I6nfdSN6maCMpqe0EzHnK8vD+6/nS8HkiAphj0UYPKGL+94j86DweAJh2prm8oVmCckTrxM8D
sgp0XpQZLOYxwHamWn3t+16+jlBgje6UEorS4FgkzpoAEq3ngIBXzSjzrMZR9uYprYQP3P7TqT2M
Dfm+JjcVC4X4b6xIQPTfW/Pxs3/JPWRtS3by3cwFXt1qD+fcqlQguzRF+NQPcHzeClNjCjHWDyqE
OcDDltSFBEwr5D/PUQ0EeAcmzFsEPxVUmK4MqajfdbSHzzLe4MjCrYSKQ4J7sXYaW5BgvESEL1qT
GN3XPNnYCVikOCwV92OMrs82OlK3O0NQza2jnHxqadNeO9O+FsVM/xEdS0beXTJldAsDFLQNKpoe
CHNvuZxWt5o/sFDyAAcem4uoXmv7A82eJ5JplAr6vpA5eMxQ2EAMZd4Qa8+JdbJy8A3IWONrvRDN
I1IBH4XmN9LB646oMY6VoChM8K/8MN/a3Gmid4qrGvWFVSspvF4L377kpw0PaMuMEdtuHbIeWVRM
P6M5Lna9otzLEDxNGZo2V10avi2gehdaO8XzTusV7I2LmKO9qJyTmDgfQCGDH8TArnm3NdRzq559
bllXRQUmnD46LvAq0cFAxX1hTzHyMsiw1ZPCE9fmYsTNbRYzfQx21a1OFwmHGM12DEIZEkNe1NEA
9PzW1y0DQOLJxlyYbvPAhytx6NCAIwiMd7IQl2B5HzuzK0grBaQUgyZrUmRdy/kK/XpAvlkzBgbI
0b0BPw2USefdGfyN/4zRRi2tPtZetKMvll7IdGPFd7Ve3qeh7C0l6RoEXYV0WoUh01svM76H9vDg
0GtApKCNSv3svvyTkm1oCOuBXAbutnUCxyX6yRegP4ein/uD/65PFm+138UrBuzvcPBFkwF6rX/a
Y//TAK2w0tO+zZDijmDYMqBYqYuhm9wElxMrfe5M+T+FVQs2d4sUhOI6oxgXb1HTsYYUTJ5ddiDb
d14oi7Ibs5SI/579o1NiLdFTf8l0PFAHuVW06+1ApW0Af7Yh48GXSZauaCy3h2NOpFH1UK5p/qKo
U95e0tXQVwfUVX7Vep/UG6E/O8bNcEmI7DmT9amlh92MvPmHalduSulGfoL3gzi6l+cY3LJIfB0u
SaIQIfTxSOypGOX6G3hItjV4m6aZ/I4plRF7RQ6bIaKgQ93WhBSZBGDGDXuJcg12oJoUp0fuBgWU
zHlxyn9HNrfnLcEZt/ySX9VlYy5tOads+Yimo/1vRf/YxbRgZLBxzmkgthHyIQbUt2/OJcU8YoVK
oIoRfkjUR0xPV1a4C6MbS8rohyk56pdNtnVbeJnAuRrz8yMDsH/AHaekgURHMdCn/YEikSuNGSQS
LLnW5D2pRHOAl/yakHKf4KstZF/asVvzETISI31cGObuFQqukmilBCDPjcBd8uDxIq2pwXkpRV69
+kL/pmZP49Xdwgjg4KHkvFEpwDeNngUyrifLXGgphTTCXTLdl2xbNrrmDUxmahKpZ80FZImkfmUK
qQ8+Vh7+OtmmF7Mimg1xWn3tVWO9MqKyI6HW/ZcDDakauF6j0kPw++088gXtNm73nGZ4JEjf8Ofp
KfmPu5r3Um3tuJz5GsJ1zkUXKhFaU1Q7jvKehJc8S/GDZiQ4x7b8SiPafY8+VOr8/5ofibFzMjd+
N8hiE/24uLG2XYtd1JuqN6mnr2ZovuzAhqeQuWVu4sxmQoPrKMzCSvaeEPRENR/sXclH1/qwEqhG
WJGafNCSO5qWTQ0mIe+cVXYzFPVXvc23Bhxz3DaQMTWloVfPu8ATCXjRCr5y7HoPU8DLT2yXycy5
szPIQF5KVhlaqaEfuq0S/M4ckJNKLhL/iqXaS0q3DRQcdTiFOSjzz96J2oCEdaVUnyw0OH5W41EQ
/1sGfkwuAqsPjbpSVohbdNqlWvZFF+HPUuM/tv418sk/FqHBh/VufOcGhbQTNDahNsb4F+Cp2G3M
lmcKlWBK0Kf17P5PezTEmDvlY8WgZcEeZS+GFQj3LJNClGceC3jbAjbEerwebPZ3suLU98MyMfap
JvBbc8zuqN27WXgUEtgp7OIiTRxD2gN7GHsgIpv2NEweznz4M+kcf9xiGojIn5huz7GfQwSNfd+c
I3fypWxMdOF4CAQEvKhXuQhzPIFp8onPkvIxzQqriEwbTbYi1AAvsDTAFNlbCUn21mKZk1YckwCd
Wl1HYv8N4PfVcpKMS7fWu5v3jjtuAuL9wQEN1hjvzJ8gd1voMPlRYhYOdh73c0ggW5E/XZ4j/aDD
Hds5Wv8L6vE/7qP5tMW/UIwQXypmmSTE+yyJrsKF7CNb3WP8/axEogYobnlQEiDzwzSzqcSiPMbq
fGP/UGVvwJGWwe5K6x8ovazo4VRc46tXhnC91G4aN/6V9hO8+EXqbMM+ZEelyH4mCpxeo9rqfBhK
Yyp9kttp1suk0Kth8m6B5k/Z/MtdRqHwcVg9Rmjpxnhq39Qwgh9BaAw3ixm0zJU+Ci8XttvMjUun
jojpU9o+XujCU/UrHgj7YrdAgsznEQrDDfyVtUH7flXDv/2Pmnj0zMy7fVTHcjUBVqB8BV063k8D
UZsDlKdIoxgICJc7d/6N1W14BAwz7cGf24oarhbIWiVqV80NIo3Ny5UX22ns4MVpvRP+WoCLQmvo
iaeIQDLVZPIEcB4OMmxCU8Xoq7PyiR5yMC2lhuKeMQcmyG0uLMSzk1T0Rfqf6Xbd8dF0Mlmtd3KE
SlgaDZaW5DJiG0Kv4ppK3QYNsXOXfCJLbleCTvLqc6CeNH5uZHAdJFzD3tR6rHe0g+d8g9aegHDU
pLqgT54t6qYxNZkxPrRDIadJwffKmlyDbOUm7To8QK+ftzWIVHH6fSAotRhQm1rGcQmBZfM/16Op
BtBcDmRiIsM9motFF3kjYxNWnCo7N0v+srBJ5Ad37No/V3KMVuALMEwrS4JMZ5GvkFXZHLfoE8OK
7lgQlNh0dUTrW90YmdjAiI0ok7+qVLg3AmPrT3+TB7rpSKflHV5PIOL9drtyIpSCMorXf9gBibtJ
GOSc7QLMn6t/KvXM83WqUJ3o8T//l90eb/gs9UO59zm400MskVLiE9zuVuR7K0HvclwaQg81qLjl
0gVC79d7tOgp3p7vCxbSUH/1IQKGsAMl692u1Bpbnbn5DOUTLfzrXwGsGXVB/9zmvyfrcxbP8fEN
bbTQEj6Mhxn1FyLLdPUI/sJ/SWNNAijk4na04O9aDLPMVGMK9YHeUyfnoxnQfkOKAZ1o7PzrHTfl
eO+gN5HPAxYzrLyc98n0r7NnakwgQBqoIpQ2oFbHzIg7R6Iq67Qfgp/mO5OspjNob1K/CeN58g+h
TkNPabKKtNXqAWw+HEYpAX+5+ICeLstxMU6BeShF1G/USBIw2Fh40On3zZ0aEN+7uv8r5QPSDgIm
F9YT/NQzeNfJLTEHLOg/hx2N5DuHC6ETIZpV/74mSe/WwjO2V/IxsJt9U1RH+6baf1YFUf2F63o5
tgaA9FadWZtM1v08uUoxnOHx6kQC7tzW8K5pZkIjY6tEkQVS1tTWun3FPVyBh4Q8C1dbcp35gEY8
ZhfINVWjKEA/KXsD3L7qY+tuMCpVi2EN9gZAusR0DFbgEOybChQclrWhk36SkFKgiamBVOrvAZTS
TbE1TfJvSBwltaBB8tgJSubkvMGsoe0eSqru0a6A85GBrwQGkLc92YGYKvaixFacDw6aNP8kUY5u
wrMiBZpjgEy9DcMMsdgVh9cb/hMBxdIcbcGq3TrrhqFSSYtMggwTBtXj5pA6c1zUUVNDIipwLNIh
S+Bg7jOQXLBrsieb4quPxT5wqL817cBRLW84z9xtTPPGtJN8+OlPU9OMaErkKbAEoA4DltXK2Is9
3XhMnMDp82dce24gt+X985ctueuMlmu/+Yegex2NBipFS2UrDrD2P+PlwvKDqTtJPHVLzqbvXNA1
E02bseJv4XDZyYp0r9vj9EEtXyQADfIb5nO+OBipZZr8tdsjhnGUnQF8gpoI+htuPeqroAZ9rNYm
0RcjtYU6QEtapl8A08ffj5UgHn2nJ257RZAY8XW7ahcfhukwUYgmIbGOgSuAk7sxVlx7/WxVwS9Z
PVjwPqelqXm2+iYe6dDZwPc+JANjXOwvGlHx+I8ITr1Q1KQALUZNDPb+ABNrtaYySyi/89ZmkRxy
Oe6Q0MOfuC+AVjIGqwmwUw8z1rJrb45a4dB4C/xm8Z9LLO0cSF+Dd6C/2g3H5xhkRF2TivzLA20B
VRILDPLF3GtVBV2yT6nBAc5YawWstEP9qNsoRFrHU/BlidkOZ/Be8wAqnQoviFYHVYc9M4Tlb6Jx
8LNtb2Cru2StZlaUJiSZ3gs4L/ZVqUaLhgo9ZXPtyQFIfYIY4Rwq7bm40oD+P9HuyCUz/X072tmG
scJI59q0MIRsC+z/pUje+1TNABZQ3hMYEtx/2lZ7jVsKIlSl13UuiybaqPaPTKwxz6Aj7VCZUxA0
R24TH4NgyTxbM2+LjiE1hL5JNcWyBGp7NlabM4DLRHOZyj9szjp4ulnlrIJGZSWqKa7sZuf4zfq5
KFgbAs18BSkNYOFM0zynkexGHdM71fuXUwICgp+Ozq2bTWTO4kguTSNgss+bz19iDo17vPwOEPqS
+tkGUqDD3vxFokOOoj39xEJLHzj8ghbmtTpDBWI9BsKrgygBenStxhsD4W7JAPMr8N0Apf6nAbdY
Qah8/R6s1vD9mlvRHHwnRb4XQkzsBdWfhI/mwDHmojmtom/FxmhIadtuR4JQ627XEh9FNBb3HkKn
RnewtWvqUrMdao0HRTE8EcD7iVEJJEbATmccjg7ogJDocgu9qwdZag3v8QiO5uU90p2LX8aI+7/L
iXzYHHJOnLIHhZY5ptl5rVaXD9EPq598jobJrBUHHw28vCZFS49jn7h08r+g1O/bCO/+Q8FwmfMi
9pJ7p3INoYZazUS5fxWqRNtC25RsI994bC7cF+oXCDa25TgOuT9q5t+kvyXhqI7zT+OV7XCPLY9K
OENQwekVBV8+Wza4FP50OeVK5XiXgi3QP5YXrWdwRSKax89oCpsJ+zxzh4DbkEb4Hg0vChcyDb1g
kJehm81Rp5VgV5IlOXfchIK/t1EJxrIN+R88NIn86IJAQd3IToQKHT2O9NnCWLg56BSbgdGLqDMZ
cXD7r1kNGNGp9fhnS9CBUYpcbAwAY7bzNQXZIKZ+hryJ70HVyfFrRLkrOh94RG66P++JJ9IKSCkc
3K+VIVaKoarbWTGtn39xZHtO6m91PaXeXa3rFeLzFXGKDD/xzu6RjfE59AV10RyCEXL39KPgc7Im
I+OYF2w3+3z7qkDdjUgU6s0Rzwx+sD/3/XTFUBu85kGiR2DfIRpl7aNYDKKjmOHL0UfQnOYOHULK
DF/a8CLvIWkzXKSpPFNFKlAzIPzZocRZBwMNMVciS+87z1c2HAtj5WvOI5UH6smm74tqo2eXMld1
UEQYW5au0VPDUhcLjTePL/DZ3sRzxrZB8X+tHeOwYPe+npeOSwV1kt3gUJ0SvYTAvQILKW40clwI
nf7VuGy2GHMorOrAqYLU7xGFUQOZDVG8TkOV4CQYub1Kn4/O6ZMDymkB6vKr0tZPY6R5SHzsdqwZ
FUiky0Pa2M6F9uLZG/4zDNYlREo0wkJ77VVzd+MdKVfS5peUOLOpVCL9QicINTxGRaZiKe49t/v5
WGIAjxVbF55jbCbSpNkPfMh5MUhjuUpjLxZ2UemFGX+lLoqBpStTKwqZHxZm5or0kDBFlkfaoeHf
QuNjQDKswjL78wnNEM82O//xTKWmjklrObpIHlZRvhEzxrm4NGN/nKAxukjNEjOXpRq7CZeRK+A3
Xr0My68T2DoRaWO4dQEt7pHXVwRhsMNIuoCPx0IazKRTyXuP2U2r7e46CkBHd1TvRcCNKU3e0Yzq
gM1iN8OWRTUQx32QFQdQC4VVVoKcTCVAclRisO+6iym8n7p6SrAW7frZpLEUtJAwYZVTMBpJO+DW
phAcScDRV3Yw4moIIewCrJ5E/dWuEYG66l27pL9ibXOhatefWK/MNeMKXI5/1oRWp1Iy5J33jKeL
uCM9I2KDwv0T2tKui9Z+o+u5Qv87c7kRSFrf3BDikI4jOtc0RyEsZ1RaLrG3e9ykF0uLpNLeZav/
hV+cRUtM7iTVdAov6Pq4iw0dtEHD7SnGqmbjyduMnOnwCBleJ5JiXpPqEoC2Uo8xaK9Hgm7CrM3x
2ZCSfJZ5A07lQk+ea3/7Y65qKEQ52Mf2Dvn8x9ZkvogS2Lj3V8jJMzxQRRg4R39Nu/kac6iWRTZ6
Gi0hewAQsA4ybAtvYPNnUBp6C3q/ZIH4j2M8MwS8rpBQ4F57d6dq2GoZYHkCxAvA4qxgrb5Y3mAA
Gj89oXP84a6HHnl3qSFEbpDmpgyZUMDTA40KOO0jft/CoJOh3nGZC0CeSKqKgmvVSsvD5tbxjqPh
87wgt+jxmNbR1zwzApz5IyDSOa0Y/a0UVnZH8mzjvdoDJqYo+gWLqtQH3S32QHAiGi5IX0DCBkWR
JBktgv+mm4/Pv7oI5YQzZKYrlEXOk/S8H5BqO57alfX/BNpgqSnkutrV/3JDeYVzB115CMiDtHT+
LUm8C3onod7WSUgvimA56TRTeO9kLaj3l8G77U2ojs9d27bYcblmTg/yCEtFHi/xKzcDGo5LQqx0
IGJTuyhcYOu4Oj9qQ5B65hIthwQYuv36AzAqS3zckMZRxcp67FiRVb2dqctG4hXP5M61SRcaKBIT
+tQxyUw+k+O8Kh0TtKA9l73VTopRzJEQK3/gDwlB+jb8vfF1LqbZvfKQ2GDgVYd5PcFdk7qfzLUL
mw9I1q5fZP81agsRe1lD8GiXyaDydFn65O+AKB5WfqUTqo55vlM7v9KLQRhDmGku1jpvPYy4TUuH
YryLbROfoTyDGIzegPsdexdFGl6fCoN4XbJT9P4dL56Ylh2tTUzhCVIyJPBBWGRnS/NDn0U6i5Pm
d8JScm0Y6NRTpE56wjwzNHyHj5r4Ke9H3y2RAs7/IjOVHlnvgTmwxEuzrco5tGKPZYFPtqWyDP6B
6pBKI1hp5du2EfiqUpqgahrujJeGmwTnxfAK1eD4azAOK3ODrJ5+xAU2aBMSdtF6saWxK8OdL6Ku
ji5Aa5MViJcWjvqHNqhNAO8u/FopPANBRCNP2z15QE+Z0XJ83HDA615tq4GcIpxMwGIXSRh5XGOe
CylHmFsfhVF3y0IyQi//YMRgRg4PiVXUD1o4FTvhsmdZ4LWhDB2hyIHRj2fzp5zhQn+QJlvat6Va
f37SHnxTzwQ6xB7S7EfNvC9tl7oxH0GVuhnLsCxaAdYLjY/inB3frTnZtwxSlxDjGtOwvcUPx8WX
tjDgCdqBYHly552yvCCZAhV5tip8dXOMaY7RyCm23DZKbr0PpSC2xuPJDb15hfYA3iAEA2rYC2Z6
GERb0fU2mgVkAyVSbauw8ZLdHb7sP/BiSibaWbITRBG9QTlysKTympmUBfifwa0ioLzkEiiakbXM
LdFCM0hXP91HvDleF7XmVWRFN5HT93eOuufYhtB/W1K0iB1YlIsYQXtPMI9HiQn5YEgZvI5q3Efd
6LsEGZ/YsGrbDrZFkJg/gR1GvpywKMiGuDnS30g9KTzF4tzUfVTZ4WcUOa67EuOMBaLixIVFXaeB
obNVOaTfAd/GrvcaE8EMQNg45EY08JhWLHtHAzAVVLhb8s736b5XwoR0R6YATfh52M34kDpv645Y
rRB+bduEx2YAZ/uC9PSzA+5nGBCJLdLNYMHoBe9KkwtaXPUPlKVyYyZBZdbt43TaPUKhtGPaXYM1
eqr2/D7J7Q7dI/yruXHmUXDaT2FMX/22gCrHNsv2qr8zAyKpOZqm2KXy2rXNyIfRylYnA+QT9Qf6
jQhGUoU4CXCFZviYJdXdWXKVlNMHcI5L5GYi0vH333mLJJCNrRmZYs1LCb3di/zDfw0ZB0YhHR7X
PfXvJh4cT+ikZmwQffS35ltxmqxi16sEprh3J1iUR1Wzm50+cmya5z5d8COs6kqB+yKgpkmbdjml
UedavmqYx7BOUSE/ZJEsSLoEmfQKAz8QCq4yG58I3WaWkNc7+MasB8kPKa0XSf4fpqiAf/oO3XiE
NGIXKSLEYWgxf6UwanIQIPXXGS3pq8PRqNSlJo4GicxmnxSWgOip2KqSSeRv5uMUYL3cWkT8P5YI
eGmaedQOaufX5pqP3B0KjtSTFUW/81cGhBuZs/IdVrBra9lc4eypgoREHxQla4HNZG1HPISsmSEL
lInIAu+VrLjYuWCvhjeZgyKoTK+fKlCVdjd32lb8/lEfhIk2bPHWCg7PBGgv5bdxG7hRVnNzfW+U
SIH4LJcIsZ+m3fmgoaEVSRygEcoVVokHhFdipZsYDV8AsFCFvFHO5lQLkyU37FpiQWEAOxiuwxxW
aBA8eZe5m8tdz7oGX9uJhnzHWTW95sc7Uzil53PXELwk2lOFjxsOEmnz9yPnOyYmbTYZUaYi7NrA
maVjU18DfGhSJZfkSnSpGefOlicYDYNuDnHuOZaWyaHnKl/w1SqVfwAXuAEKKBq57n0fuU4gT8zl
5beExnOhx+fJ+WV1ZwX/bvaXsD0sc2dgItE7yuTnxMR16qdyiBEit+sCy2BkOdeoG+oDzrnScT30
X/u+a+LYS+nmhiw5R4S+GyDoXJeERh+h9Qggwzr+YvEb2VgCbJzDRL+GuXjohRe0+rGgQCFrAvqx
D5la7fvIzVxwzqZL6SVMq+HfHUNYsPczAQ3OjXy3CeqbuXW88RN6cgzfkZIRbT8Kl2kWiK181eSZ
XRtBWIBMB6Q9c1vuWnSk03+y04WmAgYvl09zSaQm3ZddE3gsMD7rLZFgXmGbhNNhJLBKFXwvJ1MR
eHaZZMk+UpDs2i4XyGhmNacDhSHX7+70pa3A3n/TUwTnCPlU0HH9/08p5Kw00soSCWsap3EEzp1c
8w0oyGWSTRuektdlvU3MaakcGVqJVDdHbX/DCKMto3iTXlBHakYkdtE4MsQef7B+odqg2JpCiW0t
hskf1cQvy4h3K6g8vsPz+sWrOaF8OGzDoukLhbDITlzLFi2NvLuOKFaAkUXgfC5ZgxsREn/0a265
FAEF/iSCdNqtSJRV5Lzah+PU/tQWOWBHZTQG+XqVLjJEMOjDowOxArg5iqez4eLNuxU/1tgNRYrU
U24pAu9VrcFALEK8snxQ22Sdlx26tRJ3fCDKfDGsRSpMMYK0Cbl9XpWmswg/ZGYI+3H9zs6LYf3S
yQboDjuPfwF9ifQH72t/syfjsvhva0MYjdMe4PLSgDIj9jVyjFoE7rf5gecbrgM9392A4KwsAWFd
SjpflDUKFhSj1e/MnLjzsSVnlKvKvdCITc4m36nkFv0pKDRkz8fftA1F7XUpazQCsH6cLDH/Ff+X
Kri2RLifQzYI+R4yrFynyYwq9S4niQI1TGS8Jpkt4woTl2rmfqyXx8UXvKl7cciToP7tvRRv5AJI
MH60WAz6Z/maPr6h4GdHof+0jxyTkgZe1REOIfb3dpyhV2jFUlN43sUFKlSZdaEQ8m1FsyVwExSq
EcRakb4i/Yastb9IsuOXmOKFhSg/X+l3Xi+mUN1vL2tp+LsCQdZgWUDtJik22YnCsSnvChqGX5fV
c5IHFuRD1NrMNtQ0e5l8BVD2QSgUOaHbGNXDgiE+V7q4F+g/SSuD7Xbrk1RzKwe9lFm8pqZluGOn
X/9lyw4pARhsxcFiM79CLjH4KT9eWhnzzt82giu6u0DkvONT1b9f2PhTNP6rLjfhUPvxTkcfu8fZ
FRmmeCv57t++g+7rev0VbPhI6prk2zGO+KR7gs+R66Rp9PiOFFh5YnEArj8hSNM+mlYJOiA/zCTZ
otA6eRUTSL9nuMXLYfDlNKc/xd1T2c0F+yFTd17vfXkW6JC49ppo8ziOQnhW7qiwfsYb5k1Lqpep
21jhsywgsd3KjqZEijtgUTZ/LtWWHykgXb5Rhwr5SFhcjtT5Y5ENHmblR3fskqs5lrIpyuBaltbz
gTKj+KVYcvgtBzI8Ml6/eY+TCwIwyfBmH/fY8IDSnwSERUe8J1yw0tSOIuQjRRzDrtFfwT+64mw3
1rztAjEMocE4bCLU8P3x+Zj8W4H6KySL0tovT8jMmDLC67kMPDxM7jtPf6gq2RDrZ1fLzC1zjXX2
U0EQiizvU0KWsYTG8z7as3E71GjD8znrsBcnIgqwr1XAKms4/0Rn51d/gAmJGNdH/MjOz032Sb44
AqqlRFAFoITphevKkXEsQ8zi6ao7Otx2fWjuYQYyVtJE8Yw874kSv6s9rjXvuyrcg82t8t+Bzyfj
zc0BapteFjrJBL3Hr+vaWw/EscXPjgYCgsLhiCqCOk+i4DqByHgY3j8fu9evSSHY7SdwVgeX0iqo
o8po6qdWoGOh44cDVU1h/mdi7HZMYJuiK7ECKvT7i6fcY4d+4xfy7qtAx5FMKjMr7wL7F3gFayzA
/6VBamr3tC29PeSd3wTTymGPP9Ma9S1alvQE5/9mNNDoKC1vIw5IzclX1b3K5JpRDK/egLVdvozF
usJzdkXaAsbANhDAcpL9t0hJST1EPa5SVhaPBBVjCVwLoivFzLlo1A3d8QQEhLM34zvPCymtjq8L
FOyiMRDy/18i9JLTKvxVT9yCqyk2CfFUK7wKPvCyULnA4S4EWAB2lBD3z8OWaZ4eD1ZNnfIFz3tR
N5vm3p9s6FeMACJpXoKa5rqZDiXchsKOzoRnKIec/0O/+rgGYNM4+fo9EUKDCFRcS7tvvy0jEsZQ
yX0EXHX2K1ALTiDLWKOmESeLY9lfAhXihxnSQzXLhvcDS1vZiiLU3/Z0lHWNgcbEyV+fFuuzg5i4
glrh13Bud3kZoDL53hr2wAhXfMyJBuQxdfy4GjviKqch29Zvc3SAgDcqZifsWRB68oND4iE+mCp6
0AZ5FgvYIAs3ZEGJT8tL7Q/ZfH7Ebgl1sWNG4/blSDY09M99Yx1/bYslfmQ6OOwBU5CEcBLwZKZ3
NGhO6tMKahb6vKJqCZ01VsGTKKHugEOdh42DQXL9OyO7MZKAhnVm5UE0kS3QusFQ6QwDht+/o60T
aN/mfrOHhePu+TfiEhN/GWVBAC4qqKu9Vf9SmbSLV1vc03IOgpyB6hgXbC2rz1xsYl8yr7Z1lTXH
UmPa89TuXRH6fwENil4sratLls+lyqYJUpKsV656pVVWKPA/Jl9VUDeM7LUMYGscmJgRkJhiJBQK
0waeWvDF6WEm1yaMgQwyGEWRdP2UgC6cp3Jbr1VdNI1Y4QWsD6lbFH5cniNQEoKCaeAhEusvDxoD
ACB2zyH++PDKnRrEGyC7kilSmKCHGUNpfv2rorhhX7ZLQb2o9O8aTQFrJ5uRkJeBQwJ8DdpdbVMB
a51x3NYLq3CTdK+DA2ELkNvYYYDEM0H9jCZnFJV1VhGMzhifX5mSaNlIxfIyIldi0ofi398I2nnm
iqFW98TN1dQv7mKqwmImVMKvfSRAff5sJ/mC58yc92clHyrHFsuziU6OwFaEYdXvuhlynzLt0i4l
XyVgpWzbFHG4Ce7u8yG0FdrSpkhVTWJMcVxgJUA0fEiJJMexH3rIJA96mlkH47jMb/q7jhUr+zWV
6epZQJg963ymOJ7Q0nTmewSwb77NwQVw3pT5pd07C/6i9l1azPb9ZYiYQLhTwJtOjsGiHHzLElzL
QyRHWmXIzWMrUeh4fUmpeeHX+6YNba2/kfObkcSxN9hPjshJD7+1CTbY3kj8ZwYYRN3LhuzxcUUP
TlLfuG+VqDj6Vj1jOrD8kCN5cz2bX6kJT7Fj0okWvzBQKSGHYput/is8YRNE8/W86VGqAleNhlH4
crhW86HQB5VXBDPlGclOFQpU3TdwyTUqGTxmd0mSODu+OwiXsQbiLgoHjLOJ53/bmn/sUPCXwkYx
v+dbIsnRM2/65QDvdh1hHjprcc65egVTN5qiR4rr7w7nYDNPQLSRbH6dkU+LnylygMg8JHAisWFK
YWmIDz/yshNZjDqoNsPDQlQLyulIKSZTeAgR0VzDlku6qd0YjtQ5MJOHG4hl8esHwjQmUg1LH0Qs
tsycY7HkKvAsyrNYX7QjFGXpZDdEJ19dcwwrMQFVUVJO3VAvnuPPVmXHzbvXKfTBgw65GNC4Yqxe
DAcbTgbEBIhrXEDCo5zSg9jP0mvZFHOPAQ0oR0yNdD3qkrasnZxJw7x4npoXEl9zpsYP45ORiaWJ
RCvW9+ytBsNWG7hDKWsFt133hFlDtfagHuglfsEQtxmHFTGENsSyJCSNIbsr0bhjLzUmU/JnaXwq
UkfAu2wOerOJbOaE/uHb3d4FbTs1zZI5ettwBdc98wpzEIGyafxZPrZqW9HJVA245rxJwQFPXYX0
PrNw6f+opuDS8DXJHZ6RR84yBd9U8+p6PreLAwiToTQrHyCfmNljKExICAmrgKhlQHG3j72/t2Q4
1CHTryjz1GEMsaRNVPA3u0cJEAYwLECZLhs9XDMjxucAeZjqldgAz7JTffS/1sAJiH4jKFNh0FNY
oEJ+g86x7qgBq5FH4T4ue0ONfGsbIjTdq/p4XYSuOPiEbYnhV7CUOi70N9VrehUdghUlNwXUKpc2
GN092ce5xkFTKjYPghySy62KtdsVxtaA7E6aHfJ7L2RxcBzzhmmiIYVkdktUBQbLCPwKrRshwjkF
WdvJFshdmGEsYKwxUTRo7ZmqUv26evYQWvzuZ9zWaq5yZD7Trl6qtTEwkXHXspXYSJcOVx2WxjYp
aSOQaK3hwo5PEMBvPo2762AfCI9RgMJpGMbC/PSFcHFYz2qsfbSx3ZOHRFoXFIWYkePwzBUPwXGj
XEBjwLqLp7HQg2rke4QRfISSBmwaYSmmSCDII7M+bxO5xsJlx3gQqSdwUfcsfyxbCuiuagc874KV
6p/4NTeOsZOgz0bbH2ECs/asror1p8MUduG+vzuJCYDVc1c5WSOpBSHPpCmZMPUgIkV8qyiIuLDL
S5Lie7eMX0O9aPkFcWfObEDK+ECsftSD9E+OtJzgWScALmM+Wibtyi5upUlgthwfkE5Yl9BBPAld
RH2p5c8mGFPY10PteyVo1tVocj+KQzdhenOyQIiXDUgSsyQx0L/ScrNe8xTj9RHniw0CZO6OU2e6
FJOW0iPpVVq2P4D+F7m20sgEZfWpjc1hRsEoGWbtrfPWRSzv6gmAFaUC0frNYOPDui7xvEB0FmO3
RdfrQe5P1DDIcqQU1jKrq+Avctqy3jsKxuB0mbIvaJBeaC2j7EDyqpCwAJsYi2dfB9LdDweOI2G3
LdQqnMYK/KGLAl14Scp4ZT4AjLb3Rv8eYLotJj7y8I8OJ54KIssz3mxJsWz3JuWUxB1UtFU4BAyF
qkU0hq6CQ+mrKWP6uzF14Znuqgu/9Mj9pmbI0goIOrvqq9354Pm4Coa0JXsZ3EUD3AVIyZcB/bbG
BWXRtbCFUJUp+vClOAoQbTwLQuI5gcF/v6+paYucXZNxKt9wnWLcxCM8G8zgORmhEqV31xl/J6CQ
aHhGK/OjN6Ok0/U+6ivTMDZo3enbLSkghAVclJb4CDLfGsQABxVdxOSeIGRGtDOUkCuT2xS1tINz
UqnOTVynvgIFXgh1oZV6DrpNO5pd64ELXDo9iyRoMOhvab+VDtK4GBcNWLllMuC9PgbV409yTsL9
1/qoWP4ckD3eVLzquM6/nRrGTcqTYAnNnK1h5d9pyIIY5XMOziG7O7XVT4izWVSyTeh8rC0bkxpB
H5NGWpm1h/5je6wAK5C1WsWjhc2Qcpqksdys8HjRo5ywK0vYkuaGjcJMhIvCPRFjuoToln8+GWgP
myvFW2gWIP4qC06WWLKQA4hZFgsi4uljT/vq4SpWpheNe0dVcRo4QitpcRl2vC3iokrudfD5OiuS
iEzMAaCPa6H1wgwD0b4/7FQYzc/qmUkj/dosoqjqtR3gtvV8n1lKYwaM/ihmdqRdqefu7PPj448k
Ed4xT/7yOfy803GSc9KYsTG3yT/EDLJcLOEG1m+wA7Xh18On11AECd4H4VZdWMHDIYjMHkHBDHuN
GxJTVSSxb+s+zLE5YLZZE50AqvuerUiZFkhTSs55L5ECH4EEvB1LMmNkXgcs5EfE4iBphzWXpZnJ
FPR/U2T8EGcQt9qFjoGsto4oKAj7ZZjLP23yVw87YhWlXoWKhQmpnSLW0XCczbYLpK/sQPtfUiLO
O8nRL/VeBGfz2cWxmVUayL0blZeRvSKpbsq2OiHV2nAwAVgym05avg5OZM1Jh1vnFFroiwdzbXZ6
+nnAvvxYfC7+qqDRbfB7fhYxT9E/KTPuX/REoehd7W5AC7KjB6NpPrrJGtcTOfyCX+/1+mg6dpW9
Uug60Qs1vuxlw3LG7FYrSiLNQmfVUT0+zr6tpSncEV86pcxRp/DJMuU8lmEFF2cvP9b24COhnaTo
TV5qi1wk8UdrM4VGfcOw0SOOjSNXBo8YjU9/nAdopLbVYd3k2r3rHXn6gvRQZ08ZKkZ4aykxbC1S
jUilT46UPFU/+0rSYln5bborQmTXsadxhW9bxkfui6+r/6ECvCnpaJ4nVpMJxN1nZpRwqBAF2STG
9LHG/4zHdG7nJE566f4mLEfI4bs0p+UaJMLLepJ/iHCEbluoVSuiPDXJo2us45dIzKs9fm842Jnb
nYRo6NyB1/ObTWKjC5iQLRUbsjf3KnP9Eie68yRNEcUiJJrWugK9s3AAq/PVZR7OaEA9wZP21QOE
+xDky7m/b3B+UN2LJ9lq7fkwtMTSN/TadbwZDBs7RnctkF8bbgpz0Od2IcuQIHrWC98IRCq04GoI
zz+WDUS19C136N3dLGG9IAeAbxPfELyH1lw5riQ2HoEbdFcIIXYCcQ7bcCnid8pL9JR6vICTvuyM
5PkJvHz+ECnE1BbUvPNi5TSqKhloU0oPYUDl12agubXtd0dIqFO17Q8wuvU6fRFUTxdxg2s8hXPN
eBILafvfXt+94TIGGmf1QbP0XkVnNfRkYE+sW8Ps1TM0FZaNAT6Tu6GZtSl8u3tKOYBmKf/WCOAD
QdUI3pRN4mQ76LMcFa58NmOzV1Mb73PXjGEaxeN48JBEb+FVI4NduCabCvs+Y2abr1X0ZcwSnA+Y
90bQ32Nq1yEC1tdFgFZCLKHjWyKT7b5pF4RHmg3mPk0liNSHZIO4Ov8lWoKx2e7PPrBoG+QekSpe
Dksg2s+WkxwP7+cNf917G6Ek96Wz0AACUNBY4/yY87+1jftdhUtWm+yhE+YKTV5bnmLXU9eN5QnT
D4AldyOGKBaG3u1ncFHoOg+pX69hV2U3Q2glR06WfrIyZDeZ2lEwvmFl92OD6rFEuUjJTxYbYz62
DomQVdaSCUkxdIuTKbRyB/wcUGbUOyRTN/ocC6RIVr5BGfJ+elbQWVIvvYP8BMVDL1NFUKCKR2qJ
PS4Y2pUb+JXCvU5IXIngoVtiwQjhA5KA/Mnn3I5zEy4+bB9y++YJFUrFisfQQthUP8wMjczAHjzN
BHSwLdtGWCAl8oskTWh351yheaHbsutqONy1t+RapL+wu2pevO26HxJqP6b8hF6t+r9Dchy/sfPF
6ElR4dpe0QxDslgYC0Vrj5H7sArP8O9RIlwuiI9GXd6G5PQXJbvlMaNwIi1mro9TAyZFc1qA/bSq
otOmwJgmlUfObFdWUzWceRuer5scE7gxwIoU6vzwo2HmVUqNegJzHYBW5pkLxc3nccdo5GVz/2RO
jLMmExTZweTse+thstmk8fVm9MPGrE3MNPpTSsjb3gZbozLmcNEk9Ykassccey44A7LWY7aLR0Hb
XYTmZiKqSxsRIVRE4NQZagnoj7tmyG+TaYpO6iHlcT6ICrXMKK/XXIsSitq7uck9ePwLMpcaf2Bb
c71pWOZzVwjtuWBuUgOioV9b8eB1EXzGkYssvMbil4L3x4yHdvi2X4Pyjni1wmYnzmV2Zm43hXIB
sa5zPHHn0CUOW470ZQ1Ld6stxetfbMqfC9kIkz7SvBe6c4pBD79IU6v9lro6vh+NKVCqQgFHbYx+
/e8pYbt3FhuLNwXq9qgq/62nn/qjhnoVEz/T6wv13FA5mkM8aTvbKM0iyvpbolF/aMBUjJI9kOp5
lKpkFmRE7MKPNeAQrRWNPzfXz0jJCERVXQOzN7xv4aBZWSNWj4Efc8uQmvAB1HYpbKBWPMEA8siF
vOjY7dZpVmog4a1fbW1p4MyDVMQKBWiiKYQ/CRUdi+ti1BmgX+ieDLgSjV4dEeNH7Cycuyc0h9pX
qB5s79HEbcrxmsmrpgyXQdFfZ2eEi0AxtFF8dqcGbBjt4thmAA1cHJmVrF9TElHrbFP5DAIcZkQY
hEyMaY81r7nmCZxPr77r8/La5QiZiX1l6Hn6QjPK0OhHfsbTQIpouaKfcbU9dDanB7NYEYO29n5i
bUi6UsBJoggcYQX6V6Wt0TI8C0u2bjMxKq846juqAOyqod6bkFaf1/+lqYGAzNJMA8Ij1WJzH8hX
IJFVXDQiJKa0qFYOZGBjLgKeUHqwlNhQT8MohuAQws6gRQrRpz2YlsSOjiR88UQaaNRTggQwfBv+
82XuWQrscG9X/fqCDdIPPmdpGjBDYXu1SkR89tAJloH5drMvwhFrCUHC69Gh722F8nfr700kIW9A
JspXlXKedwMVBuQoxC82PkE8OoeRUNX8HQcnxSqxMsUA7M6jmk56YOxnvsVhkcFmvC1/6rAQ+Oe4
SlMizPOvxRpcoS7cM5JTNucE1naeXtuaEpQu3h+tNeoGIqR7Wn6qLzWvHtXFJA+p+dWz5mgLaj8G
qQji8w94S2uwyujGlM62bVoghrPdTLe0uArcvaCf56A1HidOiRiB4NHFHbqTQzQn/4VTzCLMEaP+
sXrI7GLRTZahrUbWB+Qd8WvCf9opk13B8nbIMWrfA4pjd9HkNGEmn1aF1GR7R3/gBuF/Ii2uNCtL
10I1+grYgAwu9tE/JV5DIHL5uC7rapIHUjZsDY+w3G/HbhrvJZAE3+jeAYfGAaqB1+oqI/VNCwlS
7RFN3HseYIPHJomlBxjvsRWKi65P/BIfb84ECfso34ZKWVuN5GP46AYDWjoS1ooRzaOosQavdSgm
ZWxhnu5g7Q462QBg75y87s6DKcbtdUKi6UEqvP+krpwWLxrUgFdy4NlO3ry9wjy0/XE5HeQbOtd2
dzpfygAykisjJYQ65EDSog6+EBgWCeoW30aNa/paDNEUbHSyIiySTHRfXd2E8wLTIt6M5jqYhOMQ
GA3CMwAnPMAXY6M3xHdCMbV3mjxnVnzuzs2dYfseohjnVocKFTLuVTXujysVZgNwE2I8ObfTOQf2
lDhwYHOLySXn2XY/OF3UZdqE2H3VT/X2MWEFewAr+L6GdTA46agI2qL/Uh78mUR23aEaLY1cG/Cx
zJRXhEPR9U6L2ONaR2UpyszeuHThIazazHWD/0jPufAOspZNKK25k8JFn+UyJ1uN89MpPGTw3BIt
+hmyKxZI5d5ZfUPMV/ua2hkDWT1O5jHDKDhZs3c1l55+4G7FaCOsDAB8PbL37LbSnIM7fmU9wKWh
66qsvr7iWuIWgHtXjwykKQT6Rrl6Yd7k0CGhw/5/3j5toC5GtFAXCohA9q98WKjJbzOfQMv3iTRr
uTQx+w8jPsRu5Z/YAPwbv67qB40OIFOIX2wuKhSmaVFj9U6ltGJKQ9vuoMrjaq1ECTxM9Q/C/ecC
gW+4rKTx8HoSnlZEw0xVbUAhmft1Myt3YS+eC/T0+UloT69M6w5owVQGroON2v73XbO9iLb8PqBK
82HpfHTV3jhwNnJco6lA8cgU3VrXE5Ar8BmmDflRWYXSkVzrNzx0J6I2MQQ9+KgyAgtIy8sKYmJN
+G4EXvSB3fU76sw+DmcKEBOvLa1LoSQMzsJaHD8PGV0gq/5a7ocZq1oL6yv2oTM92LcVZzno9VHH
Xzz6gWFSxsKKCVdXlPN1j82SBkp1eYIEi7cGSnkYacdqvPoFigQAnrOcoGAfU0GaXF1T3UC1/L+/
Oy7TcJEK+zzKE2kga2Y4hT7SlC7tL0L2yPSuz04JZmcqhczJiSTe9UzBPEch1Ii9jyyPtWbgjCyB
TnyHHD2xBBHAEejJvhlCydnHkoDy5b9hHvHKJEBzFNycTpmaMcmX3JESDcaj5zHp6/hlkeY4nPBT
FRcGFSBDtMls4t9JDhVydArjwgQsaYs52HF0g4YhsOnxGdqVpmbHHSUpNTO5DE+vrLqQ68GIg6Gc
YhowZ5UUkxZsIFgoTKB/tOmoUu7LzRBVR1gjNydYAkxHBJry0NbdnydgZXOVCXmhFZIK69PDj5tu
/MhaKke0NB5p9spTLPxVqDPaa7MMLS/CPV+iiHuzKLxckGco+w5B8wYnN558qeO6wqiAbintDk87
FlSWpnvQk1VSys1shQUHbfB01LV43hvJ9qQe9h3TWxL6vOJyqFDpv9bv9GRfT1Xi64p/nrh5PB+y
TLloFHWNmioFEi17h/frK+lYEBoPRND78UU9Fxk7DQ7uzaiTrX0q1AD6qYhhOIeBLvWczAHO7fAH
dhKMF2Mgx8VfsX3Pxqmv9OS3H/oHwIPJNp4RWWnwJCZ8yiUVBOCwDDrdUAjMWTp8pClyQxzAEl0L
4+vepUwGoSJqG5YQes44VocUeYhXY76qTvmXd5ueZR3ee6Ym+EoajKdUraiH3wqzvLfT+kzdswze
RdXmQ60vU/fLKkgVlJGQTWd/1JIN+4V2GPFOOjRwndwG8a7pUvRSST74wLUSlHzLJ3q2WA9a4qiE
nefqMh2NjVXHWapN1PuFHso4k0zFgQZDMAjxzmGkxEPJN6nOsTHHGRSyOZRSeUKyGIVWB2PIJf83
aIOvixKV+KN+ZKcp0POj82YEebuBf+a6t0LLnZc0nXhXMeNMLRuO/3k+f+Y5ef15r282jkLUVPY3
9xbBTiaGnwb+NtvrqRwvCO9JAqQ8c5FQe0UjqZVOzjw9m62heVJOJ5br55ejsWHNTtGgdwdPY5k8
2DQEzi0IuPLWb4kctVJvGTgm9kXJ0bqI5W5T6ItxNADy/VY6rvGenlRr5gDtIfIfGp30dqgj3VSG
JnD9hlxntoxUbLbMcWXLrIvr7n6jIIKhrUN2uRSRu6GcDdIYtpLoMumKS28Gz5TR14FdZjwkS1eZ
Gi8HFuidoDyX2eHY4jiUjJhhEO5ghkhBiknfCnNPIl3GwqJ2fWWT2kw9LKwJpIPSmIUSXAnBb2BT
ICvsfMOM/IiQBWyBUGR5FcyMaeI9SVslaLfVrn9+OHmqHkCJs0qd1urgOMUrE8phR1TCktf/LdWM
JZRIoz/XtSGroUs3gtWl3/2C0maqGSoGGH+Mlhj7b3Kb8nL/R73G41eXCrKvkf0xQ9iOuUcHDNtm
X5ZJL7f5jWbfBr5x1MOVSuPz/QgIBT7eh+flwN1QBYw5HFSCpmd17k7vYff8/z+hmi9HzGhCdnS5
NLglt+OhIDmyyUbDmORycZLSwibBjypePigblJCRJJ0tjUvLOHI6I3rtTTNYknFQan9u1+sMGqeB
5yOyIRMORXKTGhCLkPXj8cnUXRnjc2JP5FLDg4zdfwqRE+Rg+S1KrJn7Z7ywc8FXAPHQOuIroOBm
WifJZ6BHDbOyKRXRn9Vrz96yS3eR0hcgvr88VbJEprbZ+oAaPZ/3PtubzHMAZ95j8VElIZ5WqSRl
9UedFefHFPgE4u8lhtm+avJG8zcjWDE2+pogD7dlohjc0ZiXKQWHTvvdfvIfSIZhNszrCUJ2HUw1
K5i4nP89U0ogVfaceVbYeTXuI+6jEOh9TSloZfKWg6q4fPULyDsqFbzqT0mzzF9xTH0cVRHZ9QCP
hO3oTLhGjcLyI3THCo5ahYllbxjYtAYgtWA+Ybli48ZYXLjOXBMJODJVDOLYhXEfv14cQdLspB90
nwhpTzF4zlQjScC4dPieZOh/r5wKshf3HYxJY/EW/P4rVm16Rc4GI4t+XtmGSe9iMfKdZ41GWez2
teiVz99xINlURkpi5sRmDJ/9XzWLAbmfjTWCdl+Vzzj+oDnWi8TVPFT7D+YzwunrZSeZZhNbPThN
w4I91DWWZTlxhwUHoY0kY704Y0QJdO1PJleS1n7btbqrf+6ZOaFcZkWPO5nQm7ON/PZMcD/OV0+9
f81mxCYg5TwIdinUL2QA27w7So+4Yva+B3heUE192p6TZ8rj4Dec1Ucg5ZbTzkuOtzdHPIxheZFK
x8zATnOrovsWVw7Lkrt7hF976M3OkfqxPEnIaj0Zg3Yzn161Pt1GP5+sZxg3aLsXnxlbZ9ZMfcAH
wx0SW9+JyPb4myRvGl/hKYh32c0oFIPLTHQj/wzcy4HGJ43Av96X9dwO1l/L3F0vAhArpiCPEJ+E
Pnbu9eKDPUH653ahQ/0ewnSDzl+T/YRwdgTjz7pfmP/qoIZsFNpwrtBgO80C/6alIH4xUEKcI0Qo
znh0+j9ugW1oJKSGLXFxpf4YJuj0bSawo9edUogF+Omf+aBPGaSH33PTuTt3v1abGbjav+gprvgk
CqKiBc8bAmsn8Zj6gNwVHFryIACEO8U2AdvW1PNbKk0Psa5mnau6nJ4mc0hJMrfqV7xRZpjhmPEO
NmsdDkjXwTg/WMfFfS1x1nIiMVdyvIO7xnIFYBBnX33X6sPG6AjlS5QAfSr69qONedrfYSxcq4Sl
KyBg0Kh2lkiuV+QLC680Wzh5/q9DW+BD7sxtUaqGwnhjzT3pyd3UrscGDRtzVLXS5NukWeAvFGRr
/sE/v0xqfbHxQ49mXtBRzrU5T1Qn60d1aW4mtjkt36X3qvKydlAaulDQ06DhOC49K1N+YsTzlbcQ
f5AmMbMqUXKQjinCCrUtEAnI3lnKle9CuSbiYBS7YPH4G+krjIM4/8WlOgrZGVRH3eAk5fIEZ52n
B2aluwd0D14ui8Nt2VMh5ZE6+19WqIXRpEbd9s6RgkC+rChKyEAwMu8bOQhxSyieQeZ+thNJgq5g
gaLWqsEsDY1R6W9aZff81ZMcHE6kp4T5gBwE4e/1iYbNINZuRUaZ1tauLg2k3ed0+fw8sby1/AJT
n+3YF4oerHBtRViiXvq/enD9FN4erDjCgR1+nIV6slX5yDIZEhNcOP1z4XKa7Gs/yJqRLLb9o+yN
FrY1SSGg7DDcNW83NbieqSyt7gLO4BsUE73NUmjWxijm60NsZvlldhZfj64QGmbYR3QGIR50v8s2
mj5wuh8+2aSbM0nrTWGIhQNxOmL2zPAThNkOXyQFo/AEs4JvEyIjxQDeZtW75IwhjmI8c1zlq/Wf
23e0WD7nnlw5CQ/NkJNXuS3Nl7hmFVdMjzZiqkz3a2AcqbHR9lom/0hY+mDrIgdM1hNQG9KFG4Ct
y23wEYPYiNdV6c3cbSpc4GF9BwJMEn81sOanjAR0eQU/72ganWh6eQLop8qnJnPX0Sd8F/gG4WQk
aQO6iTXemSXUnvCv7W6fIk1TWx9XuT/m01eOvppzw850zQHmX9OGONykhI040/leH5IYbT0yEMr5
wf8KsXPZgGGscJ5VIx0VKiBVSRwHiTiqgzO3Q0t2HLbKJWX3koR1lkOO5Bus0PCw3g4vwhCNI3uY
x/1JLz3qDRS//zeXigDiVQA3CM7oQDU19abR72QqfMTmbIukZaLGvAvGRnrLs6LadRx1nQTljSnI
gMSzk5ZbdWcxdPfSXwqHlK6W8enctYiLo3UdPvXg/8S6fcMcOAjOL35Kpg5yKusCeRayQdVlEmXz
uIiLtC1fPGk/BBWWLYTAojKZCgezCEGie37G36wmUanczqf6dbWKO5apaopRt8GFp1lMBJIZB8HX
yQFJxFchoU2gAHIZ8ajtQ+54BCT+5rWUGvNTGZa3L6nJtwxB/YMmSfCd0WWAZ8ryrmTAbsmDnKd8
dfZJCrxP8t8kORRti1uCVU7BOMapJkJqCyUTQViDhSDkvT9scvPULACF9uU2EuxbTpB41ROPnM4J
J0iuKyqfHFK8HUDpZjxmI92q2Qtj6ZZ3LP1uKXuWi05+rG7tdjudhYiBWMgzyRpl6bpawyw+1VdL
0hhPCHJSFIj4mtz9r0/Xb9t5XEfLELo//A7/NUhBAzJeZxwUUPmVrNLhuRt5cJc87GgfIsXIpLxC
2At7mnjUGjouNO07eUmNBpIiDs5w4zLVKaesfwPTeDSn/Yl3bl4K3UUJmryLl1xYZjJR8GOgTnv3
WPbR04AwH2Z4cziGQ4rJHWWeJ3ts4ORNsmkpjzKfWnebWwiOELT5i7GEJWoInuJLQJHxvzuadVgy
y7IAmKO60H5zYnVN6624N3fixfMq02VDGxpAc+MxTL7DbBRiLLgYk5GtC22ErEgwTGgOGkUvfP2a
KyXqu6XyxBOD9ZS7yIMEKNVa/HhIsoXwoaXD1qXpGOh5J7xr5qG6V7BR2qR2naEdysvRqTJf0Hh+
F2E1lb/XIzHrDw0bkW3BRZoQG2ULwYV7i2cd6x9ilkas54kfEbx/6qVJzwrd9EaVzKDiTyRLji5E
S0Lup05I8kITAXuIljlE6483dxjILm5uaZy9TtcUgbtxwZeUJCAaPVV1FlOBMQrqhinXZq45vGvw
3NdqLQgPhHGyYhttRMpiZ6cbyDctZ9BQc3orpfUo9tYpQ8qfIffPjg9MK2J0RYCIcdGA5qpLWP0a
mkwbF0oPcP2revolKWqn2UB1cANlbh0DUeYg4R0R2WirIKiLAeUef3bYTdjbVoU6Wu0DxPBvIvtS
cPl1cTC5BKCDYT4t90887/Vpk1BvkjyOVitSnahBNJhG+vEk4AZt9fpH6c3MOs5tzc8cCVzt/J3l
jxZ8ZKXaI2nMxhJ246AfPUkG2bmcy037NYOa7GTkzLO1l2ST4vA44LOVPO85yvyew1bpiCdL1SI0
91aBe1QtIjwGo3NVcBWba4MRRrDxaRkYEfi7zKPOPCXC0KFrQiW+XKTMPIHtVN/1J5PUEFKOgk3o
JcK8P2zrM5KWBmiSjL1tcSPc67vznXY0SAO7N/CsVHdtdiMK/lGJ1+hNm7cVAVHKexEd6aswZ8CB
woJNOBab4MxXBxCJjWpnhO3p+i0SXVkjuyt62IEyAcw4nnBfqm39qkIs63uU/BvfveVaxO0L+jPZ
A0WRft5qXZVThoZVDgjEcdDrlrESLY0DlPmUJ/IgmgvEstT6sDt+0vikQeMIVErzlfC0IuFOdARv
L4lW8JHogieBb6vzNcmfMJkkiQbgYiNT3E9lQrGLP8TjiCjW/aXjo+2jpbjJmpDtztTWANNvktYn
FL/8AGoSsLqit4ZyihllMkRZQt9ZFtxFYTKUCSyKWeF7s3rYI/0k50TaVPeTOQ393vGLu/rg6D6p
WN9pz6BkXejuBH1YmRg9zE38T95cKkQKNXsaJqd2KXWt7VWgztDxxkSoFeD2tnhe9WqpAzb0hjtY
KGeFn5znynu8NksQHZfzOYQkmaRQ0Y9fUnHqxG0b9iSeQ/5IvibMvv0hifo8S97biNds8GyDo+JU
5IAjbz4Fr3zmyqTEKtBXY5yJcOk5szeMM2ddkrjdv8mpYvqB9hhFwMLENAk+5dtseNyMAm1Wd4Eg
KzTbpLncGUyRL/tIb1NJVbysZ26ZlZdWFZZhNq6Y7aTScZVFIOjivVw7mniAaapVzs8Bs5Mx2SnU
2WEbD+FlZL7ZPJyYm174PrIndtPeqL6OuyWCOaYhJ8GXam1D5bMBTINMhPU1tWeyu0XUqWWjSdnj
A9squJKkuUkINDRCVQxioWm4qEFnlXxOzrQmXQCfwf0vymKEtthnjGHp45K+QP1Xuu6UcTHTcPGl
C5HnqPihHMKfGkx8VDXXCNnWbLE7GDN+oOLkwozYn5ackjtM7NUi102VF7rg6f8SUNNUiIQ9Z3WS
Jpv6DE1EWihAiKBg7jaaaIoilN4AlIu3cRy/ph9qrBBcZP2ATcvwXt/5TaEdUK8jyZ/NwYABvfDx
++z9l29gOr2D7nOwggcUmcPWFgVoyn+kLfMl9kFa2HH/XM0qTMSeX4xBGa+1usigqp6L+5duyAM+
506uuPr2dmtNo5y7tlQbtZv8W9SPz5q9WT34BZTXCaI2vPF+cmSmBVotr3woq0PuyRQb+MOwnotJ
rdUPnw/ydJi2e0pKJaiNfkWnxsZ5MbswngajmCgUP8Zr9MLsXRuoJ22QFSjzHy4kP4t1vqPYA+Ly
1ehYn9PYMLesX38dF+6g6J6spjnxU+2CQ0dimmqjTeZwgmtB9cii2eRrj6PWHagbEg5I9BPzIaXS
vEvREos6LwS6Yq1+1fwKmHyDaf1IvOMMqfxnHt2KYsYCzH63U8R3Y+RXu0Ifm3Ms/ct+w+a3l3uo
51gjh96YgYik+/ku1HzO1yUjAO69p3y+OzdvohnSli3t5MhFN2naaRdo99WMsuVpe3bfDmFn5dMb
EvCqgDY3z6m1t7M7cdJA8jf+mCt07jQfxBm4haM8d+bsQfkn5XId/W1iQJT47SFN19iYs7z2/9z5
ecPnET6A+iIlz32QB1cehd4snUZswtCVNlk8LHgdKLAjU9M6rWpk/Pgxm+i3SicLYzZRKvGTJ+gX
4kHfvSYkt3Wu8J+RqVFCd8MOtdFTFrDXigaOOiRGqk+UV4izu4MP91a2XvwvdINtWYmUeoc43wB/
c/exqk3RchrFQzilK5G8F+aUpb2O/sg49f8zmlfovzr33lt+YDQab2AqnHq745rG/OnYu/iJmoNe
1JdQQ0nQFgovGPjAK9RX1+f+A7q6Wr6KwTAvbTvzkPbum+/lknvefbe/S49I9Opu3dJztK2V0do/
BT0sg3tAUoCY3YJGd/D+F/A/yVJChvYYFQCviLrjsVpzuNwBM3byevYNjKOEEBPGY4ZbdqGsu7Cg
Cpp3JeB8XcMBDxVItMMPzclvfYd2Ye5DEEk1mk4lH/zylyQYt7E/NeJXaZKi7Sgt4jlgo1yeik7m
51Ai329qiT6LLbvKtqzqkK1rBoZNFUSPWJataayvBKqJXbdyDoNoYrFI1e5ub+vgTyomRGhis3NC
LU97uB9blsugtFAmeGD7Ar3h51dihvwWa4y4/nWwsv2IGu8+VDqu804V+t12/nF40VMslvqPHBk7
A3vaj2NNCn8wA3p3WCeYSAn4wvqAYpv4cB5uv29ucAmNZXONscpjVdv6rghx7KYkONGfQXpr8QzK
1u0VMe16obxxPuxo4I9gUYPHw6Ti9DYEyjvYSIsVBeGifKwvKMJRY+QjiQhkNEpU+v4TusUbV6D2
e/rFmycnGCpz+x8j7qUwZJGOFTb+/t8EeX7vf7tzez/tJ6wjnHxFKfq7Pqhw1lC0kz+fRYwGb9Zg
kfbbnhet3vzHtoMWvJmCcasuOOEqrSzFxpKgg5Kt8AQgHAqpb6VYgXkDpGGobg3DVqOaixUIRmoS
QEfk4EIZRPr60awxAljxMRtyyYlf95wyXwKG9EG7RBnMIMjXRY0zufl15nH0qMcbNsHy8voR/Rsk
0lD4crojAJAJQJaqKx8yZBMi4SjZYqJ2I9vbDZeLT0NFmcVoAKqtu/93kfyjAQ1ftEBqz2avcktz
XUPWtfCBZhdxNnLg0i2qnJ3PF+XJpCY3VFQiGGbtEPCMLac6s4vpcHdRGtOAIQEudYmKuWn7cQ97
qXuDVVOUfL3FOMGmNenPkLKGPZFi5aLbtBQYYTyahglCTk8EY8MKc2sExbf11aELttfxvSzLUEt5
ZhIHq/JNzgg0obglVQTuUv55dwEfHkFd5lGk+c8PzykEze2/9r/xoVfOJv9bdwcJuwqj9JZ/2iqY
5EAZEylCZaZEniW7U/yoSnYvX/S015CNYsBGuIObYSygxq9gs9hcAMLEEcW9IVbqyFG9IAScXThL
KZ1gSs9hey6bD7X6sOSYawIi7YLg8NvLCfCRU1yh5kYDHEveqFChtMfmFZ5xXQeaNy2VvVa3YC7Z
RiWboT11KuscAFdZQ2bKX8MggW4UZ6TzuoQ43QShjJnowFQYlEWBSxXTimpcPWvfMD2j3052KTwL
VLelPWlgXXBHuHApj0J4katXDjok0OLZXxZdIb+Yck4c773mLi3uv8oX9EaGeXJY6Ja1ujwePvRU
5424M7XM3izdZVI7Jx3Yu2z6qCEmNKF5fy0NIwYeCBlb/g35Y8heUwnZ0ONX8iy/B3JR5NhV7RAn
8F3K43Eupv+YUFkf2AHFDnLU0vHfSjZGqN11bKEgBQ/0fI2aKABIQ8mAGmDgz6F2qvWDGxEBB5CO
3ZwkIU2SGAKDo+PuCXipVWFGWMXvO9735XeO6frQipFMArcI5J4AFN0hHrt5S6lcqgc8Qupmojx0
x+7ciuMhuENKNmapbfAqvxD/SIQaOZU//QCz6gmsZRGF93FSNZCqaGAfPf4HYQx2JWvGMMmfKTHb
dQzLsgd3ZHdIUPJVLDKJgNNhMXJzLcfwYjJKh8e/V8xvZBV/WSisUHdDr7hXRaR5IOpt8jo8zmx8
KMln3yHBteXPKalkr/XtDgMfHo8yBrMaVlZLs07rbHn7pvO66fJ/dAj8bINtrv7kzBqKOGdDYr8r
6Y096EjC3ENC+o+Vhqn1Ii2BGdbS8cjlGwBWgTUvVJBrdrnZfnDaLVrHmwu81gB0JLppCXoY4c/O
ipryioYaIf+dccQY5wFEu1MF65EzKdC7MQ6s7Q4gY7w9MWZInW/Kc8JnQlGRKNWsOH94uZN0iHod
+2YMWypHybY6fQ0fpa45Ko64fIm0BDfz6DCo34xrok+sX5k1kC9ZFdSuYrMjCb1h/Vh34RgpN5Nx
SmPGEp6b7ZCZKdTulkIQVkJpIaUahY3s9c/WXHgg14FpSUpgyE/QEzLUtwGZw4wdyex1N0knLaUa
/gkRFDMi5E9etMmzhE++hjQiMDZLxG1cUjpT6Tzw/VbgHgzb5I0njUhq+9Yoo3yaeu8RmxmPjSyg
Fu6Pc6BNoH7gUj8BJhg+vEOn8WncQxdS2l5nPw1dY8njGYEuMBvYS/tYPL+wSJGbf5CS587UybKU
NrQCjXbM288CuyqPY1ccovk7DXYDxMF/fEOrIdxRB0d1TtaThfjfeiG2mND8Daq75IyStIbKcUs/
pA4s+Ojgm4YiunDurf8E53NkpiOdoGfXn6oV54Te2UWlVvhYjGfGM/uOWoSg01AHJJf0h5qze5uz
WB3BeQqxzb70gv8wMPjyL153nvjeDHQs2BtAxmsnDqnxltT98lsx0j77RWqwnEJVDUte9tUF1sKV
azKYqZGqzjSJaIiEnUWD63T1GtaXw89hQbq1ouXN8OdmnY9oPCstmas/aILUfA3IFBzw7uHEEkbT
DHWNlg9jyVQpuajJtk7jkOYNQhOy5FGqINisFAk0ZT8NjLwUw2nLr/x5nj3wMzqB4lx7tpHE7sDR
bqVg6JgiMXJEDzkBLWE2eMkdP6xArmG1YDqp2sAzcbIQEi4pZn/dU38UtHANiu67RY2B/0tzxwZG
5nHaTxn6kNJ6afQG8O+aO48jfYjl3n2Oe0QqKr2K0w8ebZyTQcdhOalzxVMMAw12LtbQUZ/muFP+
8sGjmHSyc47HK0c6uz94n1mGIo7Yt5oAI0wNoytqQI4OXufDq74OuL0fF4LqlXJJHF0/k/JZQKIj
0cHqglV/3mYn3M8c63DzGdGKqidTJcj7uIhY47T5m3Gz4nyJxJjiq/y6cSYALQxMl1X1WgIyLfn0
K059Nw3h+L+9sDNV3m4iWiHOkOfDFsQsxbcKSBTYUbeYmZDlkh26G0FGX2Cpg1YwPqpSDSecVvrb
sbYWHm20HnPDrNpXBvJ0LSLgKre241rwkbfWGNpPev1bcbFmj/m8PKHl41ipMzARkiuie99PiHdu
nKvPEo5xRuE/OD9PiLpk853+I5NJJKu/++kS64iI8sdDziZrNRO+Mw7VTlicIClYpJDZjKVW7mYA
JUaVPUPZE73xLeKDWz8tkxj2R/7ddGk/qWQrKOVgOW1ftfTjWpNfAhBFElKoR19KLTXYEG2akus5
Sq1mwWEAN6zpn+C9/kDAz+0sjNDFSj3CSk+A0Dz2JFW5svDpBwDcN8Nd+LE3A9WRTkh1nisAfQys
Wtyb8grJH+99DTwI2JPWj+h5G1iZKkbi1wTX1IlT8gPPaYZukfqshHPMJE6HfcjU+axuQ1E0ff29
SwcM9YiEnTPxcvnrkskjoMzxH7es0C43D1b3ZtQH9P/RCkMVi6bkpqtdktaeKD4fkP1yt67xjtsm
GFkJEeulZKpfn4aRIzn7zCyIp/dts55tyZSHb4TW2WWvvHl8LA4jgmWhwAOqiWObtPyxQK3L34PM
5NssQYacjS06KtzXcoCkuY1jxjX/2Uk0QlHcCkOJLdF+dS+Pc8JEFLFlWn9qGb3Lr724Ye5LGJcO
80FR/KEg96yQBvMjPAfR6f4FSHVyCeM7OVAzlX5yGfmEHIlgb/3YI+DXk9VJBlikfAeN84Z8cV8n
K6Z5853Hoz794DRTj3kYWa3Op9YYFhn+kLaFPV/GVSZtxzNbmiJVdhYNYjR7kbi3Y+PklnpkFEct
8tVyrwmXLgJLxWp0U6XfwsHlR/9XTKdzaw8km34qFuSOtxGumxNOWB+S1oWI/fvZocMCGVPQG0k4
qdWgakw732/5Gar80XIl9ltQcgsxj1NRciu0PUc64GI6jGiWKpmFe00XqEw7SOjS40am+N6Uv+9Z
F4oOsz11+Yfw+NtrjNOme4CepoHhJRofem0M+1V3Sb48gNcBYCPP75UWVr1LGoeEUS9tQjMc2hZc
54PY/RqgHsbsV4Idq3Vu6uOfHlzd7z4QjWUWP5l4Al8z5YXG9nusKidvvDmUoqyShOFxC8pOdtbM
abf4+J9ognoU/MOMdE1QXUKxTSKD9bmgnT7KjRm2KsYA13SH7hl1wdnGyBQrJ3I7k61AjxoOqaf1
8Qd8uBfWv5NdUEuISPNWBd62RAHZ7R++fT/w9qjSPVlW4nH3M1LyyZzN7XbPLEyYEzzOM0yufZWZ
ple2dEDw7iL+foB5+gyh2LDbVjSIL8bD3wN5zBnQ8PeyyKC7KhaFHxUzNbquepQYYZnpDtrpbXxk
gmkA8Zg4H2FWZgUokokEScSjk+T7BKGOZUFGqbcP1ldp9nBmvQlsV+/uY/lUxRREQX7R9rGycB4o
vN3UBLNs50MHflIb2KYEjkBElp+Pv9Wvxr8evmEqN5FwgOZ+jL7D0vQzrY9mXukC658SDIiW1oLQ
YKCAvIPBKiEefd3oG4dci2vuYbSg4SCPGUVadO3VET6kJK1Lrkw1uYuaNX7CWmpqjCPDfFXHFEql
fHY9+SGdq2N3GLGpL0XbYqAt0jx+OcZYDCyNq5/LF1vkUKViDrfqodo5QdppI+bnj6ruuZ7pA1QA
x3iFFbtc5+bppcchRCYw2vuVA1kRdbwjheem/7QlPjf3Fsko3Vh6IZI/vgIR+MNsppNN5wV8gXz+
hvd3LLo8wJ1Bm/rGZww1KJ9WGdKLeZqv5bCf7M/Vtk8XTZf1kkfJWZHFKCr6HVCGw6ocBpzegH4P
2DSStcLFqL9kFx4MipzNnav/1tWfpyb+AG82j/TJWOEh8A8Jx6TnLD03GhGOk/nmrM4HwwBVqCVx
YCxtom7b1daKcQip/icsHt5WA2m/55EYApcTOLliWgo1WfOEWPkySlPeTKt7+GI3MD+qxF8/AD3C
t6mCmbX5NAwU3RqsHfuZv9izJLnC531bDmcjKb9+Bxg5nQQdmeEFu1FpDNMEYZ7MzZAjV/Kcrh8Y
FUf5LJK3UpHINtgRs+TFjroo+WdYc0JgVAcRZkCwLhxK3eW7toisb4O1gpfaKCtt/l+alaoXn/qx
rCvIZ0GCAIB/w6fnrMgttZxti0TsfIIt2rDYA+FOek7VjX4uyCqP8M+CPRqVrLrZIuw/FeFjFqrA
QWJ2NJ1jOVoBuLcuoQ69bdo4V+yEV0dz6DXOBtouZAhptHVon8NPxiUT1ix97c6jcqhd7og12gU6
SzuldxxQnS0ODoXeISnO36xS6vlyN7ReMzjACaDH96+p3GWc2dI/ZiMTXfhYN7VXKXB0XVzhPqh/
m64XjdmQGDMDw1lxBBjXCtWxgHQZR6GpLvyhdno0WVqgmpZX1f8BW9dS5nKOLSJdQkmZY73MjT0Z
04Wdb3kAoJwlPXJh7TDbXSIVP2wEAsMiMbuqOlSDedLTeHaT3LmJwLaOEbLOqJllxeGPOlHMutqk
4oNnbfhklwZlYBOkaDr1M5HMigo96nJufNGOLeHG7Htg/Za+kjVrBKmShk6232aRUSK/ak9MNhmK
GmI9ZX1txBWEFudvgTozOKKVeiFtKCqbD+WZ76CB6Q8pRCB/gjnzIuL+/0PU3PY/JcMh1CrqOzfe
4VFx5gX2VFk7nLWndsfDdJThgj9xQHramsjST4q46CmvqrtJL+VebqCKoDy1MxmmP7uQAM6Xqdu5
Rx473C6On2gQVCBFolx9GzpSZb0riE6IDhlIJUg44+TT/AktQQhoC7GTz0T0sA4WNzN9p9gGNoRb
2Hg6CbdunGPn0f7pzVVxWVIuzksibfQsbTrhGaSXBg1NejiAoh6rWPMO2fUDG5gfKByKrM/nZcR7
twg69Wj3c0qRKcZMfSUKvofcUesBlMFAIrj15k9++oTaAGPmrjVXfjoXKiDmtRAaNQgKiN67gBNB
K8soOe3BDMhsN80E74NRy4Fm47672AHtZqi0slrDooXo96+KOvT1R+AUeLmHwpyAczNHUO9e4cP/
RBh0Pok7uJDu1odZ8vWDt/ewRzQHaznM785qZAHMSWlTzNTn/SC1vwsvATv6YdcZV1lONbj8h4Lr
5wl6yiveRyaUwm67+ww/uAtFreUrSDA0DRZmA0maf/ajh+BTyBtWhLgYBp2V3twFU3oHKen+qlhD
ThEO/0Pmu3JCmZL8QSyqbbgzt+5R4/GpTIOzCcxt1SaLFV5JARRid6PNRBuUpp9/Y8VeysqbSN90
Odq1Cg0WmeUHDP0wPecsGPdgbZClRd3yz+S45QMWldCgg3F0vEeXGa5Dk2ESbsusmRpjn2tJhIcc
FxY+YqN/gxxdmb706glv8jG02X+k/zy8ARCnMVcFuvp2mrk+3VuFdK9VrS/SZmnerGtSKdM6oTeo
OlkZ51CAZRRxVxn9asB0Oz4ATqL1bit4vJ+azB3uecA=
`pragma protect end_protected
