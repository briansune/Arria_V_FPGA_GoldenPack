// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:21:32 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NvKvLcr086EhFjcvim/FQMCaHH2quywtYcMdtbRtG5Ph8DggbO4+StO4ZqZdTS+l
1Jy9/qCZMC647rRfpOBWRTkjb5Q9LYdnSgUi3zO09TqjLnqb8ahkgjtlMYS/bGLf
KfQrJoIOCgQCxs2fD6ZfYTEvU3JfngRIncybRjyvBH0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 59040)
QhUJfpMBsSzw0peoS7JrYAVngFbsOyao+A1l2czYTQD2l+cye6QHZAFYzisyz0kx
oj826Lfz7B4pXxqQbSbDXdFEyx4uFSOqJKyUj6ryFSk9otSCtiSt8EuX8X5xdkB8
nBm/Z+dRJvF3EoJc3c1tEXKPCc7tHZfEelJCMVvLPSN7ly9iOE0wNsq7XmbfIw+d
6a4rq8OZPvPKTWfabY4fl/YQtxeAuX3sKj2cZ23H2DedJ/99hd4GqP7Ndc05kDeM
HNmA7kyHPr8+PqB3nL6eE/pOqiRrS5OeEHhheTNc+gClFUe6XYHUxaok7nddOUjX
gxdEPiqF6pHEUWJNcwyGwVSTlifGR7hgUYE7tmlD0NN2ffHYKm7sO6o87e67QeS9
szP0YHtwNsALfbmypKJp3DZ4ypRR6yXuEqpTJHQOCw3KTyuFWzInUkPWCcOsJ5oR
3J7kb82pd7Cvo/QuQ/EAnbDYopPPFbVMWLPAqcWfPNtCtQ0P+IxGvd/GQ/lB39ET
AVHXlESo8NpdaFXKd4BXrSFu8OpWBq2TIZMKJuyaKVVyb5PnZfkPQsxOmb8aNO2Q
p8giPfZXaZuQ75bSRCZ2EWAcEswJNVC1oB9vhlwV61yBfluDz2ORc+sXVHQb2eVu
XsRBpB3uKxktWgle+H9UwMNv7RStE5df9UyxU5XBqRpZX91tiERGMTn4foZYt7P+
IvIdm/ix32JsARQsQTCkwRaODUaZvKK5at+JiHHfUIklBLZzsOTusoItWvWQg/JT
ucMT/OwDc41b9+wF70yWQJy3ClgBpci94xHb8/8344If1qS88GeBU4Mp2Vfph3O2
wYbORmtvXroK0LdiFYZO73XuP3LAfTwZAYepN8LoqbPbynWZhrQHN+6Q5th3DlqN
0Lv5ND0XyZElhM9hOKzaArhYPdSkRkZvxDekJjAoF0cNK9m0zvGgbGWa14fuEJQb
+1hXeJSHSnXRIV9enGFnZJlJt3QvjN4a/O34pOKA+em1FMrNQ+AKnyd7O203fenk
d9yVFopAUiwnmgCTESOnWfqqBz3kzS83bRddm9PU8hqoPlvDGn/pQ3G/cakj/XHA
FFISKx6XMAEGEvzrMQkOMLnOCC8XFxz0Ip/h/i9gbx6Ra6kKxAnRJBQKTDkjLuaB
sUv33hM/GYRRvOa03Ut1c76zr/5ftZgjtlFS3GnB1myGFLfV0NB50X17j9d+x2Oj
83ELh4zK74GCH2sAP0bQx8ZBAcGcHDwbuGNRufeRw+JLgnm3nPYL5+XdP4RM11eq
triWGhamO9qRtPKyptb18wUAr+oPPu3TG+cZmn6uSPWk7IouJDKs7a46iPR96TGU
Rf6XYziCnzfc3hwrUixYV47wTmdygCK2JivV2EbqIRo9mw7dA7Ob8xVKX/E5To3/
Pyx+IcgpkYOIJQsCBj3RhyUKSCxN+qSmxYBUwf/k9fBFMQaayu1s8TasM3DNdz6d
B4vKFMEW9N+cC4ZCFD33keniDKzxxYwjuWvokB/BTvbPAtPUZsChInoBVmfFjMwp
6uTNmcyXb3tOPuSYts7OhwvUIOhlUiNuIqhgRWV7uYqNcl0fIVQN1vY+cf292Sle
H5O0oOcDHAEQnXcyuIZjC12Kpr4p+HIpXz2P6PGkSOixH05TElemSyy7faUCJmKm
CHAt1e811EXwH4uUbxxBzLN1HQW5OxGDyeVFuUAIbbBoZ6IuSG3XuVMA4ZvkHqp3
IfsVTuH6fy4OuHj9g3o7AC3qCVPSe8RVICG9J5y4rGELhFLoSUWOMPuJKym4M6Ym
A9v3h7ws+v+X7K90hcSiPI+ghe1WxMmTSYbYeeQr2RrzgjUIaQ17hT3Wh3xtD2Wv
SWR7x/tE5SYq2aeVqpHiWaOJvZfc5WDRakfgQ9GvU92R1FbQU0Yqz5cPW9hDvFSH
gWxkDri5vShNeo1esaNyPgAInx8T892SQEqPca7xFZUJOXsL3x9D//bv0w0MjKE0
NQsXyXALeFUvJHpRKcJcSXPAhVJLprmnotyZlKc7PwrXdjKmthL0woxpBPjhlA2G
MwMfM15CQNgFn+wyILvyQFI/Zrb5IKdOp0mSc2AR+269l8Ky4wmzri/ds3aQPxUY
qi1JJuijE7AcwIiMk/h87xlw9OtmBcjh2RC+TS0E1do/qjVBE93UEJNEcG52ix+d
u079qo8cLabHfVk7z/xFeN3TerZSedW5l8gRSgZZgdHDkBv5IbS6rdSTKyK2yG/O
r3OjRtKbDYWDMBtvgrgEkeKMXRjEHKVoAAHclsHGQ9c6hBFq5bzKM99RMi4xQcHC
syRb7m7vy9Jgn0obIAWA8oof4NXBU8UNTBSTB3ds26NVA5yvOXGrXuYRI+gTeQYw
rF2zosJauWC18Zz1hmF7mjjmUdoTAtRSzpL8wDbtuq4042HfoyvwTZq1jZeifWZU
tJ1ml7KO0haoE3e+10/59jUGnF54X8jgOqkynyiCtWDlGHBKjcP+K7t8A3ijMXBK
2xuOvBZxSqvVzqSqQYqk32SFo7Lj3tvj7D1cvbPnoCX5TFD6med+RctXXux2ypJr
ZbsuEF2qq2adC8PedPOgxWyyS/XVCtrM8y6CfFIHXrHKqxfusEoZSOjhiw2JrpzE
lOqswKjh9RwoLW4mLM64ELUfo1hq3rvBD+xs1JAjia0QBwqRnMuPkPCtcfkoexFa
z8FBeupJaNPrx/mqz4XiDrLAhT3QaAFqt50eNG0UzS1WD1m18bFLH+kc0HFfiNBo
WCnzpuNQlT03xJ72hqff176b7FWp5oW4bGiC1y4U4Ub8lwNRNwr2ZYtLZij64fHA
l7ANonoZwq4W4ix2soNnn10P25zdO92CQb9aIaBAyh8vxr/5L3dEntYYWCe4fF9I
/RaQmYfEtPcQz7eAnaQYBcFpnsQmBCN/fno1e26jkKJgh8PLrXZK28vshT3Xs8ck
y0Upi0yaDNnHX+UwMtl5pNeJ3z1FfevwawYBhoOB0D3UwuNLZDdJ/tyyECeamcbp
roMq+AdMA6F1V1EFpHNPF6w+fty31nBT9ZrBynly/mWD4xi/69xHWTSQsYoW/Ae8
rdUEOlrQszBjI4HyArMGXvz2n2r3gp7OxtE50ktcbo6WZTRzEDLjIY2Nq8HWYngF
pNanV/cUEJCxvD4NdfeTSmpEAgg7FpmM3W0rv1mkwm0sng5jiogkQG0iR53vyQYm
tunQwR5U4eo6Os6ruvLyDZqc4NnqnHiUH61Tmpoodik/uDUwSVNvoecGRkRYUvHV
YHMlMTnKQ7SUrHsD4YICZc3/rYSij5mozdEPYL6aFdUEIZIGk6TBTfMqvqi/XmMx
l9BBAiC9pke3mLHSCDGPRCgAjZTEI1rnirpEA9DBzcEhehyClNyafu+F4fqXFvLG
tgIsC2DtsZWlb0R+/SHBWWud+d+vYrlrwfB9nqB/K3yzKy+sxT8xlK5Eh+lpudqZ
F7ESp5g1KcgZiYCvy9ch7IjL9Vcf6O45efgqDO5qfuMqDjY56H2C/zYSSO3/EwIO
Ef6MJkPzgMRHXzr7dtBJpHui6Z2vhL+xUAHsjUnU8LLebMiVRCtozlmCcBlQgpVI
Ltaehlk5fe/fLbUZ9NhNyYkNtjQuJiWYtMPGbGlCG+AJdXG1XzAlYKQyBbPQqOcn
hjZSxzmVwG8xr9C1q/2PKXXRSj6lFhmpCNDjZN+kZRRlt1PFjx7L/959N/V1pqIl
SYbv2KVHqq778GQae+1MozCtSWWhOwkMR8cJfsxLCCYMJU5uYGQzSLc/JBwglMJv
0QckBA+Iz4JO6kGjUDJ8gAJUSUvklA4MjF6kiGao5v5E+ihWgzhcQkRm1LTvujlq
ICN47Az7SMc6GKnCPVMECIrXJyMhviKS7qFrA7UjifmHxKWjRsQsWJ6Mxi8dSf7f
703z1oxqQdZtdH/klJy0iEosJA9DPDX4Q/wOVWqcQoLlbDMS0qGI47FkM6nwRDWK
6kZwZJzmUp5JbHjBmFf12r+uunibgVXh+4rObG4qCEBlOTD04xQvVVo5auwdp8Xy
N4yXHwwt6BP436+F/iCbBUzplg2ZUo6L1eO5fuTTDspM0La8i5oWVQTFrPzmkN70
uUBca2VbX+CqMOC0qLH//f9uxjbWSPaoldRjWBQXm9Ae5+wPoWzc7FAIT0nfk4Gw
ooZ5VSof+J599p5lEbExM9fODV7w6GG64yyaupnUnKbc3zneASDWVqbehvNqyTL3
KButKBN0EOGjfORvMaNBDVB8hYud8AEe+gvxrOk9BvAjsrGa4vfbPvHm0/2hJCmk
mpTQUV9GX6Ry8FJC3b34l3Wj80Eq1RQkHugiFjQW7bd++hWNRnBKboVlcLjkvHPc
fqXjur1jCENg+EOjegO/eJfnazoXvwCycggXp9xHoaxTFv56SN+7U6X5o30l+fwe
/TWfMO/VwSN85rLWZ6xxeLmjMbX8Ydwdn4HbPCZrLCVB6Fy5fwwqtsvkcWm85isI
6+aHK3cxFder8v6HEAOlGKyqvfTdxZM/LRt7r990S5rHvlpHhOKmxU8x0CQCRc3C
hcptiCxtkuXUGA3VApnCE1KHsvSFqRll/Ry5zm7NDKKRHlGGdSl9RvMjK2NClDxT
gvvbLae55aor7XL+ifU5ORvuuQP+mTsidmSl1SRC7FytswkImeWRjkoMcaGloK7J
2l6fyaEkPDl9QAEHLDt+n9/tQtr7m/YjIRHvPer3WILLId3u0+hZt9VcvvEKEuTP
FL6nKZc6flq5Sp0Tuldq402WLhIXHXSXui2OW1BtP1MBGxYxGIaLO24wSaViWo+L
6NVd4rl2BHijgDRXvGKid/LZWRv8xYOuxnI0hbwKQm2ptKqIdIdUndjd/nyt7mMH
EiJj1Ta+1G2lOt6268hYBdcHfPCg+aN1KydEH3tlpwg7EcMendkIrxSqGyEYnbT2
50exuX57uq2QjIKXJCCoO1PJNAZyPdm7VyR4v6EJhH2dch5hBsCQlfCZPJG+Rh/e
MjwlTvvVgK0YGaWS+k9bvgv4GE7Qt/qH3z8EMG99/1d8nknoPC1+qUVLvoMt8DgJ
RCRNOaQatOmkO+8kMER+jh4GN0CctufMrJILlKmRsTy00fICcgWoebyh2n9T6XUq
0KF2A+KJxbEmdiJi5Authq6VNcDt0iCg064Kv/D+mJL9xBpPWvLg9QkgN+hGs3M1
iXY3zsVX4sRo1FiGlxOlQ8pA6f64MvNGuZz42CZbv2scd7YFWsP0ZvjExIVOyZDF
vGYvS+bLjaZYl3G5sz+zupmRJhT86xVFpCoFN4IvtOmBkm4aCo9KLEFD+1o1H2+2
KeRZKmPdFxbd3ibpDmv6G7PaJRmEbufjs930bpDXPiJj7GiUJI8VAHxSERxYPqcE
54pIVnUucTkx6OjQllPIS/h0Fke6sKNAjPXJg0qQoFTBg4G6xx/vWCHnmTxMhWqo
ySH/HV/ZHDU0R6aKqwA+6VDms8q459xuDtPcGyZmUjO2oYH3w5sEquWHNxYrviZT
wNEtnrSYf/+lHipvCT5Ub0T6C7BqnJ4ny4SXyLATu9HB4fAmVmftA93yzDIaqOyY
t0qITd2k79Y5Kpm8Dz4sL6yWeQmN4Wt54BMsNS09+jLkWMGYHjUUcJrdRYVUP+xN
9PKZKr8Rfb8808vXQFEfSZUGo9Zd3UUIrwkEiRQwUsx5D4TA5eUAIvTn+ihIt2wi
QsP7OPVkSwK3it2Xd000nt293PrDmG4KmmGdhjWsvOmMyAXPXUEiKuglnmQqMB4P
aiPX/QrI0luZWO6VV/EZVDs9nIvIdMOX/cA750rtDdh/G/a4+XE4GFRn+m2pnbP/
AmGmxnAqUmizdwGFbFKq6C2+mUp5fWn5N5zlZlAPoZJ7qdMRhCoAXWq7m9egvmod
YnqhgTCQ5qW+wbBYDpYhc/Wg3C10NlipBBYp20j2PyomYXckGRFXqoATge6x8z6p
PbXrf/rptMWG8sYv8/yOgXxUAOM7uYfiWMChiPNu2szJuUfbekg+WXbFi2H2suir
7Oa9upHnzA6RE6tUFPLusXo1SvLLSATl7MO8q7tIsctITIvTEZ4lO0ppizNg87Tx
QzNHfG379U06t1ou+C1ivBioAAAYMoW4r16OypohbE4WSwUSwSUFCu8IKIBU0h3R
tVppwTq0+eKauQjo/gQipb6owJZCgPVqG16GkdLOT1aH+3uzrYmgf8tI4FXEsQeg
Y+vGcrmiq6zgUtEARdkQYICVR8OXjevuWs6q9VSdqT/4YZqXcemoPfxGO2idniWf
jPbfP4TuDKzVS4TNgPyAw56MjZCpOphncEzwB6LnQBrQpz3OpdoJU4T3ZlPsPsYc
JSBJbTrNtMqmP9wPKN05GXfoBmlCuoGdGuv5MzgyZl9Aq5BcmKbxR4M2Zv7TxhJK
4cE4Aef1dFQ+5phLJAYHly9Mx/wvn8haJJze2bX+tZFWa22z6GbXmJrLYMPeDv3V
GXMQvshLbGdxpT91LkvGFPw2F+ykh0Y/PUWdqI8P38rTuONVNQOz1WzinLmSD/Ry
P7X5py234R2R5Y9Pvew01ynwsZSZTs16kSPmG3pbsMAbjbfW+OrvPe4Q7QhJFDVp
4ve8l6dPs18eSIrXq45KM+71m1/wuMu6UWIdrdeljuN5jkSs8VcABBD0sZnmw7xT
DPudXaRXyi42aSAU+9NkP/s0nu3utMP+F8/g3vCdbkKHnfqmzNOF4BBKa+iuQK7Z
tz1mK4sWobtTd7+Wk4ANiO6zPTQlS0/BeI8+dI5zrSSQHKO0MwLY/IofCGkaIZu0
IrINU4yiGd4dYiwIZWg9vOgYZoGhGd2cVfTX/1Lo+yPNUpYPGz/XYmfIZEmJN8T9
k3e/8fkUr2ZoDMhOwGaGTBcQjbLT9A0Hy+DjjEuqTdqUM1crfhN/5FpDQI9Ptty6
rLmIcOuZRHSDrvarpwPW04t/imPZVIlSd++wZEIoQI3+tyV3t2vg0LXfVxnMmnfP
O0WT1RZxPtD6g1lOEzYKzjFg8gn2AP1tpku6hVrKugFPcojsSNBFWOTrNNdi2jeW
V4U3OoVcKWAKNToTxoavOwp8P2jS5i46tNKV0SPKgcYTb6AoaqGUgmB2Mv+CbQSE
7pHCPbiN/mk6rIbdEGgybHTijYTJXaSI35+R2o0t/w5q4F+g8ADavRQlSUrLe+Ml
CXLLiuvfdctQqZw1y30PsBeRcMpeE+LKgaLn/il/QdcLTVU3ja6MrbpYvbsLENbT
AXuvRABLL3zs+PtGhZd0MJL3A2/bpYemykJOqocwaXqI6QskhXOoS+UPE4OWHLgx
PM28FpBrjI0maWiEoRbqjhb9jTqZ2UZpK0AKDozPiqTItGJatbkY88iX5wypwsRj
q0xOCVvh5i8lFhtwHid7K2OOjXHsV021kgtBX6KzquIXQA6talL3IN5luiF++TLv
FZkUdpmHqD/Mfon7n3jWOe+HvrY9OOq+YccpYTgdmjQs3z01xe5WPATKTXP5lpkq
AgqRC1Bk0cJ6RDv4qiXvlzhOgNB7GbmE5fi5d1rnxyRCpfgCoTJrrtvic4lYGAp6
/v9dlByrCPFaAUve61cVuAUYhBgIgM1yv9TAS8h9L6ximbLuE/Ng2DTA74e3EDtB
8mPvS2P2yrNjP9Vj2OXcDwjwW24yVIOZt+4Dn6rCPFyYrufQO4fLdH25M99CcK3R
VyCb0jdaNEc4KeF6wJ4TWx6GHjlqpJsIx5ivifEq4bPTGJv1VMlJZYjeG7Qx9W/e
xSVaW9ZZu7fzTm4De65idNO4Ksic3WqTqTOhpiadVaW02BVda/TGSKtwZSmuz9ga
4ngXsAlaimG4fwavldNvlVY8zfbSF3zMZcgohhRn6tVkSMj3/YqXILkZMSPKtFVG
DIcZ1LHcyWnbgQbKJ3Wo75ASpLjIAA2kNft5IkmLNO8c+TJgWhi1YZhTR0Tg7WUK
8RT/CCCIlvW28M+LIfAKgbeGMJc/uMvDy/iCnG6spDs6Ycl/HthsqjDglQg8mB02
LsQUsVEzRoFjo9c/eJJxal16vXV1gWBc9HPzig9drAG0TB2o18NUjSKJNXUB2JsV
bRZlSQeP1r+DGDatiJRx3trLkuSvmLlnPP23mVcEOoQ8xiNIxbdBECc0oXQWIKO5
7G1/FUu1GKQWmWcFT7gO5XcjQCwZxu5sxuPyzVNvlM1tE36mWJkqVhG7W1b9KimL
I7Elt81BcstkiN8Ih7zFIfVSQ+511Js+ZNJj9WbUDzcUy1DMX2E827lsQkmp0QrS
2tRsauBnI6uu60km2lPE0etb2GkpACP+cRwRMxTs3dTmbX19Zmksyemf90Wkzkoj
DHGbGuRcd1rq6LPHfVmCIiqduprzPL6CCimIwEsmQVeE2ger+zx/sY2V0QyHEKAN
PPUXC9wGfw4TUke1rAHXwx1b8ure6L9J03KWphx8MMrb4vKLFv4Tfk791MVccByK
tGva8GUJT247PpOts4OPeOKMA+PvO3RrvNm6odJ0prAuVKhxTMhpzUX/W4AsqCM5
IoHVQfPMYVjJpaZrkNdlmu5XgKCs+5eRTaxg3sX7M3Kt/wzUdJLKtmEQKzq2+vq2
Wc/y0GxrA3OebdcJy9nGH1B0/UpikakpgXWB8/1xUGYgxLwGEv03pvB6gB/dDmfT
Ob1H+A/uXGi6SMFb9ccndeAAB9n00+2qCEM7kYdtkeFu7LM64faANrLfUVJnIQHC
+0BbCkjbX14l8Z0sct4gLXnx2J7iVbZOc9OOBNL6t/c5V8YQogLYuZFsggPK2VNb
0oaWK5sjF1JorCOT95BGUuNxL8OprfhMQ9WgSvVD1Td400bibNUtl8LPVd4d1S2V
A899tXN/TeQ5F+e+ibVigbZ1Rx51xEXTCwBc+QdtbFknYI5H7Ol1t3F6tXc6p5gb
HTSwI5CmNfQoIRHCvAfaqA1kr+h+45YGGW5nRd04wbcm9+xnqXTiBjXoK7vpog0/
Mzi6LYDc5UnWQwrb4JV56oLH2fbzyG4vLrpmKehhXeDC91VV3PhK93ZBu7nYNbmG
NRQjGlVa73BSUeFEW4KmzPlMdFFv4e7Txden7afS8oweUB50Qwp6X/sjtKlpLuCA
8rzhbTMuFMTGNGebGNkClfJeLrISf12TCo/WCszpe8iAxxlsOgRTCgIHTZAWjAkd
UY3LqRtCtWtCBd1Yzjfs3JaOMBLCUqjRx08tDjXP9gZj27avk/CWadQ7a9q/bW53
DyQI4EA1XxYNJLUW/j4I7BYOj8lChEIuZpwwiocUj1ckl2fczcYXqjRUsbAhB0On
+ChQvSeNFM1y/0LzERYKd1yZNlk1p9U9CppvRUoTs/C5wl4sNbGM54ttnLC76mur
MPKga4XWWvufAIrOyLapPWUqNJ0VzJLNr6bI3/9TcP1te3GtoFWccWsRpcj6Ahgi
Nzs3HBCrRcpLOfYUMbaEZB94+iNzedC9JRFr0VR0QEmOiLlloErraRdj8tVBi3pE
gAIPUUxeZ2s4muqUswJHEwtEkc9XZc3uF0OHzA45c/C+RYshDvqy3AmN451qmkuu
Vma7URN5Puown0kj8wF9uplNWtyZAtu3OKwQPTA/ZTNwsYElcIU1WbHLxNWF7/4T
CJ5dIAY6wbWBkjNmMSWM2xGLXOyv024b/+DqgGkcx8GKtzi49OTeiLp4L3Yjo584
p8ZvoFcW+I5gCCVRmTX7QzNc/OoedsiAT9dVQ6TpRgYR0Xi5MMezqbnGwZ7o5xVs
T9a52EdMGtORhRroLcPOlUahNhkb08lTgpDyw1OV7tDNG13xmRS3bCvBRGoi4FEf
4ZuoV/ihWPhu5v7BCqwqnfftUvUAvlzUTYrtcO7UNBQDqJsg5XesD/kJFyJrNlGo
Wu6MndxTtxG+tg1upZNr4kuvYCTL8lgaIxlgT5M/u2gkMG1aZ8RQKVZn8BiNrJgC
eQb3ArO7jsCv+LMFRPyh+N4KTIcpvpVkNnNjoYONbBncVBn8Ajbqcqhqrlax9zR1
YE40a/p29ho8u7QM1m5bgxgNt8FiX0u8bjMehD2X0Jlm7JcPl4YKt68P1KHaObHv
DJpuPzgOzc6I+cTuQybVnMzX3MVK3UBx3dic5aGXKHnT9qFNftK20y2OZPDeapfE
Bb5FhQuinoiBP5yFZBpgpxZNSSk3Pq0PV/aZbuHVGKj/7iFkadFbhLYIXLIh6Hg/
n0VvZsVeCc1dlAv+sr5MvSnVTarGWbU9fACe5wEWUS77AXuQtnnpj+8XcGm9w9Uk
Fatpl4TLj1hxsk+9Qruwgc69uJbhVa6/FScUwvqKDnEnFt8Gd6P7py7+UO9dhI9u
wW7A8p6X8lKy1eZGu2/KBjNxwntH2MyJvOTBpkc1PtXXpvz2TbHZW3RLSxjFd5rR
xXyzn8n6VT6Y/8uuy+jphAW65Y2oOUFJW+tXV+2cjl4StWQrTHSgLwNeZTCtoyDu
cuMdnoNdHiyGlgksWnI0+hwgl1rqJLwcclgD5FcFelluvz6ZebUB2MpAhC8ppXyG
ivP0X9b1HloNldFvDoyb5Mz/5zkOweKkdqhGOXH4n6gWg6XTmI1mUiQj/kEDlcxG
ESOgKqW3bB8H9ifKLFLHFwkNjjgpTTDs2j1W6K/xlNXaeWDOPUHg0Op3okrAKa1G
33FWZ06oooPVgx4jkzcjdd0fnw8Bjv9o43IE0q34PIZxH7Ayww16WmOoZWg5d26v
uZo8OgBt9U681ZHasDf9t0/ERLKeS1bwCQhxOptpCZndOgLkCaCZKo3q2oBlpYw3
FUq8zWpxqr0ZTSXuBhIlXPzf4VSmuBClgoU05MM91HHu/h/Nwt3wmgctxWPaXy4Z
7THihMMnwrCsoL38GQT1sk5sbNZcyh+S1HwkYDfU+SHbOhOSXc2V5ug3SrAa8hoy
8l0qATCbJ9d5lHdmoBkZ6++xIAMEjEovGSW9mN1E10wzAulIvQ22W9OVYumxzvv1
UeSWwq2hKnVCmBsG/8TepAblxo1HyfAAn4S7br06Frp+6xXylbSLDzUwGBSlpf4y
w2KsA/IFo2r4o51LP4JSb97fDVYw3SmwKsEvUMW+fWMECRSqZTeDVsbnO/rrnAmz
fHKOMcDhnzPVqK+btxyMTfkhX+XjsOPgvAKGLkhtYh+dizT7j4tk0OxOqCtqzx5K
QzUj08ky0auj0rC6T/2EFkr3eJq/6V3936vRsvIheA+ZH6gsezorlkH5JkYHr7ct
2X4vfzkuxt0YP7LtGkqrAoh19p5M70KDGCyvJw0BLQbpH+n8fjkJz+OWsDSZIp0g
OYdgvefAbPm71M293J33pMEqtunmLAuaDDXoOeMW3baNWZYaDue5z8Koc3/avYy+
KlJkx/TAhfhn/ClPi3+Gn1OoldW356tsLs1/XRkjQQAs4aW5//GRNFZn7lipaal/
FZxEB9785yVBdAxPDLQ8G2vzgF6ZnFr/HnOr4vK0wI/ukA/5lFj2KVPNtxEepf+G
aJynC3vJOs4Q4bXip+fsvXBHOEDSf0v2chRAZJKG9ANF2qBmrx9ih9QLOXZKdMuu
Ziy6lE+eo7B0mDEMOMn/TAOZgc5mY+Bp+18Va7x/bF1G3Lri0NcSci4Jb4vyN9UE
FbYcArLLA39YA6n6s+CGqeY0zKCwlFt8V2soMnZGnwggmuQ/Ibhk4hGDvQQdL20d
ZtjvA8Lrngs7BzuuFX3Jo0jYV6qQZ4nVTIHYYZHQECa3xxd4A5NnqXNIKbuusVPg
d6NP+suSXT/veMfBcFeB2rzXLZX9FQk+rW4ayYNsavBpF7FTIGlwelqeTPeAF1om
CFFUPlFtfQ9zWXoss1nd6uBIazOzvkXuWigfnXdYpqrmycTmntDiepWADj2tn0jc
RyB9yuRYljapJc3cRtiVE7bM2kOeVnHBLOy1jBkY4V2nAxKFgIEW2Ltv3J4NtxBt
QugLFdjfwVhOMtSk80yUWOqMLR9vQjefh2zISAANdVVWgvEHFkKXD4m5t2zNv56L
iWu93zqv7pSUixug9nrGfTVdkBn7e9uq4gEURGxYdLLW/geV7oHq3qSlA3e44u8t
iLewz82NS6Nul6UOlNY4F/p9J2GOb5eTpXJecU4EBZeGz0hRvxmqvT6a+k3Niyxv
1+FYu/VGbNcqch+DwKDgaUWiV69Oh+IxAaK17NbLcsIkzZSPod8BiBs0q0OJI33p
NMxpDGGXt+gbtlBwEXjCtjICWywa40Re4cqCG0tryUnSAQSyF5mHypTeXzRv7K/Z
bxgj719vwA7JynY636UomJ4CfZ+1bRnxsR46JWoKnVM2g6O6/r4KTBdhyfV3U6o1
J+ntpz+rmIfjp7ltPOXpEjMrbYdy4yIC3r+0K9leVYCpOnG28NZ6vJoMWQ335l3p
akt4P5vx3+z71R/Z4zgJVBNQVyLBgmQbY74Bbjk6yrXjBFL0m4DGjrF5cEvFskxM
AlUAcCvlKsWokjdvIloiNfbS3hQ9r6IOliKrz0emP7iDw+YAXqwoyqB9KwC/5qoR
aSaS7FoJZ7Weqd3/vcyR93lUjun3iHCuWo9JSBcWpivmN6AkEB/3R5FzmCnIbEtK
6u66McajUETWn8OPvuGu1zypQCxKY2ovKVr22XdAljRIvRfZZNrV+fBNKl+rDQLV
BIztv0ZLexJVncjXgoJnhVaCgKXh5cPtqINT2Vu5d/d5RMVvLWojz3AU18N2ZmTC
6IbwDVAopUPynYQ6AMrPGpq22n9fztPoqnmJI8aeeSjEsZ6oPlDD9chLA8bhl40r
CsgwFQ+CmP4toLwzHbt/HBzesiRhUy8hkg1+Uz7B0f3yBYnCV2kTwGTsvpDLZs3i
cjyvDSouflro4IP4M0KhhaBGIfJX8J6l/r3njuCs7AubDn/lH/J6cgmv28ydEsOF
lZ+UmQmAfBCY7Pju+pcTAYIskX1zCYq4mfKZq/e8B+LKsly9Ac9z2N0SSzabq08X
9YAUOKorkpiHED+EYUnR8Kla9tBSaDRS5Z0XGhqM+WxDyvVZOVpM8Wk4MXlf8i/d
gRHIBP3fzD8tA80KtqDvO38blYTcI4nauvVITwxgZpXiGFWaw29x1o6vd8yGhqRb
IaVQH9WwNh0W19cDaK87IS5PDlEXvoPZKf1/H0waDJwNK6EBrowy2SfunI5ijHKa
BZ0HoW09RgWdRt58Oigq93blxzkS9REMvI/AefB98+PR9B3SLWREqDATWPxvTkye
VVv2eS7JAzyJ8b6nTjpkb+fYzTwx365D/o9NPnolStv3Fxoy48lsKJ0RdpVCa9p3
/WjWgT3EJRh/hkxfrgER3ISaPfyrF6wf0jxwvwWFe0sVwNp/zoLtxa2x7VHnWdBL
qWvtpqi9x9lUNupSe9//O4P/GsNwSUsf/8ROJTA9KQvvu8DoWNkGKaxfym9TZefg
IKjOt/UV01K8VHFrQo9GlZUygAIOl901e44pf0XNVMYpcQCsjankW8M4eIfyu5Av
Kc9I/NCWgJy2ltCyjVMMVNrZ+gg/Mintu1dP3lQRzOg4GfROMP7b5+ZMZrLxy6tb
aY7ZA/hIoPr0dgl0cot4EJgTP+UTX/VHQ0QWwXfTf+c9ducYqFC05AQFC2LyYUKW
k9qz730GWTtpTFpahvSSxvJglwCWyqt9dWY94bA9scWokXaT8BUuMAqJ9Td1aLcL
yBGZ5PvHW51/y5Y190QMkUYMUkpkna6U/VLSKqgNO0luJ45dpvNc67/A9+9zZW4j
ApiSXy9Wuzqjp770dF+dlZ/ezWiYtvfiUjSe4NovmcR1CLP+kvrKFDXeV0VdG8C1
b+5yNlpYzhHhau7XRCiR2ke3IGlblDBJfbUHYk+Fd5YrVCalOtJioeIJeVKsM5OA
HlVx6PBotIUlVE6Tt2ko9J3kDGjHTEO78VlkL8KcZmpno+lJvsfBaKjRl+j2ZCx1
vU8uyNSkA4WX4Aezo+9Lhu66u9uSC6SsMCr8VdZ/qVtQNA0H6PLh/SWUfpRXTRhE
IYY4nfw+W50k7VPW63OrYYz07Ry53zELCjZCx/NME+Me1xVWv8Rwa6q1HKtzHo3a
HcorXhb4Gimheeezop2nri/F20jTXOgHbwoXre7jJxWCSAxTW7TOJKqswuRMXQPo
GFWlZ1wIhzAOYm/xvOst+EhlWc5uWiKmzRs9b224oaQWHP8EteiTxbpbjekDjt9i
LkH/8vgcnOvAT77g9j9F9HDmc1f1l3BHhVTXqbrGL6WOrpQRRGOKJdlHNsHCIhUv
9m/O6AD1RgUrdGTktgMDBpztreWLXt9TW94cGd2cqu9oWvNy3IflWv7nnldLjJXm
QdIVEf9aEZyyf6QasL/p6ECOKnQpvOEq051JNggmwfcFnVEYcsm6wBuSLzDgwcI7
wNq+bMQLqupqfy88BE4SBS1O0OFRU+roTXPPqQDoM5U/hdAySD/UDS46NCnxRxLB
48ZgIcYHFTvSDeJ5JyFmUwL4Z/8tPnWFbowP6dY/29PAaoNu5wcPrBgzINy4lLh0
dCTSGndWigWDuwJrHZCvJDuPglDSj45ro3bbCDceJmhNPRB0fC289sFzvj4oP6r0
OVqElB5MGJUwQsIF+i+AOP55+TJkbMhO4Cu6QDsjnaNHpI7R0ySOFi/surOevrqG
OcsrVTf+f3uyooRo9wByAUPYAuDe9n/BHbxSA+abzIynV2hVd8ADlt1Vb7RJ/I67
J2H945SnMzFRTxRJSxDPeiLDSIQejil04qVk8NigGLqC0D8xfDBOe55ZeGhLYMfI
Sl7Lww/7lp/tkO1p115oFPMKQKYWCjVHxm8SZePehaWsPuHaUy2qUQ9GKG/OQoh9
dEHsGvFAYfrX4SXbe1JSNHZodRCpVyUA865IiheuQN6SoKijGuhQezYc5Ly4rAP0
SfSBWjho7g0/12E6DBaXmZTVKFDGy5HFo3BzRihoPcN5CYEM+PVC9i6/U4NoeXUA
OMTEpNpGfhU7xktDPIsv66W0dOagk7ZK4Juaba+vjOSeiIHUKgpjDWdYEgI1rtRS
wCqBgVwkueuuikFqtLwCf+cCtZr6DvMNVZOP7OXG33ipwKgqkSRW98//aGgM/ErF
JQbaeIJdYG1YVavfM5op8L6easxl+LFxOlLeO0WbOYUyLdoOghVtmnk4q3mtq0eU
RcLOeNAQRDdMFLxGk64hJHgUoR2gvB7pxtJz4ACX7fqb9RGnTSRJrleA4hcX7GNo
fotCWWzrzuyw5zREgBzhaCwWtp00vCppNCluo5ZutCKkf1mGX7jdoN1IDOw+p2wu
fw/zj/16UqrO5Qw1Zg6A2cfSd/8hf8rKcSjVRTIILT9LiMrms5RHR0ldYlzv22H2
XwpIWp8jA68gKBJCW696jEOh0Xksd1kXBp23IWKZYHwmadVQlrJnQwod8fHaQgMo
sAj6ejYVBsvhccZM1/zc/VtNfCTSr8K8GCaZqu9j3dazP6O3+bq3+IdGbcQI2RNi
TFxU/RrJ+RJZY8xLWq3k4IF2vqz/NClqTLApIx0TUU/g+57T0mQBAV5xuwDLtW3v
OiC8PGU+pGZc8p5Dd7R5g4+whXcdX5xzlL9yc8/kci/4R9wqL6CrSHvxek5SEoeA
rr+uDsBPP5wpTVHKNDgFUWp557E/d4c6TiOQhSQ1o3YFm6HyM9Vo1f5aQDWW0me5
HCt8VNmr+TVxP4AtYurF06yoNWlMOVVeSSn8/UT+MtGaiZUcZi+3Uz633FRS0Pwj
n/WzYN6lshi47qjQ9Pj5XcGyT/DsB2gTKPSRyOzTZQ/XblmAQhah/sn2JA0rD/XT
UaVX/Ff2ju42uSfQq/lnFv1bbnRjhNovsxsJTIJxgUl17GXNsSVur0HP55hzu/6H
87pJQl5ktDCzF/9C07neYabfO0W/kSR5EdaH95OeEbsyN0eAOCClZDQimZJg4qhr
1sdlN4xubbt3b0PXRPCKOuybbnpJEMcgmzGhdAr7NJSdF4pnJPN1xQj4P+Fnn5cN
VK8crqlRgaIRQERVe6QPOh/LDcOKDlgpzuXi8/eLX0HrXy3NflG2iULOnJ0MuLQY
P210b3VwNUAK/wmwHvDw5TIfOuoZ5lbf+iO0y56tDOXSem536sr3ZEDq2y9hFdMh
FaesDUO5nj0c5KQ9Murydq2sSDtTytKNDI4gBnZSp7iXgLFhQDNZWqG61eC0yf5u
1YkKaadfM9b4o+8RtqpYOF4z6s8Xw0At/oGTqNLaddTfa45Ha3gLk+/w0w1UE/Xz
FqWtdopOVtw/He5Lv5k9Epnn6A9MiYuna82mc/AOtOgvaOefvCDGjsqrVBNC6lg7
fJQd4R95zfy6vMf9Pq+6ljlBAfDWvTTdTVU+M4XY6SMiJsHeNGw7U+sY8To/6c3x
yda+wZlkY8fVVZHwAWYj5f00bzVHh7jyC4iGDhpsLzBDowvA3KvmTFrG5HlOPKYl
X5CrktAkpNCyHj48EST8A+KFRZB+Lf2ZR/K6KiSvaLfQMQgf9Q6AEXpRKxqeew3e
U8rTiTs5OsRko8B3GfUSBzDi1esmtIhzp6y5Rm6uqVaZ7JsuedJ8feY1eNZ7IP/H
/i6XcvYOdgWBnSj4y0LR9BrJxryAvCYz45rLBbbsCJUjca1/bp5v/8AgmjiDy5XE
QaB2JAaDzr7vzjU1fIwd+5hmxNdyLtfxAj5DZz/PRKWSoa5FpNC82CpBw9ADhmOk
ajz5V83/dYDjv32gFo7KzpITIvc7NPVALb8HECnMmG1ac68r7sXakpgBjUr88A70
WerKiRieo9HGUQvsyUlBlCVxRoHkkZ6+yXVE2xWDCAds46rhFf0eP/jFpsHgNyXI
AFYTzWV01lLxhT8ndf8bSnCaiOjgXWo61mSTT/IrVu43YmLyE8Ch5Vcx0VudrUFV
RAssKDaael1S01Kb+bf7U/pysFnXgL4CdabA/2CH6EMd9+cCqAkNs/0eOXiw/0yD
OBXULmHrd5BAKtyGYCgqLup+LD4p+ediz6ZtSTohliZgyX9Og0EFSknZeI+e92qi
bDds3LrUWMq5M/B6hW5y9glMxbEO7nfl56ewX1Iuf89G8+d/Um01p4oH1MNmCnpZ
cRXtpawdb5ExeSSGwP8QVczVN3k0qtdjSJ8yJ5CIIvMtCtSwCG4IywMkDU3jG8ho
53cJ5Xqm3E6ZTOvjrJT0ww1SCFDi4vFphrwkux/Im11RnBG46+hEy0PnN1aPci3L
CiFLEQoGchtH5J0haWeo+wHSZkX40Iu60ACkBrMcAuveifwYcDZu4pQaIiirKy/K
+64128xL9HKLZkmNu9BXZUC1OS0MAnD2ASV4TW+/Vx6MNqQEFd3iBOMNoBi6dFFD
M+5fzSIAs9xRg/KvrjhpPNePidhu2Xg7N3qzW2oEckgumD9GonAsfin30STY8pow
grXjK+BKof9hd2h8CgyeIWM3S5qPvFUL7mLHFyiPx4RiV30mqHNokBp01r8ydVm4
azw8zonP9kkNsYXXgj0TncAvMzXZuPO1EGssUhsRWrCCF+0YZbCsb4W4JV9kpOiN
GbZdZKtRtLwXd10T2BVUzhvID9+Msx07LQtof6xs4+eDLFSMS/jVPL761YYHm4YV
GqICq15jrCvpwKRxAtFgzssWm5uZbqVgnbsCn8v3Gm4msIUOIq8LT5BlZx9e5AZy
vahuNJ6BD9+OOkzmlFS/SJHubkfiL9iTFJVphLK+kiDYzuLlCdpgU82qkiZuDv3B
hR5IGlgYj5d69KTIHlgdrq8VPKR/0xhEN/3Sv64AV7H4wQbfE0bgZmxPnkSABxc1
IFJIQzhK3m5IoyyP3ZyjwVbR2GvOGT38izbg1zAwin/mperPCgLYf7pioDj/AyBe
vTOPw5Ty9ffmfJ9vMLQtfnFsisA7zVBY56PckbZUFDuxETDp9109zvE5zprQU1+E
bb4NR3NYxsQ5Lvpn7/Q75ZlPJx+ee9IbCAUsVE5F69YxiqGKXdooN6MiITv5PmsI
V9GmlCUqCkn/a1kSvy6XdmlSjJkwmEDwi6bfw06cdEDf9uFrSNsqHDDK+9tGuya/
wh8drIVinMWrXzNum60Xcgsf0+906qyCGSeRBux6m/EUQAbkIohvaFD2JwNzFM0D
AuaL8ngp6hLKkHAT7IPN+l3AASvx9pQBVnymAcdUAcf0aQU3uE4JXhm+asFrxb4A
X6oxqKNZQmTcFknzAf6cRgRwR9XareTT6muCb21cy7vkW6PNeDkeLOZKnYXA4zA5
Bwou9WxTkapPOFM2USK4npYWvheraFkobt4I/TW3FkBd3u4acQqbcCZqD0zonP7J
qpq5PIaNWj0vL+FElEsGCcpC/L5vpNTUc7peg2zPn7250rsfPz0sNBqyks90sRRW
0Op7hpKLnjOMQAJmPOrpUg4Ft8d/bFkjkxmXGg8L7fWXZuXNmnoPr/BeJGHZgV97
HigghSscRbDFIhbmhwddZYErGAKhGFdnuNbRXcpPAnpBlbzQFMed2jI6L6JKEpoF
RBKYXNchRp16RpguxEqpKLQqbzwdv4K7vbTQWq4Gqganc9CgoTKsR/RRyij7+XhN
N59Ek3/j8RlLyxBgFbsJSdGZhFaT4E8hO/eDZvoxRrZMXTwGLHkTIZFAtCr0T84R
fxbIE5YFfsp/vh0I/2T/xm51NyAV4LY0oOzLljUopjc45z5T0E7kD3f9hxidrtAJ
iCusN0vYGzizbt20Q5QiMQjesofaR2sTURpmEgs7KnMtq5u9jGqye/tQwMP3NTo4
u1hiEghMhvxbNEj46xR55E/b3RdASna8M1sm/RTSZnAQcWz/Ke+FIFw1aaOCTFJZ
vkX+m/8gKDJlVgQ47+Q2bK2py8Kc8cFrIkijVbS5B3kDe66rp+mdh9rCAUex6Nbd
XP1GmDT6x+h17FrjAIiDYA6U/07fMMdlAUIqe94FBpn5uwgk2J0L1H8X8NOFQMbe
JS4cz3azOew30W+908AMMQzr8uctNlB6I2KC14S+iU8vitBcPh5SaznW0mSW2a5p
2s/EaLE1h2pf1x8A+49iGP3SmZMxZqW9AzMI7d6o/OZpVaFQjgB9D0YVTck9WMKE
CS+9Jbb71e63wAR8GBkkpoQxMfOi4D/OqgU1I2mFkF+V2EDh9HRdi7k0QKCnq5ox
jBymSyTp/VGdClKH48GwegoLvu9w0jghX2bKVs5FjAS3QDH4Vl2kQGV4RR3Af6jr
7Akr8V4FkeorY4l8VpQzsGU51OugVnzEZjSsEsFkkR6wh58mdln4awcLZecQHtRE
d4N3FIVmWhGBkc7Ld38IrVNWn6EcqAfwb2gkOpFLZtjW1xhK0F1OWKEud0OAgMXO
4IeL6eUSGgkJyzzne2z6MlZ2sq4/A8mgBpIYF13mFnEvaxH7CA7e6xQYkuoKx4Oo
c3DaniRCMygoih3dOAX4zB+BGrenchyYtotAgLi+VZgDezS8FowcvDPwO44+e6z4
vGVf5gjekkUnPXVziY9SwuyfdBek113vTPFdK0WupNCbCTVoSXCpIGFV1jKZUR97
m08ZWO+YBcu+ZQvBJzvi0n4F8HBx1rfGLpmssiqaW3DHR2BmFqYcAITtB7aJOty4
q7H9Kv/n46GYUScC4+KdmnLogufW+ghN/wvsPvHIaESNrHu5ekw/8kG9vQq0VQlE
7sEbsils926etajMSaRhQkLvNqy4aMZALREG4E/tr/uIDDYzzcUdFJ936D05RAtL
u4mmU0SNNdYf082XgO355GofNlUaSf9tuuE2w7NRXlTm5lcHXKdVz53sNo5ZuAUb
eZEQmXqjT5xFvT7NOaIXeueZW7mTow5qB3fP6xyGMZzRN9lmyYpaDQxGK0YfjJ2+
0Xr3/H+WDOtRMhm2WswLJJq7sals/NwnjFcVRSjSno3XjorY8QxP2gcSTfU0TCwl
OLEw0iBiAKTUHp63I/+lKeTvze2Ptf1hpJQ6cp9y4151wyXQo90M+k5+9+c+LULQ
5M7YeHtpe1ys/5OW1p/SmmmenJFMjee8sWSOD0k6SFEogL5HxkUHovgxfCVwvwxL
HO3ZXJhI5L7YMov87w+nhsKO7pzhB/d+jwux/OyqUVq+/M2BTlQvBqy9q0eH8kOZ
NLf96FZCyc0znfjRHpkbzAs8kY+XItkGGUCM0UbickoYKwSX4y8TIS9pjCZq9UUZ
l2EnaXGtHKjZ+y8BhpVekJrXFsHmNVvDMmeTErWKMc04rBRbul0yeS6wgJcriVCV
XzttF+Xtryzmtft/0dsl6lIvWpCAMm0omc6OitUhqDU3L81cXpbYoj77zdx3jeT+
r3ihr8lJGVCP861wK011+asOLkL4IztMz2JBleS1s80Ogc0tfl589Z/Isd+BUgQh
QAsB31JZc6W55Gr0/P4qzoOGVc9fOiNLwDvIie1nAd7F5nORq+S5ea72IqP09Rfh
dg+EdNxP0cg+PgZgmJR5N0O5TqINv6OWnZQcgMKTZcmOPx8Hw3aHXJPOJTbgI3NO
XtHdIDl+F6O44edzczojQa3CRiY8j1XpSAAuIDfCPut9SEycDBK5iNdjzd1VyvD5
LProR4lbirxBo9EBEQ8BoktKW+8psBDGhDsTUV+U8qkv0SfzZG7H9/0S8BvGASDb
wRJNKVlAssceHVS/0o1BAaOr2NShpeKXYFqevbTRmwR62g8zjvuYwkQHrtqWTmO1
OZBvDdqVHIOJgH1Jy7P8LNsTWBZe0F5qyDhAsgEKyMtHyToQsYZnrqEluVLFVmW4
i2Btf7c/eSjRPlVoym7hfuaF93/YbvlLuZYC9yTOCmP0to1oC6PSyKFuz3Y6HQEB
mgwIUXQSbcoPDX+8boPj1aasfJeZiqoQoxMYWJmKb/K/ygVXD2kEsosOwlbXd8GR
5rhcU70oO6VOWO4JiIcEGXZYHF1hUAHbs2KeIbxsXf7m/VzbliCvAmnmKTtjunvL
YNE67X4QXog2kZjkIJjlmhUngxZ5Wj+wDXWD/YeCsNETibTf0cYzAx8B6Liz9pPa
HLc8SW5FdLvGVkDJIijyTesLuZ2YRANg+GrQpdflzmug24Ffuc3azrQMIVVrIQJC
AmMN4TxhwkT1WJKoIPXEVoNBiR9QjNDxb7I+Xya4cWg7h+/BR8cx7r6+0QolYLCC
X27N2zF6TyKIkNmThH0SykFkH3PDcZU9mzWPVx5wrxyi77w+q9Bfu3WO6EOlfKew
23Av9N9Pf924mK+JgqOq+uKxfqUQNlsWAhexciOx/BsSYrQtncccScaYru88yu0Z
UO/u9LemH/PkOWGQuvDZEegwBguL/cLxJhzZYlvMj6o/a6+NUMqKuIYM1QLel8F6
XLI5KCG7C7x/1ysexgojeOd7vJ4ItoUjq45RbnfkDK9Cej1tW/VGUgR793yflNuE
M5FuVDST2ToFHY+kHhGMbk3N4cRnQwavoZoPLId17ezaoXT+MyV27aDOjuFaa2X3
2OlkzOgTJav/myarhf31qHWMX6cOqVAs49/hlRflh7zL8/kYcWUG7MjG/+LA/t/e
pAl4vRvXHUjNhbVBL4r/Zx3is0o5sOxhWPN+b94Mkc0XmDK2Ho4OVrjfgXyroDS7
ih0oUV7yvRdZQNTTzPkBziskVPKrYBFUvlG0V48CmRYjUNgdHKFVearCzZsWrW+5
tZ8aEzecyQKHYAUOTeP5a0WAM6uqMZXP11ifMjsYtQ1ps9vJKjhIamHSZePTDHpo
ybEDFlizgN76L2HPrJG33NwFouN1zk59URMeMhC4AZ2oNiEVGGG0LteKZ2Yk6djE
xPeVNcD+MQI2qEFxkT4ij427+5skWCuSg+y3PcAupgR8g+9n8Oy4TGOGSUis0BZL
ZFJkHtqq7ENEzvfa0IoNHomYqITCnyJ9+WMVadr/CH2xp6+3bjy452qyqbRKhuRq
mVn8FgBNSFp0vU+V7dq9tnVn/1a0/ZDSw0xKvftpNuLhXbSPjLPv6EJwKUc84gJY
19VBw2cvQYrYoPWJfgexGqGMqZ+PIgdeio/zlwMbs84DzFsO7DfEwICvGF11xyvI
XL+jVi5Dgt1Vikhmq4RUfB+4ndZbZq1a+4zgXYlGBQQDOZIKQhU8kJsqkd8d5mQA
xIYFrkt8cTYbQCxjcuCfMD8s6mFC3XfEG4p+gcjImZnZW2vF1Owe6ZqnJ6zxUB58
4jVKkhswVW19aGg20Bzs7r/za/HYFccxe7Q2BSiihGRyqpLoTBFYW+PzH0H/rYvi
6y5pNRukrymXnNV7lO+t0cdHcLvPpkrqVRYHac91kb58nmertefhi3oSRb1WMIYJ
+CUYPBs6peQ4psiGHGlSM/rZ7OS0dPMRjTARJ8aOR2yN5b5zxCDjjfL4Civh4Mb6
2FKmeNHUclHzcuhBbz29J6YJJslcKH544HkB5b/tVAu1vX0I1woOxS/59B8c87F0
QOyJOKaT7wmG0l+NmljDLnyMtMTXEzazq3T8cJoxLXiNv4AdVpl70XVEWjNTlqBX
b8+MlKYxhi8m+YKkXrkdyaazDAYhfkezcwAs6uClLJfJg0ungj04b1p4BHHwhUAP
4bxHpQx94M7xbXuN++RxZ7sNnxqyDDYmqWYOeYbkR8UmgMYkgkNiBcCmw7ftc/O+
f7sgqG4E/XyrMCLFGY+ZtdAUmILv5mGChPeV/42vRdxOaSUUuWO2P23HM+jam67w
mLlANQKFHKuKJ7T1vDzI4Oh1rvHcg7RFkUY0uEKKlAa9jmmq2Rw2zUtFDrWnn6Db
XUmDj30dDTzwPkBW+NahaoYzKCUc4kW3jA0rVPT4B88lI9+SN0BZq1ZpS2kClITf
nq6AkMeSAWZzVZug9AKzRul0YBCUb4EDSYaAA2hnAwMUeQbiWg2M/jsWHzjr59oM
5EmNbUJWVinZKcXZ7C/ZZammlpSOMznBlZ6j7oSCcMSaPULV/9tjXTZ++2fKPsh7
VsgQXCKrV8eyX62uJS86CTcNqhE+MJIZ5bWLtQ05cW1XuHv5qtRoXe7ZLDvn8A1V
qSy0hs5XySbbddkvHfbxo5dCr+ZG5FEHCrJwa8oT4k36bVNA8fULRLw3wZLwGsa+
BqDsYMeyIzQ3fVbVgYVEJWmeSJcC5im+oLPFGiI0opdzOne9onKuGuan1bIqr2YR
ZKbHQhJcx9FUzm4jgMnhsA3YE0Pk1B3JdhrstoadAp/6h06H0PzWMm+z9Yi9OAvm
eYjfG01iZOb5SUhZaEYbvoGuip5j1JOuwgvw+/YJjZkwhN8nnqy7rSdb/kljQp6m
CS5fDK9u39Z1IL2SLQZ+MufE0fgLxX1xdcWBGWTTwnasoBLauTEhQnay1hJ4NeJD
XlcjliFVWjwNDpPtdCSc2O1C3aVSmhMguewiEJVB10MLy8b9bd5qaIl329GwjzqU
GUVQzoCF9/eln6r6qICvxc7NcU36mNaJ0RdJ8cL/RL4bly3FQoP3XyGLMl9J0rVp
KuK/otaEkzUP6n3Ms5amK6Ea8/Nr3t6mXVPoLbVTAJ2Fcj5EwEIDCBSbhf6+/ehn
TU5eNvYZ6YZT52qeUHE2bumB5qEnlezpUQYK5P/uaPFjXmJYDGx7x1kXjaJc1DuR
Sr4oYJi8fv6zyrKsr4orJRa7+XrQBDfAECPcknaoq3WzTFAQ4ePeVD5uW5QdFu6Q
dDji2EQB0PVWpm7Mf52SqEYwcdydU4PH92cOcksZMe+rIZ3KKVKw+jp/HUgHZj4O
yDWfzyCtuhnqTXH72gHF4EsgUhGb2Yzy02kLkDC9Gl9nzJgw7Kzj5rQxUAb4yt7W
VDW+KRTI2tVB3XcMII/EocbW4HxV2bwpGL99LUQKzPXMKRaJiZJCbedDyEfGQVui
+aWkAQPkt7svH+mT0aYjUQWc1kHQ4l4/B1KFiHUQeiEIe9KYH3iYLLdnIL5IZwIV
l+Wd+JxfF7TL2KP2Efhe1o7opf4/UNbiQlHrWOlN+OjhIbgIR0opYVGZ7Zp+JTg/
6/tyCP/6+DXt9M9cuSUH0sbOWQzLe+u29Sizv5L0yCEg3AUtH3Aj1uRrh7+PTamE
S7/ZIV+mck0wHpKkHOn1oSvz3RKTUk01jdCSHb8ylSmENbON37YkNCrlasTJMi50
yATcIqJcdFf8ppaCndwid5CZzlzaYzl6u68AQhyRtvFpNzh+OmSw+2gtePjZOqiI
B52bnWfplhvw8GoCBmjcSldk/yJ5UIQZZJ34rdzw/xEPRuEccs+3v87rE8qmxMbM
iybPlKbXbz/EaDTFtC9v7j4RF8okYKCa3vPfegAU+sBPbmuqQfXi0Rr2lrAvspyB
4117LL3V/EbUBgmln25SGjaFKv2aOUV/W8DaKUk5RGw0TjYARvWSfG4u+qeuhJzH
3R59VpM3RlVKV91+DoLKGUAgKKpI1KThmXnr6eHnqstDlvApEg+W2wszbmmNp3Il
STQIIe9b6UX5xuWCfD6iNBBetQiJ+P2A5VAliwk+FBNFb5SlV9uQIppodttjuhj9
9ekHv8Phe9QQzFi44ZuJ84vbajKvCtmJQeyZb0Ea4UI3Qxbhno39JxwcGWxS6DGk
8H4Unu/PplI0nKmzcti35rwfJG+ZjQ6X4shIiMSluGxNJXJe9lQCO/aLBGZUOQui
YVmtz6c011iuU0aBSyx53uZ0+d6ezeTluHEI3FloWmhrOm4+G8gRxg1sMpyCbhoo
mOsHYWtdrE6U8wgUgEoT1+VYRu9Auzok2Okohwg2CMwKEwgkxCX+h/1enV/cCkV/
h0rpMrGesh4aDXCSUS9pq/3r47X10QsUGQ5XnJpo/6eWFaylqlFfomUXwKOiJ84c
Q+sC8sRdAufyU4RA/wa/46HadGj8U5FY7LjQc9prDDSSqPj3JwyPYIc/3QbnbwLh
YVdquFByJ0J5VHCNQ4Nqrc1pD1e+90LwuUXm8HafPjSp9Akt3tDynr6esalKg5NF
yqQ57U5OBROa7AI/vp6nDdjNQlfItI7TDubG8kwHlEXCvqPVj9ZXg9WaT+b0zYc3
Y05DS/MADillNZ/0hCDCc/5PwEnJy+xzjxq36QZuG1aorbYaJXbk4mhoXBCMuHJN
NtgUNglEO4iDGSnR6+fEvgFaRmQ1XvhgvMuFSfeBNKf/9YjgmaPRO/JsXJuzQUSr
FGvYZN6YtBU4abBaJqJ01rTCZNFhIxOSPNP69Xe9R80jPauPEqDfI1sMcMhQhdPW
1YxozkIegXmncf3YTzJp3iBnJ1vnkYuOu1sjg0lvTxWAYTSlrKvuiUV+XKENeJfG
i/VJETdZmolpGmqY7OkGqE7B/8IbJaQ65FynL732pi34xLv0MxV05HU1HvhJOaDA
xYud/09TbV+WqxE1mg3yoLxZgDBpcyF8RGYvJRdMEZu5cMoee3eFFa7nqfSTPZqs
NJwYovcLpGK6aSmsLWa4QN6iEJ00qWyTsRME9dpvy2HrVtYwRnziqXPuEV5+vwYL
KV8iQgf3EU41Il1Gq7anBn6VcNdKaRFVRrtd3CwiFibv1yvmFBXKtyJTDZ0mrxEg
i9RBLSU+mrhTztEhyOfKEd4c6vilUhDQrK5Ev6+NNJy4dqKdcSrDPRzbZl79foG1
CM0d5x+qxB7y4N1WwJDQa704M7FK45B1lPn4DI8eqnY0jI2WgFYKsEgP7OLrFmvQ
xXVecbGraP5NGzNywULJRh6frJysUkB9k/MhHWvGwk/mVHw8VKb3CWgRRTH6W5/5
3xmYYM36D2gpqv/C1o6n2VKQlnehuSxHYN1Y+O/FizYnX6moY7O6h+5kGRCHm1mV
pDFOTEFxqrkMk+JO/q0KPV8Ozqey/YIY4nhlWh25QE8IxtjH9or8OnmOBd5QI9Oo
xCLq6/sDpJEHhLewldaTzYiI+ZohQXjj1hWaJskCN2jVfcqV1rwIYp8bRHibGoEi
V1NxprRNt0gTx60AJrCvIFf7l1+fhqMVqwNsgBUpZyeDoVknfYSvbLxA98w4eDKj
YRr87ctVubWQJfgrk/kbXtZV5Kx32Q2VqUpV1rNnrRstCwzZA0r9q5cG2qbQ6kpW
7rDdp4DlG+zBY9HFZKTLPZg4jpLAeQnznZJwHF/mS0HagnUg7zEh7mjp5Ju6xn6Q
R3Wb5x5ATeZgW4oGeRNlu0V+wmmosm+J8luzXJXYhAF1eAWjsHagSZp4VUdrYFgi
qkRZwZJqSc/7WDScgqKyrmZVVfEtjtrQxHmBLnsBnzX5Q7Zv8DR6TjBmy0e30PEf
zIyjb82aoLtKhtuWTjjwYxFLoQBDtiqb8IqpTu/qpDm662hTbt7mEqpToBTdELMQ
Tx2KGGx9dK7QTcrhP/kAZ6Tj4mKAByG9UlQYa0riH4ioG9dW+IC+LdGauALVVW7a
uTrm+whWVYY6sitkeUvIydtmKncYUjmikzviB8eDs225m9w0ZNrkMvbH9L3TUiI7
MkQUE0QIPvUJ0aSl6+XTX9iKOOo8eatR7UhQP8zxrmgvs7vQ/tEfZJVYcT878Zvw
mjc+AEEAArfEASrLcvT7/IVuULkRVN+iytTAqSeeVvVv9tngtdp1qmshMrrLHs7P
cFx/+O//N8LdDmxlBylNK82or6X2wnPr/VxyvCkRjYsSMIfs6aJlHg/IPKha2NjO
VIXEACi1rPhp5ALT55b5qjSTzRDcNLH9iwFOaN5C3pv/Rrgdd9ObRii9H7yuCkpv
WjIGx68LAf+F5eopWGK1tddJcVJxJIhUXvvzIgzphK6EFAj3kWOBV0/As0auU3tv
6c+ny6/r8yB1gssJQHMqTOGC7v/B4ZPan6gzw+TRF1+SGgqaBvEL4jsieTnN80nO
Zjd9RyY12TXiwZt1pTiN/dWy+K1Wi6yjh7+zavrIP9kY+uVRSoPARqlHcvoGhbvK
A9hP9v/+7Oi6HSxdO98M+wOD81agp8q7yoyjW9n3WatgY3rSB/s4MQmLy4Ptkb92
FkOOEFgLrPyhFB3w5gPFMZvU9CAuIzra6vCcjYVc2XU/okG3dkG+ESxM5WT8MGab
YLs3jhc/ymPkq/us9bsEYlBlvnIF+WA1rMQIUDAYzcGNP/K9ZUtUs2p+ezwFr12t
8QA6oUedkgxtnaUHQW+JxGOrWCJnjEJkIGqukjnDr7DX81nJSc6Aq4wAypLB/7qW
R2C293QHv4loS/bJIkPy3ImT6FSQl1FAbJgipMWpQ59iPHtJJCMGL3TQ07QmMaw9
E58SQZxHPgNewwOZiAyWcl03idDb9hoJTTKmxJ1HF1h1yHUU3jzmMiacnUL0AWkp
UHt4dlIdiM4x7YKSppQiznEhDKnwILdHRNgFBZNTl73u+ZZp9mWkEo0I5MiAyswi
iEWIqnOQLdzANnOgtwOY1aftgqj1UvfzmMzNZsYrhrDqxu4BoCGKqJnpAHn34MUo
T13/xTL5EhAPnq0TRq66kQAZhTB3P1VakaK96p0syOWzbF5nRkm9tT5V4LpX/2d4
pt5cLAnd+OmpoewG++fd65wi6WeYKUHZMGkjR+6Oh2s2r+gSREzu6dYGz5EYrKqp
Zo106z5FfyMkciGX2E6Qg7XVDEBSI2M6UqaDr48tRPHrjgh3VVgF3KGFoYwuUbF6
K9hOdpEWHczSr2I1XvkZAmWHoUe8qq4vjQfQXhO/pj/P9qqVkEeZ2GpotEH1drDG
6Zkj159cWGBnPFyuDKZWge5pPERUh9/X45swHgPRGdHmozn1jEk6Ok0MIrEF93ZY
9FT7pw99oTblSXUb+K+MfT0NGmgMZYKKGZLvkTj3Ez23JUogzmcrrlrZfO3ydIki
F8T+Tm6LgOq43zEsw6f2SHnoomz1nWdzP829nqqPujYsQMDNAttth4HseBmqHfrQ
aWu3DuEQatlZayPzUtjGTRZbC+086ZypynUr0j7Am2eJ8mEnVRfrvFoRJ9urBq3g
+SqlWWvsdMVJGqB2e09/ELZOuMvWU/Dn4fOaYig7Ypv965fWLkmvM1Qt5kNwnVkv
yN5gXkcgL6+IFMxux2adMrQhAYAzlka+nqUlxjWWz7+KUGhln3yDqbTPI25gk9vY
0M4JxvSKM9PjPGc07qYY7Ea7KsvniEIweVmFqHLk4UZNyPAV0viZxQQ0qX1Eixqb
NjY/y30sjKd2GZi9r0szKzOQTZkrsr9UHcUHOWbbJ8rsm4+m4QsA5aDxsaxGOapI
KjT2nYaTY9U67cmPndngvbrMqVBxMZ3iBOKPGCK6amClEeKKbahbSKbU1IQTsLo3
uZRWoCwmWe7eyJDfCCDSWcr2FqGvatq273Lbyt+l6hSUo+LHz63jjIGk62MsXW12
DR83w97MC12DTamgWxC052SGVqCLdaNcLOJPt8mqy1iZhMxREoLpKrQIZtPzRIx7
fmzxg3o4w1fuInTvJZsbp9ef9jSsZIB5pl7mfWBcv9AaOuhabOzf8ysgF9byn9YA
Ts8ht2Dzmw+RxKp2BL4UvuHmjcnB44A3YxStKts0707175t60lkbHP6x1+mf17Yj
PYG+APcqMm8fBPN/b173jBAW06jznzapcEI7Oxfbpr6a5KGG/s55HPowYng5wQK/
NgVlNI99SwEdfIC6g4zU97l/jNjmKQwU90bYKGjwegeJRKHkO3bLeHaCI9w6JXmA
+IB9+mc2ykTyznpv21RLkz7JLsZZd8lwJ2kR28vY1HrjoAtdyMW7uTTqUlfkMxI9
c37qE7NMWB/JydBurGojCMmR1q/F1057A3Sp36oE0YlZKsF/rEtrzpQhX+zjJZZt
0OzB8EG7fKyLnDq4CJFgDnPIjJD2z13djnMX27inQ5Virss7shggYFOpygAmirVP
/tNsvIk49DhAaL7kC71Nac/lAD/I7FFX8WKxc6eLuKdNGgYf8wr78w9Ki8niIX1k
oqYPyMtOOCwsLm14GS3yD/00ouOCTBgLm5siE/r3cP77XsxZtCJ3wVp7tS93Ww5K
yzR3/10NR+vwRYu7Fjqbed01fUdHY0bs8oa2Bt2tWvHrg2VH+l4tB072he9JSVpw
/zMi6FggS32N9PnVadxtrJkqYhz3BpI58sq5oC925hUjkXkxAAbKacd171H8mWrD
/itwbSSlecErC2bpZNjEylcfIVg5IqNz3edjmIZxe4IJx6ZYWAjLQLAuFxYn1Es5
20hGSanY/c/rdT4ezmsphv02St8gxsd51KWTxSePusgYEdrwtljlHc4cEOPkvuqC
7Is0oCFbMIRkLTy/YAQvKFYz67eS6X2wDY98gylqKFfHCJLo8CLL9E7NebTbA8Kn
0GlOp7bjVAKCVPJoaWMv71ZhrWCdrdQQz19qiNp7GN9W5DqoPz7OzjnwlLuTsL+/
uWbfuw+lqYJlyplq41xu/0oSXFjrPNuwWwqb+oAGcVu/y16nMeh0zKRxPNLD2g2w
e1CT1d7aVsXXMO6ki8MtFnBqaKXIktprM4CQhju9+E7mtO8JRLlrPSn6aFlEKWFr
uYEEA8Ahp5TQHU/jCCdvYVdw/W4RD0oJUU3gk1pV7RAl/GYfa/PaIXBOefHmNSnx
jga1ffh7REglggdCkiKRgGMModrZ565LZ0FiOu5RwN6BAoUSRF+m7FKwXYPTReKK
B8jJXuAqBLeXyUpPfQ3097Tz0+373MTfZZ3jcrJNMNZVWgUjWudAyQfpYAsr/rHu
E+/ZCvO+1TT3/tbz6zg6i55DE56thqC48HTChVQtdCvQIbGOLjTC/oHtSwX0nSvd
Qb8uaFHlXM2LNKav5mbL/DlY0yxuUu3d/jBhbewX0Vl/kC13S0dYYq8SuW1Byu1U
+eOIbcQ47kg4sJL+kTxIhgMKTgx3xpsIjH8H4jR7SCvqmQZHOP6O8DUOnZX1KDsa
wbFzvRc9r2kP+RmIXpApRMilZzVn+fLk8S6hEAi3P9TBALNQqajBCLglgXuh9mHW
PP9JY4ltePMbFjxfPYcr1D8IC8rZA+m+vG24SbMJf56tAxksppR8R34NeZleUklt
SDUS9GRQ3E+sVAV5KNGvlicowWyG+OwQZx6xqhiJRHW+4hMruXamCgVtk09OeCYt
wEyRE6HtgOCt7G1Aq0uRkZfKLcZrIzvcH+DtgFpbPJfrJmuCOXqT6k5sTfkyDzaR
v4qv2fItqFnjanbbmu+b34hmLF6ew/oZ1U0WD/XEoPoEc3JUsxE+QA3iSoBroNB2
p6XtXZiU6Gq9Or1W7cL6xLljbmNSOJwEsXF85HjfQajhskFOmcXTxhK1IF1HA7zt
7LJ9aCP0vY43MX2nYXj56yk9rLxIi7aa/UOI94fx+qXj3lo3N7NHPhWCzFEjLjQP
5gQkUfjvW9ct/4gdEr61Z/j/37XIQxgyLu56XvKlXLaPOyOv4tPiLaQeg5RyW5N1
xDBzuK+xyJgRknJPLAY+nQcldg/YyNXNmDgbI+d97aAgaDYTjUWTcXRc8obppGQv
aXWBlZB60+Mda3UtBIqKVTkLgKRfjgSzjbrFWGHuVhXbT0V1fovDZyKlTUmP2XWH
Ina4UJ03V5fz2yFb4Iq4iqABg77u7u1iD9UjGFRmkJl2Ecr9alrhyfDLZmRIvBCE
sxYiQW0kf9ED2nJo4jwswL7iePJe541PKI0IzDDE5CaPipC54TEKKjJuoOTN45lR
EkO4S7eDZ2kBaQAvRULd0A1uHrBR8zb7PY7Xyxog6T0dM8lp0S6FEDgk67WrYmjk
Ul+qHGoeIzQm7cLV2EtqXKW/TDaGK9/p7ETzmkeqkDcWVqPXFrW558YPJTisXIRs
YxCfZnY5MAUsuc0+5kBJVSOuTPmUmcVQvpyuY3NSR/MEYmVXGgPPGEEkMOtXtUYR
yAzcIHlHq2/y+lIyHCO9/x7hlNt/vIXJwsfG8YxKCuKdVUMZMChL9cp+Jkj306TH
lMajhbF2169cuP4JOIqyeUEBSBBUc/XbusSiAGAkbpkMrKfWIhpH9Qxyjv9nOqX/
hcxs+e7UClIvgqh8/WZwoW33lbilGjDbGpu6rYbY+3Q0NS1nEzpGKyfrXKQYL8g9
2F/ygmo3FJfSC+UUonTPbzal80LEVuY/8heIEcHtuT0tbb1LJeL5+fG6XzBYCL0x
VmIY9+S8IQCstixzpV/dSh4Z24x1fa/uv3GS0jgOI0GqfZse+mAHTvcLA6/HHra9
UVDrsc2Bli6pVFu7uqRDH3XqffsXFt+8b6gd+K0svy3R3bjmtIPdBu89XzOPS4w+
ZIc4iqLWvj7+ELdk0NaaGnNKm4NgmaXDk8yJE9pVinNoGQsnthj6tQIhvewZpIgN
cXQLut78vALVqJhDTJIVObimQZ8S1AY3M8ESqme2m8Vx/2+wi1DK22wjLQ0QV8CV
QvN5i0/x3uVJ/tk3vYzY/2mKLhTxlrnzlGaCIq0DA0j6eS1zY3/OiDAe6xLkjS/U
SvpUGrqBsGMwKNPG57ejol2/doiofq26YkD8HHKkUglX50ZyrckDjb61Yug9H/bE
ipscNUj2jF3nDfcRG5j5jdyuVbMCiSJZoQ6CXuLPmzxmuXSO0ywn1IqAcMzc5sZC
v4zln7XGxPpGpPNvq1853BCHdkMk8CsewK/C/iUkx8UTvZRIrydMx73QuSHBXoMZ
r3h0kZZ3E2sV+EKhOr4IX+9GH1nabkKZD2lhe7rECz3grd8Nn/LkKSxMJhwrZS2I
JQDmR0MQI2dha5LAYDx2SReI9+uw8UbnFmCGHvvmLLpuiRFaWE+au7rhOeMtOOUO
Y04zV+cLjtwaBPjQcHef0C8sgxkpCHKIgAf4xLv7H8XahbmnY+WpcC8cYzt8vOIO
BPd/77nvMrr5NoOnp3mNFRTKkPmf4iDb/uEELBt9CdehjViHrDDYGXflkzSYf/3a
wPNHvqciyrp3kCqHlTK9SJA0+J7oFypgMiLClqgDgs2G2MM2CxFbxwvfxDJV5ECp
ajmIHIX7AaWazecq0udgZzmlG8o1N4GDkvWyJj9ju4moKTwwE6R6ljBURGF7z0Ow
AwebrIwQzsx+NSr8K2XdMkJMoWPcHjMIAIMnDKQfXUS/4UfqOM5ZIGSNmJUGPmXh
lIRNUciI/ykl3Dtwgr15Mra5fJg6Z2+AFdl4inFk2qrtg3Y9NDerOfuhSnPOpZHe
xuHBNmiZZ6VJ0PThL57OKUhHyOjk1A45Tqcbx4XpJSy8U8U26em/mRMxA12La1fY
LUsaYJIrZil/bU+p/Knw6pRWwBFtf6uKCaH8cxejCO6FawFlKsiy8IokSsbtQy+q
Fl2AFTlMa5ydlrrDwlN/1dFuhesv2ESmecG68SiurkUP3Iga/VUMQ2/sXqMiJcUE
ih+bF1NkPyyvq8ky74kMKFFTSaDNkw26e8otreTRJ5woaK8Lvc3rhg9A3hyjNfG1
F4jCjs3oJJF4sZG+B1QsMcVqhixW12HBIbGXznBO7K0foJwrmuqFIx3nsCDywFGf
25ESjt8GUYyqj+IjurY+4l+LBLOQI4dF1jLzmOEcKAmnKN+s9qhZtnlv/j3omHiJ
qMVEdHq3GWE9PZ+eI4BqJLq4ecB7nEcOOSepqtW6697quVMUsV9IhWXjE5O+d/zI
m6kbaqx3s428IhKDcpuTJO4pDJdbZ3PQcOKqlp0Eir0u4Z9DN7Wh9J5ecuXuuifI
zsZ++AP7lMaE8KqdIcQWxd2nnyKH1im4z2bnNtpWvLb4X0/QfRQ+bUMia23hG76l
F9BdAKFPLIUpFIKfpDgRv4IkVAsy65pdoD7KNF60SgKHmLkB6aBP9wNRB/tPBQs6
8eeQqA4k1CHcjZ8ERdKr0+Jds5OcpXqddqjuQCxn8n6wDMXbnz4NIjGQ3KMZgNdJ
crU23/J3BWJhbDpw4BdC/VPo5Xx2XpflqLtOynFKdF1yLgapuBCf82tvZFUVmjj/
2uxnYQAth+s3Ph4QHmtonR8s4GWoVwXrsbf/rj01FI3Etul1fBSmiZCQg57RFTg9
p0LyJ9VK9YsWdsM5NDeNv9XO4C54ELlbDsqL3LhHdg4nCziehKF5cGLcXtSkqWqz
pvCRPsPKsCukZYc3AcMotaCtnX7fp+coWUBkfRqPLtjr54lYkO7oUY7YYbS+SFVj
qiOvlW/BUiu7GcJDVoCIokV8dNKyl1squjH2h2wqu3JeEAOI1jh3R/yz9JXAdgWL
8TrwJcYl6KE5aqdpdZGQwbsa1632PwIYQ2qGwKqTwaz4ibQqpc9d4Rj481Fhrv7W
8Lqvqg6kphnqwhZKidCwkVvTSpt7b88zM82p1kTrBgJbEGBd9U/3q8cIYI9BD4+N
RCO11QaqnPdKwo21j5ulVnl+RuxNETDnYx7bVlZ1xpBJri4DNwZnLQ6h8mJNEer4
ysjSsAythCru6QFpa/tyrdyZC1KDgmD32hBHmPyEUKd0EAdumS60KzF5yFVFFlX6
+AKhMltvm9YhFXWJJ2MWfEgMdzOyA6YDb021WQpXnicW8gd8JHOrwD3ksW8IUomo
kqWOLYl50m/Me921j27SAP8bb2+YvKFS9s9grPdSCLVoQ1tRcO0msKzxDBGtqsko
mK4TphLpt7mc2YG/9zWieHug+CgHGjk+atEK6bSzsmNoU9W+KkLiXAMJRQr5/KJr
6xzk4q0tMXHOleP5AMF9ykP/KGGr/zn8Iy6gTtQGn+wi3qCfZLaTFg+lDyV5O8AV
VBHMQe/l/ZIERLBZSROQGlQjM80tIp10QIvRom0ku0pB2y8Wd+X/nUipdCv6SM6u
r95cCo/vV39BrSdcUlqz42ZeGwDyL7sAmuAMhWQPgLiy7xJbzaBoCMmiAsfv6bcx
S7NkpeZMGSwhPtUShvSDBxlrhAjSNWjwjyLixK9RoMT7CPgxm75OIYU6HDY+oKu5
1BR5VHzYMylKMHvrijAE7EQs31wWjMO2rZpA0yyAwpm/RsG5ovqcjtSpDLXnTRIg
6Oip+z+e5Bb9fIsZfY9XTp4kJtPsoTW35Q0XP4huBu+lfOJK8tXS5t57t4ceXMPj
oJPlR/hJZA37pwpGay5VQtg0uOhqQRX7CYOBtc78+kUb8FU5Jfp9ClviuBMHCq2A
y0VexSG2+yRYstaVl9QXPpqh9UnKKHTewzhAwW2tBCwBmO816zgMrVl/7vnivzZt
o4PXHvTWAA+7TN11t5WRY1Lpb8KlLMN+/PkmwpHWYNSYQ4NTWfJ6BwFP4HjL+b/P
cmSsvXiw9aI+pQ3YdVGPvfJRhuFur3Nryz5bRiCWXwwAtRVKAkXZ0kTuhDqyd2Os
D4A9YG9fXfRxk24rOzvATOZVYNiRO0xL3D0LFaMWl13lXuRBfPbaGhKnz+x73yG+
GRBfMlRbv334qWidEgasFNRCclg3ylF8DJ7gea3+S+c+4yI+3Fg4frPc9tkNhHZe
WhcnnFvsXcbyQiMl3NSNxc2F86D45iZOh/zPvGx2eJxKqbUJgg5BJNlGhS4MYYbn
6BTFz9afhKnsLT6jql0R/Tgbxkc9LDTo20VKYYcGnMN7XDF9qA+BJw0DDmnOiVq2
BkCDer1ZazeDsSiwHhpnGjPljTyLiQt+1Pcuh6PaFS5JZbByxzrpVbQAGewP6Lqg
T6IUJDQSVvdyyGIx6ha675/QHL3OmATJ0NWI+SHaRiYjDQhng9iRnOdl/eahkCEe
ZC7SHG5ZyCaG8xzZKBXpZKWpcDx+hDBrtY+gbopkPIA9ds8mFt/4/HAzcDNtOzuK
l7y6wUTFMDa4JebV3vVNwl5NutY3L/5h4jvy9me+TV3nVg7wmca7/k2jvPofkUgv
vZ4QTAgEn03W1cjZdNPNFx7NGcqJGWye9kV73nNRviJAX/x+CZgMdGLpYmioPQkU
H5NWfMLQjBFvMs5s4J45YrD/CQZY5gr/HnPgsDnJ33cLk6VlYeoTuNrY0w37zj+C
Bh3KXpiHp5tCQTwH62pH93nxE3MyQkAbw5eEMw+XkpO0yeQWWWYnWOVROOCKxpnM
254ZzIp9ah/2E4hizS88vLoxGSBVYACQR2aVUmPKdXq/1Kx0S7aWEMuphzT2IC3I
YW3SNqeJ5N/jxfRO40GGqlw949gV25A0x5VV/y88fW1VxewO2n3q2rkMls21Ds4K
tzWb9Vgm8yxszbev62JuGmHtPChW6Uoz4NUha1N3oobNpUj8b7wtXts8qVEGGhAv
01IabTeWqpG9mKx3QYUUPSL7Q4EdU+QJFLaqoYaIsxwobAKxMauFANCA6LeS8/c5
fAHWL2wBBaAhwsTbMsBqSYjqNY1YpieO7p1dEwevWi7SCJdU9y92lDeT/256UYE5
KL/Ps/XbBiQriiSLaPWfaf61SuCKxaisA02ufMd9iJylOieD/A2ZYd2lHbEdWDKt
uPjCfSykzodxoQ926s76wxkuSwjEvfAWJgeTcRpVfCO8f7derBglfwyX0niZmQEf
A8xHQoai1H6X0Z30HfAGVvVnekNmgMjOFZ6WAO+BAGv8spBSj97Q/OwYZ3LTIsh2
4HDvI0CQT1qC16VT7OhkIFHBpbXjSpL13SwwmyaMmOKOqZ3XJh3pHyC2Lg5HTjhi
1q22XDluzU47CMxtD/Usr+38LKiMEY3Sl9uEbUqkAaW9ucY9a9N/GvuKM4t/+zmz
v1eIbY3ZnuMN+OXggfo52/vuetpCSEoEvSSbeZxD0Y3zGNQtWuzUvF0hNwOQGWaR
mpq83qjRLmqiTXmGl0yFuqdHOPO7MTeYECBXpvjc5KCr7B84VjZTB2wpH4L5e6cL
WnDHzFs22wMyW/jy2zZVylfNnYIogltj/Y/icLi6WKlr7f2oVTQ1qHHdJZXwzDDO
TMhUF4nMS7Tbg5R/mmj72y5qq5liMSkL3Cukww5F+D0HTKtN+/iYxkvAQ5no+ORp
XAouZFL6DIfjCwmzkBEZ/wz/fx4uxgowst7oIFn/DImhnQ2kfWjCT6x8u6sX7Aa+
Ae0kazvq2NopFzCFPZFYNyX1Jek3PQ+mTkStHy6+fvI/VU6COkkKzpc1Fn/MB2PM
4qf2YhYKAxnAUKMjOX/efTyC561EsFZ3GaJqCs6hEYT9fcIYr7LniZmW4ewX0A1/
KBTFs8AoApALHR2Hel94S/3MXWskmVpuKzKHkJsX1W5Qfb+3WJksc1fVsbZ8b6ZN
LvQghDm6DfCY9Sn0CvQzejESrtlR35UPB8wiWKK7mgQGfnvBcUzLmkhJXPhtqlcG
3BzFMKYlR/Ycf5hKwo4Xmn5owPijNFRFT39FKnurw4bAuoqwZAYT3Lqe6/UDN/2b
Kbqk0QaUDx5QxRTYvwUPNdXSX+5U+KMIGZYfJAz/BAqfzjCM832TmXK4GQ9+C4PY
WejkWmKiouj8PVIvawNccQmfXwQrPStuehSayNB0QY1Zt74wZNbTzyVX0Nz7163K
nazA/9LgyKXCgVgjDgUtzXvQSg6JRFci9zr/vrHUZBnU8LxCHsi6yItYA7iLzaJy
i9JDFPP1YU9thSK0piNOY3Rxs2fbyD1PNHinLJNsIOErY3Ko6OOGmfvg5yJPmFp0
PJgICNvsM7aV2X/kQpD2yRI4Mef69YR04vf2deC3QQgcu/62e+Uxrn/4IVWkj16j
eQb0dNg22cCLw3mQXN7DlCEuuf2mAS90M21RToY8LFqoTIL5pqu8Eg7Kv7S9GmZS
GBhWfmm5AuR3yLt6oQbrqXzd5s2xnlaEAW4hV/wC4LYkN4+Z8gp/acfmC2Mpm49z
LkOFnlh4Bc0NmqHt0djr5Tc3L2poghFNNS6vRQXL7NcZAl9lkUHbM3d4n6gKRQIX
c30zF4oV7P3WGCxkpzxGsvrf4OqlasEZEbnljeZekdrVTHg06BU069ODnSLjLADM
CEuEmPgd9LGNFhupf4eTe5mQd4uCW2KNayW2q+1CcJvq1FbgLsdAUpidoBEk1RrJ
CVJjy7UA8MyEIveCRjx/RnDBGEpU7ooKeTKqv/ZnsiJyLMnJ0Tc/y1lb8cVjmWwS
vARYCGPMVPvAzP21tIcpgd3LycDjPmG9+VoV/lXV/ZRAHqipW7loPCWjYjxcIxHb
d+8yEVx1/upcfGoRfyFZRdlVccHDwMDpREatSXyREKXz4wBtXUve0UqvOiSqRDXc
iWhZ+zi8zxusGT2bW55yirMn57snFbOhiaLtJrI26NqENxMUeNslFgs8IItRzS3O
Yqb7Rt0S+XNc6rTwroWhTFfAytqAuZT0H4NP5MYaFx1W7t41ZYH/jO/IQCbcyrAl
nj0vLrlqD1A5JUJ3jfDQb/4QhPY1zqdc+ZvDgUCOoJYh9d03w/I60g3vWUOgwSOq
3rXD5wAZMVYW1il20zsMbXk9TW1m5STAiWSzsIuujI08Wc9p9D5lUQKAPBT5erOe
tDIlT5gpmUx3FghK9SaBaLIaoZgP7uBkscwFfmJpfeOuwtfg6NnkTo4SpRV+cZpw
90M0eJMNIeivPicW4fjMid84J5vcoSMvX9WzjX8xYwSVs1R6PsRPPzXTqr774fLL
+QSAQlYzNE9VBNKE0ET/s4lFmvBDkywF+oU3HQG7VOEEURM4CIN+tQkI7NT7D+Pb
zK721onPbdRZTt44S0lhFlaJKnU4drti0Ftksk9zTBa5cHSq2EpOwb6J5xd2j2Lz
gU08o9oiaEJ+sfq8u3cxUveGL7DjF7FQ1K38Jc2rd0isems0/0itm+DtF06N2u/c
V2sQ7V+4bANXA6v/WnILtB6C/+OfXO8PiRlCtl0DlEENhAIYbminhHR/8c1Eio+s
kOY5Wf0yhdFfxPTU10PLyLe53AGo1dS6PLOf90p2Pnllwwa+HjKe0MDw11fsC2zd
IVDfBvJCndqAmVd0pZzkiNpbQq4dhXbamjAXNOmaZlzEkRCGJot6wkcn05diIZKM
iIAvIVX3zFnuVMzd3pO3I65HWdYFJPnAho7vIvA6Hj3lkCIt1wTqEyz+p5Ki5yNr
FQwh8NZdjXTxeLuU8tuv+dUpf0TZCAt86drRpGOATubCrOUpPqWyCG1G2jZjPkkJ
2GqjOkC+aUwH8niULtPD5F5NpbEanbT8VvvPqdqumf8GriJ+BvEsgpferDyQPpOs
uGZX+JUdAPzBKlLBZSGqyV3RCbbBrsbs+Pcgy/ysiW1/WbbLyf6p+r92aJX9CDRg
eDIHD+e/AYqzBYTpzWhKQvX/CdB9J8yQsgWj1gOy3ugkJsFIK5LzAAUgbV+tlWy5
qBujgIEBScUXp2k/tkmax78jM3a9LvRJVeJ/TLUTsjtm3fDZAEbzAjYPAgqr5uc3
ObP9m8SHXBLoEIu/zeydpyaU03BaGn5FkY2ZAazOn0ZbqRrS1ovzFoS2iDX99toQ
GC2im2TlsL9Lww78TJYvHRHLPYAc5zmhAtEVPZ8FTUvoYsQ8atvuw4q67LzGE5ME
g+amIUzeFdSmuA3yO7HGATZQZm+kCKspMNlOI2WqbuLcAg0QK38sUjMhLbCG3GNK
X60gVGBZUdp8lMSKytxWPBY66LaEVbuIzgSi+yrCGXML8TgqUE6vCeCDaAdbOcFF
Q/pKt4VQc+K3Nb6XftvHjqz4EXlQuETTJ/kZr2/wKhkOSs9j7u9CE/Wssc+lRk36
ecz+jT+7jkMFryTo1vAGgmXyq3qCFpKJNuLrhczIK9wlbY9vXG9VjzUrFoK4o3Dg
QbdDYTacrdkZCTTJeWe9dX6F98Wblkwl1ynWcbOhCBA6Ew1R5LmcBaoX2PoQCaA5
7OmV6khAsTV5b/e3r5B1YX76/zT13eFTiOHWULehW6IpuD/PpGbktRg7Qy1DoKOZ
hdl+ic6tmX1bZp/YDcITU7wvfq5YLO7dsU4QNf1VY0westoIt3uiZJXr+rykFD7D
m4QaJj/dulPehGjCFEKrUqXpV79ZiLPb9qWbYxGBl8UxquuW80GoRKLMYGRi4hlV
uhj7r5X3qlONPvr+8ApZSHHpSbIfQA3SRsiD/BmTwpQc1uhzW8N93MrjlZCtqPBT
0FfxvNennXFYe719dxChJ/OA1LXX+4xJIRFMt1qI4bBVHgQV0fJXfzaPZCsGm8GZ
GfDxZG6l1+jpKQ60c44LcaxwdXq5x3Gra1MC32/plo6nMLcAlIZZC463CwbF91+G
5ehWdKg/Ds3BnxRcY05/RCdOxL0U9Vfr9QJn49S5aYjoPytgyYqmf/YkOTmYFvMb
p8AxEAS8i5mtceewx+W77kuFcukAOMcJBEpx/XttemXJCd+bQKVYXDXvNP5A3+HN
Zms6+fZtjWUcWQfJFXKKDQdpB4NDph1tNRMCWPjZrbruzbjiFHJ2l23srcireyyv
WYqxm4hgwM6SQ1P2DHS0W8g4vkdU0nG+dS43S1FXXj9e9G7DiztWXhipA2Y+JICR
PGmbUC7F2uxbz4RHFGqSwYYXZVa6McfxXPRZxESujMlFZdAU0nWjXUeOpc0rU8gv
JgU8fr+EeM/tmZfBiloNxjLm5egsP2NGkFgE8ICMdu83bhBao4+IIgVMa9B6+ZIa
WJoTFlVxwIj2jJ+xEWdXyTdqvX465n7GbqbfE9mUrwuMt4N03K6LaN+8ldU70yW2
VLoH849/dMHmowQ2IT5JCs5/Rrmw8d79RbXijjeunDDasm735YSXEypaHMhASweg
V0VYN/btI5ubURPgq0gk3wJCFTMRZaAMHysb7edYGYdd3FQJ5tW5LouSkPjV4NLb
DIwJ36kctxc/vR8sd+biZeQtQTiqMYqrui+fGExoR9SQBkmB7zygtxMLRpHLf55O
ngKn7odwJt9nlGPVMAwjSPryCjxa+eiOhjXB7/ZoG7btL9sGyO8e49i8Y7QOuVzA
8kIn8sFcZi47xIX7R+wf5ocr1A5SU58ppGQUsp1oS1xJ04ezd+VJ80SQA4gm0Z+l
mt+Qk3AetVAdXxbRz28yawhtYzExTWAxr/vU96fs5+t8Hbtl0XImgaGuQvQQYZBo
wg3ejsk2VrRUtbOTgY5D06ksE321tqSJ96g2Dl2/CVzyZZYVdHTtcrsPwgnle+hy
LnsZlZyxHGS+MKWN2nm+HZnl7zhHAw/UQBTbHIfkUEmrSG9K/r2o1CdhxmLpdlt0
UR+wNsl7MKdU3v1tk4K3UzrofYfGoEadacYYYvLYRnJA5+DEgKLQrvB4Y4AAYuJm
0hHAargZCX9dtJhSk3/rBrJnuazvB/T0+KrSO2aiKaZBHEoYuIdSFjaeaq9k6cLQ
jp/W1jo90j0zolL9HpJJ8vDUvaxTa9XcntCOJ0kq8jX3TL+WR8uqSdIHkAp2hI66
fupcPM92QHmMXvaLAF+BSz1ygMIwqQ2pbtIAigLhTKhNoR8eodxL3ALvCaUbWrCL
P4ah9VBr1axDX427629XZfSKFBZYrIqyR7Hac11ed6cXUWda0E+5xqMwMfmaqvgY
RFoU+xztxGTHTfemNSnU7JxA2EASNpyax/FtrIQMT7MPEWlZsAzIBzslZTvlIPpy
E4mQn4tARgoZWjfsOM1DJeGaHa1yp1NN6gkRdCYFGiJhmlCpxtvU2haZjNYlwbOc
AwPzRtMxYX53JMtpnegH5TnJ7AAjbhQqKzI/YX88kdJgZt7C6/Uqf8QK//awSBlr
0r9N7Uvgt648KUj1GIb6S+QMNC2c8nkUjCJwLb8Nj+y796OSc5hoJVzu0HbCxV4M
TKc0E7oqcQeJkNKTxWszwjFByeAR9KLySdUzOBdFPeaZcv9ek81vgDRv6ayPTs82
NrBfF/+g630b2QK5VCi7nbNDk5n9kuJyyf9GQy336B/Gh+Gsrv7aTafotqNNY0m3
e06+UNLEAx3rwsJziBtP4LI/5FGjz73QYScF6fo5d9I9o/yFMSEPFe2x1KdmfTXI
LqpVu/ADLt8Ja32MqI5Uemv9wRoaaO3KfdFt5K5RO/y/LKrgxj3CatpgOSn4vql7
W260FaA0cOauGM6P7yWR0ri6YXFVyQBgqMgxU1/6nu1ZytoyxH5TWKdIpOSJvn2t
kvsroIybuThiyXt2WNobMeASSeyFVlEjeSbWbinQQW7p20uJSMQ8iDPrEdgtGVX0
DDEIiekXQ8p9igaXSYhT/7VUXBGNUmzi3ThSuPFzwyQTmZRDK/gWV4ozpjdMbqBh
ybf9anSEv713Ug91WEpT43ls4SeXAAAxFwyX1yaiy15Yli5cLZtJ4gzXJAvetAto
YLTS9gLChVBoaMiyWfqSK7LKvYQX8BFf3TbRW9iwp2QUZpzJIBV0mbCIvPbfnIqt
+6QZCBAusQmdyvrL2s0zZqv8ot3VW2w93Li3paqDUSMskxYbVDeoadUWUO0w1RBK
Nsjme/wS6wsCK2Tbtvch3CEGk9/qHiGL3SGs9m0LV7yHKYuiCr3Pn1o9NOQ+pk0N
V4WBoAhTx2MjmLvC/f1q1AigDeeYXPJS2h/i08oh47k8KXzp849dvOnm+XznGOQH
aEbjpWdpovhmBFqRLAt+Iso4L4PIDLZtTIpSpkGgNQh2mSB6JZ6VqnGbekePrd6u
bN9RPjMX1RRptPtuOO8yAn8XxEvGKDk6nACNauMiHRexgGjBW3GA7QV5WHykgGxf
0KAbopNlW6Uwkx5EczPEmyF+M7ovSFnoS+/cSNdYBJDV4zTa8KQz1ogaABxiygTU
X8ONxpn+ypsrmnHa7QfnxMCwUnFcklxDN+U7YcF2MHFF+bK3JbcjDJEP33Tbg99V
9hdjYAfjtBD+9cx7jhqK/kNHmA+RYKOjBp3eIxaaZlWVmqHVXEx0dpXcryO5O2JY
+K6hrhG9C4LLP4caL4OsGcsXgb8dkW+R9G0+4yrSioECVmQS7JqYVPqPuavmzqCU
odA2m1O6L8rJ/beZvIrdQu1Fasd4ekxiN/Z7gCBmyudc1ZczTAa/d7hp+/mi6aTl
EfnDNn2C0gBpRSjl9XesuFhiDahhWZF6t3jMXxcJu4iiUclv7MitwekCPrLgqeAn
Q0TqB0HQbt+jZ/hUETtMbh/WWrQvQGSR4XoXVH1SkNR+B4j7RG7YTnLQ63eWCDCf
C8ljNMQGgueAeK6cKxZMZxvsD1st6h+YWIdp6scZkv0o1/Z1sFr/qNUp+mEb1zy0
+CRLyCo8bIkQFvcxlh/4DUn6VjI5X2D4UkSLh1HoSYFLij8/8OCPVk4UQTYk2srk
mR7Kr6J8sqmtImaHEHjIfu5uDGfItZ1RybYvhmebzBjrm6MYUK+b9GtVz1v3FsVW
xN/OsZH+lxUMFf/X1iN5I2BpD6uVryuaYTJtZfKv0N2RJrBmWZI1eEMY+dZ/Ks2Q
eMAQ0xaiaJsum7QF1sWpA6VfzCzI0rRbN3I6OkCiH0L3kCrLzBXFyUoNxgzSZYZ5
rlazlOrpDY3JdZlatjvFAorBD/GzBNwPKsSzu+tyqvQOPl2u1K1LvYtDGCtoxhQq
U2Tnz1JW6anX3/j6b8jdLmXNPenjpPw2yV2LgirqDhVlRfyAfE7c1iCmnLhtS40A
55McV3mKk5Ct5OCb3Yl10m5jHboivjnj3a+0zX7koP9Zd+fFFz0I0lClFp8icWRp
iZX8ooU/tcocUFAd5If1r/Ofrq5AfpiBp0KdzTRTZB/zuhA/dlzT47adj4Qho7Uz
9qqHBGTiDF8fwfS2db9uvfqxjr6GuaVxIoRe/NDfiOo+NAaAIjKUurR6LboOg8Hv
4sHexmE/nK1PCOeMxEhynzW/RMCrLuFFUZ2STeY1E/AX2WIuD5s8zb1E6Y+oAstJ
UcpLoZDgYOrC2URMpLVjBvwFdOZ3amHX1xngZKYr+wcXjkVFFfUQnDt04upQfrhL
YDeX9Z1oyFziT2BZDlPZSUMDBfrpi5xK/Ohb9Ef0yFHnKUBAJQSIhqN/0/R8T89B
Qub3auz10fA0kr8RzvObuhAgTOf9edYGvHofJbZKDGyYXmSo8nTOV66w5BE8t1Fr
CTb9bRW5mZQRHiuSQnDvZ8jhVDN1JmgZbSxS1ZM/ZkhWWnkb0MwNh/sCEiFjeB+p
hRgE2b1QtZHNQFL+oV/uQL/AY9UNkpt7PncCzYesoueOWvCkm5WmasxorBloYkpp
1QHkYTLeTZYuApBaSns4YikgqCEfzW8mAIldGuO02iCPHyt5QEt3xUu8SgYW/kWU
MKMQ53TFz+V4JLJjLOklfGJm+MD3ciX707KVD0pxcWTiP92MeTAL5VDVtjCIphly
V527cZ4RkKCADQzBRucLz7MboC1QMFoGajfvktpIbNA2ddvlKnE36c8gt4ybts0/
b9S3qO1phg9p6LBgmrpBy+w4FVOtg1lZzhzIXkKpQA6XdxOeNIWmkxgiUe3e66gh
4dwotKRCwpnxTtN1z1y5t21eDIWI6wcrXj2d/4T3XjweyWb7wA4FW2L6IEw8LW+n
jwbKfuowwxFcIzZpTyOFnKf/D4b47iORxd/lmZvLMojvOq7AaHeSsYWd283PNd4U
U8IHlM/Q1bmgipVkU2drtarpw9eql/xfrQJ+9KEaeKGo1Wk+++mzQFm7XsO9zI/0
1SOskQuCFObeFJD4NTg+DHQZEZbpAdJwtYjyMYguUtDC3cJNQzQexQwUXLA8uGD/
yrJYT2CQIPT3rdHBI+nDQJx0/tfWfVlBZGus/SCe+k571fJLZiH0uagLG9r2wL9G
L4MKzGiah5C2sHWA8cEsExHQU4JYwcVvzBNsORHvgFDSUCwKlyQSTpaqU5yjAvdM
i6hsFWU+E7qJlRJ3/3iSVgyxGW4hdnReGte4rwFaniahZvbn3FWEUPJLRUiBZjAR
3UVzMepQ0tLTaE/fsgOyajVSlVKhdMRqwujVmu6tJAMp56MEt7qmb2Tw81wsQBS7
ZsD82qvCJ20P78yxUnGSPn2atyjYqBzGF54M2B78oi/U37Gn7VU1tQr7YbLAcDGd
Sps4XV9Wht3INKoFotR7wYJBGOqBWNluj+i+YTYeUmeqw5wJFepn98KkYtvmVUXt
K6jRa6NXCialAl04QrBObI1hoyJYMu2p7cxW1uYfbGmDgh/5hhk9ygZT14WbYgnV
cXa/6mZ3x06w0DX6a8vIXUd7+eprqRPjKDYCcFrobfhrFwX0v+8cWLrVbgrIUZ2i
x4BH5Nm6Y6WmoJjyYuRAex7sH10V1R4Cuop+7tO+ouXcnzbiVEyLmFoFjANvQceP
IMRNnW5bn4ZI/joOCWypNTvBARoRJ9R5xzIN+R2ES4sNH01SvhOKy+mcm87PiXSs
y7zXAMB1qW2jeP32itG6B6GCcoUi+sklTJj5oVqKmmryH5SJlZew0HDu/IuupK08
/eXMUOVbIc7BHj503E5BmeP3oqkip/nREa10VXB6L/2+GfIQ5Q5tycp/nGMiTD6M
u03u1OoDlG4CEQKbPeajLSb1YJCzljgO1fq51kZrENtEtXea1hwnfRUWZY9G7ojV
fEzV+yBnWkxkUWwYteJXe5hFOk7wDioO8uyWEQB8IleLkqsLqUuJn1AxEo94JWo7
oprX0hyf+xgRFZy03KCxZS3gQSqaWTCw48VLHpz9E5znN7NpOfqZzsrJUdT2vMBx
ydWiZKE6k1fH5UWu/04wW2vRz4u+/dAsC7ZkQm9SmuWy8VeWlhBLi7F40pwVp5dV
qvLQ0CmXvOR9P8fy+2ajg+FD7lrMFa2ln+4kjG3SyG63bdxSGcZZixEwNmbpQYGL
17fEudJLh4KRVqAkS/nbzNgCHZv7MpX8TdaSTLpxRIsXNOTh74exCFgGVq9zJQJB
McZ9/JLEkGjAbuMJV+TVhhPgRt9kqXizbSar04UXxGeHgExAM/1DK/XVx4Ohdtjf
waBVgWQf5i/qLw0e7wnfsewGYyVzYGwzGBx4/JLhnhTqFGkDzF7kMCfcNnuyzzY/
wMIcg38ZMyUSJCDKTE2TLOLg1v84Ijp4pG3NlkN3HgsBM3jIGzQW9vcVCTwAGD3M
ispdQXuaYnrAqHddXTHHqVI82zxY0OxsPVVOjq7GKPvePLOrwTAXXRQs3qvef1yH
5m5uEH2QTYWMKdN63rgmuOBDx1UpiM4mnwuw3IvcMM7ZFP5lj7kMKACsAPttBA21
KP6QZDRcuP6o14FFhEvoF/aFWdSOJStTgK2/lcWU6ELqTfqfz5xTM/j1uhH91yRe
0jY1fAV0Kr+vBpUxD8S5B8f2P4ZwIWLSZ6A3Zuh+rEJSMgyIS9VfmMG4nZ3Tmc+V
6xLSSOUZqjiGQjLsGBoU4e4uyGbeXoniIjF7mq2zBA/7eiUOQzdRKLbpmV4plYLr
wFJqQoxkURt0ewit2jUN+DXuV/5GYNT/1rO6w6KmuOT5NJq/7SYQuKiBnHiFEHMO
+a1WdG19ZutxFtEHN/raVKye6yVuPNnHt5G/ob40yzJXxnl1mUSnWyLihrv3ZQLO
7OAzLl9eHTh2rs7FreEinlo2yOWqREiy+6pIurgmothmq7lL9u9xT+b6DNUPFGPz
6CU+u0j0SNVSiTy6R9NQJbdBnUwS/dA3NNYofuolj6s7IhZ65exwHz5OQmf/6GNQ
+d0OfMvN7DFA6oOoHv0aH6tZ8+LzRgvDSR/OhgrMeis/oq/VotUviOFZWFpgMDxY
Da/ZhH2M3TqA15e/eMG0tVtxDt66fu/+vPfqSZgAOc/myxiLeXQgRVU3bxSpzfig
SvhxlSJSOE+pzTukdru1Gq+dpI4DF+FnObeM8w999F6KHV4FScEBWhuZX6bmHcsN
VGqqDCe5GPgQvfbitX7khK/KlvCReAdVuUfxpylIhcTPKR+yFw4K8OLLqZ5vmlOg
41pzBECi6EVZTUooc9DzTgyBKlhC3JUdG5mkGgydj0hmZP9KDau5DyP9sAmM8GhX
P+jqGszBFOQNlzWeL6Q7xD4OlJUbOFBwlqJYLiGRTdFmRqMfO4NyYnhmHuMFupda
RTX2uNOd6Qh3aFAEP1390CcMaWxQIZs47cQNof65sKaI7uH8MJ0nJLuEL0SRfezM
nQtAKZ6BhT1QIQU/jn7aK8B305MfYuDEJazr9M7yhK8OwJhuI8TWMBxpfXyR6TEl
di8KIu3XwejGfqigcOUVwoBexAd8arI7+ebjnriPDNLrnl0iGimZ/SUYhGGJ4wQH
ywrRPu1YQLjgy2piOaW77I3PN+okFS2HQR4yG6IRbqiFMMGUeKYZVs/+tWjC+dUI
QdCV6n0Xl9qxyJ5aIgzJDSnkQT/2FYl8XMVfoL6Do6Hne6p5AK17y4yZ7J4N+Txa
9Yq/vG5tGDKdSAGBmXNX31Gsz/6CprF691D0e2lpXDeJp5txa0KULRddJrWWkSUx
UV8mVBPc9j4Vi0a/f8EHk3/00lLjOmx3JWIzMNLaDpm8UCa5STJML9z3TesNQPL5
nMOuUWsFLdqQMpZ02kHft3djmrze/t/LnSTYq7WvIPJWvy1Eampv8MHOdtAsDPWF
I0h1v2LaGHMfFVDMddB4O5AXKJV0xLnDF9661La0PHstrmNeQoHFOPWxhFcQGkoB
CSBrg30I93RrdYCnXKbvJ9cgbK415fmAuIIrmsZt/lxmgkK5UL7uCZ5AKv4yI+PT
V3tBlULJG1GMgG2pW07/WFzjQ+iiiG1ASwiqeyymb3LixP7foMn9RHpg6+1GPDrX
7c8aGN/ovr8lTF9SoEnlaqoxT65pQEgOWsLKRp4jGaFEagobSnpRbCzvXWt2XNsX
WTz80bI2V1lGMVN/NaYKMOUfDvPaOH2Dp94leojFA+SISKC7+aTMAsECRSx6EEu8
zM7gg51Em6wMpghIcGCiqyLnzkxZ111R5ZQOR0JHpX/WUFEY6rNaOutsAs8ZtUJ8
TxKAobxpkmKKc++GEXmSxfKXb8P/mVCQLWZeRAjRfTA1CKn8OhqFWsU3IKdYyXWd
r2fXVtrZX8j12Hrc1BZYWTti+PRnvo+pxdMRYE1jtCZYkny6fn0ftCPTUxq8FvTc
+G5TJBKffnaXrhybCazrVOV1Du2Ncum6ytXew9r4ILRMLj8zl74n6Mx5/Chde4Sv
maer8qqrdGi+6h0InJ22odc37DJHyCsg7hYCWHku+XX7fG8Lrp6JFRovyPH/Wq4w
VATQ9Q4Z+lvvoVsChhIjX8DLFAU7ZDwRiSGw8V57bTj+CPTNd4mN6BhNQzlBgmZP
L9PwomhmUjp6T61LxzSpf8Cy1E9/xcSFHAjsgrZBWg/swayG4o/Vx7kIMGVc1o5r
ZO2CgeCheBz8WV4BqcOaS4q/gzzJZM9zyX39QmoUb0LlI5e6v6jlC7DiLFSnK6OW
Dz+HUD0UJdPEbPC9AUf2NdtDoANY27XyxNfDXStu6NkB7koKhNN065l0RjdQ1tuG
1FE7W90FtuaCR4i+M2IqeMAcKYAXf49Jg5XJ6AEWo83KWPVhJ3Ecd4m9UPOXnS3j
LwMYCcjjZpQECvHwTfCx6732H3XQcCnklRMGwGg/kIdiJvl+x8TbB1yHS/nHiasa
EYYxD7o48EL377NSvWIok7eiJ5fObmfT9ajaKdOxvc1F7kaf5rnfvPiCuSoy16RS
ncmNcsJepVj2MjQK+jS1CXBgP6UfN5eqmYAqf+xUd6RRonhglnTMwX34NzUTdHyq
wkeG+qFOXe/qAzX0oo4fO49QlFyaqP+jvV7oHFrrPQfdZYx0TggT+w/NXDMQqoDF
vzTpGFy4NTo8GjhlysBvWbhaFWsbl24LBt9NrHHCzJdADkH64Y6GAVHDWrs3pK03
1f6dKqsuxwhiA5OfcHmIaAoHOWeBMjkKVjBPEUijcVhLAi9/9b1yJ+3dyd0hYuea
SAveB2J9ij0+UsNN7pH1WKOrPdCbIBgAO95nYOud3/YQaLEHj/BHIZqOqNTQRqIq
mfyXTeGbPDK/Z8mhGKfHt4eMXtmJ2SaNxrl787FXm/SvyPfJbBUFR13yc1SMwIj7
vFsDrFeX6d2cnJ1IXyvB4vdJ6bJG3PmVYs/89rDuqj1eLMSGIBr6QGtXCpzeGwGQ
4DQIUUCRS8CCwlyBfC6RgFV5BI+QeriP4JO9n/Akp2ZEubILIXyHLj0vYScXTmSO
AS7ue3JImTEZj58eC2nSwGx7DPVtFuX5OO4C6ZKdL6wg6vPNSR3yjUkLdDcAghzi
bW3f7f9TRCW1bQcIYnNo0uvR12IeECuxDOPzVJ8oJdnAKDNiSXw6kUrvfDoDGL7J
nf3uAx0g378XbjeZz7d98H3t8n91Aiugz1WR4iGR47jvDVzPV8t5VcWvDEnJvFnv
3GWxlET10TVvNXeM91Tp8ElppCLBPME5TxjJ765zxTnYzgDkagIU1muOWr6PeuUw
jo10GrRsUUwy4OdosKhmA7JhAFJGUD+Inc6QEnGtDii8LqLF77/1iYLKrDj3+Gkd
PJF121kPuxgz61aRg40C5G/wn5UZGNkiy/Joyl9WfGQ1IQdCaej6X1HCZK0Dl81G
8IY4Or7/lCBP6tTS8U9Us4y2Vd3vWu9WrB+6pP83yD6MWmfE4c/tKaAt4tKGkpnp
DKNzwVHa6Gt7GEdZ6vbXYTurH35/aFMZDPoG2WIrEWAI9eI84y3qq/UkiBWQfW1g
wAisqZtKazd/k5nnHDnOyJ7pxqYiQ7s25cxe33M2mS8X6WkGEa5GlbV24ApiXSao
IDZ5QT+eFxKS0SaETKeqoCpxeIxju2xUy8NY4lgEOnamSvC1olbkHrwsbi2VrPhI
kHNO/WMCayGzi+26np40zCl3mdvP6ZZsBfr/wNdN6MNScD90UrzsiQ3NLSBwXKKD
b/fVfzlgbuIPsnH4gVepm7fU/EWFyhCM7ud7NajCbPQHgYpRcATBXgaX1cVtVcFY
WJAQWAmzgA++orxirgSJUNkyv/nzD407d/01NEhDSQR5AQjGXvfNbFnWshckZGjD
m6qz0pWb41nm2uUll3clS37NJf3GrsiV4t6dMvNY8P9oxJfVZuJBXN3+IxU3/bKi
aBgp3vP7Dr9ZeA5Lb32wasHoBGMlviPiqDBGXAG2kxEzsCTp+ZGjO6cA3quexO5P
nf08Qxk6YYo3+IPZtBxRvHOaIIjo1afbIKaeABRlU5AWCV6Z141f7zL4g60bCEkV
xXT9CeTF6mlyNuvJsKdnnDL89AKa/tnOS8hJ80G2t8rfVDMatF3ZgT8/ha4MVqlS
rrJtQ/ctaKHOdpxRLbt3ug9B5EionjwhaaFNMbHF/Svgm6fQ/InGTeidaLo45+aH
NvrXfh8Zapc8QQ3TU1HFJ0Avtc2Dp0ZdeAVHs6Qoqm9e+xA/g/r3tjPhgSIJQtEy
u0pBNmvQTXljsc+T+EORQW3IXH9If9Cr1+DsKtDIIMmx+QV622eGITlPdvu2ChAw
vVCf/f8Lb4aRRVT0GHVFhovmv/+W+/C0cmFm3boSKnEuSSeTnWu5bS1F/8TaposY
JopoPVXnTrnHrRxc01F2M18orR+4DP/PHuRIwNkx9AeG3R40YQJw1NpT4CYHgTOw
fCvPvNCtgPy6f58vRBxg28jjf3ixeNog1ljAyGcKzIhlc1FC7xMAGbaqQllDAAL2
J2aZ0mywb7RkJrzILB1jjTdl1pYjBsZD4/m7p8z2uSKaYQUvjENq3GMd5Yme48/G
JioQa0XphJyeM4JY117N9/SrB5cAblrV3Akel7ClJDVMAiMgEHxMVTimUwdLZMlR
fPrdbBiHxE1c0+3PW4LvjDBtsW4bxbIupkINnVPKVJzp4qRH0FPdlEbQchMBjq8E
bbkyBVG0tZqRD40zIhfQY/sgWosSj2sHkQXf+qz8oy6nVQhMdWnrS2+a1g7tJ2pj
5ZQG99UNmGCtzjrWm8Zln6cO43X8dMXaYHC6/6jCD9l8ZtlkuqMXEppxkYHGEzaF
787cuJrcw8X56/2l1ED5ma7RLxl+ODTW+P3iwMy6UKNJQTC/W6NBgrad/8n02jxS
BzJ7Uk/kMGnzzQMdtWuGptKuYQtMZQ/QP7vOrJoWsK/LK9RO+gPHxVwh0cbLUsVW
5/MJUw+I1YUKxVE9uqfU+6zfYPyr1Qt0XsnB+394LUOFOk1uDn4wL9KG3wyYS2u7
w9sUwoaPh7WgT68vfpQKitYcHSRMhtvmnqs+emdDI35Mik4m/BVBbXy6I1CAWhNo
8ylbNIqvnassAqS9e091UmErI5kMsu8gP4sqmTzhvXEf7cRIg3HTwosbG1q+AtG5
zILwEch11ALJd84dDCqyB8qeRFKyEPG5AKtbthC4o6ng6OdzuWnYnPQ9EqjoM8aX
B12nflwKDPSOXr0dQGRwuP+0yan9DjG0g9LbWA/tJkJ03T1gEsviXWPhPwPbGwru
w+/reYaKK7lgOSnwNgrlnzj14NhurReic5Z1mMIaleHsgjnteqvbcOGmce7WRZNF
gNUEQpl+g/PUNNMSUCcnRKHnxfelVtG42OgQMdExCtAlS938Og54iyFwTIysUPlO
/LKwR+EyfuXMDT0TEnLdCWYGKPgRrCBMrkLWM7IAAUsKauC/92YbUlr4617Dlfgs
BTO8B3XDUtkKFVow9E8yV4MXdgsAcqGHFby+mKw9AbmTJRiSPUqJrtXh8C3rfbok
pTt8VZmmhWYXcxirSfq4szVLb7YIHF2jZUHYBw3B/oFyVpmRTl/7o0SQuwjBJAcA
qBshZNLzYc0VSWAsu3ueL5ams2aq7EP9AvfOhONRt3G3fOu5lsqxoVL47MQzMRAq
CLck8Ta2YeG2uMAJhClcGZmZAzNVd74WuiwE7CC9GB29jeevjbfWPuEQuh7lyp0q
NoE7ZXw6cAlWEhhsoAvK4NXIzm9HotRi9swB8u3EAtKHaup5ax7NZI1NvPUy0hmS
NIrmxzBbTEr4MlU3LC6uBlfZganJuIW+NNTvmlqjx5xzCSQRm1ML7yTvP16ZAC6v
K0S0aFW+mDWbRtq6ow7QrvozZSUU0813op8ypN2frKUtsNul7jX2LeQQCdpwHCwK
4a4oVG4ZjLq4bBRlOCGu4w31MzMZwQ7i49agtGFrbOD8cbGiESW81P8RUd5KINEc
jOJ7zbnQ5qJhz0QZNpsu0X92sX0KFoHDiKNaFdZrsf99if2DJV+pehyRnO0L+Q1E
BhLD2GP2SXlC2c9SZzH6k4Hxj0zRbZxW3Ne2grxzmRGJGr82e8Zlhd+DPNyF+KsE
jehHH3oKDcAczKH7UQMsuSxmMOTpDNQB12bJV8I10wBHN+f9IcL69h1WjHhA/W37
fbXg92WMeW2bQZUpV6jwnR3KodcR8FVZIQJPQWnREwZN9jmk4rpZ4dZV/vVc7201
G6hJUYgjWqEehK4hKL1223R/3Gty76Pu5mAse3DQ5QNgkWGmnbTgU5aApxMaw3eW
jHBu5QHxzPP4AOgEWh8XFuCW2E2bD6P1kw1gXg+zvECXL2ZfqECrY8mWWb728uKe
pVrabg4j0mYkWRhEmzVIpwEglJVpFCel2LLalGxUN3+Q/o1WY5Zs+NSguU7O27JH
VLeDffvwx70j/xFavVk0cT0qeOv0Q8eZVuucspyKFQqk7lT87+LacryzbYOsaFmX
Qet8wqzNPvMPSBCHf+ISaYOPADceycxPqVUd/xlltcAQoWdbU3DMDipxCC8ZIa0a
B2Qjd/SexdN0Bp68KYnCHJx9RKe50RklYVdZOsPMnAolxuK+/8pbf/b/zxMTbpph
VeK/KgmczMiM3XkVhhZ3HwWUeWg7hL+lieQzbuvsEugpIDDeohkOH8e5G0GBYY3K
m7Y3wIsKMEe1ZxJGWGplEHohTPQaVh5XZw0H2XzDHnFgkkTl8RapUEKJSNKYJ0u0
oeorrIpoAnFyKFsNrWvqZ+5az2yMEChqVPsE5Kg3QVQdCFHbRapruuQcd+cwv47o
rAgEp9/WwE78jtC5aJk2dg9/rup3A4V2LfknZm6EiPkqAUOvBQyXbIP5e/o0SoZo
UxE8F46aSw8OJDjZbwOTlZ4GYKGEZi6wMTG8t6P92VdygQgOad1v2CpilF/3ZEHZ
THY4XTqWMujRvw5rTfBFBAmICvXU+R8dQBCvVYk4kxJXEaHJ4zhC4pPFO7/Ukcf+
mg1m0B5whh3tR36fn9tiiLBxjJWJiEg958NuSkA38ltDktSffx3qWsvMzeuadXss
66D+ZjtOKuDkFnzh1/6Jv9Khe6BrQepVau8uwofh7lmuv71nlE722WDJASvEXF6I
SNxi/j3Pvk6a6LRW39HNgI6eAWN4tAUvQXVIzPwTdaguKDfBO3CSmpKlnh1kfgvn
ASIlmK5hrIBEqKgWz3NnbxXWq4GIH1VV5V2kaAVNHttftjTopfrRYYz+sFUnvop5
5GI3X7v8pOnNKlkFOXYIa2GTy5q6j3kWLRvJpo6xCoGwCrcfAkJ63F6429hg96sd
VueOXFyR8yI5AC2J8rKwvAK0L16dgWSUOSNseg92DsWc0pyFPdBaaXU+SNwHUe29
HnkvP574ODrX4Yu7Z41UxdmMGjq8ibQbrcXwR7OYxfmSj/pPOlzkRmk2G4o898ZY
QmEzApHUumaYFOCiR+n3ztx+EKCtp9yxlnkoVBo7HWuxxasPO/9U4dXyNQDtJOmu
hMMkBQTIGWswWcDYsigByK7U5d1gNErV8nuVQVBZLdgCzsvRwMsFHzGL95eN49UY
6t2ZbLQHXopXBW5Mk3QjW7fcvjHBUiCRztiCWvqNCZT/a8/7+cSHj8c0drIAOE85
ie8x4/u1YesGlsCdLvFB+L7iqqkQUoyHUMLXuGU7udnOsuamU8TtVJdIXVvM6CvB
vHIy69fBgAGOEsojsTo+IPOrdkFD+YL4VYjSV5FJlCLi0p0SczLWbbhyGIowSTlh
xXWK+QKuGLpDqrHBXccurA6aR1Z3+P8uNllMd+oO9UpZZs7DPR6zCLHO4wO+m1Fu
gVkW0a2obxDgy8x7ztp/qNt0rXb3oMVZeorNXu18q4NtlgQIlI7PUHWa9D3s54Ud
hvTkJshzZOxx9qHT3nj6gGlwKXfKm54hOBaN1Dm2m84pCoIZew9EZb5OZNvK02+t
SiWErGxbvlY+65Z9vK/xV7NaVhRzF7oz5lk5BaGfPXWiqPym/SzTWmwz9ekLDCch
7+mu1iBmZQdquX3XFczlbzIok/ZE+Gxb9ABhXL6lqFmHgPF9HtMTrAYbBvyaenOG
dAhQ/PpFz+1yCGr+7PMAfCIPuIlUxISBfQjSvoZmBYbCf5s04y7rFSVmrAlsDV2U
C0xXQCTo/7yF0Gp5LQz2s99f17+dNjbdm6PI3sn5w2fv2wooXy3XrupriDr2ZMRE
dZSIccicuMfLZuyfJvhc0J3kVlMMDzlgfrPlCValLfMXI9WyNfJnjkmyCUMBOgKE
r/OqWTOO8g79VwdammASpb2A6VppnGUCuJZlL8zifONA5HA0U+4xFO7MY/u3tJjd
XqIVyPPUjA/cHlE4rQlOD3O+pZwNzSpYPeUlg4G8yadnam9xvn+Dp4PLAOrtSrEh
HIBVOKeFm1vRcboohMJMEoVNYRy80qeqt7KADlkE7lVLKUZxDxr9YXJ89ACnYRR/
m1R/q8Ux84mgdy27B3PE0iS4fOIGEwIO3hnuBf4YYEEGPSEbhctVcxqFHJQnZRVi
DXkvOhdWHRHe+hd7G5k11TnTZdG4ulYOyDGsWLApP4urIo2BQvE88qlhAQD1vE1J
aagepukA4NfqEg+lH3+s8pxpVtYNP/XdVieoghFKcT0BC0qLKAYhDDpBkJBSCbnZ
nzbDit9OqhM7Lzy02AZqnkP2JwTHLlVX135Xp+v1hlAazE1fF3YwId/mLaFpc0SW
ARtuncBH1SPXdcEEIRB++JAdwO8+8r8AARJtLP8FxA15pNa4oPtYHptrEenDdV2N
QQoQJf4oryNEF5rFWMXLzoxzpWu+RdfIknR6hLhmjFS7R8llDxmB/9682pntlZta
T0UeGXG7NL5xJ+JgX3e4dP8k+I4jE86YSUZeKdvvccu9/K+dbSAp/V+PQ73UzQM1
T4iSCu9EiLUBYvlFy4A0v1yXzFv+1ZH0i/YyjxOZAVTBx6cZkdNK1RoBhCI+yZNq
HgoJ23XqZOLZOyHBiJtHXLbvUDYz2WIns66YGNpj1kMIG23XzhNp2/dOjSxmlyFW
tDeBSLFpG8wEQ4vLZ+Svw/fAjCQPUv0RBvvWPnoCKWuGthdMJYhYbMPULrWEiLBM
kRjCAUKl/VxbsqbwjU4FzHHc6XeYIWazZKnK1hkfBVYXyAi+vDHo/Ti65otKeTqa
+yQlrl/P/6jvrxlzzVB3M6HKUNRreLtIOIqt+U5/AeReNgXd5M8Kr1QJc51ZPFyz
ajpsnSs9ZE5ITknpf0xnnQbhzRPpIuKPNYGfFBaUb4u4NjVRZecsxp8kxOTjokNW
nfE/L61kgNUfc2Zn5UOzbcz9KJNv4p84YOBp+YMhlpQ3CdsedfxeGcIQkwxQLTiI
Pc/19zWYS+seoXk/lohbQlZP7CBQSfq0Oa+0M4RDagfCBU6i3UmTQ+BvV5/lB7dQ
/F47D9YE8dA2W00og9NzZsxI6OmIzo2nXWdJ83hx8nXltsXLIzGEelSijO03qZKJ
WmTU8/LDrPirDJnQHWauroQ8MRL/zAUrxOoO11cOPM8SbLlzPVJH8pSDfldBs+kP
Ei0+bpEzlvJdKf+b939lgsGXdCWWuLplv2vMLsqZ1KbbYyad7M6fc+oMWFgmZB0r
6srFTc2JBpbZxi5S9xDt+Nj7bGWSjcDR8p6d8uiDrCcnyISsKHuApGeLQ0dF5PL7
IY5tdY1NS/Fsp0GIuAbz3Ub/EP8bRruhhfohNzn8axuYVrHivsSrSg50gzX3/soj
NRKRv64iHbMl9qR47ng9ajwVeaAaLyAnPKQ28ixM87KlOT7X9XEkFAMSy7aCwqjB
leUcMNVUxc6b+H+NOxWhkFZjYfDI0AmciApxbduIS5Py7BYKeANt1CtFqvRqwNE4
A5xQiClG3QbZEGHnQlMHQC75i81ZBuA95yGcc8bfsin1NMs3OC6fdTdAdBxhT488
MTEmVNWYfV27GM4mOnwARfMO1N6l4IhiuRe+2l2RAUIZPtS63pHJ/YDfNJ1vBk6G
CtUGU5WdBBmGxuOCvIGD961PbCH9/rOVZ6r1xnqV7B9XGO5Go9YBql44x5Wi2tl4
vSQHtVb7DubYWKAGBpzfIrE109KqZCsHvfD8dClRw6nyt+MV6Mt3aD5KyPbT3Z9j
QchEW+7YEWOiXCpmPYLAJxah/5u2mvk05f57WhuS7LY4gM3GnM9f7gtI+uYTc/jh
eLPEG05iAzDwBDwAR0/85XgP8ov9okfSH67xHTZulh7QysAlZY5053egFXG+ayEm
WSZXjAqYJiPgD0BALOVGEQageuCbTTkTOk2RvoJeOsJhcXpnZjuZretMsLwckWpQ
pU8uWeFycuHxrMiO9QKiWakKZ9Adox5l1P13UcaOujMdfqKMQWCbVP9KjKbtKQTU
y49FEg/ize9628hjnCTIL8W/VBIHMI01fvjTolDg1Wj23LhnlSyOQ/uQ4WU3+6UD
1JNupKDah0t0/gpTLQ6hhMYGPgIrWJsZx1IRxCuyJB9neDT5bI+A97p1jb0OtdNM
SniZVyLKTFmd+brrVXGiBRxlsRw9AeI4j6oyueEY+KrocYtJvklhQ0spLvMVgVgK
yHC2b6uMPmquBl8y3wRHegrm0nGRskcZtrlMMnLxZpnL+Gp4oGFlYsklBybem+bv
gQOQi0g6BFOu25A88cPhyqAqIfvcF9zBkchZ2H14qR1WuqBF5rByGMBol1uN+qJJ
Wp/vDqLybkMMhQ32bXfMLFo5P3lqjlID1Hpe90H9wdDAl40HLpO+UMcIf2S7lnlA
9at5vrjNmtQEAw+b9pJTE8eOarYd1vb1AVjfq4Mz32Kc1XyUJ0EQqNQtbB6OicFh
wkB8WD3nhl2MeEWu6QeepyU7Sj6/DBmfkhEkzwe0GG74yHzBxzs5uXdqpVqytY/v
WaIwyHnppLkAmy27L/ATEcB8m0iunvFO7lVqdivD/tAuQvBCnjm9n2e13dvTsp0r
zpfyvoMwFRVqhgv1Lhe8OqXHsIUNohFsJItuB6JnYuBshuCJONrzzu7Envbk5bCt
OhcKmsIZsmDh/CV3KYeWtXL4+XOpJ6qvBMwij6mDxQjubXTqs7X2D+FNHsgNuuh6
VUcK62/v5sZtHjd1R3502I327MevjlR6oSVwzkqYCSGHr7OJ9h5dvmCM4daOnLtq
Ky4jfAKNDZcrHDl3Aj+PuomT7+3baCebU/tozN+hYkRn1Z6aTSicfzOGgbnP4MSn
6eMfxeZTtJgblPx6EwrChyNsdQm8odoOBw4xu4He1SXnP+o5sT17jt2qe1sJPfou
RVR/+J0/tmzctPXgCWmPyAigYKw3YUSIzLEruNdVA5QxPBbjF+EN6yuhkhBLTH+E
FSWAd5du/GK40XOoG76MSGFPwDpAzuYLfFII8VjkaJcI0BXMkvDgzno6B8X7iYub
BM6SBC8cLYcVAUFxdch5ubTRbkNmB/E6wwzYApt2uBqSky7IgknEnR5nD+iIGkZE
MI/sssVjTSBw0K5rnPZyPMDMJQsu1cS5y4SHGr6FVqzo1QBsGuVdpKuH23tSOIHy
yWTafQ0tWJ+K8kvxfC5cDKn6uf8LGfndQTAkYxaps0XvA4bpxVFUhQQba6Hd0aHD
zIW79CsvJY++fzVd/joiEztwoUfan7d/uNWBFKQ3wueNO3/SvWtZnOzJr1jO6w2u
aWL2T1bH4JkcvNPoy2TLj+oZmCFCxw8ZttbBqpXWpgCL7GYYkjlcBdI6CFvedZs5
LxgVxuGxjx6QJXWhzYqXCfj+xkFZnHI6Y5WBTt9/rhIecGmO7YioKXMW2VYAtojH
S2d9bm15ZBfM6gusWQ7mFDM97jOk3P5+nBxahgWqVBDBa9d3A4YJNM663KRcYa2q
dQFVJ1gp+i+oc0F80xQb2hrRiiLFkeqDToYj2wGMjz4mOszuDCEQ/KrlTF0AK0mV
PGPAECtpNoRexgbWXJD5x9fkpejTIfMD20ZIFEJKHwqUBHMLHUHVbdEiTPP2RHxR
LhwUEq6Cv4IVzilGBHNr4910jAjQ4ZFdakZegVI7RFM5WQBasa2SpTbRYnKdpZMA
2Lyj55ZfkzeUrZztv/XsHQVhBQgOXpJgAy9ZWRlzflIrP3cWjt8DcpCiayfY0ZgB
uL33YLEam1Ols//aT/9vopRvr9VMvZybcAG6rK/g3hTSCoN04+O/0BWgNpGLMxfG
NXGpkOhyuGfqvL8hwGLsTWwfcQUDwVCS6ny1qk0hLtquWAD9ai/zaIzmx2TiPX4v
T3VVbNU2akcMKAW2O2KxXlmzKhSzN7sCPWCd7LlqLRUHmD5dl3YDRF0aajX0hgdn
DfaXIRXqQ+BR8r3hgkcDOySzeEyAtwBQB2rfGpwt33jO0H0oXOkU2tATOwNjuvUP
cNoNKt/O+vE/6/I2tdJeRwUgDTpJZgNYGq9A7nn7t0A4PJZWYtUFpedYlQVv7syn
AvecnUajAQxwdIM64ZUDJZf/d8oDCkjH/U0f4REIV4kiHOIKBtxbT3uL0emY4sMN
pytCgyBbUh9dwOfdiRrcG244IMifHBKo51zZFvQ+/ar/ida1XaLoWTu5logQmJd1
+beBztkEbNzhF2IcUrYajYby2ONg6g2Py59fuzYfdNU31V0Tsw2+OQi+f4l1Kvas
Bj2SVFE0wBqz3fRKffCsyNzBmM7MREtkXlHqqxw9QjjY3XvnMYS6DwDmj634NpvD
SZhgRa922GSCjmoLRLe6LQz0qKu5l5enTW951aytZrD8WJ5YEkhtul+wmBYPI+h1
Uaq7K8Lb/zbRsaRZRZIYrFcJ5hvovQWNFx3L01GxpnbDpb402qZZgGx6Qv8llqyG
MHX9YiO8JKiBWNF6xlPFk1O31/9m7IdwstlnfXSY5piQ4oMWW6VZDDluVK5Eum85
nlzC1DCGkQvDtcaJv4ugfL0tXR2Hf5tCZAOf6yNYaukEeHLCUPO1ZKIQLi6WnZFQ
ZDhnl00vGVN2uL+iZgYQn6l9NP9VAxVQ4x3YAMo3rzD4w230UkFB/k+k9NsrcRT0
oXdNxkaaQhjk4lUo6bwDw5H2ywihUVdGkYTQVDlOlw1gOrVbrnsH+ZY7HnqUU0O8
Bacp4Jpf2L6ZJOeBn7LMmCt+Kj3hpvBVT0JmCltVowx0sA6O6j89TLuFs0WW1Q4d
yfJqFpQru4FW59UgFJCE12VDrfLOQVtUFuS3p0dITOnUiFv4l05Q4eJjfByvnV67
BH5QqlUKwRqmrJqqenzhnjKM7x1/FfMKGlWnzhVoSarkhcloe+2sH9SLAUlWey/Z
FcI8RZs4vZQ3sJOXa3aiaHInJUWzzfknIF+gCN0F5z/PgO3FIvloE4Fzv0mCPfBs
4/vaEuMY59NabMkVNrmVHrTA4UZDAzR/Q4gCfdTPDDmJF93nw99Opv7S5aRCceE7
DabtBmOqVRRmXIxwgty1/klyuLpeboHBTQPQgPieXDrkOxe7mBJnrmbzQOCtFmQ6
UJ2wzCtXpF9usuLii5YDGQIj6jNxOWZt8fK6viVYHrsg9trlpDSos3ieS6fvDRpC
eXs5bHSb5dcndppLlBoAGykSxF77Rp+50OMAEsiH4SKmVvB2axZEM/mFkX+0DQtb
GxdR0VU45bzt3HVahKxOEq7aEYFeM6vbBN8/f2EJozMS0SVkq3lzd0OmXjBX2m6q
qJdUtx9erikX8hMEDXqUlhmG9t6U9mitf0cwkVV5CYk4yNBQdv2ZwXUeHAPkA67f
o+GsVOOJRiT7POBdqOC2I6/da2kfRRxcg+BcNIWzk2PIPD/BVr/X+r2ldVgGE17T
tD4G9zncZbT8bXf3JX1uFtiPymKEpg/IkPvFcSsqAEPG5dUj2SUmb05g7N+C9I2U
BdJLQ11q6NkqR101vFifcLFrRCTiJynFYasGahLsX/tIqQh+wFYVBv4vFMwFEXhi
YbDuB/so91DZNppj1inhixvAdTqlJugNwdtoONKF1X7Kj9UWoOVKPVZWFy/cCWxJ
O7NJ66tf6I0M/eIEOVP3OJGWsYBDjZ26y01yyKbcXXnCwtFxHro4/Hv5BU8h7vT1
RG8+Ll3oXv93+Sw0L4FMxChb/o+0tXjqbrzMSLP6OSSIRl2rKrhM3nYkI1Ijdo0B
CzOMdLZ8BWwRSXgmSTRx9sOF1wuMQlwC1nOa09kDxpffg8X31Wo4qTmUuLMvccpC
DaelQzmbH6OcDkJ5bm0wxFepvNSUHyjBLOx2biHb0LQLTHBmE5VTQgBNGdlczdmb
bJUNjMcsBMSiq4rFFOMugalsRIXJVA0xQVInLmi0kHC88EZOH0bOui2M3G0HZIRA
2Ot4UFVQx6W8OEXT5waYrV+8n16C1vlngTUeWs4d3E/AyGST4lW9QhGADqu1VZFa
J8ON2Rmhd3Ka1ABUX/6drl63MBz7l5LNAawuICukQ2jIShxeVTRsV5KUkTSfGgP/
RTZo4fuCzgRjvMy2puGzLnngFcLpX4NLlCdihfXqqDymi3JOKgY5brio5DLUqpmG
zunotfgxa9gHQFUcxrzWZWRwi4Te2hwacLNeBoTGpmmCZT7abxZNBLCjB4b5RGHM
5vKwRY2H939vIuiGkn8HAy3EjYlofn9j3r7z6wy37mUtha/nNB5KDN8yvsv22BAH
j8bn8dNWYXb0HllTtJiowg2kRrxc0c5uNpF6ZOpFnQe0uuwGpinErTFkKPifAE3U
Ol5X+o/ZmGS/gpbIpM4mdIejw/u1sG2gBCXgYaly7PKiclToNxApjiylHxaYhqFO
9h2t+LdQCIdyLsMtfQqqrfn13FLXd/OVYGJSEH6h9pb4xJaUblCf1CVFmdok68mr
ytJ6Td5lo5+aKUJouhtCK4/ex2s6EkXSOa4TjkbAd8pK7TvoAjxTBTISt/NxHR7u
horKc5vSQ1yq9HOJMd2woe3p9Ll7ux9KJOUKKzBij7bUp5m9hbCoslcEQZHmEFP1
cdnNtz546S6T/L8uYsyql7luegR5WXoHazVtK51tED7rSu3Kq7bk+kWSJwlKonGH
i1P8zRHqMqZs+qD0YBwbpGiehLMshXEyrs9u5oNOv+HbEZTxxGi3WQb1uL4pkSGs
9BnFmzKQeUwA3yaY6ETZjmYkXimp526vciJfWnn4gqOgJHGIZFWS2TMKf2V8WJYD
MlI2q3O4mvVG34Eay1ZsBPvdkZhSMSUuXMvbjh4Pz4GyOeCyqrg4by3Ph/HDvi2h
q9qCEVcUqE23NViiVdLuA9k4jI2t0vx4JesQj/ZZLxCYuTZZ1HE0UfgRfxpHFrqO
CC4kn8dKfe7225v6fIOwgZ26sUK5wRs+tu9lVxMBDF1pcxqSevZtEaucbEEs36m6
5YL8WrMLb4m6I0YXu1mhSy92SjCv5Wxy3r3bAhr0gfyb3jIwleSR00s3M2V/veei
zghP1pqHKFSR8IfEME9/3AxZrjzYmt7pUI1RHmZUA5zDpuLKFbBqzfZRPBik1fxN
yRKXuShB0fOJ1RLayt0zXxIL1Uq/bAUbk24Cz5dOmCb0GNcrdmeoabKXTv4iYxia
TecTBsetr1xSPMsXiXAdWxb+4OOu5gg71KEFAfSSM18tpjGEQoFksFWwYjYMHxJB
bhMjUHgsFZwLSFwjA1QqMjPGUBiB2NfAnwxyuNtkkDOxxLgLn/+y98DNPUKd1bst
SPufhDa8L3xiAyve8r7SgYTa0y2XAtyAFdnXVKyYTIAI246DtqXsBrQ53VHMIG6D
4y0CPp8bYe18iVdLE8d+kKeLpZxhEKp0ReOOKImiX3oazJg728HFUCxMLKZcdw9H
eZbxyOO9A8N0e7kit7BeOdeXHNpsxSg7eWPDvC60POSvkGWlwvb6gYgk/cpC+Q75
YOZZKyi3ZKZA8rk7z/Y01qyq7TJX9ROQ+Kqf3WyWS4xTY0Kv9BNAg6tvIY7GhHuF
nnhwt2m8Y6OXVInDCkUCiG64NAnbpruYqEMb95uU9iIxevnXlmnaudlDxv8Nl5xp
D8ltg4IF+CzDUYqc1gyUWx6ZURUaL5y7H/OLMTXUM8FFjPgUwv5NxVPsGamUFICY
Gy4IP+gMIBAWD/RqaZaWjucFS0DJkpm1iNb1YvWOnN/uERxvEOIHi1GgpLTt0Yp/
1ZXnp71ozBD1gRBbeK/mX+jNkm2PPfK8VjmJMoKPziyaOd6bT6UM1fUAhq7Yg3i4
enMIThBc5Im61kkewPf/Q1DSHr2uTM3ylWUcYCg27j0fT8FBwUV/e19+OJ5voLQC
t6asLobREFhuxgxXqLSBuEz1Bwcz6cEOoN26HYLGhpAaPHiC5OmJZ4zhW6IPD0Xy
g9zxVy+444n0WmfyGMTmN4gWLWTFy79goyVD37z8COAiXnhqE3ByX4XEZXQgGPlf
WY3F2nLa4GcrO5xB0CggJkv2fkI4Sn2cZeyRt9PwFfyn6SA1GB28zkygVhvJA/dl
FGuQTIZrqeyhACzQMiP+j16RdaN4gcsptdSR0BuYkk83HOKE+EyJXKnvso8P2U6C
MNfvEuPiUBm0GW1+YmrEykFER6fyRMiRfT8Skthe4I91q1vkfLyz1ux9o1J8c6iL
Cr32SmabllJ+djzHBQF0ouopChtpQWZ66tNAZClSdthGL51G/8Z/q6mtfMLwWFj6
lUXbwp/AX0aT+uYVtYg6houb4A5Mkcn4R6F8O5p6+9J8PefRw5AR3Nzpy5RhenWX
tvrW8fcKW1KPE9ArXLFQFqjAOoMSwmpuBUZw5wT7DydIIcPPlAvIOApoABmuHnym
oScfYpUilE8FhEOeTY0aIbIVLGTsYfP2ISFlLD1GeGrHt1Jf1ubyIPt69gbsQiJ1
xX/pk0mxdCKeHm7ZGaurJNju4GaAmPBTbRj7ExAoDQbrzgv1d83gUCESeFlQKiFS
ld0XAp41OZsOSYtWFy51jMBXJ/gQd2oakDwz1JvjEtwe4dkK9r+4NKOJbfIWauwM
AXcKhDsK+fMX54gZcUeLC3MQwgXLa6X8Ps6wcFiQVMUzmcRXvhO7KpG+z3ovHTVy
HGUA4On9fdQHeiqREu1xJStX6OZ/tsGSk8XORKvOx2cfgGDFD2+1F/BhY6EQmxvw
7Yjtd9WEYUA3P33TkJq9t0N3mLdrcdRasCks8rfvqZTXu/2lHc4BnciUpwmFgy1n
lEi3FX5xr4sfqFQa53WMlyrXvbFWJsS6R6ffFzACY6pjxJK24pFE3xK4PhEixwjT
1SIFvDBkm1u9omyyXozeJyMdi/s0P9MY2sNrhxy+cX05Oxp0u76SQvSAJkYk8sfV
v8rI3M/UXpnVHu9fa5xp7oA4agDAeSuwMaM7g3+l9MFxneLAxEqAWv87L7Eqv5Xl
tobajJBIt16Zpt5jh75jdTQX+EiBMoTMhfcv9viqD6bU7rqyctR9Q45WU3H7wReE
BkwX9ewgh0pkt/u0sOYgXOhviRqO9LfGh6fR2IvutfYb3rG/nnsx8jOEVUnyaqIe
Dy2yqcf+YUhJ4MZVhIDg/jQ+ziFgmZ3HbevPXM7ihWk2vanLQpYl3zPAWezESrWJ
Wp6WvF+vMmCCJoUkjqaNxtzjyIeUGvE0hoki39ZxGnhvb2FZ50m0ILMBl2IDkUQy
O1yrAo2GijjEs2JoVcyMS1CwB+x7OGlgL8/Z4omQy5zY2ce6XvMo3DEc3943bVnW
G46GObe9fq36q1clSSY9CiaGm6fkYQ6faoDLKqpcrffOv7n6/30wbi07ZfD6VMjq
/ybzbcLqtKk6IJKBRSNojt4jVBw76VTjiJeG1DfyK1bcj2ABxVBxAP9pwQsncw7R
XlFlAgTJNhAK68weU40+94knnfT0+G0o3OgX3oNGQ59IAgbw+M+UR8a1zOb1HwbE
DvvtLFuNxnw91A/Sc2hmzqSqoz2xEUN/enXSBY45KXt4aTZJkbj9ACStsoMyVIbS
Sn72MpN7yDKIlaoxWA+rwE9iMZo9wPbv3hbRI2VNWm8fgxhRY1DLbIKg/nmdJwww
P4hM8l83vjFu94srDZqqATjFpLB1BmGXuFnzv4YNYvsNN3QcoVQZF0VgVpLWKNgw
tAsUpW+ZDJOq17n22AjzQQntIDQg0S/rHd2Yhw1rdWC3WkihD7hh4JqEm6freBAz
YlhHxB72wWILoI85By3IlhI4sPe3AHaNlB44VvmTKl7r32sUWzeRE2caMtd5Z2pj
z3cREr12grw1fK+yhrfklhReMFfMsbQxbFJPtQATp/Xl+WnADgC8HcOU8UGIalsk
j8sPyxDRSdi4qvnCQAHj+G3cqekisdjcU8u/i6xtSedBBmZaNNYy6qIs1tWACtnc
kdwd84xGfSMV/GddA33+lt3FRo1/4m0Sw2+zkcns5dqX+DwydlZZ0fj/GWdQD2Gv
Ptxgs5dCiB3TG4b964aZTPKoFqgp9XrK0oiXRqAzr0Xo9AN6PuepDWXDWF1StrLT
jauSefNDjBu1fxtDWGcWtE1fptBVsJxZgcCWYEqLv+k89A1PGEm0jAV8vgPWcgBs
o10Z0mYd/BvxoA3ansss/nS37b/KRjs9CkkL2GMR+8wZquH9CiD/GfhCD7VJ0vKM
SMSnyDQruKvR/zuGyeAwm/Mjbi0Y8VmJVEDyGzCnOpX4PUv4VUOuopoW0X4iocB9
efrIt/I/7y8UsZn8Tc+KI9a2ju1szRaMcSMLE4Zlo3w5jN6z+yiedgwGe69KqrDr
OLJT349YN9IOe+56I9eVbaZQaEoPYqViA1SX0Tas+n8ceDQ1BVS43v8iKK7gA0uu
crP6yC1zQ4ia2nwAS6DdAWJ3lD62pNE+8yihBvCcV3kXXq8knItR78AfMH8ACbsO
UsOZ72KvUaZs2u7shb2Vqjj8YtaJEG5QBCU6cf9yXUTuL4e5KMgsFO4a8MW8DvvY
ZUcFCqCQA1tDLYWE5JfrUuL9DYVsUc5luz07TVGsdPOczM8ZUOgAG4IDg435v23q
N8yDA1lwRngRaneDmRgGIQlQ6n+h7TIYXaWB/fDBsrAXHt+RxI4ZPtF0FTDEnHs8
rtTpwHxROrX9ZuPpmEE3DBjNo/77S+t7ZfuhZXqQNIelz8rY1z5N/A5NOd6yy4xr
fv3/sGqjZSPBaK9WMn9ohP6Orvp+mwEpblCweGS6Uy/+GrHMSBwYZpsQ5hEPBrx7
jvpAbgL8skW/lb2DsHv0hAdku1LP6JMlfTUKL6ZVoXdNsG9GgtWhaQJMzk0a9no6
sMljpgKgSfNFAPgINRjoTelOZ6/c6xv+miT9vekh10iycrKPipBT2W1MQw//TM1v
0rtAROFpbbrUC06K3f4GvuRjx6p7IFxiBaa9Wk9LlfUp78xtNmHdblFev23/LGJo
rmO6PiezwclpjdkcWyyYsZ4xXQKNLXaNs80xp8/LiydmRnSh2A+fR/vWaSD8/cVF
BxHZJ6DgSkUrJksNOEQsnmnnxQC0rFxMkEXGbz1qiJWhg3XxJS39lFZGy+Y2Yyp8
B4mEMEOJkkSLPY/VVeqUdvpVQWpmTEp9jqDmlouoRuFGr0AafgtnhNdgcSDaxUQk
DPLF8oOZ7qa7b1RaY4auqmz4HE3FjTWDfPy5PJJ2femPdnslp7Q9y48avPUyhgZ5
XoQw1Z5HcD7PNeoIb7Q4E9TiaC2A4Xce6Dto6hEGNvWT+mUm9h9GIjaSQeSSM67/
4PYJdj2SChWUMpoUrcG2Ox+4m2keZqzBQulCordG7iZxd3Qc3xxleJtXAk7j67fT
L7DF19EguX7lBthaae/qAIyqkianyXxkZ71lplfZx9V8sAJqSyRAq0Ky6wsuXFAK
ZwkNz+0klKmhhmSVEI9HG2G96fEU5IdO5/7LqU/F0j74i2KjPSzXv8eoeRi3byX6
IgaTnqiyop2ofPRsGE2QHnh6HCk1Gt8bW4Eu53MrWwgizZq6gnQdmuj4X0x+TNVJ
fpnTCCxqaAG1qHtx0qBh5KKOllivO4snA7g6g2wo16y1TdRGSvc2Ym2BMw3rAdkO
/88LHTfUVlBZa24J//Q5AXHReKaLUuK2IWWsMdwo9BLwwEMUcGL4xGNv5XmvE7Ou
K33oWjU37Zo31haCpam/O5WARdBh8GZVCOGCBlOagQXLVFYZOtD4RXnlUFow4YFD
gwF/Yq8T8JDqYrNL3gHz+3fSfMQMxWSN1pBQ53ATq6h6sT5frjPoyM8CklvLE8Pp
MWcfJTnePKGX0RbxOReAItm4TUTULkDok2YKzym17vUxrEBxl7E0BS5L4vEUyor8
GvVatNlnrFodFXX2i3yt32h2mhgpLzXr371mDSZv1wszu6Q4vyOgJt8G24cIQE0Y
aHboYzYxtcCSVlNlrJEnCASZdyd7R/Gdlbz5xhaJrJficVIxETg0V+cGwlEKEGwz
MVl/wB6dYQbchvN7uqqLi8NMobTXK3r1sEvmW56qEtVZyJg20PX8i17tNCRvDhaJ
AxIXU8edIR5tXdva3MMr8bNIoabNbfV+V2z7a/4Rnr5vtVPstFhxceNLyFInTnav
G39WK5n8o1AWHjEjX6QwDFXLv2YXdlWIhPCeh2zRA00y/OoXqtcI+CuExxYf3vqv
up2pMnJIR8n0FdJI7YNvOkTd53ivbyt8N8N8H0315JNjzvajV/nLKgy4Bfc4LUTa
Dby6ABqkC5ohVysFGB8BQgWpoPIGkn5gjqyC5e0mXnPBh4y3TZn1Yn6+ea7qw0C2
txwI9bKWC3s5zXLimBfjTylX9ypEkCoAREsXJx3wzvYvl5RDVhHTmJoNvOQG3xq2
sHtvefSqp6BAJH7CgpovybgaIMZo1nRznYH4blhHj9EuP/ObdicKAVReexIpv/y2
/2zwUTYoIiJpa5c+oUv9fDHdwpm1N4GUtoOw3GhlEr3jcrHH4W10CrcZIC+f8//C
tMwTXXE2voz+cHLvF8u0pQ9nPEsLI+aC2Wh177xO51aLkzbn1+wHQvJfC7lvcjFt
vV2djXs01lpi1KgaXAvxD3bG5fhmBiCw+p4hctNh8Fu9qPIzhZdFn0P0xCIbc7qP
tYYB+UT/UMzDIJsjlp0DfaXb7HsQS37+pBZcmDZzfit0nbZuZQzfNDpOSdm1q9Ld
xSTmv/fry1A3DzKuZ2g62a4NmhIzvgNUcHTgx+a8t+F+I0R97leqBd0k0H4ZqNhz
+F1M+qbFZLRx5f6o7YLYDHIIEQMfoD0O+6tgxtEJ59yVh17Ax3ItTohu9Fu3fM7p
buG1ivGQkDPpQ2LWUAI/QNVdYgWkRsK49zEEHFSNDBcUnirCSYfAxTeZGIEnIKs0
MTgA809rk3K76vOjUmoi+nZjCmSGM1iq6ESQEoDss9/Hc4ka/guCMI2RHB+Sc2vB
60exp4AmoQ3Xb/UdqTsdwGNYjAQ4XXmowGLbRNURHWUlf94Kux5IGtYugWlC5pdS
fuYkoJpytX5I9IRz//cMB24Zb91r1eEJnoWtdI7dSY7FuLTIkhehnyW/WfiAIlDu
996xhtcIFbuqOGfOaQxbMCqSFnOEssxbd9CVW1jlaMbwFZp2Yj/PI0TTF5kEfX45
11Li/QzaIO9+Rw8socAKFpFnEb0NV86d4jLpUXPHGqk/gFGH+LX/MFYSSI8K0YGl
LRP3HxzeI8OCEVx9HFQX/R2cgjJqjwr4vXBW/eEU9IiignjI14Ux4mYJJ16V4JQt
i1k7tvSga+2kmnpdN4rT9qFNatMMs06GTgc52YWlEqEMxCTPmy2KXWUmOhzT/JXM
EA9WHB8TVHijQr94gdH/se9Ky0HDxI9NDEzDD325jpOdC/vdsJP9onu6lG79SLqP
9/A3dvtBQ+rADAzK8BBuJB+kMA9cfWx5lssWuDZrEkuCp77jbOaw/l8JcVH+Yuah
7DOyL8YVcxIdkDsfxlyqlvv8y4nj+tnD36VfMrR72RG1u2IYx2YkRnNQc137yJDw
3X6E40ljfWBA2BRCjmtZ2+Jk3x855SssQpG98qyeNtD/KUhknV3DOkTxrTGQL+En
13fZ52zWHKglvomCL+IhvBWH138hFLUJDdI4DADxxrIT6sviWHzF5lOcneN3Vpct
nVGILP7zTpW7nB1GN/cEHgFkVHz1kiKCEwhq+0m9P4otdRnhesGBEbghH8pclWUa
G3La7DzCgkywuxeJE8YKogWaKWqHkLNLNh2QPeL0IvHD9UiwDcFF7uSJpS2AkJXh
g7ns+PVc18kifHAx1ZD1NgIiKAji15s6rSUBqZ7iiLJxm+bnBSG/OCivCWoeCzmx
w5dD+qc3F8tzlOmtMfMPvC+gjn3P1FfX9v5v8mnSB9Q54/LK8cjoAw3lLaNO/Wp1
1MRg2IzIse95vftCeIeV70hfUrJDeu+fj7nIA0lUXlE9thVwHqAlKCZcJSYVS36M
yentasT8c7pGX7AD2xiYJn02OudlfZpf3AJdrKFpdXJz/r/xAzlM/etsp2JCNEel
no6CZDtoh2v6Gs/clwzXjpsK+SAB7NEjQAYNio5v3R7YUL0vOF7YYGvTWHeoenp5
QSB7+zMLuFzZxPO4eM91+mr6GSluYj6FAEeAUrZEL9uNnlNXJkbMU9AtPQesnoVt
STewRVZ20h1VlbWnyxhzPP3qFd7WpblGnJbSkK9J1i14fd6Fu7B23sfI846LgrRf
u9Jn2MUZi5buKtIl2wXqE9hU880zr6MlGrtUvgPUMEyE7iduLYGrYDSlg6t2AI/b
N0Zsqy3QVvj1gocqBGFeRJE2xwjSKjAQUU5ZtRkAObLi0Pk2Y8AQXmA0/Rlw2X5z
DWE54Kqq/xqGhgyGitoqCBTDRmO1nazyiJZMiY0pypx2jbG+EfHaCtY6lS7/xLZ7
Rdmc6IRiMkIs/RjqII12+calAd9tk0ikhM3+hStjBKcgHxt+Frur3Lq1HhJzKeIO
HiM6+C7kTmP6zNbLXZcrJoM3S93mS8LLVpjQ+PxmLD5REKIcg6QdJJiB/cTfyR2J
mHmaI0ybQPyGRmyTddOhSVoZgxTYKmlCXaQjMT77TaauRHinmMQJ9AW9/WdnWfgq
3eSF+XefXyEzGTTXcsF6x2a3c4dLHJM1xzFqwrjWSeHYIASUrgwCxBV7uoKTYVsa
NhuzW5BmxoR6KlANEj9D0ED+gzhNTegXNLHmZSm8zsNZsyZseQmyhr++M0LSgQD0
ar9BcJWI2LBhjt6RCfcU9fmcNVsPXNLv1Inwecn4xgb62Qt0mVWzqyOw6hrP5ET6
cTvndP4CDGY9Qy9oQ4NQcNTLqn468yI+2DqtFmHfI2bPU/4pHV6MhmfNysgcz4Bp
XXV/JL8LB3ctwn327YmrAb89sn4iop5KkcWI3EgI7E85/pdrHVMOkfOy62soSU1M
8LJDeGRlRzOIq3Jxlf38/iHkIUTfZSj9zI3KzluQzfMCgxj39lyOdXl0fcm6keiF
5twdUQaUJWkI0Vy4bkf8Ybk4Kk24bjOmqqnIhCWrBd3GPrkJhZHp4V67INizYXBI
rGm7AR1RRAtVc5zKvS767Q9pnhnvKfADqcbifcUkpCvYmIHt9oBqKxiYNsZYlsyr
xwrrzIGZJceYC7Us8R8lP9bKsCt4PX75WkIXz6WLQzmutw805exGMXa6NTpB+Z5y
sqzuXypa0bo53EaaB47sCzaNDPQBZuXb3L1J7FMIpxvLvg2CuKi4TlVSJX0Yn5zG
YVAPTdMLhSN4JZUk3hCqK86w54PgPUrpweZ0ZzxaKqbdagXk4Y+xtxjt6VGHtZ/Z
ClQBLu2dmcGHRGeSmuyFBpLp99TNELyAnGpQT0jN8KqL4ACc9mnjsRJFBiBTUNOM
rHw0YDN3+R1TOMMM1/80XeTJ6z+3fGBokU9DESGAtV9R+btxaUmuET1eKiWTIHds
Ozf7rVlEYHkxPwJVxvgVHZUUSl6VSoiQjXcsw/NkhPjSdszt33/b0ofScOJ1kVr1
oHYrVuK9EZrcr03KB2wnAORD2JHeQvwdnMhu+sV+PrUcjaq2lgdV7Dd3iTNHf+7J
udEgUB5Npp618eFLQ3Dmra+f62eUmMb5c6COiTCJ6pYIaSdzu8SMNAeKNOaqDNkC
Ojs1w2gHhp+89eOFpEzz6oLenG8K20fILaUFEybmWNLxGeR4GTXrqx+B688QQCm1
4OuUzLsGNJm+ATkFYfei0M/s5Ekd7Z7yqA4Fi8skTWzJ620N/Y6YE9RxVnyrmIlO
LT+VwvKd/BH9N5pBBFS0xdqNX5r1vC+wnEulOC8d/JOQRrUOisDv9QzSFEh5kPiN
tLvtXPqWTE77jrgVGuLn8XRHcAgRFwaVcLjOqNNZUwYH+TAHnVlY7BGT4LyyZyTH
ss0USZh1uAPLE8RILWF3KiazYTO5xDatwKX50WVyrIyZshWoj6P81NSxxn2TRIbf
N0RuWGriMURbrGwviL/cGs+GLy4ttkcJd0ikCFXIHMFHX1utFGA/yb4bsjzzCwek
S0TJrqz7wMu2idksv1eJv/MxFIdlwp6/rK549YJ+WNclzFcURADrzOZzdDDTislK
ncH6RpXBt4EMvaBoEZvALHzhriyo+Dr9PNZjuaamaek/0NZsCUt7mpnZ5p2s4cSS
e3dQoKNJYg7txQ9I7ZGKPjQtDPhr7LMLQPo7ubYEzbhpvEWWeCWY7eQDWEVx9fdJ
cN7XU5lyawWQ8PXYm5el4zucwuKmf31h2NtVt5ECE2FAoHSPNJa0XhkCz7mBZKWO
l2sn0qjRJ4zLZ37qLVqH9N4xW5QNNbjAP9EQGgw5Q6jY2yR7dbPrmHkTB/fy9/u/
52BfRkm20SPcrWjZeqBQNMsPjV5/sEqSUFihXArOSRZ1+ZJiAaF6MQRxJV/OCKOx
ZSHVE7Nx48ctPi/vdicpvQ9A9AjwlZ24sOAfxwWDWTTOqSXIjg1CU6W3U/pwM801
mWOlgFApthg+WgG4ow4a5T9AA5IioxDtwonParaH3vKsPql3tuz7ohH16IQoCDAp
+hSYPX/rf5kxeKlXC9RU8OLgC6pDHORc5dhoDJgMBea00tTmK9v03lNhV3jiejo0
Bc5I0KFsojItAMqYGHLYqorquojBhvJ2Uw08zs3actxsIBzKtfmEHTzlg9l3fM7c
Qxn/LZsbf99QFtO/P6T1kSfV9PDJ3IGRWapiahsKvBMuOx9zTKw7I9cp/5qKtdlY
n1Y2V9bYlyTd2wdYwCIm2X5joWVxbpqrHUdUYkc89vEe8oVdjWfJ0wt/G1lLPZzE
HcqlYMbqjKaBcd854Lt8HTKTsn0uZFkkcGtB+9V8/15a6jQTfy3k+55UotsbDliP
qw5apPrNLynCKqEVr0TiRB10K1F6VQD8kZX1BGBw5k+L7E7ykuRIrKCW8bQem/r5
bvRnp9bmuIFW/5vpq24pOCqbEYoPQRogvfu83YuD1nKhJsrIXBASbej6nW192hXb
3V9vEGdHDgc1A6qxJDnVtj/fg+tBFvcbO/Zlsl+FBFCs/SzIq3ban5IqasNMw/MQ
LDx9iqqjI7Wdr7yVEXD/FKuoYGdgPKXq69SfKqsvpRKBD0BhrkHKZqglSpHkF1P5
7t+uuFf0vBrnSXlIwtrqytec+3jICtsthJabFx+x8yO3Vns7eb+gyHsD7wIkUsUn
eQU2DOOGSxzGz36h7icjbPzm88+c9KlbtMehWLOQbyxhgV2npLmZUd+spJ/eg6Ee
IWIHBkWFuRLY2740nPZh1+y4a3ttXUncXI6y7cFWx4Hehmy9RJEawjQGI+F1Jd2k
xtUQNH55OTmkLs4fbjezAm5UyDBvlVCzlC7y02heh1XWI3nZxXgCqvRX7Hgkxc1p
g7FL1h73h1KeRl1LmU6rf76GqeIOVlkjACdQJXPoO73dPsvQA3yhO8myqsbkyqJ5
Xtxh3USm8MBd2KtOvkdFp0RrUeqVPr44fR92SiOio1WB2bPlxsKvKupRdLN3OB70
x78wGA8Yr3wyFmkwHedMuZpwlDjXN9DlBSUY6gc5B8xshCyqfr/p1V6g7lLYI/7O
hsPUvgdm+FlpWOOgJvrLC/7DBKQ91sis/+5DfCJMzaTcaoXSsFZsdIdfZ20t1HBK
y+MSrAIF0J6m8QvRpFVFG2NZvEae4rgZmg/0ke2xrFbR09n/SQlkSNHNKIVCdtVt
ynM+ylqJhN9ksxqtUAv4KNcm8vcNT42ZlotV3b+HouKR9gvp5RNd+VouCH7VqQzB
4B2+FyzgHQeVep0RnvHBwqAE1SMTnILFtj5JdDx6vDKOE1xooXPeO+2K3c36GLPi
EXlypfX6DkpAC0tgBcuSResy8s/qLrEpR6myM5+lddy6Du3NcyhoBQeUD95rOBCk
lJ69ms18TWL77gA70HP1T9vLGaSgw9AwQ/7TQqS1zxlajQHn8JN6Kp+E7cIfINWU
jb6EqXBHJ4zyQX0mk21uuDIuxoFPpOg2CZoF3VvzHEd4pDicmjtBcAUYFViYAyzG
gdxFG4ZA984uNYoVfQ9hKST6MmrlAjzJa1B5w8rAzVtJTIR8+Tdts6iS8/tAm0O7
f2XEeJAgtkAKz7jfw7/byGJMCZ82GGMbQ/7ic8kPusxWuUvzsXfhZGUIM7qbpbcJ
s8DAcwEgKwfo0bpU2PDBywtk0K+uhjHweK9c0b2jm2pvJ23jJJR9x+plhGTib4KY
zC7ilTnH1yJxDtVVC7afc43Vbl6hRFTegVTXP+nHDlWryo/8+pj0P7lLOwHVB5Pl
reS0teaIHD5h3SZtozsl1KePXSrRIzBSQ2pA2+Ge64BRuY1wFsbzy+9PGBVYz3xA
7j3Ga0jeDcwwWT+kZUDx/Vd8OHnPrCGP9pv+FguM6LuTCb1X+GFFTG+VxLBCzUev
3bJgbO3EWw4nererRT+6kmHAiNmuV9ljZCKcwPrsiowbn4oSYo8tBKxhN6DdaLWj
N9XWsZsT0z4zzjG9PM4+vi3ivznKyQzAfl9zjivPJTMgo+JtGnM8GjgwcGjqr4UF
Dgv+6vgWlE0DrMjtqmoXgn3lY7UhzTLRRgId9PuxPpSOibgcCPZ0LZecwmE5YZJl
JaD6cVJ3Pp5HocpR/dh+Y4U8gTGcTIpMct22O/axcZuNULDmLZd0WlIEDnOimTOh
kOwDwnEHTSUR7Ydw9tfSI3otdyEREyUDgHXddyBBryBQGthS6mMb4Vr6uUDwDu3W
3mbDDxqLQlsf+1L2XmarzFHagceC0xUhwYw2IBUPKydubC4ZtCQtIDGnmhDgokEk
UTrsUWWJKdtWr8kpNNE7ZMK+1mW6xSU+NK2uivewwxTEAMNhGggm29GtTwjWtleU
MpPSdCYDM1iiZJeq6THoWOomqtY0LHl061wIQ8YjOYV4AdvK3woFylvdEBc58306
EwsN7L7RqZVaKZ0urD/2Jkxc8XDaN/BuR3jCbZjroq8XMX0aRSm5WyO1AgmwaGUK
QunuTuT8jimNzPtyUGSvuMI7kw1AO3A3wgFkOsUZXXSvq2H4X93UIzpKmKnTW9l0
RHi6PYKARU6LfU/+sscccTRWYBNL39UD+2Rw7ENhnMWcFgH83+XpJd0N7XLmRywn
K9EHb+eqc9JL2H0XGNlHlxzOiwboeWIOSwoNvzKISXTG19qXfTTG+ZtBkDV2oWPY
jZr4E9lo8ZpV6gg2CovU/eP/hVIk3cYxNXSF/QTo1lcQJ9TO2jn1gk0Xu9Ntg5qK
f2CRvRwSWpNg7NjXMVYYzsGX24ldboCPI+/M0hO2MNzhFJq3XqttvylglZmkle++
YBdW0GSWx9hO94GzcYEtCwlSArrNFYlWDTFLKtqctZ2PC8MMd/BwYt3suU13EE7o
wc2C10FP32SX1Zc/so4vRPzUHl8jEWJc44BjcJN1SB/M09blI0REVvFQ6RADppbr
OUl4gzsJz/svsarJIKJKALIkZ+DB4oKeUE6c5EpYnOb4xPhBM6U9nI5bL3d9nMmi
ujvloAfEfrao4I7TfggMF7BNactKafurKMQLeTpPiDmcx77SjhUFiIpdKkk28CKr
Uhpcl8wjdlRJhmdFAKCbHWsUvzRWv1gPkEydhn9TEUg8bCtU/Ro1S7p4jMrUwcHm
AmhmyiPjGm7F/3QkBzd0qA+fPuD426ZEpuvW/O0fEmO6A5TI1BN8DzSbe7Ny8BjZ
yXmZ4zrFPJ2t0czYrYaUn6TaqCv/LU+9iGovnYr6pOgEWi6XlDc2brATBFps8gmQ
CALxHOiuDTvQbH7Jubym5QdENWEOSPWMLOgV0QxhnBUnDFLYnfZeFrUYF2++P+Yx
EPiQTlda4JgyXDkH9a8NlZcLoqaETrsKRY+9Pzr07Q8sTZRNp8V7HGiN3hmgjGnq
fEQBM9TWAF+LjNLgmr1jn+IBXQtjO2K/BzHiHk3uS2KNAFxc4n242XAv9bLKS6Eg
q2x72Eo1U6Zb6AwzvPDtgxPiqbq+OHx1AyRvDujAKHxuQ4J/n8pG9Cjz1KphXu8K
pTwvVGrRoN6nLzdriYB/0Yl+NUJD0KC0LUmxFCtjA7G1Ns571VBbU0TW4b7y5fGc
+nsFmMFqSTNLwtxmRKICGeWoWOPKajGueCY9c9mHcUj5tvWA1p0k0BZpEDbBqnF8
qPAfttIJmKqkP0UgbfrojHUKHgaJKTFHaofUa2Ay/KyMCgtyj0rvNAAkh0g4FfbS
sHtM5PKFUXAh2VD9DcRGHjWcyJbD4xWZ4sljDuOnwFX178aWElH9tofjvqo79Z+/
bW8WTD5IuTWJgImxdTyQvc6KezCxrrLW8qh01KmDkOCr8gP3r/+JmeFzgOf9c/zR
BTWtzYs/rAhdEyFwLZa09/BJwmf94l3a7IhKZkdm27eJXfKRr0bvvjPNFeW0yUF+
EqqSKeNSyGo8ncg1bgP9Brslv4wVE/1ECcdqbCMkdnBLPk5bgyBB1kj+4/0D0Mrl
dzBr6y7ZN0R7FngpdS0W+Zo1ePaAWSPTKDAlh7IeK7FnaZldB4XxgdYKN+wnf+6N
/xXd/h9VKCjukImUKypLMK23MEsMUd214Z4NGP9Q2VXFW85T917DBaGQMH2HsB30
AgS+kgdWmVin6GxAN07CqtLxiaHBy99jjlXfB7YNv2AjIDpkfkNBavrrxbRhEC3O
E6Sy1KWYPbY0UPy2JxKV9AmnouFD1PLjo/9XrwTxd9CFCWQefRmjAyG1lN4KIan8
dUO0bPsMZ/k/tCmDU5IDp3e6xDjJn0Hn6giWKLhKz/BN7extkSHxdduO/ElfKtJr
pqLyEzJFH2kLUTSknoVd2DFj1BDQaY9BX6DOe8yoSSXMdkzvxoivY92E857FX5k4
JRpRn7cUSC5zxuBvWI1hwva3ih1Twc2TZQkIZUH7BGA6vShmN0sl+76PgnmtXCa3
yWfhYM8fZ7naCkrVJzJG/Y3noxZvFdH0b3jYSbrlmy9b0OPVqKIOPm7OUtmSFPgu
7SW6M2xnzGbe/Aiu770p8xw0r47VBRQUYaXYUqv7YixyXTvdrLaddLwqjGMlqtPK
hnI0g8KhZsrJP+bO00c/wde73et9kxy0lPBFhle0fNJeu6yMzTeQiPVLMoxI8xSK
Thtbneq1KHyvWNGcDAG8+TeScuVsWAXrIS/SVeLzXgqUE5HOoyt/PocgOqXS18BW
v0Mu8eZiePiJElejbARyZnxBc719VRqN7ktszglb7froOBDB3uhGCsleCpbGMXII
aXeFKF7HcLkRJJMNVp/dYkQvkWD1yPOYd79M/Q/pI5y5Jvcnp+DriUZmVjOnNNAV
pWRi7hwIyoalixkbcJYIFa62p5KjZcv8P/6fJiIZMQAJ63CfmJs83gr1kWu14VvS
WuWlBtvS2dRcBM5G8FiEbKDle3NRb9WlKhZVCvBeQCXFakmHGVp61RvAaTZstcbu
E+c+MnO7wCOf7LZ0VXLbySJOftFAOz5gdRV+w/6Poau6QhjA9U3p2WhX7/iHl0W4
pxpoK3hjFogId6CCmg2Vp/GNlhJbwap99Ordd72NNWRrHKG8gmk4gjy2WsBE2hei
cqJEeTQ/da2zS36N8xyYJNAYt9DT9eLCi4x7U0DgM+USM5w/mO9jzLArgMlFkcpd
PNM0uov11yCjVHlQDD0lI5AWkhlBqiZoUbDTZir+ierw9A056XGKW66MoyDq5p3y
yDo7WaCpG94cVlDU4jJG/WSFunv3gMVSESWK1oGEzOLdC+Bwnb59FNXh04symzJJ
9rXKSXZiCEPZYPIqqk1jR3E7ZGnc3AZMGfvjnjHMKt5B0TjjTBPBy1Z4/mPo4uGS
tUmj9hSq49OgqVK0YsFw8IzoMlqKlfM7bLB1YWAw1anR2ClzEuiHT7YQCAzXJZkZ
quy3EZzxFAXMu9h5kpy6pTk/Y9KHtlFbWralRxuakBcKTMm/IMQmJiggYIs6ZDRL
L8YGxRlqyjTinmhYoQUvuNLiVlej9yKsZH9ZgfdUAgTbQQRC8xkuWb5FaRV6dcc3
h+ya/lMC4ni2RXW+1fDsRkgEaDKiwZM2mzuyBOGiVsBtq9DNtpUsbLxjAKU6SLCg
289swzOM3ZcsmilH8+zsKPZdl8ixxVx++SYWYYvqyJFnmb1QXM8Z/zks6g1cMAWy
IgfO9WQYjkgbc/c6+mR+LTWM66EWkEOsqKlX0o+TUppTO01nMLCcE+qQJU806F3+
N/E0oGsZh4/Pka0x3J81UNPgv1E0c3mbctSPqJAtNDESO2yUKiIgzuSJAdc5q37B
EYNRDJ1qeNq6s76NhQY7UG/d82F4hQAe6HOvyXK57S4gSjTj4n+xa/+nOVWV3ZHV
rgBpi3+/spkk+AkS9He4fvaCfuzK0RJafOYRegk7g2BXT0RGq9cuIL+vCWm8o/Be
iij7J2HLfG2A5WaqZ1wocUugmEqjsEGik5XtDiZY+FzpFqj3B2n4BeAmyzsq2Xv/
Vhkswd+/Bn3ASy+ZvIPQjkfqdgUdDUSXg/oqtIZtZi9zw03tLSvearme+KAqKFEB
3MVIUJbCwDmJEQXW4HenbsRZbWvpYCi7Jv4y5bmD9MC82dypzoMxQrXuH46QC1Yk
A3t63uXSIH/yVNTuPyY0Vx6INU5Iwc92OJs5QiPOSTY6A95JA15hhB2rOYTI4/PT
EdPj9Y8on/QA9u0zfjNW4hu6F8khkbp1GlIErIPpZ4WjGKR+6obny+O7ZAGSivwU
lASSz86YfhFhtxU+tCsOHvLgFc9QXHI438mhnZctEjKT3sS0LEjW1ZxeE3wxsVS/
hfFV5tqmrqjpZO0cj2UnGJeCdXONjUNEpB3EYgh1QF7KopIBNXqCUKhq2oegWN4r
x3BF6HjaR2etR9WkOCUhkG25Yg5Lq2ypN1Pw0+ImX9I1DoGbDBNAP9/bym8x3nd1
Hfpstc3JplSCHG3YQCnv9Z770lPJznFCIAE0hFDenzZlTJNSQjvuKcwb4BonkC3d
bNzvlo8I+5rnT4bx9wywQ3eC9u9Dy6NDnyPPbJRnFVG6KqVoqD1kOTgCHLIZgiDD
zkRqSMFJsSEaqzeSCLir2cTgn9z5dRxsGrlDJCgztxNHtU5jStKDLK/zgMXveRSO
DRMMJj84OkYdRW9hqfR6OJcEl83rrgW0llNDjJDTFQh9BfIOOb6V4Pt8rSPr4QH/
uaaoYQ3YRkzV4TotpGTqssz9DWIH3RYQ8qHpY9lUs/TMsqU06yta5iLX16PwtD2Y
dHBMJF2hZ5itVBsCgWvtERNqtsiN5GXKFj1siJlw1q6GtunXaXtHuJFYAWLuU/XV
s1WK0UG2xFe8Z3rujth18pnfieWEOQ44GQhAFs8jj9WuvM2/m1newpUdCo8Bj/LJ
sacFIC/t1UV8ltqANqPyYWj7zb4uQ/xuQA2n191Lill9TwjGxwlFxajsa4jkG881
rFeCut8S664V8vSZFh3vdC+0XDjL5PPUk0K0k22xD+Bwd9MwqFYK7fwNN44zdghZ
6KY9SutIsg3w2y4+AmXhbWKQBfMSbG4NeZD9tMoxIJBnHborqjJm+WDbUf7aeRID
/n+PBSYeiTK840jecDcm4eeN8copipcWJ4H7LbKwhkZopCExmk8E89BHhIYx9ajP
ckeZRnmUzWWM1B5l7TtnsVgsMS8diV55/+U0w3BgKIfDOlVKXgF7O06ZT6n65RQV
Frg4deCRNbrGOr+iYjXVJn8sJdvFpb3N347UxOLyDK0NqP0DhyBeLqdSN4B1Drsc
wiiIKS5bTZk0E9j7OM6FpVO0X4CcFkEldsEZzAZDelXHvCbydiM3ofbdooNmWNUl
0gOWX83j8A4QxNV4qnR/Uhi5X8hMnU1YJGyXQ8CcrAcOK/xYUQaKib/w/z5saWsg
sNVQk+cKlWDvzKfnjkiud/kxIpveepRTsR5yskxb6jm+bhko7UuHwGHJKs3OISj8
xPUng2sEysf6EbVFlVzXzBI/B8BWprXfpMT8qe/YEdweaoVLRgZQT4jIbvC4AqM7
Gl/rha8J8DCFKZNdJGXhyihB4UqqlJhjQGOyUUwMYQQ9i7j1MNAjB2HVlKpv6m1F
8VDk66VU612a2maw8xKsSH2ZrlJzAs5RsWlq1BYYfEg6xa5yfqdW5yD0RtpNJMen
+QrdAmi3mkj0XqBJEUrtv+Y3CPmv9wsuaF/cJ8ozA9jQ3QGOehMLb74Sw3G/Xyra
A/SE3j/wB/XivB1/EG2Y0puja4pGAY/rGl5XpA9OqRDHQu6rdRxLPq1XZWiyEGTD
HtViRmtLQeGGS7iSgpUAbi6IwNa7jKHN1eN8/1sisZfKL4G0OgidUjQNRo4moTC+
IhKnogh3WFuMYLLu4WovkeZ7RYqUWcO0L0DkVM5Jgu72jRdoks65bbO3E1GU1vWm
2H+vwy/I2xRN4g4XhzbjgXRR+D8xM8Tz0wXtUPqIktzXxM+7icpMKV850YTggekx
NBRDPozq3eGL2qX2hWbO4AftRQUTKYCyUrPs054nFqdjxMeLBSi4NfyLYO6d+Iyc
AsA3ZLiTTo2nz7J17Hgiv0+qd2yHFVOqsbx43zZiM5eqcY1rD/JPjJ8iK812coga
yDM36QDFULiv6j9kHsj1bdF0JDhLL1lKtD8nYGAFjZ61Kcpqb6SFz8Ccxdyv/hjL
Y+KLXBnWEiZzwqJFHUHIl2eimpMTzuhJCwTB8dkmL2h72Wjm3vjypcZ0P78NyzFe
4xam37Iu96XH5EfKCqVnV/B1CQdWhsCkDFiAFBcl5/Q7lUDx1zJE5jYvkOqtF10z
Fm4kWegEeJYvOL1aUscb6yQWNLgjnngcyI4UjYOVtLMtnCFFBjIcBrbmEKKFydnZ
zum+Oq3GqB+45rJ4ocAgUYxfzd0Ekru5fRLtcLvTR4bja6AaMTpj4yBwYi8MuSQM
HE+TdvWrfCf3RgeykduQ6kc0mZ+umjVJq5xBgjBC0t+MVSpcR0SVLn+8P+MZf225
q/SiZDEvgYQYlyYumfTc9ZcpFk8XI7iQLws9FOTeDPoRI6gegGzy1iXUjaQMMloY
sCFSuN1s/Xxf4d43DsyWvBta106ajWrNJhVhVZLGStSU5WkOIShHxlcZe/pqp/D9
tfbCqLeUQMto34ZuaShiLt9BJigwOMgpQFxUvNQCpj9WWBBpF/4LjqpMHQEuoUGJ
zPe0NqD14NqjXLwMT7BVaobiHg5ck2TJo/4SJsrxc5Q5NAbDDZkOO6xYucsx2FLQ
jvGSIefBdZtW1mPnmfT2BXpUEMTj4X9MV+wc7uS5uhGVjO3Rl2MyiuYT8zasKita
De/IHA4tRj1LVf/B9Qv4vNYbFJHdXa5reUwjd7F0ZMPMszHT0OimLBo6h++v/63E
9TRp+ERslqQkMXxMPl/Bdw+MMJzJQLicNgnlGO4CnzU1KpCsVK6n474lP8r86ZoG
w35A+cY/LdCXiPf2PobkcN6EznJ+L8e2f++qY6jQtRP2qYBRVpqskczo0RII1Mva
vDXCLAVjh2xCSJkrhWLM+RYysdH7Lc9ItdVQvGhf47uXTLOs6m/mFIqQDtQmjHU1
kDaNEIC7Y7e1wo+GqG8T5n3H9kJnj61gm33aFcSXbj/Hgvq1VhUGDAQTQ4YbAT0N
P6DKWiOj90mXqMUP+PS15hxlMZUtlbLVGR4Y6cSgQZG1tJz+gMhIJ7Zhd6so3RL6
Zvjh/w1sGvclwO1QyUypsuDHO/uIxO9dfKd21uIlgKczYO8vaPDUSTR4aH3nRZ2w
55J5yEA9BvbVfqKWwpCZIyjO1TxwD5+dU+Va9p351OmuZMFJqxmOl1K218o9FKII
`pragma protect end_protected
