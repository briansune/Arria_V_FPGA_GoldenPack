��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t|� )���� cE�-�?��Dpy�yF�ӽw黨@� ۔A:a�t�C����>�m����y�����C ��S��������C�XF��֦��������T'��^s��w���GUV��_g����a�b���\{1ȉ�{z<���v����a�������������z��P ~;�ʮD�0xZ�7�������r$����A�"�ե������Ո^f�' YDJ>��\X���	�#8Hoxfm�����9����>W���*q����w�AY��}.I��v�ڤO���%w;m�h�>��*y(�pյ�m��DP�h��: -*�3��I>�ۘ���2;��BƖ�f�"|�5[]�9�
���^��zФt��c�7�q��Gd��<}x��vr�[�b�7����j�ˎ<L���J�^��*��O�Du���s���8�ɫsn��$kܾ�ʅ����%ܫT��)�j�6�I;���A�[�')�GT��:;bQ��A]@�hP+���E\IDw��m�nB�����B�o����Ǯ�bsn��E�q��.��|�SA��x�N��m�s# h��Y��y}0���h�P~|���E�O����;����>�]�c�Nk����,+����ϫ�L���,;e�}v��p�?c�X������ň��;2�_3��s��z�]�ANn)P�,�g@��^�@���__j�t_`^/�t�b�.�Z|�/��¦,V1)��an~B���X^gW�EZ�jg��$%��?ʖ�p�A+�q�,Mxis�l����w���q���#B�5��4%A���@�45��i]]��m?	�f1�ʮ��`���i����4�+,&���c����-k荓��w�K6��]�+���iWФv��*��Ӏ�������l_8��Ғ(���k�)��+���2��f,b;+71S�x}�}��T*�}�V�$'}�һ߳XC�6K?v�92�!T���XIN�"�������rwԁ�LRb�H�O��j�L{{T��c}���$Wzd_� ��Y)	�Cy��G��~�w��X������??׬]K�|���x�F�YH;�Y��~xA�\����]+�BR�CR�!�/�bFI��婖wv"a�X��̉�� k��1�>_T��%nu�R�e�u���vw��]$� I�ܔ�x�7�8s6O���܋� ä�/��@E��!N�2��[j ��p�b��hU͞���@۠�%E���&{[^�Y�G���p�f�',:d��5�w����v��H� ����"����qg�<P��e��)���k[�u�Tz����diӚ+〡yC�M3s�!d�h�>̼4Yjͦ��=$a�.C��'p���T��̭�vD����JXc�����렢
ۓ׎�/��^L�\��Z&f��,?�@:W���Y	t����,-�3d{7"�3���*BY����&�qL;y���I��+4����]��lu� $G���D[1|�c<ɉ��r�Dz]9GϞKy�zg:��[СH=�Gb�k<h*�]���$�cÝ��;R�<)(��sش�⩮RW	؄��:^�U�6#�h�=vX~�%��-������/F	��~M��"��OL.�/#��B��@;�N��xp��-�U9�9�eMV��v�?瘟2:I�R��Ap/5^n+���ݎ���y�w�gJC�+�k�
|{0y�q�D?�Ͽ�$־o3fK5�P����]���ͦ�Wg�"P��-���PƑ��
aV�[�3#w�IS��H���R-I��٠����LtFE6^�F���%&����b��P�ԭ�b/�=ޤ��K���\���(?��,��^��D("����X�Og! 1v�JS�؀�t��T��b�CLlA�z7Xc�ܵ(����tj�8���6�ЉiA�Lc�,���&��X�,#Ŧ�SZEam_]�������Ƙ������.D�fȲ-����1Ύ1�_=���9�J=^J|�w�i�
NR��l:�8�KwԽ�	�C��.���9P��qD��ݦn'�v����O�,�;z�D��\�ݚ��p���6�J�\���i�2U��s�}�|����<�~�4�#|^I��� t��9�ؔ}�\d���dw��������-w6�9����@/N���im'�` G{��bu7CЖ1.ٯr�=/F3���U`�)�VU�Q	�`�LpC�l��KN�qQ8�r�M�C ���Y��2��R�]����M���D@��WN����[a:���M��@�w�I"(̒��`���(c.�i��]~&LBu-I�d���{>eg��o���90��@�Z����-e♢��q�G��U�G��B����Nu{��"�
��d*Q�j�EA�H箦���9%��zk�>sf�&}>t��?w4��W@��&�{I�Ֆ�&e��2H�����j���O&q�M*8G�]�Wa�U�<����`y|�Y%�fW|k�أ���M#�ZóLI�w��Ѕ�ΡH�,y�1#.�I�#i(X;�=�D�L��u�y��+��½Q�Θ���՗������~�|p�j�B���ۍ��4�~u�F�C������q�h�F�wH��4�¹�)�#Չh�?˳9'�R�H"�Z�Dص�cL����)�4���O@��3����x��w���-f���5[H�4�H�Y+<������I"�n?�!!����Y�5y�j�� ����=8Y�zr�����-��kP���ϸg��n�)ӓ��q���f��?M�8�j'��a�/�CGN]�[l�.�L��c�F�j��TCmb(���z��[��7�D��9~y���H�4w�|��ZXV�4�̏�^�4/˨�I?���;����{���)c%=R�u2�i���$L-�#)$$p�q�f���vl88�&)��X��#�����?�,���Q�3��~ؘ��೅rC�-�uf��zU�� �tuH<"��ck	G��I&D}����B�dZ6\&JG&c��	h_�p7��0���ļ�"[oEJ�jw[W�i�]�	鋦kS��$V@���GM�v��3Xq�8�9��M�VSS\��YlE8)v�J���p��LF�m���:vAء1F�_C�;d��R8k$������v%4I�����ld���߹v����	R���ӟ^b�-��_&-g�P�Y�J�V\�p���0��솕X��a����)$�f�p__�5�U�����6w7l�Њ��#� ]-����~i��8�E�$s,6ɦ �t�T��5��� �+��\��|�z}����J���-07r����f��gk=��Q6�������e�R�J.)C�u�h��l�F��6�8�i� ꫄��V��d��v���A�fuJ����D��z���#�R���5e�QMW
 ~�G�:�W�㓗w_C��K�WwG����	ڌMMWH�