// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:54 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bxLd5pDFZNtE7bwau4N/8fz7vc49XeSeShEFjh3JxePglPaBHK83n88YdqwX2Zhf
OZ/aG85rp32oe6Oy+zo9am2N9ja+KCMSOz4kbZflMQcgA4Rls9bikSXeJMiUT3ot
pjjcjde80bj9k6kqbM12V8hS4GFIU4trCVrg964/OnI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2272)
C595XsYNNrZXwQHFljR/TwxfQGMgtkSOo0Uogg94cr9UfPCLIc3DZGv8Q8EGxgfg
VSwDz1tZNLdh7saNDzMpVo1L3WMGqZD6HNFD//JSY10ZNfXDn/bJJE1GX6uJy93H
t3deDH8gZPpKKKQ0Zg/ZbIDfpQ+OAOAndSt+3v8U8G7VCQITXkVdlW9i8Alf8YXT
eD4JItdDTa/7BvtQNEl3gEBNf43Z76/ZdXpkIQMA3+Vjnia5HJvSa6iuzdbkwn7g
wwujfDcC+LfJgzypw0p018RDVlau6+vqIcp96UXJby7ZMP0uYfBQ7++9lbTj6BDG
atP8ITl2LmMNuSI0iSfL/EuyCevozdxfJddia+QKrJ3LgqGYYv6yaq9VctsfZLfX
FDEGzL1y6sg26R8t/GHlqWRLZPPYqUDnyY50Atb2J261tQCDPNXbrLz1BOjO1Ytk
NXp6XlHNyr4XBhXdVHxOUhxcjuVeRd404YvtumN/7LKHfdmQ7KedZfPm6h1yf2g8
42BLUz/O32/LdXRtPS7tzGSJX9iKsZfjrgxF7qvxd4GcPAaKmsKBoioOrq07xjKS
zSOoDiIU3uR3BP00SjyQgr+htdH2IQ35TN22+NJCtEciVHqOswvvabXm00uIK+9Q
w/2LgdDRyA2QuKu9OoVcbdJB+LTIlN2HR7AXurPsE4bm5baJ9E/Lmf1Sr8XB54r3
hZqKXw8fnXB1Jmhs4HSphZLBTnqGG6H9JMP3zmgdet7/YNiADcW6YJ2zdH3+vkIa
v+ndz/OOk4pvbGZyJqVZL/yqYLqr7wHR1mhwjjwBGqvqndoAdRFh9FdfSKZB6Smv
ynAzFyhD5yUK+C1p9bHq/MV8DNjS8D/HUJmqDZOylfxQeMWNTmDjqVNjkos1BiWX
ZGDR1I/V2PPxnYFOpFHqXgy5K0cRH1UZmG6yM01tveBAZvH9jCe0BOZmKzDpGwyC
w6SI48dAqGiXyZaf5E9reJS6O+VdKRQ/Gm3h5ocprXUDrezHH0gALJAmySR98h3J
3fMc/7M5Hqzrr1FIOVqeTLSOoTKbV48e7cm5XmdmdC9vu5Amv9mETl0qxoNFOqL9
4Vo0yg7Vdjav9AbynkQ5ChYogX56f589hUBtxNDG6CaDeBTyLdzISR/3lJUm9xBw
+ts8owHJyKu9GMA9wWUSShencK4QX+8VwV3sS6mn6MftvPSUsoSZturn2dA80vGc
dAVIADHZZGUOy4iJObheo2hLC7n7BuII5cHRqVhCuEBz0zPgawrfrOkwn4QE1iP9
hs+6brwVLPeLlos2ZWV0HQlCK4Zd6QKRVbHC76veHJgN5ZPUk4zFu/mXjR0uQ5yH
1bEG2wyBXaTf6BnaIZAUfwGubWuVtRaPZ/AkkkhBm2AxYsOMFKkVkNfjMNCQeW0L
nRuGxyofJXkE8jWHpvQ1/KHM5Qrv23P4DMipNy3LRcPH8Z/wX8WcLoBoMCZUx4nB
ip+r8VSrgwCo/Kn1z0fu41bUODo5I0plSnuUWNHC2oqCOW8tWSRMd61tCuz3d5PC
gBHsuACkD4uXJDPm9dTvpOWsCf03/FVZEa4wTP3YMZwkf5CM/IoK246ytWNCkH78
8zxARKliWW/NKlXSszKE6KV9a4ZScXAKatbln5NUHa7iFM78LhDBvD1J9xlcE7Nb
FNvJEUdsdRtRF6bMy7Yr3ugG1mY9x+LlGvwwUBvTu5MPRQ1A+W+OsPzoDCkhZ+fM
5y728Snz98lgh+DyAE+9ReqTQPh0j6FX4hQ99pnDARqc7nCy0PgEe663gV92e7De
M1Gpv93jB6JatIPBcvrweoh9E595as3kWUC8AJDdWPDO3vUd11bf83jBpsoqt/pr
TgL4tdLARBLUOBqDnBih164pg0XspcM+02OxF4TGm72ldwtu1BGQEPUKwxMrimII
tuRyuGJ/zNFNM21zHd9ygZ4XciEikw4KM++4dsK63Axjgym+z1O4aQKlhiT6yja0
PDUQHVBkehd5LjSEmtHQHIoOT7BI+4mshLwqHt2pIHKuTaRiX+WYboSXGT3HqIij
1CMiTQnDwTFNrTNCQdy89bdSXDobr1lukmwddGqCOPPSrrKmpyqvvIdFxkqDRT9u
XY7swOSrviMgc7uhYTvHFeigKt0oGzlJ5Rw8pkuSJwPqGFma+tadaXQwbnZJRDaq
ZmnrdiLjU3SNVqw6n95PQ+rRjGPaJKYnh2dIcFUMUfp2W7gEIp6kfewfDGhTL6bm
4Cxfxk3wpoCUu19OzprLIalnxTCkGhF0g+ts32FtfHn1NVLdhlgtlp4aNkb5a05y
8WTl5jEgLkJVu/iGhb1CVzy9HDXvBSQCMfUqS8IIA7WMNxvnoaTFDUvd4gjS1NaZ
HlY0ddufE1T1Ds5gegD+/aA83gMGUGCr+xZ1uIwbDFuZEwKir6JWK5Law2Kvl3m2
ElxtrgYr+1h/SpUePgaTU5+FwBFKxrkgpQzsPZUR7Uk+sR6I+g+r7xTRbWQrSz8h
bclhZg7BwOLlIjw6h10++Qd4F0M4TtSS5M/Iw7KSUYnz1Wv9LUATeG8Yhg/CaBqL
4W/bBYIEQqzIojLeqeOA0NWYlNZvzzeCgZ6fcergujdNw/AQ2uSPygfDA9+Y3m10
rtPAXxcwbDW/cbokaj0bv+zBBYlk17kC9vL7sc9uRpCUL5oB28KaEHNvgbVK831X
jWb/4KovxcnRub+f5LdgpIXjflAIrGqXTyCONm+aHjWHF1mdqJolIj3NMI4llo2f
YB1xqbSFT1lpgM4nxvyNYkYdF8/XyZYUEGz7fPGfhNeqES5QzUdKjaba5eFgcoHH
MRyASmxyaY8NPV8eoOrxDJCMzAYwFWfGp7+KvGUuX+8Q3MgTBorJW/pZqJqohZjv
qk24XhnsAg/lNym2yHkn8HA/DOVSxoGWsVeyg+vu0BTvjUqdP0mi+1POD4kpKxO/
gVaQUFaRc2JG7Mv4JLNRrbVk6X8qqUzniTTVhQnc/scog/baWCJTkBrCV5l66Zw8
d4qz59ByL4Hd7ppHVMSCCg==
`pragma protect end_protected
