// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EiA4a9Eqi2flcGx9H1ic3zzH/Hk8PD/tMs9aTe1vaQjGALM475l++g7BRmIDHblO
leNNAK3e5+GtUf2qK553WxEvyh3AKDNhx5OYIfBSxH0vwnqlv9VPukZs1R+ugurx
u16Izf//AIV8cZxQLLgQv5Iq3s4/0bkIoWHjF0IkoUs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11312)
AcLeWv3klJ9A4BdW1Lb7277WzFrZJ92xqtFhaKrOnw00Z0AS/Q69FrXrkd9nm6s+
Zo53cBlvsRPzOPO4bA8SHk6ubZLcNWrVJ4Z20Fps06I6BROkpWuNAOG5wLil/MY9
a03GZna1c7LFERdqTNdplG+geJy/QHKogIit3nAs1wrDCp/ojvSVzJdN/zWEas0d
5TRaZOv4PYGxjfAJvuYkRwGObfGvSRMqqdeVNzWbJYmwCW/8xCmGzBceMUaYphK1
GGxjj8EpE1G0aP2gW1GsY7lGSf3KF510QnFK9CX9ngpXxehnN3S3XKeWJjabvv8O
/YrY5pdQIbUpw29V8g53rq3kf64fyiB+TKRs+Q8OIA7PmCoOmBBfjRFw+S5zLn4+
MDMi4i7t8aOFg8LEM81m4ocQpapiQTlXQXvl4cij0dioVwYbvo4QyWjKpBskNSv4
wtW4wB0cA3bmURzFcIquUZneEC0T8hPRKJ4bBiM4NO4A94UWfjctRMhX0bOKr7nF
bS3rT3JKvWXVspd4JBOKKCv9Wrl0lpjd2hlbjZeLqqO9xuE3nbT0RubHCJfRKg05
OaTFlJ8Pnmbv3sYoCUGqBp/jrS0WI1/nJ87biPwCWNmFGgWUUkKbZ+p7wy5QT8WE
/FpnivpoP6X6hetnSDqJ4XAjV/rOxTrg0KudbyxV3mMjb6pQBYMjSK91yXBgmDLM
uAT0VEeqeiQIOP5xUNhMy/oezSL8f3+67FMGCBO3eaaftI4ABMVQKq8EHAtKRkWS
0m/4eVMlUJR+Ih2RCiSWSNOAgHmpjuKW2705HZoDGCU403wrkKViXM3vqHRHXObW
fCfBIrQg2J/z6A6IHZqJVcfNxtvBDpVBFrEIgpiwvgbpO/4AOcLNvi1GZ/WUBPki
ObhuX2oXOtVjlVDV9p6U+9s4Xg8CAKr3k63FvQiqPnuNrPbmz1vsUp5PDpi1VBQv
MZUDTb07/WLsDRA2uNIjwQ/bKrG4y9Cp9UhLqorkKVfgZHoHTmo+bQESzNn+d15F
a868CzlOyk08BfND6Q2MGJ5mf9tnmQ2q/TVb4CL5IutKnEn2Qwnf0/3Ww7uftUal
XFw+bcJv9mw+luBjpJ68BrYqtzxFezdCyGyPbSUPIvDojSdYJGp5X+mqmKP+8OKI
XrJXdaXPSfFH+46qdGYuuMSlw2VO63zkBmBpiLgCAUlqH4hcvqk9rK1eKfFD02el
PzIMc/n9SyC4MAMgrK+vF7mqV7AycTZA62c7c9ZqPcXen0KMEZJcCKC3y7d86kGc
8fS7zGxaiXkjbN+MGV4qHer7iYb46o+sc/bQh5Upx3jz3ySkBVG4DZDtX2fIq/LO
lvF0k9jrcSIENiUBh0s5C+2KNOaHe0rX01r0Lf72WqpdZI7EklmG0cDpnx4PpBRw
U1aesAL10Rwz99alr1m24HODgwwr7AccfjT4OF+72knaA52jTQ7ACj48UB5qw6jL
qw3ZUat372/jwXN0tnqpnKLaFlE5IM8r4DMs19B+xdCADuL0CDavvLiO+BB568cP
GGQg8R5gKSZTifGyVdi0EfUJ5Z7UNjgJ+R2oaRp966OKGydDu6NPc2b/Z4JhA7vt
1ZG7YD5sQBetOnmEzDR47dfA2zsfyHB6UeR1RmkqmNTNaVs+lHVWq5OzqKZtKZ8u
5H33UW3RphL9m76OaF30bHfYQ6KXIqOrAYdpVUf0FwzysiD0m9xEhVvcD71EZscu
f+FtFqlTtv/xNMZu95v8IY9vyQLBR+lSq/EGNiUPiewzIBbikon0IkrWEdrxB62R
hdTE3vVCRFKhjBun75aBpflGpkFfRRYp00c8wb0pILSwxkmZWRFXbevFl6DymDb3
YLZ+8xNCJg2uFxgVBQW3h6enaHKVb7OfGuXagaXlI0rNBlrJYjDbJjF4uCbBNpAB
65A/yEgLokOsnNumm16tsgt59hCKy2UXGg/XnpmfsesysbrFB6TOGfBNzTzhI9Fy
Wn9/HD2iLv3xWG+Qkdb1cdFQ0MnJseuR7gTdzMvCGmBkD8qooaWYNZmmq5H/RMr0
D82C4grym3AxkjB93LwxTXvPDSYd1GvHvofNZBAzpHZNY9H5KIzYJ8GSKz/xfJSK
EwIsTv/PDE75+VgwzbswuPE83v0QVsTtpHbsRShxUGHYl0t4xyIBS44l3iMP8kTZ
cTrShoSt4rbbbVpBc3nydL+Axs93bWH6fdrk3BDGeitEjv+JGA1QpkLQ3ZU7ZxS+
jJVp4BXl3ynXohFTE8t4kdqGxGZFWfS53iWyow/VKY3NaFPau5/2cZJ8uVNhkHKt
wtzM0RJBKnV2MbTCH99r7bfTaucFkaGWPRthP8txQmV8Ax2stpKSmKlZ0RsUPFal
In/CIYCSL7lVB19wNMYRUAUM2bEo5IsEX1tQ71DYFEmJg6uSH4wPZTxhkQwTt/R1
AtuuuQaJbwxjl46CBEEg7RRwBgeggfeKqR/6WbR4D4oHgFYjHtZ7Y0jxwv5ndw2C
qXYzUlIoK0Z1vkgxEOzkntsPsZOGMZN+PLEoU8IBuXTr6aNmJM78bK0TXiCMWZ3Q
vAEXH3gp5sXabI15huHOzoY1q8xN8BmtixBjtcz5GSwJacL8UcXAVKEgUxQ3KWKw
bh2hIzUBkWpAH3SFJooRFVV34zmr1555cRpj2swG7gmu86vIS/b/3fQ7GYqhaYMv
Q2DPoMMtBZhUjthEXfgQDSL/IwzzeTzDHa7RsGkNMwJQ4/uhLSWt2X2R0BJrbjwm
ESN6Pa/s6kY1nxD4I1AnRRX4siLfn7QItwa/O9MY7FtuPd2oFdRDY8ms+ZstwzLq
tpeHvP3gHwITW4s18tpynmC0e15W+o/MhZJ/8J4pAJYPyy6T4wHjmtq44qN8cOa8
VTCAIpj9qhTE74tXbTMS0e8uHaj0l61LLXSnyTeRSBblggBrY7zzO4YASTsJUVwp
mPa/RC4fQiNDIlAhe0Mnzaj/8VCO8YmbY0MquQ/8W1y18V5bWDwgFDhRWj9LWiMH
hgM4NXakBccUMTLb2ahVT7cvth87qh4ZS0Q7HwAOgklBMjhAvcNQoQlJA0FM6rbu
udnHFe9I7WcixcDEzexanYi5/JP3bhuuLJUlz3LSlrbdDBH1lsgsBj3MsYt0niJK
Sr74hdatexh7/Z5Xv3vTvPO19yq2rOf7+i31gwtGPrski+xiDM4vBJsdTRMI6sAI
B09hY6JDx/WSxUjxCozBLb3U5bFC2BMFdjv56hSDe6a9tSPYWaDGjfgdysLZd4sG
xB32c2aKdEtw+L8qkfBJErQI6QzmloAu4OkJeiPmAj+bEQXg6tD/I2a/HLxqeMrU
cThvWjAc3THVYXWjmX35nQwy0yjwS/xZYNAAe+H72kpkoq1u2j8x6w/ELVzMKyRi
Jdb/Op5ePM/WVzeeMoEiy9XWJI5lj7xtqMwUigQyxVVnlkbkVvZSSV9QcJdSz/Kd
vgjI/to6qrhf4OhEBIF4qCwq584Fb8YJXjo7O2cDY0AQh4MC9G31A4u/Nl4LKP7Q
bDGr5X6/Sav+jQ0mKeSYSRuWaFBCw3KtFGmxNv6UBj0CS0LjNmsi9Xx9vTJsdbGC
6eLhlUi0a6dAEPNsTbge9dNzYfYHDDrtxjeGndnUumnBYEc6w6KY4miwjfq1qta0
fqNBaaxQt7RqsfTFIffxToH+Lg+ZvCfwu3PyFgB1BgmtE+kGUc1MjO1Rt/2gy01z
uBk29VIZoU5PvaokqjCUWI8Huh7oe02XHRnN/GkEpZGiO29oI9cLlkmqSgz2UjUB
j5/oBr3C/zqxwyi8hjmHwLhNAntxJJJsyJmmm1Nk9aa1Ef1O/b+lXIl0Itye2Lq2
hOchBHTKvNqYpq24LRNqk7VuU9Cwx4qL0/y/osU5hYE1gizTWPyLZo1a6mZhamca
GCZ4wgXFNJLn/sk9mtofsTp71wecau7iDHSBgn4DiDLB9QbZqJ4DwufjJaRXnghv
OvIiEBVx56XC7dJ7DhYHSXZwDaPIU77rya982N7D/0TaajihRdfBaBsjgBmmrEOe
6VDHHUEqEqU/JAjOHq1wyLGourEoZMmwQONmShYn9+leCQdTShtgXMLNYOOHrAad
rXWNH3ZvHE3Wk8Wb7NyQHxvoTo2LScA033ODATMXOXidfaYMysMDPjd8JLGb8gZV
IQ7Oje9ChEgVbxTXUoSd2slCDarOMSJUsIynZrdpe+Rc+SagKVu78qpDb1f7YXED
9f3Dge79M8kk5IydHScVkgbvfeShzYzMrtGhQ4QNiS+Y990TKKjTVYS1WdUK/4dg
JC50MHXA5uN7yhgrukcSVf2XxmGM7P3x8FuFcYrbNVW9nIVQpNbXaKoFtIB3cTm5
+g53zTZ/lL4+f6WvEwSJRLl2tk0H2b69XKxy7FMosyD46K6b7ynzw2rK9rHW9eWL
8PqJTjT0LxE0UwOYCA57N+g+B+C3kmmF7jJTFS0KnwJAnC5p9trpDTJeOQgVBQhC
CeFR0i9yMiI4DbbTgg8QNLNFFwFtdDlRAlDbRydCRtbPjJd3oRsMsIAFstn7SuxW
gbY7g0DuHyeYAW+f4DtlyLhcqZ8/f2jERrzcsZxwu1fgrYLUN3R/vNWoiOypEAoF
Jm/KzXA3YxqOuDSFcuEj2ZaPXYe4EjI+pLpjUQksWGCYfojHSL8NLwLrpm9XZyOL
U9iRML+ufyPynqzU7gf53TZQnu8KhzuwJXKUbtPa3qrFKDf4RE7QczMCphdVxpgY
suLWJRkbeErQUsNX+mYejMUPVbUT78gYFnL3mWGUI7enQrifStTGmveaFIr6UsE9
5Ht2tapux+UelHwgOzNCW6Q7DgsGmF3GFjuTCWzGSAF4ZeXJkV+jtPsgYEsf1kxT
4NCq+j0R6Ijsd5lS2+PnsZ4hfyecGReun0GvajMEhdYnUHA1C3ADavGW5B+5LiA7
74eZSxWuvSQpBj4GWz8eEfEBd4jLB3Pw/kZ+fzsVq6v9JhKIzazLllTrt6bIdXIs
Z8LIhJFjGTHv+0gUmlFIO1xiFfjn5YTDv0LBEUsiljSu1rrOuIUB7VtS1Y/u76cC
IeZkg6ZLu12nP8HPm+rbv350YO1uAkRXdUGSHgrJcKnrP3Cn7qh9aUpPk9JcK377
4UqyVV+mQczKSdRs1jkOEOQMFXeiuUg2Xt3sIYvRv/CFttyc8B7ZTgvFlX1zyCo3
1K813H/4xTOY4c5SyvRYpPYu4JuPsDxPGzVErOajEocta3l2BHaU765rMWeWSYh8
V6ESmyOLc12sPWBRzVTPMw8mUNLHWGpkIrVpvLqXyU9jRSK5hEWDch6Kk82Q1856
CDYqnEx+hzs0BYpDhLR0CyMRX+1k6ghUh8728RZ+reu13hWXlQdG90NZcwIVaf0Q
QXVg5p2/DdLTE9aLYNNKp2b6+UMD8g+nC7OGeZhDyT0x9Yeb7olha6ck2d0iJ+e8
uZ++Il8XlO4VEhpexNmeLen2uJxfjKUzAvXSQ11YMr0ntbkQLuEJzUNEzJ8iqmzX
+YIjETFJKgEwlG12rOKaxv21BHFNRxN0UhjtM/lxuMZIStOJ/djaxwWdSL1J09fs
qUXEq5YJeaz+CU94BnzTg5DNM2t9jg882WScYm6+sXAUj2tsHJTrf8urKwgBkXX9
90gSY58JysaFBNP0YNGL6u724VcvqeAWdpYf6eJtDlePqJEiRXTNX9O4KOKtKykw
ZppSuz+UOCHRi2yARHqp8KX0d+4n5Yf134As9C/UJYoDlIMATf9CxB2W6Juwge5s
zwAAK9SOA7CsR+GUj+KIP/3WwapHnqiEhmVpPud7RasRCtCJ+ly7p5xZbxydER+V
7+OiuelkYsGfhNndeLMhOHRVBL8A3klwWjtrDOjhXLdzlORPXCNQ9ZTWF418Lxg7
f8IC+ruq+8jFN7caBjERPDedMW98vt8o26KPbbeYQv1SPKg1yUGFu/kdWUYE4OnX
K49KEpivZYMn7TCwLmpGyWnEIIs8V5gs4cqg76r3z7aEjmPoSHX33tF/4F91Htxk
NraSHwkkysu2wmJb57STJaEl28cskTXROHs3qrSUSqDtu/gFYJrsiForR6pMiUHK
s6Ddlvf3TRhzccZ9W54AqHKph0MkD2GMdlmXL3ylYS4v8Xm6TTHcZZ1yiPpJa5Xi
UFIxhpWAcCq289tOI9zu8qz9Z1OxBsNpqrAwKiLKBzS7lCCJ9n1xAool/7f+hAsC
r8JFgIwmctoSnYDxUBkj/wj00cWH3P8EumGf3l7v4xmdP4SdeEfch//I5PLxp3Xp
zEgl8JZjMQQUkC4zPBA6ABj9x6L6DZ+vDszm1lLrpApGDn7mNHWsnJCWX8nNfujR
oL/jWAGJxnW0a6uJEmHTqtAH9sWGkURRUNh5p3VOtQaaj97U6eOqdAn4CnW9kP4S
Um1XWzPa+Us0bNh+HBwvcBXmkgK/FFMpxhZH0hf60DREy+gKxc3LvTfz9d/fMO7J
Qheh8K66KEvfWAmnRLU0RoJtdRlQg17y3T/VeqOrWE9gklAOsxIJ1jkNVmaA5bup
cLjs7ZbJQF2I6+uBQvb/j4xDAgmy8Altq8xxf97PSoJcIvkg/nf8fDiNNuAiysX0
TIdm/g+iUcokOe/LPJb1cP9L07njTyZtVMaIeyhR8MWEkPn3AkljBqoQJouIa4LX
z715ZWELmrG8H64kjTKJgQO+qUKN4F28tsTl7zb9Rud8DNZubaMO5zLwf9xMBYeu
9Varz+Pb3Z6o3Z9zRhPEZ52YAxgPWatSD3HiBs6rhBktFuEvOCi/esqvYQePMrpz
dYJoNXR/RYs8QSfxkU9LTJGejhC1xQCJQd6QJy65o+WhnvZCXO+FK54zW2Ynmb/g
exqdA2UacmZV3+a55avtpW/wUixpFDRSjyhvS/WxjXu5tpsAGcbcmI+eVdeaYt17
IMqMnfriF6N4JUrsn75YfIFckaMW2qmU9HFFxAg6Vx3oxJbuM5D1FzF/darwd7C/
wQ/VMqem1g2LUvsUfSQ0ZyyefA8NQfiwED2Vdv5K5u2SOQr3kKvcWUW/rnOjZWGG
yq5qGxY3PkfCShTDkcfvtKKmVo26OsHU9BV6laDtj2f65dOGfnoeKW66+PNIs35J
2vjc0013Tq0eYCDUhn2StRoyDtYHqODQ93kZ/RcLq+chcGQCWjc8UJleAKPu5+5D
nZruHylTa8RxOk6pneQgcyA8mgDQJiLYMR/9vlwLiwxuFSvd+aogVzW9g4qfW8Y6
BK6RUIzEN5ZTfx9r4KvjJ4V8x6B6Emjcm1R6voR2ciclEmXrlBU3WQNOpLhZUC6t
pvQ+aa0N3ZjcMnJbVmqJ6wASdW2JJQ+IWYLYmy0nfcuxHbGCFlrQPgPmTQNmlNGc
L5zCuWJ0neRHBJZAmrpluFTFPZ3ZzX0z02G8O3Xw+d6r6T6lHVlYRUeScYH4QP5d
4AD6GEcZvSMAQ79hXQxLm1yYCLnKMOJkXRiAuOIPdRcqwCsJWfg2RqdqRTV9/gzc
22ZoXrJQaZsojANd+5BKncQwvMjv9UkLHXQCPz6PHUAwxAka0rgMkyiXqR2YVrpy
+CyXGxFuyUjz7LaTmIImBlosLs4qbjNOMrQ6nLfPuUHEvnCs/vGRHhsMx4q+zRmd
8SE+MdtCY5t/X6MtAOOAnsgUy1t/rpnynI2StC+KukZeBpaK3BAuR4OLIFcUxMyD
OfMqg4n7OYvCTXWx45P4GpHjYfNVtFAlmBia7bMxhv0gpT1wJUEJd/IVIyQWo4BS
/7jL6jLbgV5yd9vX7K+fD2BTVLb/KtFxKRZHiodUA57YDUeUxRr8Hh8uEZTsUqwE
+omKBXDnXpbMDz9bMTLwiCtir1MKsbPQ8O9B4uMgnZzoARppko9CDCDi8Eb9oZMg
eMq0i1Fnks+Mvk/+cPpUZJy3NeMBVAZIH7cVyft8uxdI11NrgWEI+kJYcHrk4P9s
sCIBycsWLtyNHka4J7TfiRpFDa37H7E6bHAVdL9aShk7R/Gi+03zDXTOqkYCMrIA
6l9aLNIu0YxSPpVlRGWsY3z9GBQpfeXhvv3twIUu2TcV+DCqN5uv7FK/V4oVuoPj
NoTa3ggDIchPvxtpdWibpoLoCUnrTDfpcZhg05KSR3v3vvzRZ4jyuISFz15KNLGZ
c1JrSqRsNeL6tqfFhs6PH5YVzcZuArB9xCf6wonStuZsaPl7ynsPc2OfVS9Hs1pX
e6FBREDmMB6B0H0kM6eXDJyOCwybEPyg6yiJj0fZNOI1u8cpZqODhAe+gg0edlM+
8O06pOxM8Fr0hU1ubuImQy6CmPFOL6ZHZksAIvTJtSXOZaqWdu0LoG7rquK3j5fR
5IvncLRTBdK4R6VMMLEKlxJ+tVcUR/Q8+N0YgNA0lm6HI8urmzkdsnoZAPK3rfrC
G7GLYG0leQDMNxsW4xuo8pWDCnq5ci3c4m280QVSTUKY/XFcmuEMTN368aH2Ft9r
f9KbA4xuXVn7IPHh/o3pyHj6O8SkokTHgp4W2rrkOLS+HKunUa5uMcUfQabwSgsC
wy+JomsoG3a0pze5SE9TSsSsoU156gzmvShb3thmHIj/MF9LhANbNefT/439XfVf
4JBu6CwXJ1s+IlTKykPoCw4eG2DWmsx1YD+BwLInaf8EGNxI/aauVAdqkZRt7X0R
T9SFkj1Ze5NUmGT+cJfVbjlVwG3z89of7rxISiCh31qfK6d37xEAVLKBI5NwaO4k
p+sFNolTifVwrmIDjPEeyru14xjRdsIAyASP7sYVSdynYzp0slhCbsLNwwGl9Ewm
LudDZw7daWnT/u9rjOH66jKNTW43VgIhioeptHbbhxdSiN8pExDgbF6MPm9v3v0S
+g8Yb6sana6BNzrIKxceGOJI8RGHAe0dR7zjxY6h2Pny9noJ86ksAkVY+Xq3wCpe
iV5UUsvTs14SfmyIf9Jjazi6v54pg9S/URPgM53Zhk0pXDiIqj1DRm5PeERj4yMs
P+ds0d3yVlVF5Ha83d/3Q3GrCqBygSSMzuOFcUQbrcN6DVgGgUbO+jY++TOis2yv
muLwCdpuB0zC1XJNnvvTF8jQN2Id8tloR4Xr3KKlQiuHy2oFCyEgGWe4+hkRZNRb
4NZ7a5YVoAo9GsLgydW7edZsmtT8BSuU3Od4bVsypVLcOhhxpMO/IARJldjIUzr3
stDOIOaoZ/MReEM6LfgLEv5+qyMlb1FZFhCO35XCUyKQC2MWBSC19hyLZujM7zJ6
141nXoqjmRkdlr4ZOPc5m7zlX5rpmYlvO4ucC9BOQRT/FlhvpzG7BzygXJ5oFgl9
b9DtJpKaOLrRmAB3+HJEkpY1A3xTRxnFF1dhrwWc7G95aovK24HUaabRYvDCclA3
LDDIsOqMQsxvtkxNSivgDCLmkRN13yuNpTmmgdS/RDRyvO639YSt/ksJ2BZKQtJ9
EUj1ZD36MQftAnTKNjx/nUTBSjJOO3cbcAMkhzHLVt96bUc/XEFsalSbNUcs9SJX
hii8vtVAGuVQhWoRSi0KkeGajdpyVqY7JgrccKdkImealhleMefMTnUQGHFt/ndi
rTUE5BWwp50oBf8FfsGNWSugHGqOoJEDSGeDSIYCwHOBhBaSDgURmCJ3JRMPp/IH
BQnshG7h8iY9ZB0XW1RDnAn27BJo0txfpqp8uHlipIi1SQyz3ZlhWCwTAhJDu5AW
idBu0+/4F7WPRNQItqayE3roMussEG1Ri94/8mFXrRNRgOmowma7LLfnrFkifVGO
lkR0GUxK5FzHlKeLMeLQ1pISOg4epa2B8tC7V75izAzoSNElNfPQR+YmpWJ1ZQvU
8Vi7nSjNFHYOvOxbWFiu4LSSW98Y9uTXAlOfqAHuxSGNVbE9QNMLJJSONbYp9MFb
ERNoBgpYjkY1Js6+tn8RZQnNPNbL4+tu/HJU0jpdQ8R7+ESwYYtM70DEZ3NydRws
eaw9NtZnDF39FuSn73QpGRQPBo1n1cz4ToJD2ygBuIGbx9RdkJA9NliRH3Xqt9oH
fv/VlzNs+dY/CYQRz23/UaTYiBONlxj5HpSWIN+9ESYqPuYtJaJVTcsTQNH6E8xR
6u91uE8TahLsXFjFGSAMkuGXOW3thEL04CbHDNkU6Z6aa2cDmUckOveaGe6HePK7
9ZXsAk6tIvnyTVl/xuWWIYP+rXqxtkCX2iZcCRTZKseVcj3BOrnKKJ31OBnWdNl1
EUXGC2M2EOFdPHH00tPcCL5c3MhPP8QSAaBNf9iydzDVJBQKei2tU/CnKJ7fFwRI
PgtkVulGPUC/TVCpuXK4ip9UWOmuxXQ8vcsTMGgjtTiTVkDXDAs1/pBsclq2GKnv
w59A5GfOxpRtA7BqjHTXIqGLNv7dsfsTN6n7rQ9utPcCXJv6Qb6q8j9I0MBtgy0f
ZlSK6WIlfmr2/sgfMcxtqkE91a6nfRbSIjXZI6RNB1DeLNnVnazATGlDTXNaXvY6
8WskYq+zFAEh+KxYAPD/omNEWBMRpclsCFX6g0dbIUao8jbqtVKLzBjFAlax+Npt
F9X6yGhDJyPOhEq3BxIVwWUjS86BRIF4BHQ8LoD99Ew2dQC5n9DdhVjJKAFPhTeD
2LjyLNKqI2SS6K0FpBjTMLprVwK3apJBX9SGt/ZYRHBCurDyJJcNfhtaEsp4MwDs
MmDpyb5YYhAKctjPjdGdMaXGKm64jEaKyu0sDpAHhvXX7vSED3822PrYT0yX03Jd
HYDEqUdj1n5PLZuqn23M7VWcBp03d787TBE9e5sHzu4guKwSBF+Tdmly7OLmWV7J
jEDAVA1qKPZY3aF641s4LZPU4Wuwhg3Idq7ENlvhnFqaXOYmI9yeQSqQH1tsYaiM
YBt3nPn8iMGTsC5Pn9KS2zoGlIP4NAzkLfi410UoVkV+tJ5s5N+YZdDWwtVPdzNs
Ohfhno74Wnp9dNMuW3xIUg8EC1EIY2Bj/8zF1mmc0+m/dubBbSLbCodWDXDbmQLI
NYKqpMvtPK7KzOHBPLrG6eLukvErtc1tO9U+/VOXbpZhZAMrQe8/0WihlOQO4UWF
kCTTaY63MYy/cJxIwRM6phdGfPQeKYA+Cq7kYQjrEUD3Cj9LY5h7FJWwW5yLwtW4
QGvubDkJL5ZuNDI+f5l+Sr12hTteee0KOmsyovrzNWA0tvzoHptd5v1srG6Vg1l+
O3PbEpzp3UHgSJeaBLZh/cJ5xioXQ5sFX9Cn9sedTphFO5Q+fN2OSAo5A+q2QIfv
ItzWB+19H4xWtlijLbl+3I7z8l6fGUOi2HS1OoKoDeuGq5eBbRRlRygLNXZnNd1S
KVV9Sl1YqVYhZtV1gp2z3CcCjyvUAfOGuExrPcnYSOO/K3mksNpHgYqV7WZBKvfq
mI/cLqA2VOmu7sYZPCklaU/km031qu7EDmbF0YwPw+O0HXUzBXWZ0CP6N2WTqIXs
S7+nsHJDumNJQvb/FXxA+7ljMDoe4Bwapc1+FT2HgaPkK8tbL30h1b/GQCjjH+uw
3YA8L+7phlo9C0Xq+KXAeNzxNt4l2Kdb43FfgIvz0yaW0s8WpZ47aofKoQMtTSRp
6JEe1u6e+l1SAgxWGfs4b4NB+bLt2UvrA6EVCOce7Z39rnAuE4VibLYFyx4SLe1I
3Kbkmip1CcYSLQGDk64TAIkxGF5YMfiVO671mgez6rhjfhPs6RQhYVqY8tGS0Td8
nfs3Fv2fkd2Zt8MRs99Rk6udW75Ayn1siG07l9+jHz7kJ5/0I1XWwpkUQyS3hzb2
t/euDX+cK+KgOKtuOyiUJ6aDpDsJnh4oVQklyPqALvcas/SmLr3AG2G+K6XvvOLT
5NhMGPyy6qf2Z1cSOLlxELgw+tohzQxPq5Q+7CoPvQK/Zf5RSiAcQzjN+OuKe2R5
izBG0L4t2ml/76w6zf+yJBTR4fYzsoEi//Tp3nDcz+Qx2bh/nc8uOllHzOpYhP8f
h1LFguxYXPkYdDxPf7TA4tb0JetmoShSJ817TAoqXNsnmKqCtpG+46Sguphj0RZD
BXkVB5IhuUUStICNflQre6GuNmBXfkVml4+pgM8hcncId8Ujh4bx0F6MYauKRlVZ
R4wGyNyGk8RPTB4CfUc5JBj3oD7n1dAV3UIN+cTf+LkVXtp2RGg7onXUot+Sr7F1
qMlbUW6JLNhkHOtkKd4xgY1pA1nUny7ILPuD2uGICLzqtBqazGre9EwyHe+N3Mo+
GijOyZoxBUG8e4T4hRfoxhuWcHpOf5PvJ73AxaP5HCY4uzOGSxFta0q7IjRsz2bQ
SY0+mASxsskm8WnBqOBSuADGxedVV4LoUm9n6xJpMgNk3qb/uIvTei3YDw8REHye
xFC7rQGJOz1sFp7NfVaY5lIrJJQ7+CmIP18Y6Z8N9wA6U1dQ0XcJz6Phflt5Tg9u
ZbzoqA2P0mi9TEypQImkwfvB0uKNiRPMD6Z//p+iobp6z5siaGKINMjXPK2KAvfa
e4NumHZ3tIysdEccfZHYMhUcYzVJCBUlikPKqVJ5kB4kknJUGb0jyc4Sm2C8Cv7e
aHKYcxi9baRu3eu7zzDMTXEWb+uiidiRxSp8pxEnadBMbz7H3b9NaeEQAQBbEJfa
amcb/jc66MIQIcuxGwWBhRYgQd2NyfNute70vcWb8svwPJvo6fwXpyDOPyHhST+i
YTFn8W9JM4No5mgAvK+bOUs8mZLcxqY3aIoJtemJP06uimri3aqo9Bg9uSBQ78wt
jaHwkaEFdgIjzKAGfO/+h2RrQzmMJ9ixhpLy9HA9eDN1vUPR1CtMPsxVrt0GhczS
LUeyplZWB57g1q6k7cA/xRZnWl1fliaaMmBHJH5nUTOn8/IEOU4a39X4VTLtb7kT
/vEE/yLH7csCdlcQj50v7Tx/0tYDNltIf9RdikktC+xVTxY9J83w5AtrQ2vWBiYd
uXYeEn0I4lyeom4uPIBBCzHuBf5tyCk5vAa+t0K6TZ0g6awLgZHjTOguRsWOq0cp
hMWemmpCPMooAvweYT80C6RKxqE0nmJgn7KqKOMM2NoKaf341IDOkDq6qs1TZcFZ
08d1kACBoR+Mxn6GIcWS3OhSY7nfrKOp/eApTkDzFlygj9oIbkERRQK/31YTkd36
CvKjlewBKbKopCngBZ1Fuyeltm89C3tYbB9NsWoT0HoCfF7rcxqf1aXFLIlyRQDU
Zp4VT5Gmgv6SALw4lE8Nd9GHgE8C1mKv049t6kOzH8o2mOxJ5mhcSxZrJ9jTzn6q
EunFPcdoRXC79m2Pz2VuRJeDYCz4+VmhQXPKnOWhxOJpU3h9aTnte6CWwcYJxVNw
UccONSHChC8zYPbbbeaAX91uCsAvV4mGruOk7JNz0fGGbWSAr9RR/al/J75L+28u
KliH1NWnwrvJ1SdwTiEOgCrP863k8rCc6d7QUWQc7b1SGNgwSyDLLjBeWtbtmJtu
H9cMjxzj6Ofp2eJ96w0mCHTBV0wvp09ssdvdVZokhe8dv4ss/3FDSjHmtJp0J8Sc
pxqj+NHzx486i1noPWAfR9OKKelPrGLTxlaEj6X5NH2Yceu+4MyyVjZtSiv1s3Yh
m2D4dyQVYjX835x7rRJW/yRtek5dbx2heh0hudc9N/M15/gs08hMr7gXhCOT4qFC
Okn0HDDbggTbJuP/I/qO17wHMhBCi8iVbphSVr1oEgi/K4qRUK4mcchCkzF+UMPG
ZiAVZeziQWfrpLUm4DZkHZvuZjqQ327wV4/WXnDi7Xsxj1KwkJepMm17oG2K2zda
uqvhZ7PaihLvCoJP6TC4ylrljCa0tDF5WYZOzkNv+W10/i2CsxKveTHpa52Asxsb
yDOnOC564ruGuOaUXIvZuM1+bzugC3L2gSBjBYEsWoYtBga6k4OIOzdfHLfWTUX2
fle+n26o5ahpZV2eX3ZN3r+Nr/txxjLjfiMXkpglrXyQZ5c3m5lvMxo4H5he+/5j
8lm7L7PNhSulbh4uN2oBDWiutA9N982oFWR4K+RIS7bnsgmnCxO1TSB6CH+bjP98
+BThAIMKmY+rbDzXcSpEVk6IJzheXfT2/SLd3FyAXR5AhRDsyVSvIZMF0vl2UILR
fCgDw2/rfpbR3+oeOizIhHHUjHhNgqGYcbID6P43th/3JWi11JJfu32PPo4ibNFs
BdQCRmcngZvaxQNRJVTFlVyWMEBc3hMCS7hXaQTJL66T9ZbD3XdnjrLy1Tzr9qif
SzJYgNBUHpCQzxyIocdwMX7zWbD+h28pe1KGeTrsQ+MvwiopLeMh5rfmNCyts1dj
PmioTgNNlsFzvhA5me/TYii1txS1O8jjxjiV1bRpOouW0Td9uBXOYoDnFqWuNIQa
E4RRlVZ7M2K0ZBXv+c6/f2byrFbJq+IisN6CKVvtFwO0w96gC7ex1+GxrhLxK8Ul
nFnPPRSAIgjvOMyEHBVrqBhtTJnrqR2mgqA/4EGvKWEgJ4nr/NpN++DpKETXLpA8
j+Ubylzl+PvX0y2XpXf0WhWe525w5ea2J5mspfBooI9qRkGbkgpmqsqBM3Td6D6Q
D9pVDK9WjmOVy3OBSKL7L/mNRA6hpr/aGzITjHCSd5IRboc6IzyuYgrq6ajHszfl
ogV6jvnWU2UXg3Gpx096MphCRBBSs7JytwxebA0SGi/WheYk/Y/wrH65tNZjaRjZ
Hy9FZdj4mmZzkOsQwhVSKDeg41qpP8psiVLsiVNcHeZFnyb+LIKAn7C8HXamcUJl
sB9wCI7+HB3vbc8cG3KTi5JG7rImTbo23FjiFeXmiqL+QUXthSQaFSe55160tI7C
59HFQwX3f+w6snZb5lJ8296RGJ4gZxk2mxN74YREJSK/wrUoftK8NEA0sZXsnwcJ
DLGT44osAbwT5TTXOGnlAkiUtNEudNn6fqfx2riwrP8wfrHPD6N3fCzTbZDcRqXv
UZojKfQGRKygKTQ0J1oZihQSbJcK4I/Hq9dOOXflEV+qvy4P8OIlZTlZTlVv+bt7
ADOToZkUeUStZeZ3U+ZY9WADHH8p6E67YAUag99H50ubiEYyYTQ26OHQWviQ6olX
8cxPp/7kwvrCxtcfCZuoKXZbndqb2MAYhejh1PF6xkaZ7ME+4wFj7GeGMpNBSpoT
QwEQgP8K4JCapljVCOiuj8VAG4y0vXFI5hLPveJwlHc=
`pragma protect end_protected
