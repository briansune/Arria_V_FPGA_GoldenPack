// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:19 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jZkEsbrzcWMimRLk4jQA1iWjz75tQZT9SQBsnAapx9+RzznOrYqGzJHfNyiVmBD7
ZJ6I58hc/Salym0vdvXz7i1dIgsOKQLtye8+40mqsM/bvs5m3WruYWipvQDNSJDm
rjWx8zn+tfudCmqDDrcFpAuvHyCYVLpxMnY/YvIlJaY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
Ygs6skgsNZwccIKS80MwyJwoO1pympIZ20OXki4wP8ThwdVLa6LkGaIi3pio53PM
X5uKYG8cSgmrqrPndeGBzS1wPIKKTIOekvkDNc1oaEZQQ2+TeqFMczXhra41vPP4
MSA7gUZ0PIJZsL4x8HuS1EF3C9uN0MSGNxioqpr6r7GroLfTwh7smcScewdjAD3q
8f8kgCvM7jebBBYnPRd1ECo2CCt6c4SJnR+RLcoeppVLXn5K/pVoJlJXnhEm4uHN
cC7Bhyqca5yE8c1GDkEkfg9oem8yW/a7zSNbnsj46FbuSsQGaoDKw2uwxatjgKx/
5wVefIieUAQg2uZWOrCIhJ3FLQPFB3VpL6fjRzbTQ9ISpBRU7mcvL+CxZOdgPSYV
UaL2ReOGHsimxyICdD2KbX+BojnCqYpglj57vVeR1G8T9J3JZR7ggUc9r7ZYTU+J
x0wsMqZ6phFHHymrQSolVtdYbFl82/msmhvHHD5VqM0K/jtH0pyxH2+qC5SozV2U
Zufi8UGhrX02sCrnt2fRC0O/uv+GED6vmIfPUIYq2HYVUB7e41CgXyY/0GQ+caYc
FUm8lBVWJD2GHNAH5xuLA9m6VsD7+xAKxih4bbYAKyovta8ncmA3FNK3kse5E7vc
Pf0urn0x07qP5x9QadjyCt7gt38z/Dn9ozIplboz1c5W/He7sIoSR7gOoTGZAmHs
7ReZvBR/RbE550kk9JI/bwq7GpD3f9VHB21OjKokZUWKsS4Bxvwr3OTKLo5obPA+
UMeSopgujWoJle53xYtwQ6531Pfwdi2lLBKEyHiphufQyCJ9P2VJQKFy8468xk7Y
Ue6ocr1HuMLylk97WRNainbQ85Hd+lrC5flILTODpW4HQwS4kSneZoXw7YSaW8sV
Swaaqh/zg2vPVojHO2fCpJ5DG7qpKc3kB1c4H7WvCtJgUcJtRobYdy7H6XfH/P+S
0HLDWF6LiRtX9vLlCP6/Ocs02iLuoygeJX1ZlkIgWOVVRBNKHDdyZvs05GLFnUst
ZGni4DZz6BmMYynqS0/9wMyavG0whi2MhuS7O5qF96tna7PBxvhWyKuw+GKQ/985
6pxL8RChdbw8U0sP6/zv69yMUGbq15K+efkeIz4eB3T1ibsURSeRWlhWqvazSDc6
rmQyUqc0r1WuK5i78VjFPFDm/JbTatJxt3Oi1+sKIojKYR7kDuVf2bv2vjpuAd9Z
rerdGAHacZf/E3dLrwzUNL4WXsNJo0WcePDBEYFvBImHDEnrVll0SbL9K8sFXIfe
Y6DiT4XTrttMl3mTummlRXP3h6Hyoqn7xKmE6vvIZJdSmrAKrv0qP8z27mq6eYvu
96R8nIrt1P/uxNrPDuLG7Ji5mIiTgxZTB9UXG8KVvYzGWeuSt+Tf0zPK+GqbeJrq
YzHi4MxALU5xKq31sUk3pXjMUdfV8Lur/vFfK9YUzYt0bTCKVFvmrbi4G4vOnjI8
HWc3aFpqn7yXcUMHoGfospN4i2/v0kgheq1UjPL3+i3ipwXxBwyhbU0XdkIGvhV4
Gl0wxg2g8wsVdEdw1wCFEfLnLCszuND8vABy2NVR6be7IrgAc5TWobdSq5SmAnHb
RRoPq6KsDnbrB9IuYYWIwwoiswLBvaDfxc0E+A+U5VolHawOO6OU3BhMBsRRcRqa
WZ7h4dzwGPVxUA5Lo52RzfiMddKAjjO+O6bsgfQJfH1p0ol7q8D+TtAWzVqtF6BT
81ZU9FoePVbZLBnSh/7SCT8RmZ+jxUrucqDOh8n9hJxLdlt3ISnfA6026OmmxhDc
9J7w4KZby3zY2K4ab7eZ1TtQ1TAEHXsjOJJWz373ZARFkJ7/gDHeps0I773CpC9k
hRqUM5bMFujZBfRUFItqsROK/xsg5fYx4mq7IElNQYL40mNvUViy8yQkOWg9Iu/7
msTAlrkfsqUvYWUjkBQ9K4FRoroIsjV+rFCI0khG9uZ1KMucfq9+o598T1q+2wrE
OAd3qko/4czeb814SpRVOGmr3tWwe3s2Rf1XJjl7PVm5zdccJQYUwbzLbaMGZ6Rz
GOD9Es31QWHsdhixNr5a1MHtQOcH4WpEOkYWlxW3p29gk9sMT7X0hUaraFFj/Ziq
B63XX5hsvpc+ikjvsf9HMjP/XNYo1U+2VnHSKI0XFxEIOxSNjk9Z57aYCfOgQcz/
7f3EF0OKF+NAKL7yKaYfyn1LrSLuq1SFa4jUMTTN9faGQMpkV8EjdBLKD3SGth1Z
1nGwAL+lPRg3GZs00BHm1WDCQywsjFH1M53R+9lcELAzVHZiY7LfBLUs3eH0/WZO
XSQIiEE6cYrQzbs1TBOX7hSTyVAVELa7yAhDXWf6RsO1tGSQIkWsdaLYAIKpXEak
li0KK68F8h54XBvkhQDEQxrABI7vxvk01Q0Vl/zy71y6dDkEo0BMB6oNStLCLK5o
g6Swg9sHkheWy5GHrjYPCpk6cYLGn7GLV9oRbzGJh2SKvQVj3E3SzDL6e7vXOLgl
R7B5mJPaAp4qG54JY7D7Q+CA+kTZXc7rf0vTVQf08mpbz9c8FkZEnRI/Br+qd55O
GVTfkCgMGsTQy7SaiosI2J9HnPzw+4/gY8Z1rZu7bTQUPMY6VOyY682k5UB87I7E
MA4vE09lTaHgI2c1ThSwe5c3ObVuIXMYuk7+oDjpW4Z0uKeD7b3i+vg6/BKyyFna
0Bx/BrrEZ6tbQzhrhTfLVSmumSHKjokdSS1oHxi5MIRJw5Drf4dAADTs52//fx5D
FU8+gkhprwX6Z/cSrsVOoSql3LTcNvomV8PJGLDkjqPxRUf1hnuMLhKMzPEfCIg3
4qQyA3jDaim4Lz6mZ3JT4Ws7wjCrRJzPsw4ysQJuyCb2ZRV4f3B6w1llErsnZRTP
+M0V768xBD+1NcboTmdEpkGpWFLNtcNHtcFExY75lkpgxh4B3g5OQX9OSdGNKX6n
EgGlYeHqfvVuOhC2ryxiMKtKETv/NNh461kuqCWb/HAN7eC8Ps5gcz3Wl1nRWCPV
e4TQ4OzsLrLW25oHPwPVi7oMtm5BdsyFdv0aGfRovzAjLKRVG4Ec4tBx9AzlvCPA
bP38hxZFHVeVz0MHJn3EUlRxvUX3+sGmuTSIgJNUThUAmn8xD76UlVFiEIiunXlM
nimQF1tRLeZiszYAQ3oFxP+/1Vs/nScJ5WEGn8/f/xQwI/Zbevz4OK0x+fBAJCug
/iC3CWqE8D3icEpxZZkdTU16v32rYqdV0t6DHXrUaqLgNufsi9ysgltf7ooJGC4G
jad+MHkdmgFMIRITipgR7F+ym0frMW2tcvluuKN98e7zjE+nqbk+GPco0uXUooI1
wbRyNexnWjo0QfAHHTKqwq9WkqGwncJQNz/RjvXdbsexk/dDoIMtzotggtAMs3/z
AoB+m3L8bxO+uJTrWD4AnBCE18nqWalLCUuKmvV0PLnO+MUtCsZZIaK1s+l35k/o
ldwenErI9Lt4VhBYTOb2yEuMdF+wVHS7Ic297+7un4xifN88VjWK0qCV7Ucx/oym
nxczUj3HcESGZNnZZRhW4EmSoGZdA3kQdjOZLVWzwzQETeFBpWZuzWNszqPd6hp0
kzGA0s39GXes0Da5x5CH96CaKDcgTd43+ome22TkUOOAdQDkM+qTilxeaC9R5h8a
SuBTVIg9V4SjcWiOZGQdzLCeo+G2kAdAmcdVFOLmOOc3N1oOF/UCZczU+lDHrDPg
Z8mXXSKVZn5Epm0xkiuT4I05zVz1WJi6B4lzEWVj9YtsGAy7AuqCVuj3LarNRQsM
hKnjaHO18ya4QMDgJTVxux/tA9GO1y/Z4eofcYclV+G39hR0yJHfrSMT2q4WTMod
/UaycxGHm5E37l93E1S7xDmGBiAWKXMotSuYGl7XTSrzujOQfhtqoYEf+XLZIk6T
jvtT/8XoLDuwMJejybSTv/D62mt2bFeL/BoIBFq4ByT1IGWdt8N9lOybzU/XAQhi
aTPdvoee1NaijrZdWm6QOzzJzk7a1XBfbWMEp1s4ySlCn2PCLPukcEmkpmIpa9Xa
8mJOCz9XhfmdR2o/tXzloLXqB+CznGkK8wosxuQZF1UZVXj/B60Ifet307ZCW5dy
ATSgPKmBn3MUo/UCEm8sYkVD0MUlDz5FjnGP96OEY9j9YnpElSkK6DM3H/izpD/u
5WShA1rarF5OylNZgF2jxZSME+xD820Krkhy19ptve3Etcp9rh0sJMTgf4p5lodM
haQc0o53/QheM3TMp/NsqsCdtaIL53olDvKeG+F32aSQEMgfwQ3QKtbNPqY1DEQo
8+wKsS7JXy7/AR4Pjd3keXU+HmysK2rKfoV2zTOP2mrPHbgatYR0OcO72NGD8rkI
1Tj0NT1ea1f1ncpquYCSM0PS+bR/h4gctA+G3so3J79xoP11mtJdKcriwW9bX/pW
+BoLwDvKxYgIBmgoWEFLm1q9vrCbBEJwwZH5oKJAOtTRzEFtaqaj30POKDzPKjMD
DpTW5t7wMp2yn3OywbDo4TrjhPSSk0ebxwYgGeAtY4jSAfrRPkTXy9loJMHn7A1I
UHMVPcxLKmwhdu4T4EVkME1nIdEPRnSRPaq4kEyvMBNQaz4KSCc7+kErey3JeHJ0
3Ve7UARRHqdgdT2xyzjJHlMPmrnikTEULXiQbdJHiR8LwJTmprDgKTQnOKN7U+CK
TtKPa//YglqY9qVnIXxktsSglSIPlJ97W7I/lEck0DWfkpE9QKRq1ypzSPcf5hgk
ksbnPQtOsHlR3qQ08J/ZQBk3XpMPuRaL4WuHEJELFM9HZjodYpsQ+MVBpYaDGOMA
L7rJTMY04p+Ehn/HqR/cqfF2OYf5RosIQxbTe1Vyz/2jAdUFGzKt/mXBz3KzKqMY
CM5HbvDCYA6nK8PKO+NNXO4Oao5hDh84YmQ2cX1VgJNRll/Hlja2YzAQsmkEK2Z9
ggxv9dcDY7tsdmssZg65ozKwpJQQ/14wrhL6XigaWcBR40TTPD7h5Qz0qrIzJV0L
CT8NIvMBlnfAyoZiEuxqrJWhW6vcUbTwXw4MMdAS5QqU2QGgInnCtYdmm0MAJc2D
azDdUX23bMcCeHswRNM9O87o5U4bXU6K3+e8EDWTrQ8fQ4hh8T4YimmspumYJyWL
KsL0sWOfrDhbUXjx0Voj29oE4FM+gwiEluRxoM7BHJvN4kpn+Mot7XW5KV6ePmDk
sSpoM7uL+94zlasdUSSc6nWpmRhzvqK0nqnTzUvbn8yalFLIUkG/JCVF/cVWKfYp
KsjEz4jIdsZdae6OfrKTwhyCT9TNbnkJ7ZnhzfDUFwdtrUmN+LLCPQTNmjL6Z+d1
Lw5rLTmrVgfvl6J5TlVVdn1eESXR4FuXw09hwQ1bvTuU/8qKzGjpzU41ZW0XXjCi
G5weMiIkmIP/T2RvZBnhP1xGbLCNUw8r9+Sl1mwKHmTHnRiIE8bKoKN6Atlrwz9b
GPt6cVmSGbq75a6OBehWlliUD8EfImZ3uUgeFLOWVoWfLltUZyzGEltAy0CxYcp5
vwbSjAPaKrq0U/yCrtDYiEWhjUUz6ycPuupxKfCLZeS0rCaQ9NFL6ApJkNC4W4RQ
WLZs/x2zzkZ3vTlulo6OyOL077S0BSJJFRqIOeVZYZH8eQ9KdFZsn8tz7iY59Z1v
9CrPIrvefGBgzn97aFHvD4xWtXbsmEMyr1a0UdpbkdxgVS8rNbJ5ykvk31PIwb9k
uUaSSYQFW0tfIRGzsVrpOGsBzGaP72MwhyYBPwxV2ezrTFCr/BGMUk1FCXGr9pud
+ZCAsa16NA9ZXaNInDqbrtcX+137VerMNaEB/dbMgIaM50mJ4d6ZAjYIzMKaUZgO
ypMNlsEh+7IP3UxGiCvOaPgJjrRbeEiTiYIutPlg0ptw1t1vo9YJDDyRP4J/GE1/
IdeWv4/mbPjoNK0KJJbU6yNEdDN11HWxfPA1KfJagTBa2E+OPWVAM1pB39ZqweMJ
hDF34Hs0kP7PktTvr6RjA5QSp2YvwbQkD52mAUmDweC2Hj/CBjPWHd0obVyoKpNf
DIiKWgTxPR8xTqf+BZ2Zag5pfEz/YJ420wcIj4NjPa+fgeh+b3VPL5b48jm8G8R1
ZSxDUVOiucApNaRyDCmWESmBqQV/njeQBRMBBSFlhZPiYB6M2EmkyKNWshpijT3u
n+CM9BbgaKLwXLSVaikUkX9vb5e/72gGrwwU9jlKeBq2RZxM/zzqr4PY47yFri9H
F3iYcAiNopV6UfQ1lJCoUn+Ty5E9MjgKv6Z4jQesdpch0BEAd8HpeFjOnGp/ivZI
nlJ8v50QmT7fkGA1bWAgHWqhn/YESvk3YTvJRebYZ1Y8NXWxNN42f0trPb+gDuvu
JRp2tyMgEb1iGePedQXVZhmIzR7/VOi5X2zXX7VINe2Vck4LEs+evYDOaAVYSya7
C0yjbiT24g/ag31xF3mMbrvgr3fzxa2sj8YE22qOeydCEXp5I7zazPnseQAmzWXs
dDxSNYR5wq+xcFq1mR4BkMA438YNWr+teecwv8jwHK6HPrFwYpIpr6Vsj3SFsMMX
sHuFvE1lhaHc/CxNSDup9zT25+b1LzfE+9wu245Fpe5Ych/RMxH2ESug1pePS8k/
RaUawf76lLI+Zh1VlmZ2Pdy9FvFG14rN95FTU4lw6SJQRqcarE5ZTrDcZ9ZyrFZr
qr5+2Rd/cJAoJqM2LC9F033sIAwSOxpEve8ab5AnqT1tPnyl+adi9XMUKYPdPquM
eWxe0ZvF08/WBt4sY1yM5ZvUX6TMny7rjOEksHpDRoEpvmJb7D6v/3Esaf0MVgfj
CeRyHj1Psrjb/q7CIgz2Eec4yzAnVNf+WqZlb77ihd3aaD+sHluFOlsBcvhgs8QW
CE6kZRIuaIo59GbDtsH6GqfE1kENVKUSR9B8Nf9LeFlrhGJJCwFIVFh0ga7wK6wH
jDqiTHfWLOhNuvl4d/vWkuwBL4cqxILcOry8EYwZV0hOeVuS/KzTqQKvwMufJJVo
51qNA31Mr5p3cFhWm9dAEM06CbNkKpznO4v2W1jF5aGSCg2SXYRkmRnDUP+pFfud
rkyBMo9EuqCfQEcp3vuSlrcC+nM47nMRkUqWYg+OXIUJvfwRwykKAYBDyGJDa59E
e/EfX1i/YyNx8IF6noQJVqW9bTTxSKvY5uVAOKBE6LdKD7zqtwoHO2504yBo5hVn
Da/pD5+XKdS4uQr7k8074tXVBv3xDy37RuKfV+OeDUAMm7cqpQCfUOBlrUWmrOG0
J9PmeS99RwwTy5Xps9948Whb8ww3qbcowNbHEEZ7f5tkR9BpvWxUeDlyTfoCEoJo
fYP+WhBasei0ztltO6DbRF82Ps4yZ5vTLGqWs588R8rj6wLIecQRM4AjyZ+v6oXB
+DUHPqbFpyyMY8n/rhmfeHZiaAgTkTYbeTnSukJR0BRrK6Ee/0pc1lYoJPufw2VM
uFrFg7A7CumkXaVuQT4T6StVCeVFRmR+sh+jWZYUDOdqObCTSOc6rnuGF1PaP7qF
ZwlAvbsU8UtFPNYAZikzmg4V7JUzoGDYsz6kiHbQLhcZY22mNWignIu7C8LqgYPU
ZomTBmxJo2CKicdAwUrRNJgu9b3Nv3/JfqorfRqdaPyiqpC+Kz/3JwtrDyVTJUj5
vbDztz/Dxd1+aLzvySlRmUkpPNs00GuWBxxcG4egYmITLOjd+LrLZrLzFZH+5E1o
TK847/VASk6aE7sezgFY4zRsk47vawN2mp+4kjUv/bfVaJUVt/2QnBosQ5oPFjZ2
X5LkvHsP9JWAsFeFRF4hSCx+wlITZBhM/LkMKYEviXoMU7D0NcEQQfBCI1QwA5sb
MdXWjNz6XOy7AsuCGYeXdMgx8iysNeqidN8geWIrqqF2M69cyuezmDXwnxkNpyMi
t6HIYUaPxINaZshtmJ24EXsNFKc8lLmFEfJC8xhjurz07zbDknDTzvdZUkrDcPyu
usRIN0ZBSLkXuvSE0KpJrLyrWyLJ3fA2eoU1PQSet/lRMfkGU/71oQFyoUaCIPtq
aLyTqxR2mooQPICl/7rtvectirrAxMKE67L4RKPUEdmtuBsHs2VfvBCxyhQ49HTS
XWyMUqv47siuYM9R5rTfPubK2gdGNSes7n/NXvQ2Lhv+qBJW/mlIL68bcH4Dg1DP
kMUwlJchlqzKOR9n16qCVHiAkZs46ZmlD9ubYuzrvupRYfMiSLsMwV/QNjjmuYv/
F/mf0G5X+fmda3qD0TrtbAaaAIy3GUxmhmnONv0wel107RW72jy/ojoIIC8ne5vN
RjKchWcLIZsa/S/tjhTdJFtHesPc0L2U/UE7ynhEuKiMrvtBiGF5Z/QLLdwpE21X
b+AXTkM9crBso/qtwvIyLuJ+1jZdYb+M6QoaSVkMUXek0oaVUckpCqQ0vcqk3nwd
KzvLcuQQFy9Iyi1Q/keB+SDW7KH8p5hJnJBTh0OywTqoy4KgagABsFPnD6uEUfoJ
sJRWS8tIKKcYWbpygJmoSq+Ty9tO9Auwt51hVPPPkob4Ogw7BWAPilZxpM9dEXCX
8b5004FvqPkyFy0FAafyCY+pYZ5KFpretvpHjQeF/gLqQbzozVr0VdWFaslqku20
ksMMNJumJ7Uppry7moWUV6xrF4P9mYexnv09S9yFj+B9nifrntJYPx2y+ZqClOcw
cZrs823xrHoMf6BEDJHfEMhFug9RDN0TyZJ1kmxzGuCXVmjn60cAqyCWhbbOpeun
WoixK+e0ly4KZWCNuWVd3u7KQUhJuOk4b4VDenfhNJb1WN0iCrLZC59zu2Y3rfh2
ezAD6bFl9N8H8rLhuREbp2saup8nvMIaYihl6Uf5IRaQsBws5ImM5gey5uGnCV4Q
7fPieiDMyWYWqo1iIdIHsTUxGIFp2kNMRvI4en3xM6YGHzqfMI5EvtyYQgPRBBSE
TQ1U9PM2z/NsoDz/wq/vDwAxGcX5qGEDN6tYohVweRdDFvdNLYHUlbH2+u86EBPs
0KaiOfsdzc903B4HmoQDPOz88k0PImb8QHj3sXpAELw4/ATJO9kcSbI7WkpaKxFI
dO2ttRBJAAzLVB4SvLqt4YK2YyF1sFG6hgXz6+bhF+MIPnkM4j07Qo1yxZsWcN1o
qryIMOROre7OShXzfnrZHkBX3XZ7LVVC75OlJvJTnbPN0Kwe8SThGqfQ++K2FNke
Oy4SZmk7Tz3Xqi2/HCNCBDoz1kaH6/LKnQxpEEHb3ukNr8M2hHZlUyuzcgj4tpOz
KVcLGqpbvikvZDUjk89sWtOSt+oP1V7fZKWyh1IQpWb8qIVrIl4irMw42nKVmjbt
KyVT+4vJREk8zJ3ZL9eXBgDRVovuNhPLov8vPR/1ulggJDfU9r5W74XDZPv6SgvW
YQpxeeLqQnpOPab6v3JhPr51xNQJZtJOLFpHR7S5NiCIvrEXxHIxUNDi4ywcdSMX
av0b9pDn2cC1Sb16LHReuMweGwDnb6JsfqkO4yXtb8rgV7zFTFdbIZgUQD90z5mE
Ef9209xRYFqJhiGyLvfg/dH13Ly7nD6gBJkIbzWftkNtMlbSe8vLjloOb+E6cld/
PZU/1Wzr2VkINwA3TqRaOHqS0SqBftzU0+sL1DaFzWFKy06Psro05+dEZXhA7UBW
6N3IFGI/0cY18OynRoycJMEZ8dzEQvaAD6Vn7j+MmRwfqVGdlU3dxE00bfBKhOIw
e87/urCrH1gDI022illRG9LgCGcR/80HDd/6Ey1RrijBx+TiED2chVDS8X4K9Ixg
xRe4a3eJVool/vw+jP4uZl3OKuSN4A6ZQhZZABCQg2GAHLyjO9oGjVVqYCgb0/SL
u6VHvnm34y/j6Xg0ZnBynXzNSbls1aadZslE7veMmEADqbyliUWLp8q3OO18SIQT
OmBgDJIyDY60A7SooEE5obMMRLOWlBfVny97em5tohGc48x98mzI5HPmVf+2d/48
v7IX7Exh32mj2l9DnqLPlfl2dkF2H6lpRtHtAmTYrFChpe5SktKPDnuWwIoaV+55
b9sy4nv6eDBrLpVrYjaxUhwMmWXW3Vt16lhUbMCnc7DoNVrJ2y/V0+0O13aVwmG9
UyjoGIfbpSpH8tpRPJaZVLHGShLvQw2un67j1LdHmEvpyjkes8jGPpXjinPHdwfK
98zZWckdiE9ytn53Zi/+Bg0rlk5bkyEG9/e1i1eqYcK4plVkHvYZUkDDQWmIMqJp
i9f2zo5lJIR6OjW2tv7nGfs12iEKteILoA/ruv9rvU477Mc6/manzBJJLKm5EmTR
5F+9MKoOsuKxeah3xzEQUzsQ2Tk1R6OB1wHnpCT1kajDpgxqy45QrdJupyRoDzqr
JtqWy65hBcYkBAwY7tYph627rFEQV56s1TbQn+RESe2JHhfuMAaopyiy1aHsqtJh
TnuuzsMo37jpYRa1LsfuPXXCVQBR9Q1QnMA08Wb5YDQxY4KfaPcNOcFUAJeaTXiC
WZ6c30cHYFRxKL8ezEif0aRYxTsi91xNDAGz+O9dBZI6tvnzrk0DDmGuX9ihKqnJ
ybmxGVeJ6bcZczrpEBBxtI5l3uJEQHV67eosBTkykjul9TZkoyUIJFGaiBYX0Lah
JdKwOBL9X2z2c7f5ren7WfN+jIWKx1DWGe3xER/UrB8b12dhh910VAJeinBcXL1d
NoXWcBMvjWSFTfgft9+v3tlegt2m38mYmy0Lx4aqBIfzhB5umE2OFQu8qZ6r3+hj
20SuoofHXol56YkTVZQk2qFlPcox0Sf/TXn8Lc76l/RwNpq8hGjKt/eL8vOwYFQt
n39hHxCG2+evTxksJdH4F5GloyJ73/VqIqMIkaar8UNBfbXX2TcWH0h2Q47nSh0W
Bz3h+0+ESXvzKjKA5yPzOgTuQI+leR1LTsJOeP3/3OGBeomRzv5oAuUMR3PMpAkK
XLWDu4DM+SS1zYe8BQAmd6KBNq9byAsl4F0GTT8u6kwXYqQQXKFHeRqx55Iq51p/
tTaxSMt40PjCihbrFeyrA6HLyXftKyrTANLreaFy8earG2k9epjkFU7tQKQRgQ/H
Ul3AtQgi3DcLTvV8XvRobE0MKG4wET80ctdsKz+nfbfeQU9MyIOeWD8I4BXua6kR
h6LU10VIxhk3l6a7pDw7hOw3jg2/38yIcpCSSBmB8pE7NBE7qTxD2ICFUMxlZtbl
LKgYiJ7QfqGKRUP2/dG3gjMhPiSjPBAbzMdF7BZcFTFZYx9xJ9VARfKq6pMvJXFy
YsH2LF3xz4Ewl+MOyCLglNWpHtOgvjLEZ1FaAjqZfPQ2Px4x1moTHPdt3bU9dqeA
rWq+ypWx+eBb2PlMNB396RATQpKu4/WQO78aDb3NuS5T6fH214Nzisv1eJHA4j4F
evCFJwflnjQ+DQm0TBzz6bBC4xrt6elxspnxsC+edP/gYUmhPali7bW8GlfqgEjm
7QPeLSFBnRlORHyH2rg/HNxujjicl+3vX4THMD9++I5LqE8LRxM8lbQbdLuts/Hw
vwLprk1xtFBNDQMh/+ao+s9TJxn/DLJ7P2PjSeHY+uKtjDgLFMZoFIrzHeh3heHf
FEP0zc5o8eLANlojl5SbMCBlPGDwUb9o5/tdGEPtzz8WKLyQ9os9f6iMQnTzgZoH
3mV0g5vvWPulJpxrHdU9B/DHD5ONCSIXIWccw+B72YlGMC3J3ZkSjceGmrvaD4MI
Lk0Joe4Bojz+7NB5D3hx7aiS4gO2nkmO/3HIwc1jkkr1KZZdzMRn+4MJdsDfu6tv
jTjy42viZoMV5BOudoPeIt8dKmcEJnlXDRM+l1OzvCP/QEcWCNbaK2T+I4jquXkG
5gZ+ERmh+98EAT+Z8Bmx4G8mDflYSwTlOICJULlA/EjQQtkOavNlkdrMwbIc1cVb
gKW1p6bm8AVn03jc3w8ymoO9DIDn9fVdGaTQ10k3/CpDdqJ8MA+/b0cP8vVjlSpX
7s52P8sqzPeCfnK46a70aLFWD0EQ5+EYnmRmbmJSrWFEVdtodKADj1i0bUrvkXgc
DM6mBHTfh/72jpJEecxCDk9yWF5EpMjGOEVEarNZA2PCk2EdH1ix6plvR7zRKJa3
k6jzjXoyc3kdvuYpWBcEV9HbIUe92In/8z8Hqf9JQ7FCxA6ksi0V+AirozuUYzFT
0Sq2WBCqiXyAzQlPnve2ZB5uFysQfQf6jWYIgFc9BM+6cHLrmz/Q6/lURsmiUiha
oUsdTLNekvICYAUNo8Cps4mXt0Q40GPN8yPidKvu05CHRejvciib/jp7/i7Q1dsx
Am5tcclt7XLr5uO+3RIQg+QLVe3k2O7GYLTFoGzAhwaBvL5dsmT8J1XpAkLuR1Hc
J9VEHO+jmD8cpT1TUk8BSEs0maBTHl1Z4+msN9FWuabMu0Js8/2JL3TQob1C+re6
SvZMRbKXRc2i4j9ICiE+uROu8YVnoRBJb2PnX0qgHXuOwQVgpvzpPCX4cN2YHQCO
FqTes04gQ/WfF0uwPGZe7BEjfwQsZJX0/V1z5x/vgRb/xizFDJmCNY/iKrRzbeIE
6R7EdfyHvUWBb/MyJo2FhFjA2T7NqaeRix70xSzGMVzxl8t96b8EcP2uqnGvT6H2
/Ff94eSOYm4UwBXD/JYeqPG/6QIDaR7N+O4BoJ/9OLqQkTKFK19T5Bgsr9b3VWt7
CwZdHS4fGRCzYLyxQXjGxwzhhvRRkh6K7mCMp0AY3t88h2ddidlAqHMBxIhGSTQb
/JYKUZ49N1GD1FicLBgz6N/hLKmMBIKf6vSI/4Ef945+2yv50cyRcxHcvZG80Bxq
1kyme2MgC/PH00tUg3etGns+SIyqJ6OKu3ltpM1a6cZLB71IEN/vqjoWUtXkXsRV
V1iaTmspI0YJlgV9wn8lKtSCZCe6AlTd7qwqX5DJNBBkZs82vzhRzCzJH+xIJ4YM
UT0XZpX030l+2I36+6XBhPWCmS+pIbSI2qUQ1sOQNypAK5EOQuX6rqkzGg1Ff33y
pIbZKoowpYN9u7l/MUkOQeAx4DZc+HGTyxxE3ZsjALlMdBObpNmrVHBKVCLlx+9L
NKMOJANkhMgZ5W8BPNhmExZqBUC5HQaYzgG4SuBcxM2Tfd0HLErSU3dxrGL1GCg0
15H6EUWCRzhP5nmyNSEmpySTKG5spW+EOJZphwNV+iq2v+v5owmZUHpmIHybwme9
5GFgEpSmJzBEumXIwYI3tStDLAX8nVmqok5ut3sk4SdIrTIlwpBuW01MF7ktjTFE
sBpkyexydJwUAxSXttmAE5OnEuA094ugGnNfwMvAtae34yuovjry+qcRLleCe+Ir
qeGdqb7oAGah5wiOp5JwJ5vAFINs0JQSrskMxTkG1SnB2usgT3qCMmlPmcpp2zGp
Y/ZNiO0Usil4VZke+o0ojMQhtOa2DK9EhNdXiQAytcEorIDyzhs8X/memGy6HfPy
SlcHMTE+pqwZNDZ5s7M5DS+t67jMzfkLWaMFlkE6scsesEt0V+b0tLqwthoPSbyb
OFxGWEFRY+WwBi1uLyH+q3tB2EkgtRVyTLyluxznhBuKM7e2+Z7Co2vF2ui47ULG
ZRXhDv/ljzjG/BhMY9AN2skhpSNtwxg2/jh862wDcVYveC9sP96qBK8Hb0swhJw6
mEDtVExUstfWqWvVOIg/esTlIrE/LcNr79cTc+YkhIis3yzfryt36jv02dIq5p8O
buhmR9Urp0F8iWm/A5GS6VriBa95wWWnALTp7ltOV8ciBAjh9mP87pRCLihLqo9u
9Br13Nkue2ERvcDIYIFGcBBpYvBwy0w26umFqBn3iljLmCAr1awujVun/SZt4oR/
brayqQex+lZn5/2/g93XyIhUpVlPQko0PmvSAgGLZry5+lj6CDR2qPEED/9hw5mc
bbS4OZvJ/Ym+zlYV660tBd8rA4xgtGxh8d0dtqOpB77ekGYpegILXTr6v3VfOSzz
RghvnITpWz7BDz5MatvZvd8pLAxQdDc+pu8G7Bj1rwGT90FSChIRxjYWny1R1o3n
FPpNyWQDfgFGJpkuJAHkjC1nzNRKPzfJhgzmgIenVC6yyuQ6lkdFWyBvxfHDgWz2
39QmcL7iNLRgz6UquZfwbc2ZRXxcK1NLEXtr79aegzNKxldDq+tZSrJ4eIID8RF8
h2udm3TUz0sK73aPOhZjH9MTzcMt7l9MbK6qeEaLkKc5W2BB5khENpM0xfSvAfqs
unQU1yD3AF63meFDX6MFlf01iNiF77IKFpMtTSwy95NgUyzDigL1ecCQZ8+FxkUJ
JFcU7SjgqjKz3l8NlZ+z0QCkouAMUAPuz88/kiR6G6lr1BIoRiEs4yM/uGMXzBdL
HbKj9OnDrUJJtsCCyg9sXy19Tq9jDMO1Mx7mcWW0IKgvN4nJ503UI1VTsgC3rjAC
615PW0S2QgbS98DyPq8tLTbqfMXOgB2bKWUHBphBoL1vWLgmQAKmBtoTgOegObnV
hSYTVaus6tkTgidrfa7v6txQhG2O0frpkZexiaunlaliWp/MlyWdnfOnrjOWNFBl
jiPRqmZCaA2CvweHOjS1EXtBeiq9irmLmflifwvITeyJkbraOUJ/nZxX+sQpEiS/
TH2LE6k8J/nR1h0GvTL678HB+YKU18omsa8O67oVrgGd63mm9TgrxhU389tHlVuS
p/Tqa+FIRTW9nXzWm48wJ7TKn8p7m+NAbcpfARSd3J9eREH+KhQxCO20hjVPuh7H
RninBwsPOlqkLQFez1M6dhNKm4JBpAGjN1DSTxVg2O4c3RjtwLolhSAaDTRNCeHl
4+Qun2m6vKMDKgLGmy8RWjn6d3t7aPCDvb9hthC3TbyuZ9fYdeztEUiJW/IgX7YV
HGl2lYKuNb5SiqHITZLE1Sorjsem0PrbwVXe1jIyF2oyB9Rbs44IjgS7Kq90A1vU
D1qDBph69UpwwOGLjuxlhuMTxN0bXSC88kA4euhlQMJbeI+zT7XEtHIDX2G8byfG
FEDON0V53+dT5wVHu3DZCeOusU6Uo1Z5Bhd/rkEi0kAuX7Ri6/1m7XSh7HL/HRfE
sInnOSSAASibg6RHbhLpizdRGk8jz/hegIeadWRzWr7gWgbR40bnXCF+cPIf3f4b
agFv2LzbPHNNC+lj+xjkqDoxY5HVlGZgqmyqV6PD0C5p/4sCRldB5wzWhQ1AcjeK
9zyh7eTgB2nFIku5MjyF4g3KbX4oMnsYm3PcFHr+8jjNVreVF3SYlplk+aZXjZfO
DyGv1SnPNOmzhHPXTeL+um+PSvJ6NB1vN6PDa9i8vR89AcOSEVDmTuDozPA6Uhhv
tcqla20WchBwR9UQlMgZEJpud8IOZKcRzU4+ndkXlJ/6yxlgRrI43JjS9fD7sWJN
vODNHB65pBL3Zbx2QBEUnSUuLWgFWacUlr2NYznxqTvUczzAVsQtkCilUZ0/QkVG
UTTspUzz8XRv/H5iimsHu/m1z4P1eCoWQvSBSuydSPRyrrPEU/bR145v5zvOmBJb
SmJzYRxLEgrY2s2XPhTCMzvY6yBh+toYWdQPeL2Rob2OoWacJ+/m/VkokMlSvYSS
SwDpSdisxN4TCNqNWW08sTGG0DQSh6eI4W0EwR9w4HdTu13KmPNDnHNJi0KseOhd
PlrGx03Tcm6Psuok/E3zk3i6EEz0pkeeb0UU8ddIKW1yX6YUijYC1wqOqnO4em1n
+mmaqe5Aq4+5DRs0dKoHNjOnbF2aCGvKLv+LbMLyxRqLauvqSS7SsfzxlQa2UrXV
jM0Bsgn15LnuaZcyQiw84eUpyDl7E3S3IFFO/o/zu8xT+iwtph7skfGk149a7X9b
TmwNEH6TpV7Nhr1rbsr/hRMRPky7uGqY/hTCsw8/EurSZmoJVrYPmmPjuQDMDpWz
ArpDn8orL36XpUrmPlPjGzvQapjlvhGfX3YeP4hxB7nmyBoIKU7ddRwlX8kWEfqw
oy2TdiFy354/uNv2FqC3ON3p8zCnJNJfV8UsqDVMdce6ClclGNK4DFsFQEKvaEmK
eQyiC6pUh3FFIj03hQBluO3uEM+t1zCNsv+1C3xCO8Oqg7px7Lw1MDU1yAs5qWiB
POqnJBm82Rmh3ABo3SZdIABd+tUEFkxXJUvU2/Szy2Wiahq6ilumVm5IzL0kgKyb
TJ95+/OLSIrj4pmq4mAkt7TVn8ACQFbj/PQm2uAC7jtyXBqY5FirYLRqZHGVQTjs
Wu2V20Hgyqhnmy6RuAXBlZLg194Pk5plVdU5P/oMCkzfMKWCtyMd8LxqYVlYfJ8G
YHCsfRn+RSVBy6/cPlU9UPebAOopQmyCsQoUjP4dH0D0ZYn+2nHFObdotD9ZXiDL
/IWli+w39mc3QIAFJjrcskFVBEKkzzizMsH10eWtFpPVAYZAbB7tEXLrIpH9pAK8
qe4PC0ZX6vCKiTNRXw5bPTLYMQeofIOrz1B0PyEa1RV/e8gupZhC5dKWWfuIJuHm
stEbgCrx+aIBIrscWT6w1I2tllL8v7Xj4ljOuObPPEsdt7hiyZV9V33z2oYsuMxI
3iYRAuEKWUfWiLylnouUyOwkfFiArSG5NRaeBWmrgAN3/qRpiQOyW9O2h5NB3HEm
7SnXCPvTPX5Hanskh+GNM1tKuR9S24BG7foPL748V+/H+pbSQo72IvpE8iQE1aCl
VzVEpPjAkQtjvUfan7uFDJi2A8oiR7vrCFtfQDf8m+aGILk3I14KlUsoDWaufKtj
hZd4vzoSfCk87+GYtdH5k/XV4SrEUFmbqDP9jqwo7dUbvMJ9ejZuNRSsYwXxfm4E
zHcjwnkQCxOnvMAD+ck9jStYYCS2tXRNYgqG+cFoIaujzgb3LSmh+obIzwHL096q
XR1vyYs5xbetxdV25rGK6mR4mO1wWiTXzOfvxYPbBq7iL8yw8MKaa3V3FuaKs568
yH15jGh4VlnWXMuwIWDwvdYlYbH7pGQFQ182Uodsu35ykRDRx8EsiRMyZA4mZyhG
yaEIrFo24wuo4XxEscercoFLZCMlBNisKvskXTfW3CuoHxFsxxuWbyF2OAKwppOO
NtiSrtN/P6n3JXvR6Foa+ktbTIwc4eabg1BLwibmxYNDsDAgVFYL/2idraiOKits
OkwrlDIQJjkIiaAOAPPTlcU0qP7KfbAiwqz6z56rjYaKx3GZjqAYyhZC1+J9h7Ff
TwCbAFRVy/KbTzFg0ILHOSi+FY+8HYe8TYmOdTvmUNyPJLxsMZr4ITeZbZHdTVRZ
u+Jx9R4w01la8PzoHH+DOtEBlrsM9MTjyeYcClnvCjhlILrTeGWcud9SR7q9/cmm
4TXB52/2lHwqF3ZOIg5LkhCmUarfLII5UT+c14i8G/RmUe7S+N+oc0Yaxiq31K5x
G2YPtJZs+PxKT2le9cUgh+0ulopjzBUnzf1/CGb8CV99aCD69jfMiyWey85/ZECz
l/Q3g9+TFL93e9sGxvB4Gv4K3hXEqaOa1Gi2x8EhPHQSyX+oDCb2eUQbnNqbVKY/
TwiNIMeRWufbrxuXhBOplBf3FuipKrgFFo3tyOU04zLzlAJlkCQ4WwOarMWO/DRD
BEfrtkvfeM3g+OLI8tCk5mX8FSgkEN62fvh4iGvBI0TL5PxBkfk2svZw4L1lDica
ydBsGUc/klr09Qh8eX7A9KzSnt40+JpHi3xYFCxgsqKV0pFvsHoQ8kJmdzm7VADm
Sj/FF/ojfV2aurh97iKIQMVia211REiJZj4ZAoX79UXxotKDy38NT2/VJaF77kQI
NK0I+vcmF3rMbZpj+bhneuzn3IMT6tcDcTBIaqYE8pqtpEkBwFIoo/fCxnNP0vHQ
0moq8pb6Mo7gbG9Wtg9OjnQNPdtf6ir+7PSgK8C8vzw/bs3KJ9GzFs0hPLYE9+US
UEvT8lgTgZlc5n3/7uHeect5X23V6mT+dqngqAAv7yPy+UmF7K++ShS3ichD7PAO
8ZZzVtmfO2+VbvtRCoqxYKdkvdsJa2nPgemPxjMnRs0+Fw5p1aiudQB4ToI6B1vM
yckms+ylhyV5NwWl15qnof9+alxt8FhUIvLMZQcTfNS9M/tPmbeVmzUegrqM8KRY
mWoOyf4i5mk/xHCE5NhresT9BhzwGy634K79cqRnpejAxBU6TWwlhfuBG7mtygSO
4PLZyGQbFfIrCvKgObbgg+GZ1Bocayzsq3kPFR3E5/f1W1UkEHV7qvIzk48zynBU
UxMSyO/O3mO8rzwpP5X5xoMU1mtvJpyi4Q9/CUm0TrZdTrPNPEVkCYUoVhX45avT
t2mUKjBBtRhQKSUPMmn1kQWF1ETAHutEatMAa5cfL/jLuxGPMszuk0Km4dHedgID
IuvLsCOayn7I8hvYgqis9RroX45tJaAxSlDmku4OrAwu4xsaNMVVrRzrB35Ghtge
F0Xf8KaOzCDN7tZotR9sQc/Z1PkG89+YK34GZ3rLGt1HkKE7iTSMY77D+c+7eKn3
O/UdRDlklU7wJVUqaqNaa3W2tI7nOu2oR47tZl8MEz0N9rE21E07q2t5nuAZbUp/
MkJ2F8dzeLozBzCrlNriY7fPRFXNdVyDgmUM6EO+Uj7yvSCliB1RlFf1ODIbb7Rc
HB6psxMxEVo7avRMNW5HOK2g80ufaW4Ezpk03vrkuZkGsagijwBqWpkLbBJyaQMk
+aVqvY/q0wqZT+ecwOHHF1iVzvjFjaQI8pERsCsYSxOmLyZf+XhFpMn9wuJ3bnjk
uQJsZCdjAkgQLEsD5TFdbAtSeUa3kMIV6YSKdf7pXNBWKmeA8sjWPvG8vpmUGDuE
JOnfQHM0csnV73tONU5O+LRGDJiYCgnH9SpElB2JkccIZEasROKtsnEBpAwyPPSZ
sZ5k2EsZRwiLLMdgB2Jm6NLU9rZcxKIpZCY8IG6V91baV3vn0Petzh46z4rkXwHW
JBfjkNqMhyeOHgNLWHaceJLVzSF7BPBUI/jHXtXxHuy7Y4+RjaR+H9k/kx7//sdo
FW4BGF2yu+canEcIpLttrhilpR5xEM2p5pg2wJkFv1q0HlGl0RzDzfZfizTEY2Ti
72zOG458J3Le15rxKAXQp/m9tUw7yVXU2JPOx94Sz3DM31HrQWjd5OjkmX4z2EdX
uT/q7SGM0ME2nE5nJ8H9Wijscph2AR+zVnnGJMN+qY/NjTSzAw0DprUI91ART8Iv
2WyC28ofl64x1x2XiucwRXgfNnyASQQ9CUyKpImr+D9ZB+LOCUS1BYkDltPQH0ro
RSTSr385dn5lD0dEJGH0z5A8k1EQUz316+anGj354j7mQbbyTP0lfKvTtrOgPlz/
KI0eSIw9eVapdlKH87dFp/6D+s03NlD4UUzgxmR6uC0lF1BpUV5gX045RIyclJMZ
GCbcJw/En9QtV0MwwJ2rKzEan51qkyuW4N6md/250QhTxxj/Fi7WBHCTzinzrSao
oLqOTGuQFbX3eLmFNzQahvAAQ+6Ptr9/gyda37+RlGGdRI1Cr2/Rsjpo6STXKaoA
htmS1B+Jqo9lzWCY+Fqjwzo0QdnL4DeF0z9CqVyIhLsz0/XdjKi+1fpa/AdYKPHX
C0bvjMLbAyyRMQPCpTubapcT5i+QhpI+NhuhUHAYnC0LOUoxZZXJpdWdGPdUg41N
2rzKWDxG8wZykV88ywwlI0MNuCzKQQiS9bb1olzW37+q82wXm3HgVDppdyki20Zb
8arZP3fbcxh0d4yVMGUIZMuvg1k9n76UWkrRfwJCKp31qmnSQ6vs8Tjq6oomp8H/
ntnhtySLGsqPMQLaucmTqKXwOVx88WSWLFkyRwq2V+zhY/S8R2NxWlg7uGCFvRDL
uHDQePjNQrBsC7BbgR5k6gULxYczU4RpcoN7urf4fZddbW36nBKbr6meK4UwkW7S
2WYbgc/AsBuNOjFJUD6iljkpoQSJF6C8l256a+1+eiyzpiNP4Yb6L3ejISdM3xos
UqWbUqh2ECshYay4un3Atm1TAaAuwBoLvqaC2ejdu12ptoD9pd5D2gHZvstsT58b
EiSBqvmfZxvCGli8VOFEdpQdZmgpROQUcjXVJFXDYZ1J2qVYJfhDeekeGQAtl45u
1pb2RNnNn6ITgRufb49aypfU45TJxByRT/bL2sqevPW3zpDEXdzbJ45HBzpASErF
jwvWsKsvDOcivmwnMxRtBzXa4RW/rpoERyczsAHkpR9nIO5ppLPFNLYwPpY+PaPD
idGd/zQHFJicATFNRPHJy7MSKTRUl+PnHtjrGFVRObA30wIIfvfdQOfS8ux3NBGc
6fp+HDHE2W5tn421DBefPKQmOY8nwH5EPBfIz+oF2gq297xZLSqQuPpDJuo1V2+U
EvrQg4+2nianjl2uwYzLixzJADigbkgCKIqWlCEFCTLsnjy6d1XHHjMK/pIJDYr+
YzwXQRy1qawxsBFCQaqZBgNAGiPivn4m4VcEad6fqdOAWMhn8BH5kG76p7cFTg69
P3c7rlQ7+liSSexyie7GVsIwcBxZX6AS6XvJxYlvOyJ7+Nm14SRjDUpx7uXU3uRE
7Bjh1qS7wQhs+uHpJ3AmyYUUfItCHJtSAMa5PG3dKNDYakQvLQcv9mDA2MMrwmJi
3HO1t8RfBbT5HeEjmiSJQls+txB0IvdesFXrqZltAnvQidR48dDXwoh2TNTHZ69e
WQ1XJ6X2Na3XdhscHiBslzAkc12hrJMT6gVxgK4iWiWPobIzmRrZcVoDC2x8syw9
DqT0e7WRvqn1V5IRNS+QlptagGFCYOlyYbclRDtK9t406BbC1BY15icMRwSrFSGn
zA2lhhkVkBU90XpOkhWTbV4/3/gW2GYRLMCoJU6cC26taK4BPqkUC6I5FeqCdikb
HJ+y0vYNJZirhROKJSAK6N74KcK0cW0fBzsvZ7RsYj65bKF2jOkav53oCKHSXfh9
Hmyn7OEs2fjaAyROeVK4uf7eADSouymtSZBG798OG/BXc2HorlxOL62Z51CZtvJ7
1dPvOHCJPyK+2LveSELgNhVNktvoP6SmrYCRjjXPWZx2pg+PVUa6rUHOrz3YBv4s
S0HAbmivzhejO7IwvjVaNyaWqt1QwaI6lF5xGYrgQWe8oV04VDyxhYhWBY8Cs55E
RFGVUG8mn/hiSNW3QXyyJQUxH4jy7UHV2ebUImg4APZE9tB25oVehEOasVTW4s8B
TktsLNDxp2SQwhIbSpcr9nVfGlIlDLyZ7e8t9gThcn9Pnz0cukvailUsroDgeqBd
+u21MA11FC6YkNFIWyjeP/1xLs6UaaN7fd1bYa3nAeAUTzXt4PUS9U1hGUoQl0Ab
SKgk66ZEYzSIPoV3mBk9mxvDxTW13JE6XjcCRIQhSiMBsJqrnniF1la/FeNzAMda
u3K2rtgNDVPt4+u1MkHXP3c4bJkHdl1zHK9nnf21ik7gwFwCMwEyu5yw565Y7eLw
jfIZGy5HXMYh809dJtwcMNIGdr5oLw8mzfJCWhVQr69iFM92v9LtxS+qNikIwLEi
ve+NVm6le7xFP9CDTDStVyVUtKRyUdJ/E6PPIlWG7Foj96kxyy0tEzrWj61X89yL
qg9ScDQkPlhTh1uT5lIWiEFuBzrJLK6FLHR4g2Itf8HK35Wnc+ATXqaHMHCAbyTF
MfpcI57VIXA9fyPyCkGZQkz0Rbgrp0G/M0QCrT2mf0UoaMVCqRM1O6+5losmjuVc
dVcZBcx7lFtM6ab590UVImOGIsCGVcf4qCUQsS3kss1wiiYWkDdZOnoH+2nKVRVQ
Xezn3QQPzDEP8M6J41Qq0FV5uoGIw7TGNzPCDQRgUVKH+WNtvHyy5upNvPN42OBl
KvN2nxesv+f4VldOKuW9g4P1mWreMNyPKOitCWnfxo2xDTM51O/6cCiUlkuoR80j
9qmIKP1q5jxWc+R3jj4KEAOZEI42VQG3KHM/UNAJdATjTP6jfL3unJbxuBwyjx1I
eZ1/8otglgxMed4dPGP3JCrTCMB50dSVAsf2SXkE5NCBF9A4CTwc0TlVLXXuzixf
luaJw+5QiBHcpjGgtoqF1BiTnjfF5ZcX96PiipDcU6VIh6SkwN21FAInntCSK2g8
nqBwEnUjU/xO2yYPCvWQbVQ2FBO8zDKZU8LVdFY3s+goqNnvUhEiWtEvV4xG9SZn
lcL0tiLr7SuHykApzWhk1v8xALGFu2zBpOJjTIEIz84CvEbldQ3/DsCgVdkjq/b4
EjSPTiRFV+h/nUqKVxsFTCRLUcA3RvHFCADRMFRGnrMScgr+waP0WDmKb+KC0UWo
PAuPYJRAIcitzFehK3kS7L/d0QTsHGk4GhH3OC7Pvvdag9vjLCrlOTZbmu3O1aL+
2UpIiy6pKVrCLxdSxbp1CWIBjmYuufw3rF8hkWAafhkHdDb4zVvkTrZbOZ9YXDLu
+f+6Ka++b4vyYRxJghJ+mwFEcELBxdXireBxRPHFAv/mwY9qo/Bnb4rxT9Q06UL9
He18+CCLavDd8fFAPngrXPeJhKxqxaF6+100w5rODC89ojams4TBQp45zS8mVb19
oURVs2oFGsY0j++v6Gd+b1rspJL/pR/vdiE0OAyzcCK71pk2HxEN/SZL+DWbLI5v
EWrXicW+JO42c7lUc61p45BULJ07KzNTDSCGjwCMmrya9V3TRVxlAjKXpaoh2Kuq
x0eObs/YuFJAXOPge8kpPMzo2LuSFP4D8iNdnpQJvMSZHUXrnnXmp5OUNkgafzYo
4dlS2UkRU5xLkuVA6qnZztEUl1tqhSCGxWYm763bE0mw8Wzvrq2cqi7XmhECrLD5
CHR7opMJFwDB6A0jUdxa6Doexz6tfxZzHLxd4kovnr0/64b24YqXd2jabDyS4cPc
HzvrGzIQIKGYMhIOdeMH5W7rn9TyUJXJRlPE8IbJ+GGH86swJNMkDke76TM/+aOo
5pZ5FEt31uM8T5u1rGyTkLeST2EfnLoxgZX0WbCect8MMbd3DsWT+DPBixaXvKnR
IP182iF8NOwZNrpCLhO026EGdb+dm1yYYPAjRiXcqv05QjKiPJACD/ntyI0JXgYU
ax5JBytAbg18IT0P7KL56WOeHP6/vIoTQeImf1nXDQvmVFGqxsIEFj01WLEHzYV3
Om4Sp7zBMrkn8WjQxIA0FgWwioNKFTUCAoWuJC/8ypTx+oBtAYt4xLfIWwhKBKvx
K5UcCxsrY31mAzs8jHFWzvo0R7FinbGnJ8why7CNCwDneLJxZF21URBkTwv3vMY4
8z5g1j3BkpOiFFAKcqJAVdsQOCgqLWN/TVVvs6L/6MuCbQDvB9Qdx0D9p05sNPNn
N8Z4TrcvhCe4Si/HvHKtHr2VqlC5E5EL97GaEly9RTX53VQogE50zQHuS9+R8JPD
2kUsxJlmSCkYA/7rMxFHrRK0bHkpNKr/Ux8lssiKCeQSrn3QfGXaESii0zqzM8Yp
Mn46+z1tmKiQeJwzvzXqhpaxJuCnJdLsOBtMSiL0IE7SCrxWKD2uIv0btItOL1Ke
51Aa5gcKDUH2olOuijr05rHH/QgS9bOCr/FgI5OL6SzNn3EdKIlcpRB9J0k6ydmh
z8y34Uw1AWPcdc+lBRkQqd5lyz9HQFrMKxt4ovPHw9uJZ3k4PfE7sNwB1IV5Ue2W
05qRx07Hk/GOD+HMx2Djd9oP0agvTIoLel3xQC9gIWOYdBsGgr7gtjXayUu1grZY
0SsmUk9WMnb5zcuPIDLUzI1oXaW1iZLf9rXLloTzboFem8jimPGV77SNCN7uc+0n
14oIdhzNcv1lvWfjhIDqrpdOeS4d5J7fvBnyOCIQVg8O3tTbH3ztQdrfgAyMHr2w
JZckfT/N9OcAojiT4W5mOpkiWx6juq3N52TnKrBL5WGM6IxCGndkx//ynBofkU+t
sLB0bL+xj22/6bdPRs9h1UTwrHKUPt8PU6vXnukmu1uhuoFG16lYnPsP8W8FLBQk
1A4GNixvVHOgUK8TnKuMCUF9mHzIQA+yG5TUnnyxXjMVm5Yysl9JAZ2vdxDlbCrb
tMawNcn4qWb2A3KFRldKB//afndTlilzKBcUrJI7cmpCsBoD3wwHzR6QvkOTOrMH
z+qYKo8dymnuH+bs0Upal0GbARCzNCtIGKJhshq9Jkm8SAF06Oz4OP0ZG8xN0Q5l
0ntq6GeqCZ5+SgZALgv9KV1Capb3QT9YYqUKDBxvvIReHC+hBTYN+XBILaqciQ+k
tiTc6PvJMGFHH9fEWNcBWTvL+GukrIvDijXY0sLSqKWSO+kLfLozswUoJegBrZ8G
e1DDD3Xt2HhJ1HsvWYIR5lhO2JejS1msO5PXeUkvfaQ0+gShGRvkz9gLJ6z3iZIJ
PaTsJS3nyOlSXeoD0JIXvvLSDY5jSnwzkA2jKlfSAbHsu5y7yfuaUEvBQ3ER1cYH
/W/+e0SunwSvG3RZyEfF9Aqv0TiFvF6bPWytKptauQk8RLyBYYXZoT1kEECFHOAO
5UCCltQECLfG8K9xDGtncOr3Y4xC6tESsQg1Tno/Jz3BqDBvHCAIrGZy5mUhNPQO
yN8utOJmUckuBOLAp9RjCenAGh9H0bAnUxatIU82mdx6oaBeTJ2ij1RrYKmg1W7Q
+i59wph0ChTjt62881lnr6TFWpzblD0TZhj78FbRqBY=
`pragma protect end_protected
