// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mFc9B2TD1ri1+4ne+ii97OEFVgfCnAogWYEDevG9YStgr52lIB2Bz3PekPmDE/au
2jqtyTSAHzk9/MKj0iM0gtZSyo6QF2bNyEYD/iCPR5fvyGqwW4kuE5whcCu551Tm
Nzz1QEX0nIJaLkaN0XPplMNZKpGKqm8yhIDU9zI0QPo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13568)
FcITImiHFjCa/+OKE8XaZlUteC/gerNAUb7t0h1fvb3mJlDVn+wB7LZ2CNRQ8RtP
tcin6ptbWLZFJ+/Wb0EMxxtkxD79Y/rsHnf+Xgf/PboBJYP9w5h6892AGd0L1LRM
UN55llip15ZNrRMlOopEVi0xWv+CxCovP2rOLheQuSCxHvxQrriLyOaKzQ7di3bG
MM/9rGq4+gDaAHXg98vFZ+mSwpjQsW5OXXc57/qWqSwvP4fTLMJkPR0jLoPLJwHE
sSN4EOfou30MRu3D1yzbBAmWT+BRNgvV4ISZrLUJR9gp99+dgJzlgwrHs5z2v0LT
yVqz5bQzzHhO1ccBqM/V1e3H2mDrM/gB9QqbRFsODxHLpDQltA2PImVZyKGtDyti
X3BLE1nX/JsH3LkaPqrYYh/asJjHFIOTijMxvlzEETxZJabKITGEIJJhWRqIfSKP
PfeKVvPYWo9zD1FD0MjHJGG5mWatap6FRnxKnHHxZcSdQyKxhmypM0AH9Ep+1zkw
5AYNATcOmDfvDql2fswn9lYCOT8YXYiJvXNmlpzG6lp28/ESh6IT6Z3jurWmyjZD
7B+LQQ1D9KUgdG2vBqG2V7F8hHQgkNXfeMUqP9Ry0YUB25In0fkvb+0lve/GO20M
/X8eSDALsn/PpssN5WBVOJXzSbYioCR7XZuYPeECuymqWJDMSVPRh4exWLtDI8Of
BykBTKl8K/AwxNM/D2KyyfEOXr7iyC5CiX5ZkLO8Hv3VkSCTcAvuhxePHMvWf5Ij
0RRncK4A4xY3v+C+M9Yi3r/g06X4jy3+1Rl7daaf42t0vQQ47EY2iIGvTeHD+tHi
C8zkiBDRkyD/zgflHtz8uh28672a+ICG/lBT6PUgaTEQXbpSWrWCVV89bbdTg4sk
KINHvaoAmfhEI1Hro5yjKyPth56JyH2FUSHuWcFvKfXJvMy4yefkms9+nmJc45OP
dVV3RhzNBVS1RMurnfmeIi3JWcI9ErDpd8EV65yRY58O7crGmsQySAD1IGZ+qeln
rDdxpANzJZ50bnKyLvLfHYP8+wvOK+DDS0KdPG0g/u4NuL9B5NWhdylDH+qV/CVJ
Dn2jRSAund9gtjWGpGLgXoxYAOHMp6nKVve8E4WjmiVNuuuR2XFGj6JmLkXuZqzL
xHxIQZnOsEkGAdjRFYsJhoQPuWvvwQ9SWGLSrG7kqsQraSwmD4p/cHeEDY/w2/XV
As33YAr8VoQzaA1iDIAiB9WxanRWrKs3OWxFZRhespRcvzoYEbnsM0mp67MZBM/z
+1TzjHYsXU27gpusRI2Sf93gODQd34G/4AKIS7v4EuHzXMA5YQhwP2jMTqAhjYJR
Yh6a/1shUEnR/BqVr8feK54eE6lyaH7Ps3Hq44mvc+63Q2UG9ClWdy68c3yM1mh0
I/tVn+mq3A+ShJ2mk4zGazHvqJOxC7zmS106GH+Auf9xx3RS6sCnY6GtnGlWxStS
KxjZjHFkHU0RLItw/IEWJ21bSi2/NzZ3VsPZbuRjzK9F/u7+lKOSBSo8ArnGJWJz
AMvuMtPyhRiMKF2XaqU7J/2WexD5/c3/0HKvk9n3xYedkj5W1vvk5oU55jYzJYg6
j4J0mkeSK0DmP7oeWB1ClWwPGAnB2aMgHZN/xp3DDZk3ZjHXE0J7n696FayfDtGY
Nt8oc8CD7za6VYHZa9gQOLWAEkbC1g0yFHkdwl1wt/EDgJnvU/FoWKz2cGwVmiRn
Hd6J1J0332366QQ/DOFbv3U6bPWwpBCb7IHKvYKP5/JSs0aP9GsD07VaWjXGlGtG
WrxL0c71tHBkuIe7mrC7dJKx6hjknUWEh+EJFVhGZcXXd/QmFYbzlRyhkWn8YdhP
R6AUEuJ9UOzeoZDeAWJ3K/Zt6Y/sd34GeLEy2QlH9l3H4wxlpTVKuZuosQ+qkjUN
k4U9i4qIq+RSFbhQchO/ubvNUyxvLBIDb8O5Z4Z9iSOHjVWPfEjtYdj4IXJhOOjb
pFD2m4g5wGuer+Ady1+WbwsIFBT/NWhFUPtCdaXdLhLT3TcqJqj4QD/1qtxB5ohl
vjG9dkDJlPn2lkPGYopdcXjYspp5U5Pp7QdJ39lEmEH96MYPKOGxLbSbKbbaNQek
2vAVkdiS0TBbeVBcES4SDTLlZsF6EXhzrMbqtNEaJ4LxCOATnMrwm3tJBYJApast
8adlcgkkomnUtEeZj0y/aelkDE+IwuAhFvoe3UUrmYs3OVxFMqdcz1zPit7HqUZV
8lKpXsCkehFAeW+bpi3YzD6Ym8AGyjp4oyvBGpdKdpXE/CrBKs9fkK3gT/QDMWMT
g/nyP4WJ66XpRC2oMIA/uHpZ0Gy6+UbV1pFdaRhJ5YzOBCYcgM7jPNm1vq/zB8yJ
bWrvvgkHZl8ZZj3/L9omtJLa4icckyt1Qzaj0+tL0do+Tm3rwHVEZQNKYSKpbKoc
sqf4vRhq6OMYKOFtkkioxmGhUQ59csPOc+q1fmiXL+3v0IWMyDwFCdmjfAE4vHnr
YEGoxvp0lnw1YELAUGpFXVo/0YibL4hP578gMcGi/22/AwLj6jm+yqoMGMEAtSCX
KFEBDuYGWknZcAM/mWGT42l+J1EHrIcFNnckL9IL5csm/5e5ZDT88jbVRkH9OXc3
pcK7zeTMzyefQ9k5PLgQAHFzDFP8lpG34K/rzjm3Nuz5g02ZaEF3fo7KFlqfIA7a
5zPEofUWUHgkowVS4MYRqiRAt2R+6aLCUR5uoUSLopSCwE+BVr/2dLAVnPquOP4T
LSw/2lQsDuadySIyjlwFzEntmoe+KU6MWC8eRvYA2ieDqeXLDoC8diOaqhl2a8cj
DPqsSfCo8j6DmtgU3w+YlZzzOhDPrL2BX0fsTaOBcQkeXxqcJ4a3k9I0vvJy/ZWN
mi3WfQc1Gqns4Rf8tCkk/Yh9lyWEYRxy44ML+GFp7thRqULQ814e6aEOJy4aMYrj
q6HY3Pe/rOpBE8/xeXsJXshd2UXppMZeJL1lMK8wbyB9+US7wF//pY2bXTVEhBAM
0+GyV50hCghS98KgmVQ8tJ2Gx8Yq5cVFr2LyaClZxB8x91AxScdFxpx2K9AcaTA1
GMIhvElpLh7EiWARBsSIMSVhbBi5okMrQ8/HmssSKUUSYFwRx878eBc6dSVeiwrH
pCs11he7YvRSnFRR5DNBYHk+hg8JCtg836nB/FtAj+M4lZrGhSL8WKKkSURNVTpV
MaWQxvvbGf8YFcbVvSIReVTH4WGT1jV8GOFal7c2oF+xn/oopPTb3L8hSzOSmb5D
xJchzaOQxAH5ikjRkPD4HUeRFUSbxlZKCyCkbA8Sp1I5xSg1URX4vO9L+H6mkAZd
PSWZ0l7p7U5dHI8Y/MU0zjpoWLZj+ofSZ3af2UHnqf4jKK09QmKCDG0c2Lcxkqhq
6Vgmd8UnggM1FTUTs/wB0CLB3BooBDVMaXKQWuYYbBu3aLDIqxIZYWQ/Q3ZvFcyk
pEZd5co+hOsRnImssHaBLYHPTEKKSoaG3lsaSRYVonnwAPyEdHkBtDNHOfV06FET
WdOK9WR6NyJ6eGOYeDFZNjmstWMn5i34orYSHUAAl//l734iUnmIsT8VVEXVfDZ/
NszTM/QR0sQyy/uhkAlP3FMThV+qWJfw+5ERaB7u7FMeADBepYoFx4hr/r56i9XI
rd8bn6eh7/RT7Kp1jY5YQe8c9d+uN3DEIjboh04O8qWLBE4+cn7qgLL4ThhVogyf
ocqtMJFrsVF58CfQyhcjFFUwpcRFwhAzEp+sgTDS8t8+9GaXQ79LWWAHVPYGjfqS
ary6qY1ETZrMH3AyRyw//7+hyht5KODr0SPd0aoVHdugoJNzV1TxsR8qdy28IORg
fAcHnZnrv0p3LSu5odt+oxNp8mVXdf/JVu5WPm5+Dk36EsqWsySE7bu9bquRFupu
Wwmwgx5ob22+OsKxGH2qm5wVEWD3DGKiD1ZEuhiHtFX5+mKAH6PQcq7EIOyB8RMY
MxK87wZLfSd7slJZanYSUtz/K4ILhdl5W3JVEV804H9CxFjkdkilti2UMmBQ8F2m
QgStA/DKkBBZmmIv8U2yL4YUAwVW2AitZuC8QZn+IxF2wvDt10guwKY8z9wprKI2
m/ln77ccXO3g/xoIYS0/Mf092JXOIq2vCV1lo6Ksua3iS+zT24G7JhLqazxCGceJ
EqsVX4Fi90oVWigMf5JNQ4CuCbGVHmSPEHdnDS4lcLQf0gzHgXOLAMwtEKkmfRQI
oCfzNHv4YUM1lYTYwFV3pmb74+DVN96NkJQAaxYcz5hA7Ur2+9TfUC1AssFA3LPN
MnS3vsBwKgZuu46HOOe9IvR3bQyQobqUoOiV3LgMUvKa9NxE25UTFHdS2IsPmK3j
IQaav1oCMBRH1IAAM2t0xcjTa0l289Ds26mgXI9FUd02Bo1xUk30W2H3o1kiJjAh
vMx15jIAc2DEzmBxuL6ABmAjarXVZ/m2h8hbOeO5zH9PNvY+Bn6RHtdIHRIRzaYH
B/rjRfRgdHsjmKpd296EpR6JYh08VKNQ8NQlMTZrL/pUS29DJl0jMt/WeBcuXKdV
BUrWavY2ecIDH1DRqzLCUE66UvV4CwS5mIBxRP8iR/Y5p0/3R7KvAushgloRi2Ox
cL4ZLwX7p1k9snXXOMI/yEj9ULkYZyzrPeP3LcrfJZE7QEcQax3ODrAGPRh01ruz
Lss5JZr43RL9FVHrZMdyr/JvxnnzLp/9ugxUVQB4DtLwy8liB+WLKdOE7AWbk83g
xW19jnx7kdytBDsUixX3sqqtVUqRNjmOAenHXn8zPJ6LwNW4/E609IRrklpGpHxD
l7GqllOfqp79qtVdkFr/dBrfDka9A8V+OnWAiiy6INXgUPTHin9LpzAQitkbCdSW
Bl/yQ7MnasruCBxKnJ3PWPmfuwDrWuCvyvpITcNut0CrWPsxyTneJ9eH6xth+KAs
ZzzhlfGhIypE8iOeVSIDhRJJz2xFvYs85vtHjV7O8HR2u8zgz+Y37uGT3PEvRiH2
Ux6jOiMS1VeODq/eCkDCCD535hIEvdUOISSIdTqe46017rLY+ezAMtnJQNkJ/b1o
6E2sxaofyuSf54Vi+mdL4nSkWexC45Kt0C275P7DNd+39+ixFJbZfn9iUmOLeS99
JbbFyeOsNCRETtTDgTRAoDDbeS2UrVZg42dvKaEsENMc2mNaSY0990UeciL3shWt
JN3ucKJJqtajtSDQIOh1oHOyt/Hdq4eioQa2PdDP9uYNfPt5PItG7Cq7eywThoK+
ibblitBpNLSBu+xhk/vt64Y8bFdDpAfYA3ogGi6SkHOqv2H8i05xqIs2eQZLJJzj
E4t4nlOy25teeAYsvXpbvBmYZEBatiyyJY5mwvAVK0c4yEtwH+t97E2c8fbHzjsm
CThIbwp+OnC0q0HtqDzlQ+BdrRSm5aG3i4lg9ROCxUBs68zUCojVxzrD/f+Ee0EQ
UKMgslynJhyWER33H8OOs3sSVS7WcjwyXUCHrEX4bqJO38+a3Di2V6puqsIOLye1
t50gy4hXrsWlEpAn/Vqx87abcCenXVnNFu6EoYhVMM6cCDgv6LFOEpHeDDp7HUpE
N3l/FrrLhwYS+qyZzz1g9tuILgF2qT2hNu3WjixOnoMGV3r3Vrvy5OzuZ6q2qrgC
M6zpKv0TRLFcSVPYfz71t5SY6tHZs7HYZdM7D2y4d4QKCVEztLgU3445RqMHGFIj
k586/vfCF53mlcIPwu/erukQFvYycR2bnr+z+ZQtNTppNC7jh701oAEyCxV3nAbr
2czG8nxa8jOFhNOa55op2/4hgpj6fv1st3jv/uq1f+V/xgIBdEM8QhWxh1fB5Pbw
mOqxFP1+anVRizQePU+nIIcb936gLPcR9Z3FSZsIfvDim2z1TFZdkGVLRArTwnxY
eDj+7gXjF6a+PPO2Ut/WUAAl+89Y5IF099DiRtNhI7Od15K0Ibr1q9g9UNy+cOLz
IWoKdt+8CXkzh3p8BhvjPu4Nl07Cpay+zmbMFYeOprzeofzYP8tXtBQmJpuPDQPF
DwhtDQcerzKuqlnNuLs0tC0NUuP/OkMAMRVoChTEUYdkw/M7U3/Huo7pauZHejx9
6Hfzx0xLnKe+pXixbol3ukSbzBLt9ivA+dxEorucTb2NanxzM9Bn+L2FFxSAg+oA
97UlrADxYHkWWGrYYaqVUFBNJQovH3lyxLA/uAm+kMqOUC1hKdQuHuEQG1rmJWbA
9F0+pQL8uK2QCCn9cVmMYwu2dGof7FGXRejK3o2y+OaCuugEFJLi3HD0b+Fth5Ue
IQ1yshDYC1vccoZKR995cEFfBa1vlupRjgjfb+veUAhnlTHaTy8s/cPT6h7HAp+k
BCm8bjkGU/ewhK262tHBNzmScgzEY6wgZ0mSulELL3RMh5ZkFtAXAY3coUgHTYah
5WEUPnYM0ugDoYZwedkdyPw03E/DhHIytAuZS0+ZyKlilPo3pcCIA/j2PYLts6/R
wmx7KB/CBiMDh3w/KZ9YXrEGS50Q0/nG2tY86UPtl9Dq+92U74z1njql+jlSq7eJ
DatVhua2q79cfmiIkPekZS8C+iQHCSmDUsKLd6+XPhjJ9gksWgotJ60/j2HlQD6Y
AQ5ESJP4x5QvaIHPf3lO33Ty0U8v2HrQiUk/757wESOUhCYDCgIldAVX1hCwL+2X
AHmTYIabqc59H/7748bZ889CaC9Ytvp7UJdItqzxPBNkQsCLXvduqnPO424LQQa1
nrRPQFqPi1B9DfenbdhpPdWmOWlGXN2x0Q+qSA0Fng1qY5aEIrjZE+kgz3KNuZAJ
05jhyRKd5QOAgc77aadQDPWvH1hx93msHM9Pz1SB+dK054P6X6+bqPOm6Q51fBw1
yu+yPrz2RMKxxa21f09zrHHsTe0Qmu/jfOue8hPeN44XHb3oCPnYiGFkI/w3OOf0
yevHnGnhRul9Y+Rh7+BSCmslgzNp5a3uZroumrrMRtPPNqzT0oQ+hHM/k5gocAFR
5I/nlgL806Igf29uWV+qJ2dldM5irvlsUgeA+MGK+ByjV3tIoffsQ8s56LScdHdF
ZsGqUKT3JiN8fu8EyOEkEaFaZU+ZfxGtceG4wkrOrPKkBiwZMgtue72uLZWa2bDh
9Tff5h+ZFZ1BsPBSdMSle9eNQLCAg/I/5jI5aYtYkje/IZwXFGw61EZWbgNDzUF8
wZjwj8ehJcIx52I0p0p1z2S99aS5JlBvQDtCV2iyIcx5HN6uUX6NENyUNnO03LNn
cKdS9Kr6G8ADhU1cESbhkUlCErtq96xfwrCO4rvdMSW4NyHJrA5/6YjiEgmw5eup
C7DHTZkdVc2Tdm2zMEd4a0TIJUsWj/Im69rIol4a3MHnN0pFE6TGl6IImAevUcsM
iNEHjWoFtSGfw43enUSXzNtbP/ten203IOMV3prBn/VNHonOFhx3JeS8XD9Xf1hs
WX/74wEjX5TugdhLjMxEvMoQ93Z2uTdq3oxH1PUmgPBjmmKQE/SC+OtTf4EwvWGR
9zj5oJ1XfFGmRU6TnSK1W9X2FMFaD3KZmaYdJdblGfjoF2/mcPFv0qxfTNwVME8L
5uvWxnKK3e256od43m2fbCHGlT6mB7ocSmERV9Q/61N1sAFrJr+aIuXCHhvGuy7P
Or1JJX/hVs3/5B1SfQ9q/jv5Rps+ubkafEVBU0zeLfw92LIfDlBvyYr9Nt1eaHf6
bYA2qzH+EStQfeW+p3RzDpmsqF5i4GO//jZksl3ABcnD2ndLwQRRL+2sNqjqUSVc
7bJhnRaVtr4e6NGSAPH8XDrPwZH/FuYniMICZypwBy1Mih2JJE4BQoJqBb+UkLGN
T1krMu4pvfenLJQR4gjOkl8l9ZhupltSF536awzYlhfDVFSODPu6aBY/v4KvSu5u
M6mYMvHirlfe9G5qvJqwawDKCpoYJFe7ZA9sv6IGehvvqxGn6sX5dh7oWjHD3AD5
BNP4cBXYsXkvgiRenwYPP3C83nHlVcU0OHm1iBmUzuDB7vG10KV44ZkYNvxhLsOV
QvfN8it+rH6B5iC18zfz5d6KbZWLzeQdF8kuQHgSKT2gofk3jJIaQprZEK7MKtux
wIWwN/LE3juntkqXdml0Ww/zjCSQSc959DAEG1FJ8op72mkjKP8gwo2DqczczdqJ
1H9UdiRS6IdprSecsZVZSQq1AxVPSk8BWUinTsUXC9kOkKWynd2RI2NDgkunrIz+
SikTdVJ47wmByfZB09lE7GmWY/3ICOGsLWw9wYJDbtGf90VVzmXunCUVurT5+WJA
H2oUFyOrxnczujc2cVSL+YHz/GqUee8ZAEvdds8Fl2wV4AtmDtVFDg3Ua0LBpE+T
D9MR6L6GsdY3a0Df3ZlYln3B8XENJqIkajOahqeCuaNxsFSsanrqV59Fr3U9G1xc
UdAp79c8+c7NqKjWncC2EkNZB+YWcysfauTvwPd3NwClD86POwqnmIwbOIkForVC
xVS8xljjr1sMcPcC9TQQdYlPFY9cuLUaC5MJt6uo3DRo1mwf8pX/LXMy7NqA06bC
hVeczs7MhkAbfD9PvFrOA8GHtviXNMKFQyWjyE9OFfciJTEWO2uoohHBSdI9HuQ3
e7zwU9AdZ2afVQGG1JrL9gg+xSD5GM4zWKpg7ZJ1fobpP5FYfTbC4C/O+nQzoeWG
oLHKNSDDRpjASOg1XIwfEHppUfV6WpFHle8X55xf9tRgYAmRsQsNClPjEtfE1CL0
xFcJ83LmTuIxSNYejm5TKFdNqv9a2tANDYW28BsmEcN7+B3QUlrHmyl0eW3U0GlP
ypvE596Hb1P1qY+J3lRFjV8LvRXUmeV/USIl9hiRZ5IorKZpkjSwzd3rlGmodzf1
RUps01uk45XFClt3Cp5LzaKYoE8rhd+lFfeLNkN5gHr1YJPxgP3mWFmtFFWTGSew
5mRubZsqpzQBqX+yAu89UyX56cNZJZcM8PVCU9NzOpBoe4C9ONdRWRX4VGvHuTcg
tuqcwu16GCwOtOKqxHKittZ1OBkhxbSaEZEZsN3SWhK6kRDCdOvdtlg4gUE1e9iw
fue+EqPE1OFzj8IVgig5PCkgg9vD691K4u1qVKss2cuQKi8A8ODSMLXgCfoEnxEW
S9JymVSj9okoSNqHyf0mJ+fOicYxna+yJXT1jvDItXYWzviloQheV5UoatWkdrPb
V2UMqeCKltu9Bzw282phyDTtZgti+mOG71tm9WReX20Ff9Xz/Smk50yun1+sko0e
e27spJXy7AsyPNxA6DozVcVitbrTYio5C3Oc3PbaMMiqOXa5CVcEM8DBFgjrcoTl
l5ERH/w1UCtXgZFnbt7cPVk5AuLIrAQfXEvtc0snP8BjwRwTDSUBech68hMCWkS/
SgDYiIxUCLY3FbO88N8Hm9/lsA3xtRu1LnEW8eHKNbtcdWuSlUslA15Pce9DDLlo
gLX/OSchfabG+NrUgWinYTGo7KcaY8VIaHExS5w1+DwHoqd/NIBMi2PD1i9eTsly
HY8lrnXFbfRLx6Xi7569vtDC/ydfElS9Gp1WqEH/wQJK4hzM9LterSU823V5Dqer
lREub8S4JfINUJ7itLuPGjca+th8+thzG0ZSDVQK8pqp/gd0gqA84kXgN9UNQA5N
ak2Ymn3liBLlHWi6AidmPm8ZbWq5ucaObF94AWU+03vE8XGmZ6BrVSyvyCzyTgoc
qj0xG4VGIeABD477I3qj/2QRP26ndKB4UbXzEOsEfTAzFz/ezhQmqq7Z6jnNCx8G
oXel+xSs6Rh7yuGXj+1BO9TLrkq29+QwtWZiv3RwXFIt/dKxEeQWE2YTV5Izkgzl
VEmkPjQMOCNm77QGJB0ibzdg6b4nFeEDz7QxlG2IlJlaWbcC/5vEVNsxieAvGYZX
1CnhAqk0AjHxv8MgbYxYHo3ZPR/sTqSn8E6UeRqh8wS8QaIUWd/3nrqsqfioUACu
34yqhqjJe8qZZw0Gf9fSC9A7LD5e3xet2iOW/uRLOaIxeAXxQZcr38/ZLfnjnI/H
uetqGvnyUYbG2ixrzB6Lk79ZpsNbp8F9EVxhyRzoNbs3PJOCbaeB/kD4ThDAlIzg
ZV7+u7uzgf7kunGMafR0Aqw4uN0vNr75SuJ/KB3QyWb2w3l8ncjly1dFAIji4Iul
pDO0HU9bbr8x1d2ChJellO1i7loV2QCcRbq+2iQfpaXgUyzRpTO1Zz6zTp6Kdpfs
ZhPaPg1i1z8YKGr3bNu/bLdXSk0Rx10ajP4ejiPicdHYU2+GqA01kG6uZBXVNEKH
1JzwFnchklSKPbIm55J90I+YbvWxTQVvxCEFMGCyeDDRRLFRhUFSzXw7bwShpSew
0YDO+5TW3CWr0R/njOWxY3COmY4vTMCSKK6p+ZNoHWsEO9I6zF93Aeu0Imlywjm7
xw38mdqfGPNg/ZN6b/jTnnoUStevBrjLt8Msur0ywTAHFmw1gpTPnU685V84fIK+
djeg60LZoTS7EzvJhhwIFcexSLZlQHlS6CeO+kBY0mYzqP4KtRSZV6aVlh+GwSlz
dfmgJDzo1EbidaTDnkx1l5EMr1lJDS/Wpmvzwoqt9BqJBZbMM4Jpwp2aLcArKrz7
HSPEz++4wIyoI6IHXVs2+1Lps7KIPAQaLei3Ao/tLzkgDrNX5U2wVAWKm2E8KKXS
3LXrU6V/EplCZYeRK5jw4J/w/FWjjjqdpels49xqByCHCKtfMxmexNysvhk4753p
bDk50bCx/7dca1AhZSgp2IUrM+GEsq83iQuk8SfckW2fyHA3i9+lXLttDAaRfXrV
kzeW6FOX/canJGDrAUU30UgxVMzdz0DNGyXCoMQL651g3RDIJcJbA9dPumKabJM8
ylsWyQHiJxW8rV1Eh6lxFk9ehRsHDOB7kFbv1gAnfR0aDsF/tLZJcRHA0mKJe0G8
NERAKF7nVG1KD6mX7nCCiE8dE2mNYutJwubYzopSuBElXW9RJOWG/bHqpvOL7qM8
yM5GMZRw4cLy7UMI5QgUtPrGDDJ4BiTk7OzOkg96JNL0/tXnVqtxCJqQkX2ZcEUR
Cq/JDuwCvhMh3J65ZPfwAJSKw73PZnz6NQ6p33/3FnsJ6a65izvfmcnAnY3CLkD8
FTFLD/6qbthLGT9i6fLVLwN6/4eZ98Xfwn0y+uFVcH0vkwXGKjhcOyULvToCi93I
US5YuZa5zzGgTLSY3F6mhmn3carXtE1VwsZ8ZY+MUfxC5pWqS8b/VuoFV7eSQr61
QtSg3F2l90VszajoDdTZTEKtWDIEBBUSDWjGwa1A3GyheOWnSFUEkOI67kv8Koib
dL3+0QYdGxwvwx2it2FehyK1/T//li85BclNwALgWVyXp7U05yQ0xAShNGc4LAFn
MiHx+EgOG/3q97w3voHjaOR3cV4otYhYVuynqlkQGWjxBwbriyxKc3RYTmLBhSmZ
xLKt9ly1O9A4uewb66cda2dY/nSLWnXavqrPeUfMUxTNI2igBT+ne+jdDxFFq99M
4EicU2ijEQdjHfOUV/kva/okYpahEu7nZX7GY0HkidXuA7EKJ7ME5UlvPzqL3zx8
UGhjJf84lUzSVf025gPSKJWG/TQ+XSbRPbmB7lSGDiRD4T2QgVjmtiCaHTiym2A8
Twm0OWaooYv8idGAuMKG7wYSdqMEf+UO+TbGvyxlUasoIyF+VyhPbzRwXPm7D1B9
L/+X+U6hY9ZZ6pU+T0zd0rzWxNaVX1TfSJ0qhQgpPsbMbZQbwKSGsYpziyyawyLQ
7+uzWF9TAAn/TEhF43VXocYe27uImdrOaNej7dQxZopkg2DweHRnuf6MupwrX2+A
3z64+tO5DAfvPzIC36rVXTp52L8gXp1l1/yoGfUIujuEbJGxIkHdCtpr1bCeeeCt
rqV9D3rwA5XKissfHPnk/sRq7qY+2sZ7ans25/nzdsyURYL3gL6nq2oWRKlDc7nt
MqFFdvys8qA+XwtDPrqqPLaQ5lUxb1uC3N72JBHOBrjoXNq+OcF2ugS41vTKg0Lp
r7GXT03Wlivce7d/zrb8OaM3PRD1MBCnNTkGjlMHJdf7Bh6GAJoaHAN0YbAO+ntF
6aK3R942dq3WroxhHynpMB0Iyao8a793R3NnM3pGXn1SIic6PhSudv6RKtR7vcu3
XPcpffjIyQJ1yyxO3UJr0EH2PSQ554R4PRjppAmIi//AhTLV/CitJb4S7Y7+OkUV
m6iLYa9d5GsXo+/5MrTPUVleuzMFchynnLSKZYz1359YyE6jgO/Qwm9rbyvVNiZ5
+e9DsxicPP+jnpK0aApFWMQ2ZgQmI44xGtqCC/QI5tlcfuO3+TXhclPrjS73XRZa
LXaZ76zsZGnQQJmSgbJep8GtvFZx/7vH2yX/AblhrjmqiZY871xCi0CEUZJLTsFL
HmpQNEAhdn30bdKq9HoSU7NTd1gvGdJgMFO7hRu5baDekPP6m25Zina4jqqgZVdG
CKHbvre3Am1uZAWgLwFibYCex7nvdhVQQAeCuU7E0YaJv4a1jMcUcOI0a9Kkzk7W
yrIXqg6X1RDv8Xde5CasCk6xu7VfwflflZvXNCUvew6CPIqX0OM7HE7mZUBuAhPU
xWZ+VM50APLOQeVzWH3Y3ijfjOELMSYl3tRB7KYZaN37XMbVhc8Z/xvoeEF1B04/
qwp19yLKrDYY/CuQa647q/S7zTtovZYrktnALPrClixbJRh4ogRox563WopWNr7N
oGeM75PffgLuhpY64GPvBdhJkTPOCE7Ug0a+xPF7sqO+OCPv8an47XTUP36KxsLt
6dKLGTS4BqQbmvGSpKPv8pYBEqpT8c+SxRcuxrfq3nVql0zEnUGz6YVMec/NS9pt
vuErMymMI5MXz7+7yCVxrX3eJidkNL6TdDaqar1tOhbRxl8Fj5BB+LyObE0hmuRP
u4IuMC7yJaBAY3GIvsrafXgvSFyajkonK4tLgONDe/mtkpxcVdnU70wd/wAEO5cX
Hjd99dX8sQ1sLBe6NxK3zc369rBdU7bh73W4zDpK5kUUsCMbC59qm2Eq0us9Ae7n
bM7LRuR4FHqink7w9Kv5yiYIWnez+sdoLc69SdOjWyQtD8ms/b4yo9Z8DYQ2vQNm
TwvscDGI3BsxCtsV/HoecA1x3gTUAdB5ieaDlK5Lrb/zExy6S7W9e9FnKGOYBgm1
KVFB0jTVjJNhtxOlANbgkEAn6E+COJVqu6NMDJzovuj4Fca1GK1oi4TXXCZYa2qk
AoGW95VqYtOBIj0lU4D3l6hynDpytqyAvU4oT83xOOLMZ+EyJ27tn6zgC3onHG+C
CcPZVfrNK0wkJ896GiDymOtfeJZM3hx++K6kR7CzlcHsPJIpPbuVO+qIao1lu4se
ZL10dBRF0k4bFcVgYHdzjGG3iUyzJR/Bn61qaYdvTf9+KRWsnJloXg73LpPFRsPW
gNYnF6NNgQo93nQVyzpmszVd/MSO20HccQfAYWw2Ufu2VwAPuR1oHeouFzsHtcZT
jxLDtE06gjyUO8Ndv2TxG5riDGVEE38WApJ6Sz3xGil0RXG27TiBPUMQC+cNjlHa
EXlOI5qLVMiSiAb75MqxClAYEFavliS3Mz05huKZLBWdHg4ZjltXyURORJNd1Y/S
XwfX12gp0r3rkUYM8calnxspA09xyTYEIvviYE/F/cuWyEf6Nf41V8AervQi9gdZ
dgq/JWCwz2xDgPaHbhBnlXMLr6Vipdt2NuhtWs9ZtHtaHkmmc5Wwbn9VxkHBjG3l
GTqIi6Asfe2v2i1/Vi04Ov6PLZsbbXGdIaFDjFg696YRgb6uY8sln5O5SINbWFAr
kpTAZZ7SG609kMhyJsSBBYApC4gfqTRi+mOpLspM+R74efsdPoaswM24pRbfkWbk
+Rw6hLrvRHcK9rU38LEbVLY4T3Q4d/wEaxsLTRlW5ncujo577Whv4f5uQmlTwawM
ughVA2rHVfTZX3J4dVMmgMPTtnCFJ19rGolsJbJfYNihu/+X4Dm7YMMjzrpCdE08
PBGG9TUeNXRM19lW3WV1O3zyC/NIw+Shph7SOU9aR/Itkduk34DXmVxTTdD7JRL1
q/10M9Cr7YqeeAbDPPupguhkS1VP0ip+/T4m/kIjHUZjGi2xhl0Abp3woiTF78Oe
c4H3pw5pnxbV9Xo9RQcwwRogGoewtaFVQRnatkEay4MxBDdLzExKrezUs9fgMIle
QR0WD3Nz5tO99l5Z7NnfDLUB5dbbmVw60AniHfO+4Z7Y4YnrfTl28+zmdF5qWo88
2pJzuo6/j2rZZnr9vCtWKwIosWf1D39gueM1CF2DE7xbfkhOAI1oa7818kZsgZBp
LPjrNPHVyZJHkIzs16tQPzvvv7brlvl0JVd03Z9l0ekWl8sL9UbXXMPcBgpHuJjC
tg5elzConKGkiKsg2ZWEFk9GIs3UKWex6Jo5i/I1TdwJqPBUGF4Y5Xq4gKHvWtZP
yLd5VMyXNUuRNi1bE5sBbIyTXn/EnNWYI7nwcqjLD9I9zwvC/v2AhGWY8Al/2rO6
Z/TB3ZmB2ixw1DMp7L8XK75wGhbq1WB1IQGqZvyhizaelPFbWOi0fID8EWIC/PrH
xfpDzrZuod7t5uW07VteUfdW9umGVqqcTiW+WivVlHnd+ql4vkLG7Y3XDEcs762E
mqYeaCnxGWJiZp6ZsRLrM59hGaoYWgSm3wzNbpcQoeS1Nfx2KQD8YUNxQmhYSDY/
Jm57uwCKTqQFanxrd4Ubkq2hM0IR4L/e6BFhPH9eXEpnbXNWzag5Xn/dhxk0NbYo
4xaBY/RMTwLSDn108n0F0MMWZQrRSRLlFWyTZm5Hz0ec4SN4+sLmnZiZLjFis3cW
syQpkfrkd+EpRDGDc6/TwtvJQwGvk8GBg6NUJWNVkGUJVR6S1Tcf0xzjOh0pTg16
xQN89QY7xrYlPGUBP35HpXpsnZvRpSI6fH+huEiBzZnULXW7RK+NYICjClc66oov
dBRkE0hMJ7w9fStBKmJP3mvIwH5ZF98CgXe4gLHuOG5OtJUxTdpq+Uel9Nk/jEzC
KGJa5R43D3y6cRtTaXj4hZylYFhxZmLlS18e9sTlDQJW78V8Ew1YOpUdCGkyWQKS
0Oc1j7HDKRcVlJzpA2gSyfnZCuEPpsvP1vvUZLJ+71Kfc9QxL8A2X8NXDUKmWmSR
0vR4Xx/l1vc4++cMkSp9AWrkyQ87Kjhv6klN5M5Lw9Y45jtC+/e8gR/Uqz3TQlqQ
rxidsTCeM3s+X3GtxOhqVSiif23k5iVOyiW/4vcpx1XhAIViAOex5SP4aAs6x3tF
CU3oTlhXFdfr9JHMPSQ/q49k4B52ilHwknvZtLfoYYLOho0qPsaVdAKCYFnuGKfd
VkfhUwHdsRm5zPTrFH0Zyart02214+s6OZt3YO1BTjLovG5DSMVDB5mbShSc0cQX
LA/9MWbHUH8DiMhW2HWCj5j1OZo8mozY2P+FRWxSWMzUhW29ynX18Rv8uLVUX6G2
emdgfoBDSHww3dBLbLyYbcbl8DN7usZ5cyZM1uK7z9GKszQtHrICU5SA8PhYL7EM
977ETKIslnkTDJY2RBeQeLGrVrqcxPjNqI+e9f86cq2ahBaVftTZzuwN2yT9jICw
sqWMWSChkb9JmKnqy82UxyOe9OIzsP5WwGq/7gmIKnNHWVe4v4nENn7RSlNumlcR
0YZ3rwftBYhlvaO2Efjl0zG+1KOvoVTMfdN49Qakqogh7uI84y0asxOk0PiKrEMG
09vTPISFhJMyU7u/CMRoKn9UeusskNGe8QOvddeHVljiZmWK4O9gTVBd3lwsDHwW
DKObaHFfn9ZOeIc3bDlzdQ98Dy5F7TFZhbzb7VjFU/ALD9z9ZyAsDXSlqx2mfTn0
ETAPycMEVly3cPFQMzZ8ut5a66qVP66MDBPfI1+R0sVopG9cYpdk+878hr+0STH/
PeWQLGQoyIL8o1p+di7xDykTQzw2sY28BCAnE9fjoOpgtNLzZ4DJSQo2DSF/gPdI
BjhjoBkLwo2t9lT95BmXn0NxNH2mm+u/9SE5IHLaKBV61Yo7PZvfaGEonyA9DGQv
RT6UiNfNqwH0DsFs5Pslinh5kEZTesTk/s7UgRSvPqDY1HUV1/w33s/bwXw4fFkk
MzNr+XZ+fIb+UrCbaVQaqqN5tUbYWkruZx7M7nOd6tjlSwD8e0tWIX6riffpaDSF
H5cHQoFoWk5pYPaBRVgcVQHQeXyOQXsleO6tmOO9jar5o9RiweayYfuZkw24Q4An
fU3cSCLs0SEiAgpFMZVO62Q1aoyjiijGa/Mz+fm4/xBW4sRIHakef/BWLLFSezTz
m8QNQTqgZZapOHJPq8IhC4RB+5Zpm+mXYFWk6ZMAb1trAh2vgqtOEQ8gWpf2n5rY
GBUFC1tsidduBZwTtJxNAIPhe2MnhHyIT1S4Y+3la063NDHjnSY3fK40/GMeIf/S
XxDDQ82G9iSmCRFHG1SCm14MtUPhy064eOhwKABRytiabL8yjbaxgzKu6fAdPqzk
CuJxAvfxJmRfTrz6oZHF/IFRMiMHpiPzt1wrEF1VfoMAe//IXrwbFBqZAQHrwfb6
rH/w0NXO4cqk4+stjhSHGFJk4Sv1g3MntIyz0QlkAXO4ut39m/5A2jgktZ1uyi1E
s/g4gvY1WxTVHURLKaeX8MYKR9czDBTY2s7ADEuc10JWlrhEHr+G1OvuGtZHZeSL
2PYBxHb99V14KmNzvK/y2ERvU8ZYuN7S3SI2GXg2m4cV48eYwgOBNhq7rCXzUG9C
XHT6iWE8mRj+idunrzdhrquIvYjZ8nakMk1+KAaOmY+cOQgpvHd1qxM68j+nNhya
obo25UV0VG/EBXoSEfvP8Sf/dvlvIwT9fmrTUwmma8kdjeTIhpefkrPka1kVSMaL
9GodSlwE6HZfhRBmtYzdW/81+gQldNX3zevoDBr/QasU38xgdYH9T3/XtjOsbngf
WQP4rHxqX+8RnJmxevIeX2aBgqo1LKmZHb1uiNVLNMlivWyemwbMoqFdojFEXLbo
g5bQ6vzuP40Ce/JBZDR3YBhG2TuzSjr6Yd49vq6lKJLjSDUJXCjB4eDhBl3ENI/G
tuRkGLroI42f6uRwWDU5PP0t+fzYA1wdATjaiYyNt+lBHEgHP2q42hvKXVUHqhlp
586nNxsVtSpr4iqteXxK6cvTz2NksMEu8ELJSNeO0Kgs6Lstwd4PF8xhFOg3BHA9
a+yI1cpLZ25hPIdNHk52/0eSrHQI/putyEppQUf8bLG8KVQNObWJifgkhZW015Dl
fxyGFmT3MNgw0Kd/ED6FPjltdt7ZyjovQmYZXvj8RLtjYzN/d5OQ2ilniyixQ1Qy
rbAfM5+mRSyT3fBIyAFmCakdIpev0ziemg84JfD96q3KMIoK9fj4teLX3qPcH+PJ
t5E3Ys1Wu5PLAf22v7Y54GuP+gVY8JdtDNFE+2bqocekGZVi3uA5zWxzLSh4VFmI
UVer05QShQZv5JTouf1vKM8QHoyl9c37giHdsnFza4DYq5+ZD537gX8nVvT95LxI
MOm2lN/cj3bCpAY0dlmEpjSVuX7LXtblDAWg2NlwyYnxodJdqE5c80JIqX7DdAcP
0MVb1xrHaAOP7JsMLVkUYkiwS/vS3zSi/g1aojpfhqXMFDGOYUHTi4vNgkry8Ijx
M8SLIrzP67ULcRfF5ENU+0lQrALHODhXrYFCf+xJJJFhwlWE/Q8rRhEqh/7O6fC1
t5XLcise9h6nU1ZdP806QN6edaHGGSG4YQBywP/oLPCRY1GLgoUvUdIukQH4iL6r
lbwQ4S/Vx08Lal54G/+4Vx7jj4d328Oj+ig4Q/SfuStpVfMT7lOwztgfDgNwYvQF
Ew7OkT8otdB6zO04SSfZjFIUHgDBtbhfdZ6iFK3b8TcmnqjPH5i/8LLSf0werwLh
bade2mhGUQSauv+xMiAJZPNPr8UpY/3c1zoKDb65X3hOusG/5zHbfGY7XUJNLbQa
0GrZciuio1dlSn//JiK6sTkvaVxMmApRh8MsQQQ7lbEZVKdDvbMG0mViIZvwUjHG
YGR7cRkIQc0pAfMqzs7DISDtCikg1mXNQReIl1FGMWuf3oReNVo18TtwrB4TFz9I
3Yxc4C1TF6glP0jSyCHfwBlKpJ6X8yiOWlXJFFeTkiA=
`pragma protect end_protected
