��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t�ꎜD���O�9	/��H�ž�_����p��#~�g�7�5� c8�WL�M��ͣ"c�k;5_�E��PǯR����� ̝ �����ܡR�6נ�Gr�a6���[M�}��[8��,ő��� AǠ'sQ�JR�-���zY/���TIR��W�#�n<�b���{#�Ս�]I�n���Q��b��� 㩼�u.�����R����zR��M���{*��,������qM��ui�2�Z9&����)C^�c�3C��]��S�!햋��:���%A=m6���)�se���~�y�m�s%��^bx�'a�p��� �;�{��6@Y��UL���.4��H�:9����[Lj�4U��6�������%K}Z�S͔M��βH��[�nIx|��1�CR��� ��=g�&�鉶���yv����F�T��#�p@��ґ�pC,)��k���������G��}ofԟ��Jk�:�[e�f}�=�rs\X�Xu���)M6�Ki�4p゙�[����9�UN��i��ڨ=4̯�x�܅;-�!HՎb�$��x��L��]��5�d�M��C���ċwS0���~�4��4ShpP��Fs%^ަ+��sr����ctP��;�?+M2*�t�82#�U��&}��G�S|`��j��}�����Ұ���}X��r�?��RF���t�I�3��/��Ze���T)�����ا��AOH��Xz�G̀�oq`[o>�+�X�c���8U5 `_������a+B�|(&�t8
��w�z�lFx_�����$D�q!"o����O~#�a�ݖ�����0�R0H{��w�c�OiHְ�êU�Y���W�$Y0�.@�oK+�Et�Q�=��j$�ļ���"7�e�ZM�����B�x�J��E�!w���.v�yjU����ҋ��Y�����%�|�٤J"�o41*2���|? WO�3��2M��տ0)���j�es2ثnɾ���+]�	��qi-��� ������刍9ݼה���=-��rXa������K3��x�^���UAʼ��M����,*̘5"(�c�5�ġ͐8=�o��Ρ����"|��<3�΋���B���U�@q-�%����>h���2ܙ��I�4�$pݙ��PW;(��^_n��tG6;���a�ut`��
���0pP8��o�����q�F&�^Sz9��o�V$8޻u���L���z0Ǚ��Q��YS�*7e�[J#�[2�-I�B�[�9h|v D��a�m�a�L�Y�����](��n�,���"���� ���,s�!��F�aV�=o�K6%���x�x�%y���ٙ�U�oY��Κ�Ћ^����Ä\4��ĽO�}rb5�� �q�d�Cɷ��`w>ee��P����~�k����y��W��������=:��b�V�r�uk��^	K<�{&���N���1�O�͝n��
�I{�1���Ru���=�SZ�`��7/����' �INٿs�=�����R�)�J���� ���K�l�TYSp3H��Q�q����� }����2f��(#���lD̀XԎϠgW�����4\ѡ '�vY%����ai1JV���!$OA�O�x�2q�$��+�7�$��n��Φ�n� ��ӹQ�6����_߳��֢Ǔ�>ow-XR�=�2��x9���.s�K��,ܪ���f��kE�̓�����E����C,��2FUH��9_�o5 �V��nd�B����T��($�"p|�j�؎KU��l樵X^��e���+^���1W"��$ ��]�=�%��`iU��+P�WlE8?��6�S�M��}8GqeSZ��黸���J)o�޹_�26���N#D�]q��n�h�qw/d�'폞��__!���A	pt�:A�ۛ��� Tx,[v�\[���7���'��e�t���̾�«pOF�\�L��x3�rz�nTx�i��2�!�C�΢_ê[O$�� �{��C<m6���D�P�Q�[��y�xu���� C���:�{ɺ��v5��p1�h��U����P_}7�'�n5�aj��1T=�M�E���wJ[Ѡ'D?�����M]�����&?��qWع+X�QЌ��.��%0Q��C���o��RY�L�����8�x���T�o&-� �����M�B��]��FN����QHe?#�Kb`Y*}�w\lhs�R�Y��Ǥ��(t紝�7��u��_�f������}jM˜s
�n"��Q	:��J��.5��&p���$oU�9��Dv�-�ʞ?�4��OƔ���1iiޮa�äm��)P����P��1��M4����Md�k@(�/2ƙ]i9�g@%/�of�@��͒�a��Q�_pXGި=�Y2m{�Dt-ڿs�;��:˙G���?n,4IPCxe\Gy�o�֊zJ����[~�ù��[D(}��扳�^�n�K!�m���Z�8�6�Q6l�<$(b'֒��E����J�_����@-V�U�;Sr�j��S׮9/ƛA��;:��^?�2)�n��dݮͶ�c"�N�o��6��u��R�E�݀��7m����b����c�.^���8�fX}7<��pn�����#��R���-R�Gq5��/K��jXmvhl���ʓ�u���=?����Ӌ�+����MV`EԘ^'���k��n����a�W��?��Tr,����s��U0�l��d(�i�h�d��#XG	��u�l��$9�aB-W~�G~s���\K�G�h!8����B��_�h��g��L�~���
���bLP^G8�����+���!H����6�C*�bd�Oh����9^Y�|��
4x��'�DM�zN�`1�x���:���%O�G�ֆ&j{����O��C��nb6sj$�@3�^�Z�%-F?x���Y�r�0�4�6T���Y�{�L�L5��s[�J�"v6����g}/��*C�L	?b,5��C��L4�~��Լ�m���f��E^/����2~�����k(�b27�<�a\���mŎ��F����'�a�z�A﷝�zk���3\�`�޺�8�1CQ'ːa�q8�p���mVX�Hh�V[��~wP^��6�]8��5֏,���X�Mیy�Y>�� a?|ئ0.��i6'T~��s�m��[�ʞoC[�$Y�x���)x��Y��tȫ,,w��ѐ6����aߵR��W�B
�oG�)��%>���]���"q��(N�ǿ ׮�l�S���P\aK���a�����}��)Ns?#6���i��v�U��պ,8W3�aK��TB8C��P�Y��[Ye�$T=��õ&:�dނ�g�h�(2
Hk�UC�j�3���Xc8d�%�gw���F�6����6ȧ	�@�܅ގ��b�)};�����p�e�B���4��7^��(B��t���������G�NRZ��Y���/d
ɹ`5r&�;ʣu ⋲��Nb^ͺis��)�!<aAçXj�Hs��J����?�Pz���H�Sl��`h9L��p�ޠ�@pn��8��d� i���"n�c�R�o�%ɂn�f�qg��z7�O���`J�s�'����Y,j�E�v�Eg��"k�")R������S9ɽc`J�4;��gn������hn��,$M���/��r6��Va��߅[�:H@�n`���_�uZSIu�O�=����8Fܰ������9�;�PFf�^��6�w�ě��rb��-��}��s�H��m �R��_�Q�C�q���;�3[��b]o��+j$	4��E͒�'rp+��yC�&e�Jq'x�)�]$=�(���JT��i�'��A����]�8B���Oe ����4)��V3�p�wcgH��>��n8���苙І�.t��ߘq����Y*+��'�����P=KO�2�ȱ�ؼ�4)�N
��c�J����e#8d�4��Z��C��T�2qAdT̈́������*�`�@H.�_t�Q���C_��;����t�Dn�b8!ʿՄڝ�#���j0P���zï'�Y�n�DH��r���Y�.^9��^�u6 dK����_�e���h�w}_;��.���O��,O9Ŏng���_����|_�؍Q'�[�Gs,<�QS'&��4��ࢃ�W��z����#;�e	�[x�=��������4�e�p!}���� v�d~��7���
�W���B |g���ۣ�CC�����R�C)s?( �+���"��W	�,����R��:�p�j�z'�N�)=x(�tLA �b��Iݦ�J�����������F<��a��xe:q�%�J��gp��W+v�B	��[�y��0�nw��>��ʣ'�C��� 3�]��䄣�m	FG+L:	 � �;��"�܁��ގbv3E.̟ۇ���x�Z����|��\��z���<��>+�A^��3��W)]��������&�3��mF��X�*k��mQ�;D�X����Ѥ �WQ���C�R����'WIn%�{���2�N�������(�ӱ�$�DL>�lz}=��z{��(0DF�#uG`զ��[e���
�:Mhh��l�ĦzW�&E�#|h�M�y=W�iY�]@�Q�^	J�n�r�My��4SN�#�6I��A���|s��o.�@�}�qW_|x��6gW�9-EQ#6Y�Y$��
vb��}���Kh�w���h�]�ِ�C_���B*�*j��pM �3)v)�ƽ���(mQ{���G��\ji`"�,�5�/ ׁ(��ۑ�ת����I�?���=#j�ȴ�;�!�k������P�E�Z�]���Vo2�Ik��j����9�ֈ\�%a���=�*x̎%��B�����=4��n*�jR��?SRC���=��(tm����և3���j;]�}�9�(g�Ȧ�Q[22�gcç�H�S�sـ�ɸ	gлA�� ��br�%��̛��`�
��Wafm�;/���'͉͑�ly����i8�u컯�[9��"kKRa�7��MJ�8���q����4[��	����<0� ��,�#��y�Z��8Gk&�H�ۚ�s��YJv<���m��Z'�DY^����L}�Z��%ɸ��~��S�4�4X�n��S�����$��]�r�vgB�Xl���Ȫ�<��!2��\��F��*?N�gL?P����2�#�U_-���6{r� �m���~�[��j0��xI͵}����]wJT��54`�ض�$�ƤV�U�@���/���:��P��hzX�\-�h��j�Z���X٦5��|�6�	�28��ʈ�@|0$���fB�*����u�O�x�#X�*�}W4�L�|��8������w��T�¨�?�@��*ux��eF� DmlZHW{�� ��	�[p��Z`�Z�u��"�f��ڿg���v��TO��!�m�G�k��X������]�j�&xtx9�rlM����FHe)����ifXf-l�EkF�������eŒ�3�5�ݝ	���62�����֌#4�>�����`���Cy�S�d�%�i��c��ͧ(}�1��?��˸Q� OL*�N�wF�~�xt΋з�)G��2�C`(ڍ��g��_ȫ���� s|�۲�7���3T��X`�8�CNYǒ֡���{:����-��qR�7i³=�Ϙª����~}�[�"��W{�Aa���^Nh�4fR�J��ک��v�ȸ-2귮��f�0	��;4��G���b�������C����G�e3��#��I�E|5���`b�Z��.�Ԧ,��f}A��-�����=>��5�r9��O7�mx4Qf�P�	|B��]�S�r����+`�k4�O`��ݲ	��GV����Dk�p��♒+�cL�K�D��n��)ch����N�-KW4�����M��r""S�;��,�3~��!N/,l�SG�=��k��44�0U�Ȓt�k�ZS=~�-�L���)��<VÚ�݉ԭ|ny�sq"Tu_���_�b���d�ƞ�y�f̧�D��J���ĩ^qW�`��(��Tmfi�IQ��
K�X�)r�DN^q�O���s�;5+rd�1D�-�S�62�����j��%?�>Zw�4ޖަh��|a����������Xj6��Q��9�J�ny7`��Gu4�� S��:,��F2��<����H��1