// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:26 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e7o4GmurOXethxerWC/3W8pwETunAdghP18RU26TElXxusXr8ychgjn5r5B6kszK
mw+f2XkfkWksJteNCh6F+ogQu9KxhwPiWOMOZCnXJzQVvGGvqbCipM+twwWNb8QV
oVnRt+Kqsc3j5sCSKu/i9bALIt29DkUpxXoJfVJIzWU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28208)
mcJnuvgbdV4sFluh1wNH7Sjn5qe6KIzJBcZONlNk5pfAFwn1GkiLkv+HrNRCsxAB
RVVjCXdsyJBMj5vgXP/9VvrBv9btVQVHSu5gXusZMhyHm/mUfCQXYC5wwC9hA3Dw
Z+lB1hxm9oDMpem2kluSI0sERsS+5wfU03d0t/JXZQKbcqIa6SbPACiKRsD59c+d
lOOY5lBIDydV6cag1oiI53YjeeniBpEJGmGOf6bE2C8Ujpewdt7ZV5Bbb3WFaznG
AjuSUyDO3uC0yJ+wLtVZQG+4pF2Snkp7SpxrKfA1T5NmG3NcAJpACeMt5iT2xH9e
przWmZZIyaUTLo8WIXdrwOWIHUc+RwGBkim1QdcfFbhupSyVCjI/0rZZ7K2qsEHQ
qxxQE/Etdrw6uJ1a3QEXf4jEzdmPGdS0JfIschcrq4hYFZWM3nuqwRdPQ+8DN09c
iXNS2MOUnKICXuEY5fMKRlajpdwG9m7Wxudy48+ncvF/UPKJWIrk5xqtNeJAUX5z
InVtjNg53cK6uqHuz5sv0dZdJRkXalWWHJ5qQmx8sD1xMLSrlfLSbyRz5+FqqyHH
IITXHjtGMlrJ0lFPDGgyOkLbyy/HOED17pN8zUZQgGjVFVYqmd1ZrBbayqmVHy5D
KvgO4IMGuljFW9GZ3RXrKXKYN/TdDO1ST+/qy/xifAs609NRu9hW3QIbUiX6V6kC
bEi2028T/hkjEOH7iRg6ucZAqEpAYeKvTG8xUKo57GieFeodLlDRmWB89uVPHrTr
MorlF2Frhy/UEHMLyFLx5M5VZFGLpuTnGYZTWf/6ioOxto4vSM20P3O7gaCxayz1
P4o6wzLpIDyQ9XBoHT7h5R/IBAJmZ6tNKE2rFhCWKM4g1VA5Zxk0QTGzCNpHrqEt
sCkdGjgQFl/Ceeo24+qS+hkUGfy9uS12fKQy6NQh7mVJVY+l+NqSx3uI3IUB9Sgc
8vxo9lgpdL5vywRhDElDTlN0AZd9iuazgC0WN8zm25LnkrU1qSgJzbmdA80pnSEG
bYFHwfPQ7hD9iQRDRqb4h+9c3fg0PeRnkPEmmUw/FP1Q3/dEyNYOb7I8awGT92dH
zCMg/62b5V6ypOcogDHALpR+gmn8tKF9Keq1KRmltOcWQ+fijEb2DQ3VB95eSTj8
uyqhLaN0RHiP5YSvipW2LkR0MSfVBRO2dO0k4klpYtt9tKFHBVU+G+QQijlsJR88
Ff5Db/EYXj/0PTDcHo42YDYqiKhxoWEu6G4m4iXpYK3yCT2MyGvwm4uem7oOmPun
7vv8QopDpBMX2xTfKNqQmG0jOcAwimvlM7Li4tOA5issFmFzZ6WAU/5S0YsFkL8d
f+rVUgP6Jccw0KIc27c9nRbV0L9vU2V7HE6MYtXp7u6joJvDF7OpL0vCs9wGiwx4
l1Yefmp7FhywvHtjbc3fUuZFoO8j+Wxl68vTLqXxnsMv31oNe6UT4TrQpsLvA7uz
UUxVlfpq6pLiz5JYDIBoW398BQ4YVKYZquSHtfTQa4K+TCIj/IVx9oCXRgz4jV8T
ogzwLdwaIJhhOqzzFHxCwmIcv9zTHVHDNzApYiNJufwB/hGJqZY/dk1e7PA1HTBI
rB+/vdsBtjwnkcTT3H6KfpOiMkIQ6ew1pPYMCXZ15bnK8c8d1zI1+09mLV3okNJA
U/QMvf+pTbn7gY6ZN4eGDTCwVRZ8oTrg9kHroLQGnGl326zboAMIAEU18Q39km0t
QHWIm1QXwpkuXIWMUGPiVJWoR4zqezPUUyiVKXOxY/c8PRw+OcwD7P+RLDrKXb3Y
530sqADAVyOIyftHfU2nXvzAEo62Y8OQuHh19DiXOdRUFhhYHZ++ymRg+9qUio3a
lHfuktknBT0spvEmJezNRuhibpublCVS9LfVoEKAvQmSMLI8jXsOw6sVa4/mc+e7
ceogyADyB6DMH9XaYGfSgZZjigvnGZN8GwAO2tu4rTZVKFFyRtbJeafbf0JTWCyG
ECqdizAzSzjse+dXVmpWRp7y1AMvaGG4SYjy8FmHyLTrCrYETm4ffPGjDWeQ5zSC
rD8bVVHcQl51VECmzawv4beoLnsg7IuIJfFHPkl/x18eHqOgH1asewaJDG2QTYaS
48tTDMEr4RJfYlX+yY4Ou0wOBgbubzWQpUs6HbHfHDlReK+kmPHU1I1G+/WjBMrC
1sJO8XehhirUGA+eB5M8bWXP2Rp8+gj5ZEnCuA9AbRhu6bZJoNjG7I4DIIl4dail
/qQBYOAaBoiSjIBlFhe+fPPR/pL5uC8n15VPIaj9Yjj5TPUGLcBEhpaU/0cObRqk
2JFZdBr9G3UVWyJTcQ9qJCejnWweltlDXwJhPqN1z1DoQidWstDg9x61VUoxYkk4
ouhUybqcVPS1f89Le5rzuwApFEVi9/YLPG/zglddWi+u8RmWymteoBKXCJ9RCSmh
4RPZUxcrKRxtHWkC0ybfknNwNsT0R5r5rdN6Au2WKD63SGgeYK5c0f049G8GH1Jm
46eQk6sADFV7bIopkjy+QrIZlAfW8Otw+iEoO0+vvBGBlvIHxJ2ibHkrDoFI5JZp
jQTmzsUlslDHEA9i+oyCx9xHk70hhD9YkpJTcBsnv82zbB2joULOtQXwf2lswYoT
iaRU+ZpuhugkFtU+e2LoY4iFQzfAbYbUEThAWzUKrJxH2shxx8k2UF15kpwDP5UL
jaODDTglnGokxvNVB/oNcOETw/WKbnkihgdBW7szHD5Gcxwb3u3zKgH9Lt3lTKOI
fXiic+vvwRp5bf6vSwlWaHNlZQyKLAbcmhDCGsgGI9N5MJN5w5H03NuaTlZ4AkYV
Vvqu6UJ56fhVYyI+CXIscEnDMxSwcGgKT/m3j57Nu8nA5kQ88WhH60sVZ6bRoZL7
sYmggnSB6bIKKJZ7LHIpUl0ae9n7NgtxazDV/faqMIwicu23jHOTT+iuqPP1lnqY
DlPeCOjxVW8P7dBPSC9HZQNYk6c9+K1dq/yjQgTa/fSxKk+lLV3tone3RCVkX7yr
H0WGWIN8oiQVfI9NvWiTM8jKiVi4VGgBGEklEkwk3d9d6mXxKyG7RmPU+SYY96ey
BD5vTUyPjqXa/K2CswfSHj33TEEo30Yyb5gINlsbv74KmNgBDJf19x8UHnifFYgx
5xgU5ULDHo5p+cRUQa48Nii+5rxm8GMLC0BITu1IBvHUDiwyZgxraUsmROkHQgsB
XTW2Ct4SwlGNwbNe1AmrWTqR/BvlDjEl3G06wFkS4MxEFw/2Av5VgYuQNaS98JSf
ZVZDhvRmQ3LlM2tAt9Owr+9KVkDOxHHCJgPcY8ZaMp+d3IXjteTAWzbnLE7SSK0h
ICBbYkE6uipVUio8J+t7MafpZpTJsGt2exvKZfF11k5uAUacuIKhQBOePnYhn4W3
IKX+Y1eyub+h0//vJ5/KG+ruxnB1dixBZdNS4x4foeRcAB66inRB3gGP1jvGY495
AbffSRLe05ytIQo7EdL+yih/wFCbOhK6AL/CBm0vkeS2pBCjzfwWEYbDkWUwhFOa
q2gafgMjorNl8l+MHE9bl9CRtwAaNLF/yDxBqZ0LB568MJPVaS3SpPXJzM67L1Zk
/AcABqLkMpjHWT2iRcL2a/pZoeVQ8QSv0ZR3x8v1IP0mwHKDx/a54vXZiFBY0WtO
mfMJxZ83NEhgDd0FAtpNk4lixnXUndzLUvM/VJAMLObchzF9kfufnyOzecLaod+J
oEq/2MDwY5oXrqBSDqrWjQb4h+0iXvKyxQm53+Xs/XPrwvONLXQ2HpdvhU7zqebm
aPjPhjdNmuOO3Exl1eQ6c0Kooyehe7I2+jVfjqis6XF5deVJHBmHVq1Q9/fqPr7G
Sfk5rK5a1RO2KeGmU/BLCXN8G7boOzYyrZaVrgHjxRwTkbo7N4bBuO9mpdxTe5x/
IQyJL8Jxy3AnrFM7T1hqISA60p84tM4QR/9zjPx41Z1NXzb6jBRipe7UbzFjGEp1
cufYBshD/P6sLthajba7zhOUegrtAfxBdF9IQRiEXS0ttx+a77fcJxVPj4EarkTx
IHU4l5Qd1LtbK+Erb9WPjIFmn2PEhi/3iQz5gjR2ktn50Wc98AdMOIBuAqF09SSJ
4vUjTPodf3epXQfiTROdAPeUixp/dib6ffD0jlCDA6Kv/rpaVdOS+z6DKMSn/9wE
Q3LN0QsXOnuYF7VBQmc2SyyyU7dnjuCGehaC0+GmekQLIi4r9G/ZM5Nq3rB/HbcP
342UsySkCqfok8t2LlCKHCgKUcUC3uBcri4G1pkA6F4xdndZ4ILvRDPPTEqZmCMf
QpZc2Doe8x6fg2BrK6SFiRmNHWQjB6gaJkknPg75cAja3CBeYKNW8j4CKn4d5nqg
lUZKUiDqv50rA1H1FjOCdY3Mf/lcx6g+2pi+g6VHps51szsi3xUX2sDGVIMGxKSE
Wea4ryENMuselM2KmMNbGsH3RYtnj4u/N2H3FeCE4dZ68UU3tkmHaOlWaO4bw8PR
W8RBzc6tYcS6QWzK33EhHZjz4bmDL8Oyz5FeSIVsivhpo6CHHOoEf70k3Zwbv23r
i05HW3v9pvhXoOl/tgN+7Lk1UaP0HY3njUeGEvu9Gwu3PpiUtLYvD6CMlueZrq6x
T6if2gPXbwt4uN+q0iwDRkoP4FlYTrCYucc5inEy/4U1Igt58eLdUDVKq1t1ZKB/
lErYjQUM0137ey/O2050RvThDJBRyC8RQHersGQlebuUMMvuVcHkmpvdsrqgO9HZ
nuxZVVBki/0uxIJjRMJvcWJx29pn0D1PPnAccsy6CPjzO3TbfC/3Pw1ybKs9Rs7F
JsvPGPlKXODayLTK6TkI8BFioi2gmNpqaunXTApRkEfFnyz2ZK+mTiZa84L7M6pU
XBAT6L4pV5ULUsy1MgoKbFiDOW11DT7fyqqQxgyq7johS/aFPjPc0tyVZk9g3Bj+
aZ4yKcTGsQjYXWAwwGq0F2tJ0xCMZ1gVB9G8iAuURh8OHOOVCqMwjz5XcJu+6OVf
iAB04nsksL139xv7yxcFcRdi8hMIVKsbVgXS7KhWwqYm85vKc6477omT6g0vPFfZ
xd48nnLILEWhbL3BzXWv770CyB6XXcwXjaL+VEe7/3fk6StuR6k3NQNZJJJ+zDUv
uyB4yQaYwZFBwtjAa2qVn1jYUtP4pwaXMkcnOzCe34QVeA+S6eCF3npeNkZ06Sqj
/qDaZ/u+k1lvPpUxVXUeq3ObObwNA3UPhf11n9JdlZ1iOuLmqv3nLhJeh7QtzhJv
dm+hVOSlY7uEDc3I8vWs2ku6uNCCm9LDMVYwIfYFR8Qrp6Vrz5IdNMJbXMYPqpwL
4ud3/6yIfNOg/SqA0Algj5Y1N8LxH7frwxanI2Q01LS7OPRLV+VSs4OLwOZFQnnR
3qjWHXU+/E+HVRxOpkqQB+ABD6/8rfMmXZRZ1KdPUW64WT63u+lBirsk9o59LOLs
fP8RKBhHPiHoTAZRQDYPULCWWP1DEUTUEej9thgMi/JxlLRPglvFiDs7NNYzKoc/
fF2hj9R162/a3CNGusj4yLSa518zb00BeOSrWDhnJYRxAdq0MRXPgro4BQGSoeIn
KvbgC8YB7Sn5y1b0ktOgQ6aL8rcS2Y/y72MnZJ23dyrdQsiDFZCzaUibHbIYSRmT
CuySCccjzEBjHMgOCcKxMcjuTnbWluUqLrFP3FIc2rOAICAIPIASVwHPJ+uZtPel
sJ39k0UDyOvuDEbJOcwrL5ZPJO5+DVlP0w897ZYb6oJMyZ8MRTHk0DEDbEw1wC/f
ievpcnptlZDa+LFflbc5NYzh0A2hoO1S5/jXYPxVmO7qkeAwqya5eFrXs8OGRwdE
hrg4vaVkTxCfwC78AEsCWPibpZE6E1RUVyVt/iwNUw8uOInjztLJlKCF9bXb5rzn
/FjQU6foJN8jJThdngniECLKm4q0NUtzvWLF9f9tGUGeemTcMd+RKyqpw1TrpLSA
sZIww1RhE2f2I25YVwkOaOAWPzXhMp3MG2ORK7RkibOQU2/2nctoa0DlE3+FHLe2
7NQQyzGCIpo4fvYgXQBM/LLSHz+kUeFauIknG4nT6iYEE8DAr6GXqwyF734AaZRn
VkyP33Rm+jK2Kvme1rWvoaQHxEKv/5yWESfoiDMBZwlQUupaiowKyuTKvMjO/7mz
CRj0aNbN9AfUYSkI/rBYUUPheI2KbEbrwL0uzxDgqKVUzMOv2nOxmIv0k70q+r+U
XySHMiCWajMhIepPsZEvv8j9Qzs7VVYSfmdTHZX+vwOa3q+PUc0kb9ESyqJGcHbK
4TFheDDyKmwLELANg3qF1vu8JmufOa7NP6kTEuCwHOfjt2nU13mbRS9BKXTysCeV
t8nw6PqRrIRGc5vhg1Dd3cBZEhBAbCQPy+WFiMsUHVl0IHBx+AB/liaJ/HN85+4Y
Zo6kVh5Ej+/psQx0UoKT8qAtRst/LYSu8yc16iWL9huJ9mObby+eHZ2a3xjxxuHF
dGEWAGfYqhFEV94Z0fZmbE4e0iaIk6+nYvKW0Nqt9Gd5ISo5bIonxihiP+zM0R9P
P8gaD626NclFbuw9UcBvVG0TNGbW2PsysAnl4FZnLjAgY/1zvk9g/AxDK9egwy/G
7gyLQpZUEHfif6H/Q5I0regV6WmNpocREUCjxA8XX9h1fzCLq+NWgUlu60vLjwvL
AFBGF4r4vhA8ddcN0UAaa8vxXHGdVGvs+hWIiJ+WzDNd/yBjTlOkvYYqFMYXl9yT
hzdyu6ikwH/w4vdnhdwPaAWihnZqjosPuMBKYst3jU2ohF4qsZpzagOhOWEDpLo/
I88ks3iZLvx7oSTowiYwUnDNfLiy44CTlrdbZBXKytT1sCO8y5drDrooy3W1iMvX
wW8QDUnOUFKALrzdH3Z8ZcUJYB189iaIvDTgXqgq1K7p4PctU6JZ3WloV37Ahqao
VgwSl1P48iVSIGehNv5O2U764F4WzgEeiJXC1xZABr0B/AdpHRox7tB9Gp6uotjH
mtnzIXE/SivbdE/wb3LFvxdM7/OAHR8fUQWPypN2dTuo3Yn8xrfmIPHk86pBRRMv
5Ovpd+mvihQDQT4Ur3RaHt5Fel1HkaqbG+28TIJw6N+oSJdK/HFRNoxlZJTGLVLw
T0JLphJNLxzpxHY+qFDlyP/av56Ejaz5jFdoYWPWwXaJcNyUYmx+RBelkPs58Ms+
cuDwgAbH1hAL96KkgoqCZ6MXULLKoy4L+GLMV8pcZdxbgoaGZFMV8yd+mW62bDaG
WZF3DGPCbX/eSLBbfz+8qVnNRXjfnMw/bqhPfV1Q23j3de0qrHacabxrOGHWIL+A
sxQ401qDXQ555hrUs4Ls/SsfJmr8Ub+ylIW0wGI8mI7u99lPetXS9eiLFAQj+1oG
WbBezAy772vZ0wubnL2wcneSnx1MR23N2v6rJSf4QQVcs4xF059J7+OfHQZYeYYr
QWlzOhZN0R7Jq185ZNXSPm32t8itDuBCJ7MoZfJcsNhkSM5GTaAFPCKsPS4ahG/O
/Jc+oLxOCUFm3SkUQibxi7gt8RIg7XOBeyjtzYxDGzN1w8zHLE/5124xa5wSZt27
6vQjKokr1cvT9xIenIAddinDzx/WaqM4mKTyNNfIKIl5/bXYwP9/YkQur+lsN0pW
uFx6LUOb8VqsQY1lOyWFaqSe1+9U+g72zI1UkQP0ftreCzHzHK4D3xBXyfeeEEz3
4TYz/OJi//lTYP2hRlEOcQW/AMm5reaftHEQ8j8V8IN4Qq6xW3X+0WfL8VTiTwGd
ht/yvh4qpM7oKJaCrW7TI9WVjaWpSXWtWpGng9AbhFH4bNiKhgIhzXOLd6rKWYC3
oml3vxf9Ci0h6JSSNvAK3RNnG+mpSErdIKT+pGb2LqUaRMFR22z2zLtgP5K/5Caj
xFanbwi83SOvVGDTxOx8BN1nwWjtHKqHHueDRkDJJCU7ZhEluhsFiRkdQpXDtSEH
f0lPBjmJFSwUvmqssy6dZNc7ne7ZoJsvW0grxy7h1/HodZr7ZHIt9lnq0Kvi8gzn
sZhNzUP92zDNUyjTeKCxCOCuICDPeges3oI9GYwjkGF2OKf3288jNZuPZOy2oMjS
YiAx7VZvuaeTKNxXJYMn0muZtEhTgq2PXmAucLumK8VNkaJar7Yg8STvN83XuGEs
Meyaa3ijkQpBiPVKyF3cLUMa57rw3SSEVumm7+xobGD+ve9M/WDeE7ens2kaFSVa
Y1fa2a9wbNQVXmAcjYwck9WgLVTLC4K+72wSsNQ7r5p/yZmB0wE0NSElQMfEJLau
WLnggtj31c7wqBFqn209eUC9Ldn5J/J8WUcvdtBVSbalsT2jmFRdy2fx3fLlJpqM
2vFn9Mpz9TcQKk69r23b6Chuo3EDWglBSKSZw3W/ozetoEBg36K/7HrQhPH6v4TE
J5f8uWYshkHX1hh2ji1OPLsb8KLLEtectihB0eUHLmBS5+URC/2Dsjx0yP01cIx2
mpsflo7EKuqrT6Zr3bkA9bqEOLrtPZVPbaFuXFxMn4ISO8Utrj7VGCL8ReERzHAi
aeMe293oIfzmlwPEeB1ZMifptjh4payJcoxI288qhZBYZCjujrXbiqy4D+F3FjLk
8b1gtUVLKNoxSK9yKxxrAMLGutbqKDNSMiFw87OM8Vlxn1RR+MStSkelcqululuF
7dP5RdHUrMuJPD7kzUlQTrbWYNIuLzdMY0O62l9gj51eE9FnLGpU+VT6QiieSCJ/
jfAvY57JxNDoGQMs77x4UcbpcR5gX0i6vBBRN+utO3aWxIYLqKg2CTIIOOZM/Bdj
n7Vif6tsne7BDIqCROxkTym2NX2XjoCjGYnt/OvlSFz9C2Ovq5n4MbFa7Ey8VAlw
Z/KOrU81rBYt3WWxU6FBbwQN4+dfyYEQFktWVuAkiNkVITjEOp3xUvH/oQhv33SJ
1JNkeuo9IBPr1ZOZG6YqgPpBVu1aITdaYBlL02svZlIltwpXwYqioLl/G3lYAc0y
TNDK/VKPd06iLkrFQTVFsqfXI0Ou9WTd9xvY/QVXAjpFi80jPR611Cgliv8acKVY
qMQYqtMSdvbBYli6CeZ3kDVDirzlieF18yVMVhp2VOHx1IYL67rDoWjlvgTEdf/U
FrbU7JqFAG3SKVRFr/ORscRATNDiuo7JBhpfnERf5VBK8wMWN79nCqT2kiTxu3hL
NbCQqwGCO3LbQnVlb/zH8WqO69155EklELnupKTNc9RAkPLYAq+c/wCifRgya6gU
gt7ZKG4QjUYUEzv3irOsB2ryTCwZEBllxP72tb+CzkqS4vsEDwZuDEMyByEIuoqa
U70B3k3Ff7UT9YkmhXNBwQ1gdMbRyQNBOLom1TdVBH/5y1/03D0vxU2CwiYAOFcM
VJq1cDzWHIDuDlLWoj+1lbpk+eRZRDQ8oalWiclT+x85jflfPpd8fBvrL98h2StC
VaeQsxdh2WRYhYzR0MQiry/4xLRej3Dp5Ai4Ucub6gmv9lTph3MpeWqDMl4UZNzV
Usm3D+9WH4khE9n8JrHFmHVSsEkROHIyN1HrUZUVskfJuJsV/8Q/p2uZqa1hxM5Q
l679liqXJJAvFjkRMVonB+xF8El5ANAQD+jx+JvzIOg9aBLE/sVvtoOP5hLjK9cI
zgCjd5iq+fFoKdsFEpqAf4kx+hFG//HiKCahfBMqbHufhKoC/eFs7T9a2jp08tWi
sfmqdeOMZJSlCK6UZ/Jafl/KC1i5tBERSyP+JRXXuOhQRgj4HZVU74XVID7ERqTz
cNyBCEGXKu/YgCQG5CFkb8qXjK5dh4VrpxDmoHL41Cs95Glqw2sLhsl7FMvs21iW
ZFz3DuZm7Yz0CjpBrKrApWY3DtRb2iV5/hN1dUsk8Q5HS0i4+FvA2PD+F4EA0Wqi
Ddb82ksco3C4impvyfi9aOb/RRQaIhts8bt4GVvGS8Ta651Lq9Prrbd38ncm8Lwh
0DtU9BZzjyl+ezpTVNljUojTmY5fA/6kmV/WDttOrlDn6tirugzt2fr756GvYKlj
mkMymTKFtl4pmyYQ3i4Cgm1YspHq4dWYfFftXOw8DANC2/Eiq6fnvJHdbR71fEmx
jjf3tSXISM/r7xwRq6zz6zvEmtXcxJNBYoiK8z0cI0lccBByM8+JXi+tYHVZTHOp
DIra8xvNFQ/aQ+QnkFd4xRmBG9pT63VUb7tpFBMwJGz7JY0Q2s2vXxsbwN42ozas
00kdDOcLRDM6LIJrZE1tD42GY9DmSnDThxqQLE+HIPdb46rp5fqqhmZelIaZpl+v
2/Xk3D0d+qyHrLS3JesUYywhlvItYmd3MSwex/67ETTrIWNXK0clQ52XEPmxb+Th
qt4VyoACWOaVwjjHqH54L8TyrBDfu76WSUaUW1BswbfFuC92N+80/jDZXfzEpBEq
w8NSUe5ytdi93HaYiroz3Syre9pZYDSKfFSh2CBtAp0EXrt+hKVa9IJ5Zq9tI+Ex
NajxeoWhM9yGWfkLH5FbnfZKvEaZeCYCTzAoARBf6cg/dQ3F66/uSQSRNgotLM96
XAXYyxml/UactZl2gAf4LoAgAE52huPF4iAoMzJ8LjBJfzk6CWhd9dbHN4O1A5Nu
QemMfr482z5RlNGAud6itSstzPVnZeDitbH0FzrloueZdjjqBUsqlxfwe+zNxnQ8
kASi/bdKEtKe1mNYFDSmn0GrCgnzSp0f2UQ7OeWE6zLUh70ZWACCudWsgfWoY4V5
9inpvzrFDxTuKaRsfL4a2ly8gGgwrUkxff1lCNQTP+ClSJfdEcTTGa+tk1eBO2t2
ehA+6G/h7K0K2LiXx/j2rWYvy9xyIWHK0BEVLZY72aY/Lo+EynIPq6DKBmvWSYFe
HDV8+c++Ut9zN0zY+bCT1cEeCywj+aPWeUCXqctIpwXpfGuHFpUj0w6F7g5l8IEy
O5BiGuKWWCMCxEHvN7BTkspeo4YVtCS7+fS23rrG9sGu9hVX6K59KZpmOGd+wVSb
5obMeNfIei7k6NVqfBAOY82/L0jw5ba91sCxXDq9zTeBsM8eHxG1/ZC0MSKTekGX
ept0r3f21kFAO517VMvNvZEwzsTAC4sWLjQ1OJFxX/yd0c9AOG5FXZgiTypCMBdn
ywkR4fCsZvGfYzfuI16eOUPQIPrtZwIMPEpgYQS8g1z0cjFGhbeb5RAWq5KNp7CL
YdhNZXQ27r2I2CIbHWmzWsw+z7gSZdJb66E2luM7tgLnj1vgFculX28pa9LYEzos
RVBSh12/31Kcx24DHxNaOQfwkqunUyxPqRuR9fwDtRoiAod4aG54LJDpoT3HAkYv
acjXvq+AP5edjo70GQvTkAVPCbyVHNqfNZKIfiM+KaEr7wfB6RJvnWi3e1jWwaU3
VPVtV6sV0sAi8APAMsUENbEbw93wTenIVNe4y5x4/T7ksuv2md/o5ZDj8t0yillP
X1wfgH9YnWQ+Il/k/gwMhXyNr9fly54cKoPeTwkRDnjYlmZyDuRyKJ2T4WsGHisq
kFWaYx9NogrEjlD6EYjpx8XUUe9PjqhzBX8PAER1cOwcydhu0pfzV4+N16df7m1x
2o0OOuC9qjei//Uq2bOrzFQ++gZR1lrkQK6ouxWq4gN/PPAj9NKMsI3hJ6WjhTCC
vdhqonY7yOfV+heCjtZmHdQhXm6MykFshmyBU0XmYVGqoZ79TCY2vSTPIGW4btFV
jR2APcWJjOSlUosXFFMjjxgocHNMFHdaQAlPjIV3Cj2FiBT5ooIkC2im50d0gRYI
1wwSaSKLwdjKT6h6/0dL/KopAlcZ3fkKU9oGvbocQDZ3VWw4ShwEtMAJ3a894781
xmSJ+MltjOGNSP76gFZ9zXVjd/UzoRJO5IhQCyA4usOWYdi/HNndOxzYWZ5cIUci
bLuJ4h/kECRqNer/CHCE5yQpRGq7GWC+WT7ZLEuPJ+lya9MD8Buw8vhje7m98KMp
R+dECXVnlDite/ssf698tvIE5KU3hoXgCA2wPQKC5cbTithDZesEl90dRoVlEN7l
0bqsCd4p5FORI4GGr8DMw7KXkyZMintDOKcEb4FVrwQ66k7kR3uRKJrnMFaMrR7a
mHWN6Hth3Q017dXt8pV/XRZRHbe2KGQMf6Kz4psDmOlfE2hWgVLQvlZ80y9arE3w
wn0vTYj46gk+b4Kjnk7/OBHQLgEH9IdjAK+bT9mzaeF8C5sJkIy+qLPJKTmA3NHr
AVMCB8Sh3+18PvOkzV0Lg6+aVuvR06W4yD6Mv3g11L/TX+1NK76H8H5KnUHdhZdS
pAZL+0U+sbEdpfFXE8jtzjw2xgR6/Uix0vvpn74AuwwsmFO5DakoP3CpauGoGvnm
+08QRSoFNjmvytIt57ydXySh/EVuS2EheD5MbI3X+57SD6E2KD/2wEZMs5AdAlw9
J1cMfuq63nPmHCljK16iVK/NbKT3wKPgfyzRW7rkLsLb90HTQk5f4MfkV6ji76Ot
8OA2zay0w8O19mrJl9fkQiCIFdAXUE86lHxdiybGWiteFlU4BHcG1Nl7YvhmYOC/
oe+8Dvk5hbBXtlOszi+YoSRpDEHPgBo0d9etT/S1W5F2oAOj42Yvo9bX4thDeMWI
BnqnZwiUGPVubo4/yLFVTIH88O1exPg90GZbfIvDanhqyVN4ABnjnkCYQLk+AmWD
F2anMMN25R677UlwnMB7xv1IMcXn7JR3g5ZzMvRn+RKXKin4y5uVFrnpE+QTX4bq
LZ5oUU200Yvz9GoXfFWt3D9+OnGXBmrkY3aIbKTLuJUTQ2zv5mv+R1njG0w9XtNk
vRd9vklWEQcSPTCy0c2LN7EAcTPdiB1jwkHchrK8DzwvKJRgBKc61pJl+LCfE7Xl
mN4eCFKEStE1gW98lzwuyHEwIifNtW0Buygu1bu+IGhLeV5hvc19HmRtlpyAMqRh
mrdYa58sf+KHd9PA7vpXm5DO8rmUqmPbYPiGlGcfn7nqxJcqzU/2HnV53qxd1FoL
dmlHow3ALisfnUtVXF1n1QTkJ0khPsQwy5G6V6wAt7IZ7hbZ0TEmqbgUZcjpmYVF
hQKLN1Ngz0oyBjawY3BYcOT+3j3OPcFOlMOKYFTk+hmybbqIuSpaCSUiYkK3bNxo
yJXj6iVvVmagyB7ClciS77yCPLoXguvcrAWlxcaHXoCgJAYhJp1JoBdy6Ds7tTrn
2OH4EghqOVxw5GWm433USFpx+zEwhWRPJlNIR2HYtCHKEaYE6PI+MRAtBKmHjVri
xUsxM7kqrsYvCGSJsAtMeZ4OMz/m2PQW66scWL8tIGTtOQyBftxmk2YNqOTYW/qF
eMgUT0cncIxmuYFf1/12euvpQHx39dVJsSUe5sBO8W1zx86J3AwXK4BtxSYgQdOd
MVWTIsOlm3bzz22fd+PDAKsJlzn1xj95j26KP5B6RqTGHzyVFyF+z6FZbw+7sUjG
f1oOe0tNiqptNTsSs739ggGUCk6JukOlNeUc1DL6VxzTUuNFAc1B3RjoaQTFEg7C
gftLKlH5SOcErBS5HG1ydjAmatNwBEwMRYrZZfMXaM6z1fEyUYVevBgUV23RImd1
HdPFk/ZlNvs9d54XopHsUcjSCwtdlRU5i9SJnJOOWc4DW8iafVPE61b0Wr++2/X8
oRsjqi73YvL3wXeWdyswttIk2pH2FRnpKpZ0P+7xqi0tPMq8rWpLzJaDCwRrSzbw
NSs1L6+dZAWs/MGLavwXVI1VVvbTzAH9FZdvyuPeM1TrR98ZV63MlW6hJa8HKExY
RD6wUJlzJtQmXUEySKeL/w+TIqgwX/UxCnWZ2gzw2eTUKbLZacROkHawDFX3DWRz
6fcm+NYEmhx12FrmcbFKoPFHkILTS3fRqV/IiCU+s6JB6WousN1CNR9ycgJJgfAi
JCBI+T1x01pOvdqWZ6pfTL/NqMVEpql76aTiaU55ciYyz61EKjugDwjHlU+HzrS+
RwrtZfFWLDVdVJTNQX3QU305dyfly8Ul1Q+6esKS91sYV1cd8FmENAlGBfjW54xH
i1xQ0zKYFIl2Z13FjvcuXqi0qpCRxhkicgMTgoJuuaOMxTBqksfj1l2LUtiSw3mJ
Vb70+1tQ1wjGBeH52vVGyRJyVkoPJmbssBPEYiGoMc2VMwTG9l5J+pqJRalkE+fz
5OpbNinuICIYdZ42SPHVcLncOXggWEWbhGhWRSgRgO/OssRD4RnDl6FXg5i/GQrd
DHwbgj2sl4IS0k0QeNZQmzancY+CMwF7qvyRrL04Ddq2XCwJT4q5h/ZvQhVUqmdn
G2eCxCsb+PpVIyr1I/C8y+1I6EuQBaz29QjZUW3LjlBdk9iCkXTxswxTkyFInli4
pu8tnla8oquee2z5GL5yVVDAcMD/6p0tvBWnS6WMzJ+k5U8aFhbxqpETLhCJoNc6
BWHk1KMMfYeMyA4YmzzPxcmHdqfXHx5Y6EpX8ErEY3r/obfSQeZjFJZfnIgsPo1i
bayxH/WtzKe/YFE3nlLllr4gttxiVA42Th55GkR4pHlmvExhTJdm+iU0muu2teXI
fRWS/28TuEYOM2PRgyoGU/dYGEX7rp4hdGhaL1jcFaQAQ2Pz6cNf2+T6AVMOzsDS
lh+McHlbtvu0fZ18oVtSAGsFBL9L3gEjISXS09RMPiv0wWO9eqGxr9T0Dml69BXV
3XywQlO5S4ikEQcKUr0PLGzk2Q6b1EEIxiFDob/QPuqI/V7eyh9zfCVmaG3rald7
9PCscuoRfguVuFxaCS0HTrUaeT9fGFeQj9a/gy3V/lM4aMtSvjD/lPO0JPC+h5BO
0nai4dKfDZOo7Ks0Bxh1HsyUz7zWizVY663tDhQhX9Qo1wEFFulDfrwzfohix29D
IVVImqu1MZA9YNLPJZzjWXan8+uiM0P88ll3ccB40ko1R4UW+mvT78NwbuEsISAU
OY94DGic3wTNwZdLY1pTwP2Tr0OdJn0EVTetjGInDu1RQ/f3ViFtAoS1qeamQ5y1
VXrh4uy0rHKR6xexoneVa/B6zSEpZ8uE1Ebb8V4bFtlrYN4+UiH6DeUxJN/2cBdw
T1pS+66i6qpY3pq1T8wGxqZqXLuJ7NLMxnXEyTBDr+UwlbDhKa8sU2gd8jcdS8kf
bmtxLev2U50wuQ6F8r18FpUgO/a27iDeoDXAzxzZZbVOSGWt26HRniFXtZCMgOZZ
EWL8U0qjWA1kwMutpeql1lMrHM/xbWVcGMngcONUd2rGpaHMmPgzosTtNkiCFbsa
N2yxHu2Aicp8F+kUEeP08kKLJE6D1wRhnHEeyPbx6NqQ1l88CapzTAp6kjukjjzy
Fl7qoS8PSgDT7OQM2RIzNutKzK2ujUdZn7PzWmxQ2Z2xrmWByv8S39RypB6XfoZO
ui/stjubfRNCW5LzU+OEfMaSgFxrDtaESGQ+xh/3ZXZRx4BkvxjtpGm7LR0xJvie
LRhq8FBrZ8ZP1BmmRMUcQrpVFb7KZAMR6/EsqpLcvzNEKDuoh0xlL7kuKxUCivXK
msC76xsDoCBxHahVf0Ct8syDatQjGxZg7TaN1eibXV/tIM6D6mmmatkGOLnxQIgu
hteheFCbujed3rBvPkaZubLAjpIs0dcuCRkrPywVx46kw/Vocs8Ku6uWfBu99WQg
tVPoyhvSQXlvIRzTEYJwG6VDF4srgGUB0xoelwHMoEfaJg4wvQF459rsd4AbxY7w
kiVlE3r4NRLkOBFDQT5dHSSDirQa+aCOdsvMGnsrZOJawxI/NdaG8ALWZVQ1gnIg
VoDA2av528xYLZgFG6POCh7ymSGz7x6BZbflXccjd/bp6iwBJT7u6n7O4lMRvrIB
G8/LeTTbBnZmGKOvTj2bEZMHz2WmEkjrxCFNk5x+ONotY96NPE+rN02pKiTDHkcm
DR6AKldnuBMADDZlY+BqcTokzXGPi03VGSkL4XVuocEHTz1xemcnKnpOl2TV8eY8
6HbNJ0gdrOyFOXt6+TL6WA4GgtsQ+tTcEef8Gn81UV7zzuPAYwI/5HH2y0W0odLO
g0f/u/4X9D7HMVwE8NPHH4XwdvKHRtkeOWkkLs5uw4btQNeclbfbymaxqg+7xNqW
UiCRCwaGofw1NbLBOmiaHWNa+J8WP/sYhOp8HHkoqLm181JGh5L5RHzE+/MvrM+8
vxl+7BqCsY4FcuPC6gHBNOUGMbIfDysjzmxht9tUy19txBDPHJBzVB8u3vjy7Ow7
fumvI2bNppJnXhojY579OdVS71P+yi7/kif4L5l6oJ/fSexUYffdEd4FhPvU695P
0xqE8V5UXumftqNQI9nzB6zkjG4uqx9MWeH4niXOq/WAJI0SaRAsQdSvUav2iga8
VQESqtupnS6P9d8U1Q7l+ED+OaR1ffEvxodubsdMfEqbqfe0dACQiWWq7uHK4N3k
dtkFZPtPW2ThZvDyBzUZw6QvqQfkAZOVqZe7w9u69AenuUCjdceOD60WX2K745vs
QeLaXdWArE72pvMcQPT/G/EWKLm5PxbW0321Q5TI0biLxOuHxOEryeIJVNjubrNJ
sQaWfQyRDChywtkW7HFld2x3k9Qjr4J+ofiST5Ep96o521x4QFUUsTZqFMo7pqKg
Tvt1HacxAv//RyBBJOlnY3BHkXHlsIVTrFA7+uMlUJbBW4MYCpScyhKN8rxw8Dng
5ONSfpFMRTIex5rlRXzgWx4/cR225lRQJR5xg9EB9KtAFOGR07XzI8i0gcotBmkJ
sVa3P3VtAd4VgGjo/gdVE1XoBNf9dhJ6OZRiOU77EbPYWuEec4TFiwFTjHo52ZST
gK7Go/Ty0WXa045BJiQXpuItS9UzuHqbbwnG6rlilcEswAzNb1eSyMdHSGjEWjcK
K2tW81NXxerrI6+jPDaYW8n/PayBcBKrBXte5UDVTtxAuoIzIX39RMt6Kiec+Skv
6ruP1ipWdILmd5BQtktxkfsViGqKQs/oxRfh/ecAa7GK2/4z753OnH9GWoTpX04c
+vlNkOuiCqmNYkxYX06/x9N+HmMYCJ5Qm7H35rJMWsDkkJ2fqsf4yJX8dcgy0pOE
a5N380fG6PXvtiG10EJqnf8/ximXgkN6N6QwwS6YCzUanhIQ/2zMRhx64VWYZzs5
Zfh5BvxZWVgC5iWUX4AiptXZQcXacunU39GmtCPTiBMshTt1L4JZ8zbKqaLnPt//
ynHCMQixOq1tOIKTJBfwvYIVxzYC1JZ42uiaawn5xQy6fxtY0nh7SpQAruJh64gp
BV0NncfSD8NKUz9ZnNhckx8yQdD3viwOgDwpNuPVbOMQActaunIquKeNpKGTRQ9w
yOkIYVsiw/0tT98+tg9POfva/kPX4SPBZGySiaYSDAS6UneRmUx2sQUVYC899rUS
gArMYbV+/1EU4W8ZFxIHf97/fwJOu3CwOc3L5o3CDOjSLNHcMsQsJn6xqp0i9YLp
78Ti6hRPkvN6dCiK51XSdqjXo4TmgT2SdQH0G39cwpUq6VST7MIjoq2Ix+009owA
Cx7hEUyq+Dl/eA9E6aKL4OsqKg+xEll0/e0sI3yjtuBpSz549s8NikBQsEKQh2Lk
4TfgnNeQApv7T2W5xdN0ONvbSxBsVlEhe/LhvjjhAQBZnPkn4gt3AMdLIWzGJzLI
yheMrA1/5wcbI6nC8hdeO7+jgn61SMDMhHPs+G7oZ/6AOspoYpkC5Q2rn1TK66Z7
jg+1nBhhIyAVovywkD52sBPiO/KrslvRbEDCY3/vyE0QrY9bhg6+AG1mdd7TIpR0
WbYOjqWbd5d+ikdAwihgAJOdlG46UVX6kxSaOZoZHSdq3Svp1caU6uwlWulgTnGx
8EC35N7JhNye3YREILMoATLI8hE9ULvpVF4iOYwERS9tk1Dhk76gnObOsnnLXEdz
vBbpDgLRXGKSyPdNJIE0grv/RZQzcpWlWOehzpAws+lETjv+dy+fFU2QfFux5Khi
3Xt1x4DmrlL8LGS8Mg5x/1venuR8hKGd8+HuoeHEER8lj9QaEuCAGEF7G5ecHH+R
SIN2EKROrQm4GAIxO5smmTrcvTj4JSPf+YE9HvJYxkwudQLUl032RZ6f/vyBPsXJ
N8EpSwdXS11hkJyaGreZ3DfwO9ykssLGqzZq26S7imfQ5LPmMuqKPM7/etCAUK8K
/ifPk9MrOCuQroC1sqlEuaZN0YrfKHP5iT8i2z1hZDsf6zw+P+jCEuBoNCzHKJ2v
w3LmQTDwItyIRQof+oUBb1g+oxnoN0kav9jAFSEyZmKHXHA7W026zlzaFeaNCwNx
75Fm+sWu4ju7LJ9hTSkJnqcK5IzCjVuqbKjtwr3lJM2irZcNk8lytlHJLvj2ILjP
V4R1zsZlWtQ0jrk9q/iUBwoA9JTRmzkM6A9lFMMA/KUPoxsbIiRdIF3C8rfgF69v
GfHoi3P6unl0grRoDZYUiYjcZ9+S5OK1HRYSBos4ZxvRacWenZrdKuHkTSD5F/pu
DbzGzxZvt/kGPwxT1nWM6ilhZfesMPYRJhzbdZYTTM1W4S3108xO2XMTp6xXnulL
sHJvDCI2665asZv8wPqNMuj4oXpVAJS+T/Fr+5uumpfpI63UjoQqjnKWpHsxtt3O
MlSFR/zepQSe9T3tMHbMCGiLAY70CKVA2tfb9p+HVF1B1JYuzEqdJx7dw1sj/12o
4GM1ReMoO0A8yR9ozkp/v5qGc6fpi0OUdQ2qwpzmYK44aRVYY3D26p+V5L5nvpc5
mQSziLa9ZfXa0AhKDbcixaPGvN+ziGxH0L2iM52Sbbx44sFtzLp9/uXaczH4VwiC
t6DIXpom4CsumQLjdBZ0pGIKSNI6XNSduSyn2gpVXQU8b8kOeCE+6eXiON3GU9j5
t9BEskHm+8V1my7dzoZVfFt+W1N1ewg/xHlVb4sALd2+RIkYAJXyWknkev1YPbvU
BM37JqJyZA77HK0AktQTtqIXRAa5PSC3s44wCYzoYGtEf7V6yGkwKYqAmqgH/FX6
JnPW6csjMeuphlYAJ2kGoi516i4i3XTmCBjV5EMpxpKSGb2H4XIgFmaXuijKiCfq
unBadoSvo5z6LfOc5ByIiLDQDP4pJsv7g3+pBSPc0UboIsGPjARBbf7wkbrX5x5E
oGfEJgI/Pnwz9UhjY4svv2dgxyIiuscRCHxnlf5ok3rqdY/copy2CqMjGAhycnu0
C8/nDQwVnY8Tb/6doysqKSQL7YyrCIW3GiXrNYY6keqVU9Xf4hqdwbzB5SWp54rC
/BSx0JADk3oHaM700yAh01V96gXT+2w1PnAwxeAqj5Rglky+7ovKC32kEJgmSb5P
FDR0O6SW2WRX87xJpiC/mCA+yRTlGKwx8ulWYNtAgDzPqhG4dS8XGndAQjhklH7I
2wudQrkNClkRp7k46mIrPM9S7V3l8BegyJmFJ3PEiIAHlkCbTP+cgdJnTPPckYMW
P9Ya6LwxAqJZBPHHGQF2mrWR7ZtGm0dkhFjNxQAFeFGzPcQgUJEKzU+xgM3s9cme
a8ZZKRKD2K+4IXmeS7BIRpCkGFbvpbJ5kyQU+wCzyRLHyBh3Y1v7UDYKVtTSn75M
6bscag0ELcXNpca33NzV4DNvV67hNu7GN09umbP9o6+wh5Vi4sJpfE26dFbZuDAG
i4sKxkV0ai//ZyCBTB4KWZ6b8NBSAQJnv+cwA476Tk8CGYsI0D+ti9OwQE+db6Re
d7XAxqwdwKEEmIAuVSAgYY+NUw+L5BG2xteLGRV7J+qXYOgBIJVvCkXHR9XQffCi
98aboV50JAFHXetVj+jby9SnAdlwhM4S/G5EBdQ4BdKeMX9XMu+AgFZ0kCINYsNe
bIKqKd6uxLsL8u6SHNjeHZAj+HqF+NZ+lwlDfcie1gKhOFgXwRRK0ySZfYU2rah1
dWKBppYiBOviZCtV/QFM/4gWMik0p4FwfQE+7MiihhoVirW7VjgiYF2Et/Dx/22c
I2PdRTRsNWshH41XQBveh3JBYeSzYSsdwpnwBIStXM3LSWz+e8mnWbSZTD4V5u3h
hjoVD+jkh0e9Lb23t9Z31ySJTIzEgjFawIClLoX58/LyXR3nnJy5vqLkpcz8uAQV
WolbvYU0XcfHw+kdpMoQ8AP21fQFqwO6WoSbgbY6WU3maeLyKzqjvgvCHoX3sTvx
SxGkek5pJbfujz4z61VYqSTL7N+6KxNyxUnRpWX4KJEjiUf+v0M2F+rJuzwn8lhp
Uri8P7gZ3AdkodQQIUaMei9uox5047iuqNrLVG3KQEJylndPPOqLcD2W1ZZLDqWy
ciXaWJseLixnvKullkeFYxK2NskoVuI6kLjGyGW+yg7YCjMIzbpOV+WOJPbKjB6w
iBAnoX/stCtawIGQXXVIaOiaFtdlHgsjuEj9iSGImo4vuj8uqpuilD+9VbAe01f8
pcd1Zos3oa12k+2StTCsPtFEekUdbeNmjwEmMdehSQlpywbfDuEvnhSzLGDXLuBC
zv8M3TMRJpu5BpTCL7mtCyMGD5n8jnCnyIaBpMmDVOz2fc9zlIJfkljaVy19067s
3YdWuGLVYnZSPJ1gNifot7eyoS/JfbmLD4m1feoSSMjs1eqR0C1YtqohLi1JxopJ
soBEXDD6/TR+kU+E7KqPZrI3xm93KMW7kT6A0sGmFbnjXinwtq301XZ7chutDH6n
uGzytPmRP/AmfefdsGD6x09CMYiD9dC4mnER/g7JQyIDK13Q6tv+zjCoGyoNYEV1
rMe1o4rswe2bLXiXrXXDrWarr3Dw1UtYXXg35sRGUJ8KL4aQ5aPw6BIWm2wuLPgQ
G5ENNxS+w6dDZMbIE88gzhHxwmD5CTFuemMMXlCwqKENVWn93GiOw3VejQ5DMSo8
DmYuayfzmFyaWphbHBw8jgTiQ9bHieZHemis3YE5QU3sB9nFBOgmXOH4QJBguYQM
Y7cPpZcEymys99VWF3cI7XvVcncxx9UUHoWH9lTydkK27oHMFcg2YRdAJcIQxbKB
Cpimj+3DqGju0+V+t3jaoMC3di1voUhbvJ75Grq40t3tzWkz8YVagVFwkej9t405
i/NdovaB5rgiSc5ESZb3eKfoganZSPV8LzWzOdvLevYk2jXETVW5IEYh1uUNWMeH
5VjIBVAXLdn38m50tIfYdLCwsTR5Nmo1f+Us4VPi1kGKBDZbQvclkEdxutSKkV8j
efUAODD45ZIXSFCqXBn9eNJ517NB9wTdYFEY8VTeBMVM0K/mfCibhbS0RkQw/pZD
XBAqoYvHitRAZb9rVbIscTzh8RhjUlFaNqhPszDiS8KMF4ib09D5spfFESCwQ/kO
gbmaWmc8TAJ+IkCdm7Wf/bvTYBQqunigJRj70EqYLf5MVY/actt5yONK4W/PgRr4
E14hZeqWdrsEj8vpmp9Mwy8UydOl9a48Jj/53iu287MCAhjyqimBMdAMEbWueE/g
vPrBNpueGXyhz4O4o74cQurlfW8JzGlDoJdsxZ6rjdI4x4uoHUgJX6GfIDjx8RnA
hu4zH+BQwKp2rbz6UKMMrm3PVFE2BLkQMwboHsPsdx/3WLkiCtVTuSQZtSDTXREt
AAKfpv1K6XOSCKhy9p6g+htgXkmktFlftLXKhoR/px8V7HvjtKaXOfGcpNXPGCDN
NYpKhtdQ5fMC0/9g61yT/XAmJG8Bi4vJ975vhyfTE8SpmSOV1mpEsGxC9LpYYrSF
CvnIFC6DeJcyjKFLYgPOEf2b7dc5ydG6t08fOykO17EiUrz3VnKvth/BqOk8GRsm
6QzCcw6gI2t5wc0qQQmSBG9xjPLcxLw+DTZFGMtPLVyapboHUjTedBRoMESVdyiC
rNPA4yL40iy17qzDAVyOGAQy28V6Ms3CxwokvXLFrga9p+xCbskVt+tDVtVLmREM
sRxZ2YBLGRMbr+yf/rvs5gIivEVTsSMcs0coqrcIDcPkaqCOny4GTNkXe52Dgl/8
bYdYv8/HZs7mHdAPYKPa4Cyg6WakzeG1F2XYsvSke/EMUkKo8/uZ1yavWn2vi5Fg
Jw9fsoLOdYGNEFZqpRnVWEgJ4Ydv+h36RZ4+bNK2PAsf7e1SsUnd4M9s/G/AUbZC
yw3WeaWR3IJ0YcGmyQNe8jTN6eXYb6a1hZbdLZE1mXd96zOu+qDGR3xZUQMKU+Lk
LjG1QnzncZmwKw2E2UhRiOBULFhXsxQT1mCDKs/hr2ggeZ+6GaY/yqimuedv3Vfd
/SMl6dsyFS6JlmgzT6ivbmZB1dnfAfVcW6pUU38ZLtroCHcBsDfo8nhkOYfOHykV
XG6Xxcp8K2EqL4DDKe0Lo0bFJfeSdJthne2a4dsEmHHCmQwSO1k/Xn4fNJ8Gq05U
flml+ZpdbT/AZQYhkxBHEXbPnJYDa8rBcC30B4eNyAvq6svVB7vbRo3Uf+09ZeZv
m/NhzDD9DoPvlyxgXVcAqVUr3gSfQ30f57iNMHYBko5TQq5E5zfoyASVZYaNOzri
JALQUiug+ZlZrmah7asZb0vxEfuw81FX7fmFk3bt7lBsOZ0Lh7UzPRSWY/E8WhTG
zVfEsrDywWgGQOkBLWfMzolMdhXUXy0z6sCH/dU98wjYACc1m0GxPwCIGojKcklw
/3JkeBIH4e+LTJ+UIH42LHDVurOjYxWfbUmFjTJrKqw9Ssr/U1p9cvmXlTik3qpR
4tN75JGFuKQz3cDAcZvVtbXRwUH1jezSc9hHXVv2nesEL6t3J7oIZqKWEkwhaSZw
43E+Q/JeE1vN5WcIh3PdbX/7xOxZXzc+vhM7KUEW1XZv7Z0zmuLn8TVfpkBYXXOY
nOBjN17rYPQUIB5OQO8/T55BXyjNxm4bykdYw18S92+aXL0Ze1rkwtvp9V9Hmd1i
eXx7ApTbe979t5uWrmdaLzc3/Y7iHcFHYpy1bwHFMg1iZmEsSw8P8tInGYeFVHA/
5fL5JM1J+YxDBd2RLMuFgp3ZlBscLuGxqx/Oaw4HihM1eoV7y14C49jIK+6JFDP/
NvQ2yvKyTY7nyzoofYe430NS7HE/xiDGTgiyIIhMPxWfPfPUo35qnII7uGOdADyg
h1/YLjrz4yN6sfYYtQJJa2FJPXYLriaMBws7iG9rkXeKI2Havj/dUmZK1pRZPCus
UV4WYy7ABrI0iFY17L8zt5cW+7Rb4f9w4FEYsc54NtBbadtVkIeR6i99T2Pq+ZaA
AvjAlvYvY1ppw/98IeGJeB7wBc9b/hHcbygK0Nn+wn5a9eBA6czTQf+gliTtiXCf
zrYHjWcNThHp6JJOe1TD3n+UlfMvaMXcpVO+Q/T3jxbgBUuujIlmmki491OPTv66
Zy1l6cHMu1Huh7BezQq7WYBJiCmnfbNi7eH8vHF0ZDUwQpIXQW733fqmwO84hhXF
IFSeJVEmlPjnFMvNpdN41wCghHcygQ1c0xDKP54oYkkP+TQ+T4g3JUNBt+Xqp3pz
aQd6VjAJzGfsnnSr0GpCzSu8Y+7xiGK8r/prs7KI2l6M+dm6bkT1C3IYGbOohJUm
wJZNOroiz/OS7iqJUO1AcISOAyai4ElBjhetDJA75837Cur+hs98lUIJiVLjpfi4
AZYAWrWR7d9hRk2ZkjT9aXIjXCC5PhcYV2X0/Uu6eTU3ZarZ7YpbM6Cino/P/SEn
BW1bXFDJCBmDe2waNgsxK5/EGAEzItIvF8LViH9BRd8EqE6zY1SedFD1FIHqBcfv
86rJI/Va02V3y8vbF9Ceb6AloFfiN4i2Bq2JlRXNCSXR8d1rz/H22o8WYs3c6W3k
FfPQXtpxTXd9GjmF5Gtzgrz9/4iiv48gLWKXwGPYqwiHa3fvZM7ldrSBnnJiSn56
6ZH1nCpBbnALuKuQ+vtIcT2gPbou2Z3o0pPFl2YypzeZrWtenuzDBCFXBpO1Hk2S
Mldg9wxc1ZnlSkEvfO9F/Yhz3DbjTB2BFzY/jJi2wF9cDgtQtXMdh0ghZI0UsplR
6Tg0mF7blUfln/z1Sef5K15/EwdFAN9VUoGXj0nbH6dTXfDPTBozOgo0rwrmzuH6
Sw9hjxiX4cWDB2vr+8TFsuq0dLqTTAt7BMEt9g+iJUthhKEBPbHLhftOrJRATPcX
bQJyFq0fvOzyAnfRyM6NXnagPeaSNeJtCiEQB5vsGkksc1p08xL2Oq7bCUR69jmq
mjCHb0Gte+NPYgWUf/UhmoXhRSCvYlULwh7DyMF54BL3jxZjuK74DbPXdiCnYpGC
cYOoCzjBMSU/mmcAhGThmYa5yA/A06ET+YrDEZosQbveQRL528ZapFeL5qnncDEr
y3e7IteWF//p+50FoC/gWQpNjjDCfX2mrOTIHuA2TRdtg9x9vaU/UOrCRviTP/LT
j7WvoD02oREN/5fKa+Bcbjl+NP7q8ir+sYSYEW1ftVB8Aig1+1VhV69NDPxFhder
poGk9kX7H1Ddo56UebauXS4d0rzAHcLML75byIl/j6Xq7nM15tYXLyLBKK3M4xMP
il8z9NjRRB6P/wbCiW88bY5UqA7Bip2mDlowm7cLXGqZWpzU0SdE8B3zddFwQuWb
8hyk14Uz4CGjVwu/OG6YaaDoe6FNXlbmcUVgnEVTFGSafKa/8DYHn6WbC267L+bQ
JwS+JxjSWQHr7XfFGyxFGqU94q01ZG1RPWKH07rOmOpIHHeX9PkwT9uH6SirWfAZ
1bbod3Xdr/3Fw0OPmuZx3ItkugJdq7C6/6QeD87xbWuhzbQKfHsuI6k8TYQCoHM+
3eWeU6a+xuJF7PeZCJq4N0OwyN79JI4WEXcFs6uN5vYAT1bK8DnGE2JEeske4OU5
GS91ADjuomuW3CPdttlPHoHMyNaZMd50mJCL5pZtMYX3oqX1nsgKrTnt4a5ccUm1
8pgVg2tVgqblXac+C1fLfmxfgWpZblGVPmxWNHpkiT2EOKC8muSsSuufmWrujvnC
glpbiNh40hnAzNJtbNxzaXu4FaJTXYzpJvZA/FW4D3ZlbYm95/hE7sw6TBev6Sbn
kI1VKDJ6JMOBUyIDD9S6RiwfK179rZ32RG89hVlGSoLLE8t8VQwHRj7+lU3ijA97
UiHvjhIHwphk/8IbkMFM2KyhlRCDqkiI347bCwyYGQ9ut5SgdrD+RrX654jFTLaH
o4WeJjb2tjpnYAJ1FpTYRvWYNUC3spdpz3yvuWcqJo1fLLUsF5D3Ousd8haGCwbK
3jvYm7A/18yBxqsYaSmUw6CzrDdpL/HXyiCppy/x7KiCI5FIRTJs+a6U/OOmpIcG
ja2QY604Nij+d8oRx/LogZ4J++7+JfeAuMawAfeNs2gFOM+qS3r/aKxHwn/ZhUNO
YVdzGk9uLgGiZ1GG54TxHtU1SbL7zFgL2oc3CaI4UVnAR4obQFPj6b7pmRTE818M
YwIB/C4TXfi+GFgzfBenANhbuYoSN7L6FX8Gd4JW5vYypUgyrnuoN2VzhmaJebap
+x1AVWmZDKBla9r1y4tfUKDzqMfHCfNGAk8Run5972XJQC8YR2cmLOe1izgNSp1e
/lapTd8ETC4ml6Zuv/Se4D+nGjQLrIc+IQhEeGsPOdRf+SbXz60lszJW+xZ7aVvk
UTeIdLbrSq/ujVb6+aHGEu5vo7Ulk/EVabU56goCSQQ5e1lmGIKs7S33tn3aqLpL
WQII/cJRDQs/5a2lk5i3RHF4VdLFlIb4pEQxKMpXvn1lLareDQy3ubHa2amVYTn4
qJvWB7t9rSSS+iqZ3ZCM72LXrjxKA7SYqr4YwO5O4e5q5OTa54gkU+l0As2xz1zR
gTurFQuscYlviRvKKDZ2ayxVHA1tRBO3tTGWJACv7vJoLlOG028P4PC0YIP3q576
hImMXNJ0THMnDji2Xo68pDkycNPMfkvnqsHyXUAnQ1Fe9ua0qM53yaNca2zjPH/x
UbL0f6U/2d45zSo3y9uNgp64Jao779FyVfOj2Zd6V6uZKJ4RCId4qQByhYOMCVR7
NtY8XOsskmvypKiEo7u2mSou6t57iaeCY/78ZqtWi5n1IPz6cen9xq20lfVvOYty
shasZ8Qu2h+hGu/Fp6sALu4HaypxOMAxr7mfd9vD6lPxk8i/99CzZK0YyiQzvwhP
U0P9AbfjLTvYOoXgUbwDA8nQ8Ja23Ion8AuwUaMggSxCxCOO0Cxb90OfWQ0ri6Rx
v7F0p8PfgvL7wB7SevDfhXP1lIjwdzFDqbai6ReJlXIdwn2S3D8zhrs+4EEYe6hS
VDsTWn3KQglgxYr+2ZqU4bII43cxL7n9eDKuolboUMyq5Jhw1h4R6SgEo1lieeKQ
MgVjcsTgGxDVO4NNXuqNU0X+CfgT749lcU5iMGndq2TEedwno6a27keC0vP4m3Ih
qh/0R+5T2doZ4G0JiBh0+pzB07GguXoUj0GaBgxPiumQRo3bT5dDVt40J/qZwXc+
nU42A2Vj6fl1PsDHeQcWl6zvzKo02ICMhRCuihPlPAJgx6qmdJWRA9P5x+EKPVhH
0LEacag+TwDuGE6bQ746ujDu3vgKWw5LoEefHb3JtB2TlzH+SohjCmadvmkSGe3B
0F0IznK8qVfRBejf+3NvezDVDE4riXJn+hyTDN+3RHuAVcTfEHeFZiERGIW2l7nV
lUkIjQGLRzUquwol42xPrRuaJZ5XQ136ruvUzEfi/fO00jQGC475g6dFfMud6UJ4
+BuHEPQmhE3DPyBaw9r0dKqdYprd6zDTbUACdEN5RZO55ssGcaJjamApklIsLHIE
meo2eN2LvXNgMiDHZvbzZbmOfHoti/zFymO9NbXs4wWG/enzCUBthKDJU7fgDHL7
iQHjlkIO0o5imPJsutGx6Diyij2X/LmewJXt0QAA402Pt1gas/vCxtkXBT3o8ykd
sLAT4L6dpYJS5wsW0EFrDTJYhsvp1cGhUBYTMAWxOoyeBscpCeIF5p6c99dI/7Fm
hYLgFK2TueWZSC6TvsZ0Ff+khyYTX6w/jrvT1zigkmpeBMkK9gpOh9rtnpq7i5PN
7NDyV1DAI+UN1TD3b8PKHA23mCU8+PR5CFsZD+faaU3JfeUHYGpD487OBjbD5O2z
QqyitdcAJlSVB9xTdBycpmQwpN0IoVz8bvEMPW1jei6FAxSWBSNIciX+ijJWTseX
HQw6CsI6mdL+zbJARHTizo34J6ANiYJmmV2j4xu1+sIMg6cvFSLFxZsg/0QjqOMw
v1M9ovlZ8ESqHym2rWaA8wJ8ZnCYjsQV/XxqtntLx8OrLYgG8n8XFQnqwzWtCfal
gDSuTLIGYqnCBfnHb5sH7QpHzn9b6RjUir7SXU8CKQFdOgxFTgsAA36n5ofKZAUu
fEz//7+YqF+/rpmDURJdjCbx7gbB/H3G+EI51u7bmHSyOwZ+rXyZjyvHJBibiATK
/CKLQTEENeAVldimJj64VKVfp08nFzOfOct2/d+BVPImeueTZ3kOYkoRFssyWGoM
XM/F/ZW2iTXiNWEDGPEDt9Yyyw0d3Jh7ZoUW20StmR7p8xrw3cQiimkTHNxrMoCP
bPlLimZVW2xc2L1b5+B30PqPKYcTuNR1FlJthpRcxJ0J3smT2Tho+GJ/pi7LFXQP
0cPJ8Fu6TJpm2/GiHH2q+bMuy7V70NHbRPZBc9uFGjaXdSHDiqk7w51+GNCXbkpB
nxRN+6J0+CcCaRqXn2xdWfZ7Ty0m37vOE+TGwTutsN8LKy/te1Pw0lSA6tHlASoY
RQZ1Tr8tCL0oXVTNM2S/mn13ALB0Z3pFHbm0IQb7W+SMaNBBETCPkQWqp3PspeGY
Bfbcauj5nn+Ttmt4Bgd9X3yVhxSJNK233PLVl1I08nDSp/xWY+XV7iPafE3d1KWo
NP4IY7vH1OrZ87p3ZX8mi1CQAnikWOaq99ATCTNBvqCVq3ipUofe9ESWfetqd2SQ
21CNpBMgoUa6ubDh39KXRvuQxeOg/vik+mAVkaEJ9ZuB0ouOxv763LFeBCs6V9+h
9Qdzhn5oOaCW3KxkhW1bY5j5LRkwcOuJwAVCjNX6eTCKG0sqhW4AACSv80IgrKmW
cB5yAFrj09yzuxM4LiA0h8f6ZDkeIn7pkkgnNgmlCwQjnH0htSmoh7XEbRY9Tj3H
h8UkWljWEiRf75Ii6pu3TEfjIAlOrIVqus9axYqHn5KZMhYCb0M6zaExU6Z5S9in
QBK67+0+B7d/XQfw3agl6wGpzjndq7TKheVb4sD382p/oPZd3SQIZTLkG1iaGQ1R
6CFOk5+b5E5Std1Olm9TJ4MRuOf9vT+NfaEujKE9Pf37K9OpUfWLV62RZ/Ay50XE
VZ0cIZjTra7HHqaj1Tlb4RqBaRV/eVU0la2XuBU6b+v8phjUhgRVkzZWVBnONRbg
DI+jv4lLUGT1dPH2kZ+BoPn0ZEGmFue9M3AoJhmzN404gunVrYs4dMClY/4DyWvs
b5eE1VM8jRvObqve8aojR4qu0KxuQSEztZg0TdJbOJs3cqbMAq0p+a0GlBIaVq2K
9ebn1jDo66a74lrbwEZSf5o6fWUTXlXrRndphwJ5n4yui6iXQ22toblu7woobHUn
8wskjNN9FaxLqjVZWH0e/m7zgUZoUtqpSiBBl74z3WdTxvJPvVUPFxm9qPoZ//eo
blk8vu/orivAw/GfdR6Hu9ewMEwNlao7ECFpg1PBqi9khAZtEyv2GCfgAW8IQI3s
L82eI1tz7SmvBLPPAP5AgoP6eNt74zl/AauoRNZBiLw3t9GfxRrncHzO3+wqMDQA
JOnE95D7wMxmHMrM4JRWvQR7dWXzqSZ6gc/Kye/2rWYkd3qmzY8Lq5JkRxMmy8Cz
H3Kaobt75ve8dbovJ6lVC71/A2pPwx4oDJ36PbsIwBa8G0LTkKdn6oOozjyomVcU
CWWK3UZNSnuqRQ6X1sX4qvQlhorAHp7xLl0+GPn1dxruXBIu40K+q9s0Vwh/IPoF
o5NJthHrb9Br50R1GUcd4AE4xz/7OnKpEOXDze/wigWMTI9kRjMbXCGWscFsPizu
WIQWPokZ/jPzyF+ZLsBqgJIgryDdU0un5bs/gSi4WrgorACnmIhCdYbMnKNWgpxV
ZotxBMRMtOjky4YQeK9YqrgUmCW5YdcpBiGJX9RLgKjb88ifGSf9YZBOdiGf5zOw
hSOT1IiBaADtJ+jyIiWYdBazUIF05xIOd8cz5VrSwVPGstX+FNqLFr7KTFpUVlVe
WEplw/QUEsU7ddI3IrvZKT+pj2QII4jW2+13RIk2CPHU+jPKjhRwKXLbtPjsykWf
fJ439DQ4+1T1x3Jfep+z9WH+WhVwtLpcifdLgzCunX1zFr7YncyNnZdJCZZDVJ2R
3U01iGfIwHm+w67Vm5PWy4bzL4wYXCx4iEbdSd/f9DWrSgiCtYZm789oeynTHgTH
qfVziwkxYt+TBsUAXTLJKBGFvXSHjH+2eBT3ipyc5Fr2IFZ2tnn/jqc4zmL+tS2n
owzIY3lMLzYv++ekvW4gGkAl/y3dEMEP6L1/xNMSDKhk8VZ9zD0Tb7D8jlhXmO7f
DLmvVB9tsvxXSuFEFXyzlXI8cA+aF6fm8u+yoT2crMcOCCICLvizSSRSOmP4Pf4U
5Ky2YocWDW4x1xRt885u9W48yaDy2cggq5VagmgHlKANmYapZmq7QH2mNIV67zgX
XtcGACLZZiAIiVPBSGXlDT2KmB7f8CSQVtSLQgq/Vv47mbsU20D4AxwOxNKME5tW
MxMelU1Eq9qRJluHxeA2aajCILnJPT4KDmXQF2NdPa5fFVEZ/SlPjXFreXjgtAg0
BDVvodAQOEMtWScXNjbx8gNA+ovN5yW9EcLz5Vd+Og1y3YYY1VKAh5XBHUh17dT1
44rH6CU/WqR+zbdhDg/LzFLU+ezEGVxNshoz5MUQNydPAaPvcsMFQCzTT/X/kv9b
76P/dES4hhpDHlzf0yDAwo+onvTQ4326hOP1fgeaPqzt1gfMWlFXFf4kB/TuJzRo
78MIKL10iI6/I0SOAVPCFW0gllCa3i0wtNiVrZ970p4Z0NbjuqbIcXRq3XolxyLU
NfuzoPntAqy6wgkVzaBEYP19V08+EReGKDvtAln6me95I4k6E6CtlCP+DgU8wTrM
obHQ1p/uC+TEvpXCzB0JztMx5vZvUxGALCCGChpxhG7RI0hk9IQQ/8alSc0totUV
RXVUOpGtFg1IahblWrn6dcvaophLH16zijV0Sg/hhPZcU1HV7BXYln5RJTTggUYn
gHFYT2s1maSK2qmtNePqantfc7+jQVgpNasENI5BmQOM9k8OxbjBfc4TpvbiQQrV
xyOTpecNPRUh1FphpOE49rBPEBsoCvrdzDMpJovnW/BfFM9QIaYTkIDtQ9iHbPsH
YbXA3N7ug4Q7O79NQLADfi+8sJhVBXQxFXkiU7Sw+g5TQXlwXBa9eGfcGaBuHHm3
+1BxDjfja8DMPoSiZkNsCFyjXQfdk4jT4rpEyM8FsaP5ohfv5aYuymoO/wMo3aA1
0lC0T/TVAD7QWjDHvK0YhhozfCnDt6ifXm4o3cuMGAU3f5bAmhBSHeLsO+kym1Kc
nmyF0HvPiE2yBVnnJxZyeQArmW+5Ju51pVcvPxrm9A+yx7ydZEGe6YVfB5+EyWZi
riQ9XoBsHnHdeHWAiQQ9wxgsOrvQ0iyFAZROvqU5LcEcEWL96uM2330Wh+tilsN3
0mpdHpdFlMNyLbAHm6/0jIigDzcmw9c8s/jSUc3efjKdJ3LhUPtXd5CzidtdYe8c
l22n9bjekbiZ7tm6mm3+306qr9jJB8zIF6bnAcxk5fFXfdwz5ppF10zZYwfBKzzh
a8tNXH3ZnXC1wVoP9oXtQ5KhOhzqUIxle9dy4mtYT0hAdPQaDbvDOBdt1vyPmDTh
NPZYwTT1KBnplhKg+8608aFR6SeV0wognlAH3VmdljPqnJwVDz5EIxlpySzxvn7M
qw4Y+QZOFSqt/MUHnWXXhdyq4PqLA1qiEo9XslG7lKmBOhQVbkMOGygoAmmwIya8
3RMHXSTqsRAJizrpMrEo+GoEGstnfNuQi6Uv+argF4YVMz8WHE7giMiZKIJ5texB
wshsrxndmwKHjxFkzCo1cNzqq5bzorJq+iPSl/ctTwB2k0hXTvCxoEeqmP3ifBb+
BPyQdakOR56Huttsc3d4Qb49HwyONA5R0Nk+GQF6HRbGApFpYspL6W4zDX5Kknvn
vcg5v7StA+X7g73Cux7h5aRZfq1vY/uIsMutHu5keXxFD4UNmL3MlAq4hvXvwv8C
xi4Hr5OzjlBToZlxMebvn3pEsmRioAAVpSU1jnpIirZYl0cfBOtm0ucObYUlCHhg
ma6SdSi4E3sLtKmFsUHus8iqGTkHuyzG19XpQh1eyLsdBOuvk4TZxnJh/Jvr2PxQ
sYFDDD7+IxkQa2Dmtec2969jC8ORxiQxTfCBewUCabPzXMcBiGVcvbheasM58xMZ
YGCwkw6IoSgNXEXHUevg/pyV1r6Hnbe/xsyhrClaUV6oQU7YLSNfdk4upFbnZJf5
ro6Xo3EqdCSRDIH7AizsK8V4MQlmJEAiHULQFmOPohOCi0qQeOZtf0icyBW2PoUL
LYbcXTzACH2tdmAqh6o9j3mlBboQrgAUfJyWneCsczFao2Nb/4uRnXeXumtC1kNg
SVr0/Pf1NOO3Lf/Fv+OXv49sa6Lij3t2+axup/UIj6w/H9RHnjndzfzTs8OrxK7l
xW173zkUOorsNKJneF0ovX9jLdKBzJdV1Vf7iq026Fbu2a6xY1XBPYA2I8lU8qaf
2Bk8wX5xmJdThSQTGsQ8ln/QncSenn9PrvYtiVGm0065GYg3I+BPD4lsRPJcyAqy
pBSTxsmlusT+ZdIJIxsdP9PcuOfsdnoUmgythKd88y+Uj7PKYg6zCgkinid6eS51
6oh50jSZd2PZHHgC230nlqMa9pAyB7suGBuWQ1QP83rd84LGTeQo2+MIil2M+evG
o9zZo6pRFcEh4B7aLe9x2MjaOlVkRTjlks2Rl6+IOv8aGwg/aRXf+SOlrO1LAFNB
cIylyiQtifhYNrWVdtt2/Clk4AXTWNdrEDYeXxMuHyuurc21VHHpvpNgRkfaE+vD
MoJiq1mo945Y4fmtt8Gyqdd9KD4iKMd5mhFEZAhkL4Zdb9ZlG6o89WXnj2wh8kj+
vi/bgdCApBQHPIj+OVsIxpl001rSDZYMsZkHuwmdU6xcRclYpGgyX5aJYI8Y0XYG
w2/bKXbWowcAc60ypOcuhS4QM5f9YRRTa8nz2xPDCVZNYyKweR6odRIDFcC+TKAC
cHulM/GiAzafyw+nYeTSMUSEhU13SCo9zj19ykvN6JNUSRPB70lVzSdi8KhHRbqI
IwibvkiP3OQidbmTLoMMIwkE2FKiCuNWZ+llqgR+nkOnSe+GIqU/GF7Y6Y69rAa+
HzmXQjCWjiLYDNQbVIKsQPV8Cv9xGUIOkLRk8vIP1B2Hb349JA5zMReRn881nTFS
R9T9QRvgMgrKXkbIYk2tI/h9hQKalZpFi4v7J1dbcrhzD9+tiSfS1eefAp4cYptm
epzZlBpczNLdIv0D6wbldt8xKKwhVmkB26gt3DODEzFf+SJBdTKGAG1RK/nnGVwT
d72nAb5qaae5mQojFbNSGV7v69oHvxtDmczWKBU1LtTZdOEgMYhznFd1wgrnLsPa
la5mX9gxxDrZcflSf/0fdomYKCTdEkI9nJEkL/R+jmV9dCHt2X/kOIO4phMS2p5/
DdluUV2lWw61y9Nhz+5vg4vZqUFjjMJJr0YZLzKAEStmcRDyLosicmmwsY01CsO2
lUDPkvWHEj+OV+zSO1gmQ/2j8g82AyVJvRYfhaDW+qkIZ5E/Awf9FsKBBQ3J2Z/U
ophC1CIBsWLIqmUkrzSrIsTcyGM913W83YNRTcxuTNIhYSbvXC2UCfV2B4Gx0Nez
P9A1HdnKYmJhOFU65VxggmYjAOyPMMDK4cJeosdtjLzKvo3x7PfcUY+vC/73M3td
bkB5fY/6PvosaF3VdOtID3g/vrzItTlYXMU3szW4CHs81W7UwuMuPFUaIRSoN6s7
o9O8N4OkMJx26hDS5Qj8ekpMQbalsGmZGHUVAnc6HJJxV+uTs/r0QTD3xwqQo/NJ
qjjOr0fMwnYsS3106C8d22qFry1AutYuH+kVO4rJZGMjg0ikjjgA/VxLPqLWCQ9M
LfEt+DbVffP43dqi7ZHqbxoOZl2BgT3zWpMj/f0NhGwG2uTnXb8GtAT8NhrRixkN
B+SVCSZKZOBJKfJc3cu8S5WgjlWX6iYZPGpLQSfOXMw4OXqPvl9P2PYzEfzBqkUy
55vhfpHjktJ7cNjLrfYJlW8BX3pzzS+1K5zKHKfn0LjbfZQgtv/uVmChGdwK2QMM
c3dY32pMuMXURu9O+PmFA7Qa3Pvb0UyaOOMPAk+L/BzwaAjqjGjvC2etH1TGu2Hn
GFab3Bw9Ip2p3m+hGJTamwtQAqyjTCmEihVkyX0wP4y+ri4JdYwAYVrwOODsTJj5
wEj9nG21xcBwbb4POHdF5Nwa4YjHi6dXrkKYcnmjA3oCj06s4DiFyN8xkMLVlyAK
lqFQWi5VquOGxCG3xMtZ7kDG1vqL7Aa4hEw8PeqRalcegeqY/Q3cksl0TbCW/Vkp
pZa1mOhI4EhAvB2YVP9Vv3cLKWmrTM5s69j7xFMZ0yfEASJZChpdYQ2AbZvZDn6Q
/6cLPYCA9bx0FCZxCVccXuCAW5vLc1syU1rHgb0wN6D1WfU2+8/YDRsI7EjDvsKq
o0ypASLZB/pC0sk1tQTkCahcI5+8cdg+E73UAS9oW0sayJUhyDr3m3thqSgSiaTX
YLOy3EiL9WTwE8zXy3csBgNoroyehm1t9Hu5oWPysq37uf9iXGMIxjs78rM0ar5+
Tc3c7l3ip5pg5nQvSnhnwptXxTyHLIqIZXTzTwidnhP7UcvOjbt3nDJVsxOsy7/n
Q8iRrSG0rNOLere32ykxCrCb2VNOeESAlqq4JV9PRHZvEkwAiXamZq9hUeg0W1Zi
Etpe9hSgzRe7F+iOsRTDr9/D1+5ff8bvchLXuKwUSoHJL7rh8DBues3vHUl9mZDy
vA7i0N60GF/R4Pz8hG7jytZxD2+N01UVOamxrIALfG6YajTwKMCWfsx/ViV41rPl
HCKDwXg2pZHJGU/o4i6HC4q/7Ud8+O1zn2joN0MxPbPJV+/MhJosEMCu3hfz/maO
gIj0Dn1ydqQRVuM3UI5zI56QCvTyAxZGcBhEE6xazoHfiX+FmMwuKl7peTIgqvxf
jMswd2GSAQp3LvvhFw+ZldZEd2MhbfKEFKdfMeoWvEeZL1lOVdlceuWa8rOyfSOg
2cXy+JmqDG/8yznbIS2pkv6/peb/lKskCl11yrFS+nXxV68lpKFvPphRNlgpV2uo
OVPpUpm5vwgilMyzlUJ0cWA2d5X967556fJQ0h7sjIuk23f6g+ZFifOZPXEt+eaD
kxGdajhH4tbyfMchCRjofwjaOwM1WfW6YKOBXT+7bAsa06oRN46wF3xEgojKjbhX
ljafBwwp8gAYY0XCZVme9tUtVtVXJDds+OldMILJCX9Ch/OFfAH5Vu5Li5tzTfh6
eCLTOrLNkgZgCl4uz+FeuGlfZV5OBv7CvRv9nAnH9MkHmO58YfC2cbCTTdm4/qYh
d1PFTGj+nomIO3QO9Ql1pJ2cQy0MLnlaP9OOe6Kvt+7zDpdqeaCOL0oTOSS61Jf3
7SsOhgObuqhEnivhLguph86x351MMRKcmawGUApt+76yK/woZpxx+x61jJc/1uh8
ubxaL+t+/o570N+6erBm7XnPgUeTLQRWByCyzAhMDlG/WVLh5Uqv/M6YvCLApuDQ
mPtK9Mv+yhPbKBt5el1r1K8++ugi5uaZ0ip/OJURP02CH/D1DkdqUEdnSG2N8ckI
TyDIYvZvAx8ZwEN6pjb+JYvzB/G/bNbW4E5rifJum6vDip6zUOp81YPUpqjJFA9Q
zYf37mtsRCmn3OsoU5jVPTc1xPH/tdqyEIrYY1VuuPvIehsMcsNJ/lBX0WSK8soP
lAl7PE4crgEaPx2DuLFkB7w3msTPdt1xJdeCZZIBV3eHxZVUp7dfm0/pVUToomMW
ba4FP3JB5pPWPhJbOieYsHwy0K/Osg4lDJ8p12qiGDhGVGaZFiKRmaiFIu4UsRbK
yt4ofMYgqI7IsTAi2iLyXLvV1Bb++R7f1olGdKtskrb2zbPFm7fqjNnZmLS6ZB2x
wFHLN7UJs8x6kXD2zidSE94B9vUlTYFyY86pMO/5YWkCUaEnfUJoPIBjd1thV6re
M3jDTLRkAHVh5Q2vIz8Q4htxjUvCZ7ty2hi3brHUBt73UBGKMnYdEIoQH3Xrjc/O
cxQMu9K00pXLkxQFxDNtLc+qwakOQhcVL105vkolAW2n5SHY2tBJMMkPpcMPSoyd
qdQcS2EzscVQjN53PbFC1QYilpspB7pTBCMXUh9hPxtmlgaZMY4M9Y11Vxgkbv+3
Js3SIPFdxaNKr4tCqw0ih3a62x9YaOvBJ/Bf1sK3wRrLr6Wkr5w5VN5kNqbPGrUJ
SWSGyi5kUU3v7IhghrFU8vsIL3uGQ2J8KfEWH/Nm8q2WKqShaf5H5miVuxKzL8U3
Uwb3m0FiKInhFNFcXaW3ufS9eExexwPA9BGgD2vzRZ87C3p67aOcJ8a4tNGXi00o
MqAA4Ah5iGf8OqGrQ6u652CPSE8xv8fRHHxsbqUplitp3s3SYEzXjJXQfxkTB2aS
xJObjucb+YuOeXBQdQK61l2Xe6fiVKVtRRkFov2exRgmGQBql+eVJosQjNnfL85e
JLJyKaCelKBLN8DP4Gfd2Vbw5LqaNm5SsldSlftE/Klgt05kv0FZJMae6J1Vpt7W
/RLtfjbQ+xa3PaVmzpB1cQfUukLJlTtJ+NzjavbM/fZcjqGoWprKJfFLQ3791PsU
mrJI15ej3k4Jq3XCvkMwSQwRAXgkgy7HwV2l7xG0o3fu5h958YAAPF0LOrOF7lyE
CjxaGe74rswrYfrMEf1UoXbRWKF29CufpOOEthIdf1lRfRq39YLZhuHyYpe1SHsY
JylAM9PweLkWM9A930XGynXR/XPNfxYApsk6jpGRL/244OEoApHTTXwYEjylCLtr
qLONbCJcY34uYaE7O2RTJbWGEdS5jxiKJPXi+8dyAmi8iiPaeKussp0AYaXdRvCR
rV68LN8Ii//yDlINaM9uCwaU8hr5UTBn9Bvv/dBcFBm02VgXU9I45f7+hTRHidHV
zJEBDIBWLt3GuEh5o7LCVLL+QVPQ1Dck7y/PIR+izBuW8mzeN/2RYUPJLSTPw/q9
PfMlKTPpW/2YyOkPbtYl4pIXw0w3I35uEiQwGpND5jsz/m8owMRrMaOvi31p3djL
VTMqevgrNSqW5uKxs6TUYSWG965ZElV/f8+ALxlGYsxHA7tSKWtYgU5ZZpreWt/F
pG2ejNEqLCeYC8hUPVxF/EE1Q55CtheUajA43R9XjuwgYjSEZIzNzNywvKBBnFgn
7hopzZZPmxoWgAQV5dIG378JatQj5Ll+FC11URjYHSfwwCLHmu4IUxer+Q7nCmnK
pW3rEtaj8LzMErDH/4YbvLKKVv3ru0yR+esWgGitHe3GshRotVMsnsepPQ3/nHxT
dFI13jxtC1H2aN/i4twuxoOjbPlS33Ei9m8mpp/LACm/i81DpXOU3NxWkhwr9WxT
kJiMYZNJwUMLYcNaq5o5IcSlwjdkgQbEnPoV3+24GUsrbwM8N3Tr04eQqjKq/JlX
M7PcZ83ym6mHrYtoW6jmpWEnh2djLWFpq9ue503RF7XHPYDXei/ufjYD4mHZnz0B
3ikN4mdteHL8H+XBs/dDp+TNPoHetw9LY+GCfy62V5GQqxzuv0f49bc/YWbY0b7M
yzEfwIsPZJWiTM+UhW6dI9ugO+Wuydk2F65RERLDHakEMcLJ52JevEAYmyy7NXX9
HOy8DwqLfyns0OdPbCi9BWtYSBqk4xsp514J9FhbRu1Swo8cevhilZFqf2WkfDoc
7NCtCCwIeoc8yJWaJcR7xzSdYVJ2/8lYO4fd3+P4OGOruT07yWIhD4JxmE9jaLpv
esBu1BhRHIs/EknDTUlz+DGYrem9eHk02bT+ye6P6Qe436yCQp0SuxgGmYZ+Vfl7
H95epQT6awZxY/6kYkytGMnTzkcyF/ba8KYlqRFPu3nIr4NxqF/VPV76s2B8hrNK
yNSKJwgu2162QUxAIw7yazeIlXrkxWEg2ukoPqiwL9oq3g46Uep7C8dAZfCy7Rg5
CI2soHk17/sk1G/IyX8USfB/T8Q1YloTM8QhtwkQITxWVu2O9c/ISUw5tk3h7etO
QyFQ/tE353AcL8tQ6rZasroVvuityyqqREC7tep3hIfUuXxjpfSPHMUf1bZmNDpq
hGERnK5ytUr6IN0RMMXglBRwYSsiNs+t0OFSDK5PuM+wzzVHZ+B4vFSwIvrTlqw+
RmA5Kv4ZCze5+z5Db4jTMOEY5FuyfEz6QscQAkqMweQXCZZBErGi20n1GEsFouxu
1SozFeTH4uM8Y3n309xi1GPbvPvME+9hh4/ya914voScX3NJxbylyRI228Bj/dKE
St7MSqLj1gvIZuFjb/LTjuCqIDv12CJi7iXcPNAn71QFlaw/Y5BK91vrr1VyyLI8
pDASN3NKaSVCoGX4EI6XosQESDatxWCDbhF70+0c+waICbnUzJiiCnOSbE6VSfgN
07+Xgt8yFnRjhxfTbc4dKkb10afAkCYoNtH7sVOqri6SKZSiVGCncZ1M1Gh69GMy
m3x/0pbSJMJkFfNFGpmpBI7wGZF9wEPABoK+fiDRDAw=
`pragma protect end_protected
