��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)���vG4��NB*v�^%��_�rG�v�2�H!�W��
���1�c��J��5��Ż��Y�c��j��R��ua����U�T����#2������D&��H�d�o��9�4R\��W�g��1$�W
b��g�
@�6G�U_���Hૹا�*��j�r�	�˴��ϩ:a��<b
NpxL�i����8�VD�ʏ�P�
@���M<(��ă6��j,�_���_��˛��a�ӝ�6�cU�B	��ϻ�#��=/8zժ3U�j�{*4ٞ��t�RX����]��c/b@@�� XĪj��4��i��]-1���}zYk/�߳�(`�s�d�R��H׍;Z��C�Y��O�.�,��@׷�%�Q��C�9%�W���`ed�P���3�_���c�m�-��g���n�&�H�ƍ�X��V�����]5���`�[�I�E`�P��>���l����*P��7G�o��q  h�B����K!j��}lW�ώ?��Vĉma^?Ur���Rf|�~����v"i�����E�ݧ����W׍+3���3���,oBK��!b���0�������'�{���á��Ó2��I�e����9�m�:`n��>^��J�')��5����E�T����T	392���~�;�?�����Z�ܹE��N-v��d��;nϓNԖz�V���������>W�r G��mFJ�����`&XRC���)�t�n�Xģ�Ƴ?u����������;Cݬ����*<u�˱���N�	��!��m�7���� ��$M��T���6�+���7�>l�����I�<N���qw��޸�9���	i�|�I���!�(Wr�����|�]g�E
�nB�5Hw+��w9��ec�%��%��e(�2���p7�·��*m�9J@<�ߗ�*0&�����x�S�[FRV�����&����X�F7������u���MYK����L|3�����*H�WS�RO��b`�q�0�ɐ�6�p��q�����u��T����|.V��m���Ѻ��r^��I�p�!����}"A�!?f��������᭲���+�б�o�IA�ጏKA�q���tP�g\Κ� �+<vj�!�&-,1+Di�D=��l�a�����	<��QC�[���
�.�3�BՍS?���r5�p���-Cb�xM�u��:�X��#�1��{WR��$�%X;4Jxy��ê���n!�'^�����n����=Rh��	���ڣ���=�P�_��v<����{m햫
������=i�:�F�}A�K�΀u89��0�ց����=B���7?볬���e*�>c���w��?�E�~�\���u掔�p̍G̫6�̳�f�T$�]h��+�<B�hH���4�K��L��)M�Xގ$.(i:�&�k<����Tma�<���JCvDԨ�Dn��edT�^4l�+:��[h7�vG-�PՐ.x-�N��[��xo��֊�e��_�c�16�?�����9�1u��W|�t���G:'~C�f�ʏ�ha��haɘ�����-}��-@���l�m>Ny���/Bi����k].�c����u�%;�R���H��n�-�>�VA�P#���/{��Ɍd�DBl�W{l����ixaqr�]��`���s���$���1cp�

�)��2�'�o��s��f��?����6��] ��s����,�����&] ��O%ߘ��`Ik���z*V��@���R'_)겾H���]�o�=ȃ����E�	�g��+�a�]��<��!������atU�Q�Ѐ��K�49��fyx�"�,��f��.J?oe|���%GnbŪ��~f {gND"-�oȢ����3Z�<0�V	T/!� �ʐ�h<r�LR^_|32�z�<
gd�*&��S��UD�����Kٻ�����1��?d�@��9�m��w	�MK�]*8U�����M�5�7�Rrg�x�r�WW.��-$�R�k�W)>�;�^�+\����&i �`&��r�)9eS7���Hɻ�;
�-��&�XM$+����<d�/7�1���I��uI���l��J��qq�u����n�Y��;I��i���K[��&e�c�����S��Ş)~���Q����pcI��p]��Z�6:��D��"C����%µ "w>�|�n�����jY7�'~�(�#��g��$�̦��~k�A�y��Pz�Έ�kay<�������׭U�K��p�ݚm���>"��Dl�`G�f^O4�c�M�
�.$63$�(�!��3�����L�Lس��.Thc�<Nv�;�g���4�劗䐼|�~����gkKܷ�W $�f=f��tě2����tn��R���xr?�WE@�c������Z��z>z8�C�%�Xi�dx��G�'�CN~ݠ�� 1h�V�=�B���)�D�K(��4�O]|LyL��rꔌ|���^H4A�C�x}�������P����_wt��f^^���Fv �	�>F��S+I��w�1y
��	րHu��K�%�c�.����8Y�F?�k��x����=�tN��<�Jm4��[����~�Ɇ?�BB��>���hI�^���b������U���O�v(考�l��_4�I~����\���X~�O��޾��j������9�̣� X��˽0���k~��(�d<���9Q7�(��-Yi�S�5<��ѯ|���;��嫬��l�`��Ւ\4��#-��ޟ�x6�/�8�G7~kc̢�t�x"c�����3j��UT������Ӭ}�ϣ&��&l|�?k�W��`�b�{�A�R���z9�L7��"�s)}5F���Gjl��0OOD�d�UW�5B< �ze���Z��5DD͓��Ӿ1�n��[.뿾m�R2c��J4�ռ��t�O����{-����7�o��p��Mr���������n$B���+J�G�l��˦�'Rw_joĦ�!g1NՒ��<纆?���j�
�U0Ut�KDI�Jf��o�� ���O칼�t�T��F�ܷCU-����B��XA�"��bɽ��� a�dF�a��w���ms�B����3���O����X��$��(!�1��Mļ�5�/�no�wk[w�Nd�2O��A�;U�����<Bm,�G��XVO�h� Gw�6�wF.��Q�^O��>G
��+{.#��+e�HX���G,͠��b��1��l����p��Ae4%IN�����2��B]���l?dO��.�쐙��m+}��R�~��Y�%Iq��k�o>�6_�˞�WB�W�!�۾B�ӽ���q��Z���� ��2�Lۏ��E$�2c�l���F�B�����wz���oMF	Q��z�U,��n�$X�D�	KVa��0��"2븝MZ��*��S��w7�W���k�����m� �EDc�
B� ��HADt�כ���i��p��2b��ԯP�����cfN�_�1@9]�'��~��^q�wJ(�zt�F,���V�v�'���j"�J1��B���/�޹r'����_#�c�'�y�w)'�{����b4$_ͻ��n~|޵�7X�V�S҅��ۈ�[�b��`�T��JC��D�=�D$�M�����VF�}�Ex�0�f����y^җʮؤ��XZ�FE��������MFW��m �3�nG�W������b��y�	�}B#��*�}�ϲ�ó��L�S)�Wd�,�l�?�#m����Q{�U��jh�d+Z��ύe0Tq����P�l�-��PO[~$��8�}ګ^�r��S�1�#�"�j�q_j�rg0�۵�@��Dy�Y��*��M[ԧ��9yM��P%����o��}?$]l�R@�$�Q�j�׾��
:A��vT	Q�6vW�����$�!}:��v,�Jz̘(�c41�n��N��kB?�s�K�py:,��O��ه��=3�*mI��5Aa8��h�z31��ax��d�g�E�	2d�aFH���x���g����/̣V��Sb�)L|M�%���;M�U�}`�?l�n����*��{�|���JskJ!G)2�ɫ�sIk=���B����$Ɗ�f��T��$�Q��fR�2~T�/&i�?�a��SL!���G�ѴZ'ͪG9E���|Ԕ��`�@��_����4�v8���MCb���q)5�+��l�_���^���'��D��D���� ��j���W���W�
��G�w�C�L@���X���/M=�q��~�mG�x5�z��g�,���������O��M��3f�H���O�F��1m�N+��2<�z ����ea�X���z⻺��g���y���qee��o��Z�8�Y�-�6|��?�=�F�歍"ь�������i0��\�/�ҝ�]o@i.�PFq�I90c�Ł<��w���?ٿ氓����"�n�Pg7,����2aý�\��1X5�������� �c�]�C�jru��-S�lΘ'x/b����a5�].�JX
��
�=�����!W�18%!f��5��C��J����-X `%��iymq6��^ӵZ�U�$R�!+�Q�!<��w�i�P˶��郪g6�t��q��|lV�=�l@�޹�ޤd�v�GqjF�)�&����$D�!~וB,�iX��x��#E4�V	�_6&�-J��Ծ{pw�%F�؝����H�.��Z�w�y`!T�_�����̈	�8�9�'�o���%�r�R$�¸�j�I�u��-ӧ	�"&㮔'RSd�`�lK�v(Rm�c�e��6�K۵�t�lفݾ�Ȏ>�wga^����I|���}� ���Mu6^8
�QiG�Ru��VW�]{���g}R��]��C�u��dP]*j'��KB4:7���x���#e��<8LW�q�%�щ��mG3=ʅY�MLSw���>����:d
��p�ХZ��*�8R�:"������� �=D�r�������.N`�),TkQ��\aA��'M�}i�7=a�K��&�b[ӑ]k/Qv6�o�֙�SV7��]W���&��`ˍ�!q�#��B�E�,�ɿ�`J��� ����C۳J��B�*�&���c��v�@��v��c�ˑ�"~1�MmIg����G�l0,�E��F�������g��7^���/4�CtQ�eI+�Li�����@mGB��72��\�DO,T��R�~d=F�(��� 64�_C�;;�i��援	���j�F�	l{��zNij�y�AE�S�m�O�.��-�\�Dr��<�f5�Dc)���zPt3K�~���M!�r�+��<�F�Qrq����TY�C��hĥ!|�Q��V�h��*g�=W�4�2�qA�_�WA�zl�:|dIln�g�'^7���.H�W�?R����,�X���v��ݡ8��]fu���d�����L?~���D9N;2p�'8�΅lN$��3o|G��oNE\G�"�=�_M�>;F4Tŷ7�D2��r Y��>ś��nym}I�~�yoh��6��f�� ����[`$�Z���|ֿRòRK2'"f������p��w ��<��7&���1+0ָ2�	�`���Tߵ$$�p���̓kRf��h��#�b��>��?�G2�kQ����⛂sލ�&��a� Ӣ�`���2�1Qmx�%��!����_�*h�$����WcNH���O*E1�(DR���P��&�ܰo��%#�%m��~y�|	���%�Ѧ��1��|�=����#%���N���\��-��#f-i�*0�����P�&�V�}z�p��Z�M�{��������Ѿ���������G5I���7�\�-51:�����E���������)��͘R�K�p=�A�?ƃ�~k�O�\�a���B�դ9}m}�'pz����r�ݽG��_�aޭ���܅ o��*!dWQ��uO=�Pn|�s�V\���ƴ��m3�:�
�|��np̽Z�-=L}�F��d"5��u?�i�{P�o����*��4ԝ5�_���HH�S�+��x���6�:�B�s;�O�_!E�6��� ��e^�s\߃�ב��-�<���|%%O·�TR�Z`�5n�Sa ���xv�j%�͇�W��CF��<�ja���P�Q����)]&
�_��v�5dP���|����*BB+�FQeI|j�7f����]�$s4>za��@h�x��=څ2���X)T|p������Q�^�6�Ԡ�\�QLO�˺Q��/�K��ԕ���4���z����e�*S�*F4ٕ}�Ps��.$"�����?�Z�ɹ�ٓ�K���p 9X�t3x4`�8���_/�̩h���M�^-Y�B}��Ivɜ�Փ�z=��uqR��W㾐�~�F3��m:��;ml=������}B�� ��IF����<&wn�>�16i�~Mu�4�Gk|���k�f�f:5Po�N'}���i��I�b$'J]jֈ�� ޡS!�gU��WI<ವ�0C(�@l��"D�6��4��\���BY�٤��u�4���H�l��R��'����o�3�O4�U7�|U�����4��g��U�5Z~ən���{b9|ȃ�AT7�b��C��JnB*w�74<���Bcd��� �g)
S{��D�kyl�nt%�ON���eh�����BO�r��v:�U�-I���#3G6�J9_��62'֔�G�����y�F�_����+��#t6��y�������Y�ƈϒQH'Ւ��MA�P�e��3m��~ǽ�2>H�t��bw12uM�\�yV��ϔ#��_r%3|��!%���,U�
Y�����ܮd�Q�!�E'E3H�zỞH�ϙD!�еvy��ky��U�Yq ������̐�v�X5���Ar:�J����+KI���}�Ӆ	��O�&�`?\-Rx-���7�&���dΊ�$��N��ˬ�0N��4[�����1)��x�H~���L\5 ��L�7���d�p�U�9@[M��,�bn�g��-�f�u��&�J�j=��v!��&\��1@ �������m�Y1JX�dv�A�1�c���0h[�K��Qcu��oX���运9��%J��8~���VC�����jh��
����
�����Ĕ��`�V��D��R�ʇ � ���w�_"��%D�%������v�ڥ��������H}�Dc������[6�c(�'�:�m�`�)X$j0�e�ɛ¶�8
4��ß�O�g�#k9G~f�_�=9˼�<|��AK��t���,d���!�#䨵P_�0%$��,����f��+]w"�l�z���fa��	���i:(�t:ì�xľi�ԋ6��C��*Ы��U�7��6م$�A���/@�L�wz]�<0�0-�G�}�;�6�?n�0��1�H��pS#1�ɻ�d�?�2�5��y�E�Ⱦ��/� 9Ao߯b%�9<f���仗/i�10�)��|��s�oi��Y#�;�g����Q@��2���xD��A�mZ2Wb}GNi�?���ǥ3Fsy�X3,B�~E'�B!L�A�Nhm��-���?���	��'Q��2�(D$�~�s�f��.�r���|�sN�����hM�~\�|���'��:�P0�)S�c���Odg�59쎁`"��F��=D-xM�5�"m�-H���N�ݙR��p級��
5�I��y�j����]�����p���A�A�q��p�=���7E��(�����C�YPHJ �e�/��	���Cŋ7�u5S���7�'ڱօ! EV��!��6�dn@6��+�.T��ri=ˣ����ë��b�X}+�7O-�^�
�;nȄ��8)��
6{1}�U*�mpmP2_��	P�t�C��$f����`b�YZՕ�~��o�LA�+���m=����$9ΐ���B��ۧ�x2��iﶚ�!�����RJ�����8.��yi�,�^b���J�J��z{�9�$kη�Wphg,��W@H�b���lOS�(��ū|{n���gN�G�%^Q�rC�T�N��q�C�a�A����p�_�w3��Gk\2P�%\:����T