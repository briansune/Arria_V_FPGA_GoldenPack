// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:08 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HoA+WWl458reFMu/LL1VnI98x18WSwO30Nn2sSn5W+qdiBjNM32a+WDcu2h5Y44g
cRLot0FeDkoRPrrM5rAu9TnBSA17BXrux/7wF+OWQBdcH2MQ0NbXk5ggx+r2XXYH
yFLYNk+MsAcAXO/RoLLk/CEEioMfbotMIeipk8Jv9+Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49312)
aP29sSmC71tp2ohut9qWb3DocTeiy3mpSgZ6G48qAz3pQ+fsMhpuP0YJ5NFtqQlF
DcEEzf70p+4nwZsH4DsILmckX112+QldV0SUBZHbwt7qxgfBNSfDhoIO3zhNG3oG
S1UHm/DhW3lRhpKNMiWytzWenD+RfpgvXcQ0nUBIzfu4Mgg/9kEqTabkMOeKuFWD
EqRY7f8i9Veo64yyPb5X58pbPcUXMxx1yWhQbNcVtLL+rRy6a8sqLdmUf3rbMpch
vlKKmaX/5QFcxxd3SaeYjoYGNqBratXSRcWxxVRylE+i0uqJpRk5gH5fTkii/616
pnqrryPaOG7nlLodwdEcv+ubkqXOssO4vRus6J0p41JVIH6P+duqsM1dXbJS+2vx
5cvoM3KeE12Zm21mOeF7X+yKkhzsUhY/EbIdoHtBB2N2FXVoAhep94O3GYBJPnj5
eFgiP6QutznV2SLWQjGXs1Faw9T6Bh29wJpsksNT2Al/DcQQVHx5d4b1o0Pw5bEF
TiQoro7mbxM6Jk7cU19NyV41Jol1usJYg0vnGCCXCEvMyBmsEdAMLGAxJI0yDSqo
lXUBaIDnLTRL9+ynsS90KebIFh67k1r+yHAbos0cKf9J678S2c2wxWVj5we/JmO/
je06buJwDtuge4lsaaesDE8Yq0bErm/bC7gB0llH8d9QS6QsDrIvFjScJabR1d+x
5sEgsstIfkptm6qAdr9MfX64PMxNLXuIe26rlhwmg3jYAw+jiVUUe0p0hRvd+/om
nYfqDRKiOMNlRackiNojmcz1Fmpv0juXy52OOzpiVFap5WJu+S6ccsBdLKmijyss
YiC/CNH38jjDYhlTDTSOmsgyRhPpSBxch3TKEDqQc4JnJKjp44sWik/Fm0YpxoOh
DPyseoCWDeVzi3ON9edjK+liOgzrk/BxpaUKUevFh9JQK3a2G5o2Dajg9708s5vZ
/rh+i3So1GKFXc2vnTZ6WniFDHmQAnQESOmse/vczlynACHtgqchFHrxECylWmZc
DdO5M+TBZym7rKjFksopYdpURGmvD8mQLVQWZPIBtaKYeE1rCc7zXmKfrfEGNA1/
WVxH8rojaXFoeN594XPJqal2sLqe2UfC0n7uxQzr1bJOssxF7WW8lEsWMFkxCLW4
I+WFOJ6h9zy9rEqXv8VpdrNeyGg9XZ4n+jDRj66qzIA2lECJEHdHD+GTy3SEbXkT
flzAd6l5c1buu7x5UYhp0HNV7IP37cUN4svM/l6x5CMgC4gUcun8BkknLZoCl7ZP
aUJXMZ7drGqHCuHPUPAMxr1YfHvxqsghVVAOxfyjW8Vm4SpVuZQZ7S1plWAcOpuR
7gArovf2ICqKJ21mlbm5uTZWnhsftEh1CGPon/nnvhZIYNI1a2nOENWPiYPPmey4
FxbWjjev2sREpLQ72PYMGPAVJ+cB/xVLyzmEXn0/5FUGyMtwsSpWXmzVLWsJMpvn
B3qaRK3g42kwuUchzlmbWmXjAJkAVvN2Zo4X8xXUrn0xpJriuHKeYyuZzSTOHO03
KMn/qr24KYrH17kR1aNsQRmc49qbvhimowGg4dTo6WphLdVL7gWI09LgSpwntOFU
ikx0QLsF77ocXlL6/f+cTowFYo8Bb7Z1SF+gGyX4NP5iyMoh82cDLUGTQdUIR+Zn
XToXL2XXW69pzfFgnCZWjt05ynyxK349IF6xxstVIo1t6gxEp65tSCTKB9v33UpE
aZj3DirEDSjYAojdK5+0Y8TcfKyI+eQY2ASFhhcstyDdSMMheZtK/uJBdVyj0Vsy
5ARMh633CcMHuf9ha5OIMiEANvkeNw0GFlmTTHjnj3FzkZLcMf2p05wtCwTYuikO
51hejs1FIRqpda17W0nE/YFeBdWIabO21McDde+DldSqzOGbrZMKnWT7s8rGpF88
PrU/BiuXGSuiAY5RmhsgHq3dByEvYXh4w9yJ1FtUretytm0/N+zdRZOLgTLoxZKy
5gOw49CftvvMDmqQafTUeliKZZbmn9vQxxJXhjNkU+Aww9YDc4TFIOA+RBgF/lU8
bK4zsRbpvu18iYqD35hJkBH1T1pAmPShL41KCTsGNrbShkBMa9AWHZggi9DuZP9E
O575MdUzJ2g7PKFvskfZpsbwzJZbJc91CFmLyShydZ1ASusrwmOj2VK+VuX87C0l
8IRs1N3KXREcz089oQEGYz5D22cuhfuvwjk34SdholUF2NP3AMMIZySY/J5nT1hG
O72ivBuSMB+MbugHVoGAvwVmV7tNs4ymFzM541qrc9YEn1EZLbULgX5HH+J/AgGy
8CNKaUcbWk/DV+Z1MIoSuNMdZkfUR4tX+mXktLh7i+O6KMR6+TlL0iUzbKK9jZRh
kUO6YJO/m3KDa6fshKmdNYwlWKGaGU2kC/QipxnEDsjM8zZQl9EKlgSVEkUAnFSo
9HqunHyVVZOlujoqJd32dDuSBcKqV0m7lCNQCSaWPLJGt3qiOxHNkC5MESnQFXVh
wtOqLCawLgnQ6Fsz79pZ84oR56h4xd0jJYn4R1w2LsLgogGXy6zANP/A3taPxGaO
gjOXaJPfxTbmwylgOC+f3yZTkENeHUPhFMbGpYEpZoZlxIw/N/CRqZw2KzVrEvgO
w5EmjmTjH/8n+8tAE5BkYu3xvd0wIjFqiPdYbwoNjxtMz+XA1+R4f5h6zPwt+vxd
jaMD1yM8JwV3QBo8kDIHezEv6BwltuvVznRudRvyZvV8BPsyC21F8RkpLcIXnppX
VZ7GHgGdRkUC4A7uKzkB+EYR382Xu4MlmLDAP3Bjy0tCyqqGZcuvuyQ78yPWDVBX
MzcQsUmSrOK001HwBD+S2MXIsOGuLjhD6N2M5Tl3T2N13vFjZ740i5b0EzUyaByQ
6AXiDOfBD3ET6D3liwML4cDNzzG9b73jRpMfIwHx6Tb3kaTRS/a1SAtuVpkcxTEX
m0lKt/y55PFDVERGeo4AQ0aMNxMajMA1zMZZQ1z3UwFJWrmadDXajn6EZEwM5YKM
R55DtrqGq1XuzoK+TW9yW3aFkBc8WRgqWVSvEVlf8RWgEyUVvlkcpNzhfWAh8hlg
nyTjcLz6GFTxbMBq42+IXfIUTHVe3mdQanZxvBTzE3kNOFfbWFt0f++RGSs+lH+p
1YX59XkfirSa4DO3u9WmX3/sJZeMlvIG01UeGORvjsDBSL6M9ZCeZmc3a5nk/4V7
iSR+qxftFQAWNRTJOy5xapNRZJVDkNBNMPr0gEXlcn/or3XWUZJ3Neuyjib2rjp+
fWmVAl6TQWv0AsY68hgjhXPx/98xzoCduL9zoEE92CQu9SDu2ixKg6v01atm8K+W
Ks0Rx5KGfrkz/TQWcyVu2nh6kPBzl580YYM5XQaosSVOOEA1JwUlUBHxZXE+A6lh
3WXif3fDGHdMMcsIFawaF0avMDJef9C5tzRKsp8/EXbcDo/2eK3HkTWWcNjznlcY
ajy5eRKFeZ7UgwYwNVFWgkH4ol9HTefAa9sEPnV8FKbFNykID+X/dr5GutOn7Rpr
cDi8HwUbdMm0xNhuTR4ls/w8D48F/llKNtB4wK5t6Dt0uvwwsLzanURU0DgtaJJY
6WmKj8JDxpBLn2D/+yWmnCWXX6+2DgZ9yVnlQXKi8OzSuab5ikm4x+3opmx7eNGL
OCJdOLiMGPO8n0GHZdPaFJdeZeDaey6t3ZpZ4UfHoLNCxoBVT5dSt1HAiOMdGAlb
BTois4gz3+bVYZfz/uiuefrp5viabolJQIaUWBtP4ZUbbcc+U6hzSJj7PLGMZyEb
VqwpMNZoOSdSR4S6x7pV8R39DOkEekEZ9xiZOIAppS6rRo/I+Y3v/x9JJVPv152L
HcAoeBhsJm6MqwwHC1slu1QZ7Ke+nyuId4QruwkAF+ohdWU5D2EZvFrWn4RreDLt
L+vOEYYaZNfYZKD66JV1i2OqEseeiYjyMy9BLF0m8adq9509Yo/Nuaud57EtrpvS
+lhXqNWAyTYnY63SfeVwdh833BfNPNUWsS0ktLxjGucUv34g4uTwGIVDTi94SdY8
eg9grN8WJcRXuuyv1BpgWShiFdR3b7x/7nrJN5+N6KTM59/hJmKCMMDAY61l9toq
1rHf1iCzqDqEKs6XLCLXMizUZOqxXYXCoyME8eHC0uvekkjjQvFFjmWiSwdvPx9p
apHbN2Hdce7o5E4kUMQT4m/cECp46ltxiIDoZcLDbcLsb88XalFn67pNGoISZRU3
jX7vzc99s112aqPzmGLUge/pwyUCMlsOWhvED35J5l8dPIy3QgZUlJsYzn/fsqll
sLAurKc6DCJen2RsfACosgPmOyF/Qiovavp7xBYN86tf8vzOY1hvNl6tb9Bg6qsQ
+Vvm+3Tha0cxsmhUT7n7fpQSCcKLy++JNu98yQwWTk5hPKrDfQPm7irZEhwFyWGK
J7aNWKEcXWdUafddCMdz9Pmn4wSEgp3HPDQqUxaBZ1fAWqaKTyM1LtaEtF7PVIRZ
EPf+habBWuDUFuDMp8mw9RPEyp/V3xtB9xh+EVwPrKgjiLxsr35AZpj0R3TVVuox
88VhjmkBK+pWS/XZuDO8Sf0mM+jrV4ZeyuzBYgnoXxs4eb/iU7fU/Opf8dfEoLAX
Bt58hxRxk1e1kJa2Qf+rYcnGFd926utPj8kKdsicUHm2jXpB3lhPEkUUfSnRjCkf
pMiOybIL1KbWfgTF3SGdzbb3j/IwZ2p7vqXgXkkuS4NFi8kHuJxUcOXARBDr+A+X
DzdSd9F1QFO/LgGFyzXJeEgCiNxTzLVPLfw5betorMRHU/87vS0c6QPE+TEwZQxW
a0eVKDDDRWNpwI3dnWn9+8Qc9oi8uD9xwLO6wB3yNXjWRznfZ1wC7Ry+qNkzhFFX
T8VG7juZ8kzVcjEsUVcCOlGJYgBWJSb93lkvudcIt4QO1brkJ4tZlx/RcpadD8Ck
TBY+JT3GJnKwpCcUxFWmK7eZbtwam8uI/2n60UTGtxwWVWKj156LZd862gdBlWxj
OBLX/ijTgyc9hlN0d1qdUNg+D3CgsRvyji1g1HhXvpMaN0Iy9ek4EApCz7an1rFN
x6z/uH3vlgpfw3ct4cb8HPJdAsELBelhkUoYDXfTbbMyys6n2kFECTmNiRBFFz3+
Vd+3crigLA3qLlfGLLFi4V9FdXmr4uL1LdZ3V0hIrVMNzyOMzgzcM8qMHlV8NQ3y
gKezddocrmKYBKCt8JnSxgOwl1WA/P19ClMMqJQLvyAf1R5olqu0DgrPhCgj/h7Y
+s/ySgNYRkKP1DL+76gFJ55u0banyjygbF/x+caVAV0Ypy8r2xkdvUAq43MHDfO4
2ZpI5sX8e+qaNUePEzAkUqJvHohYLXBb58dfLK1RsVOZSDnrh+sxbh3ONvYITSWM
ykw0BNyXNTq6OFroQ/grbdGyowVf/RrpfRHQOiZPjLrsGt9ZqjwBKJlRJl9SduYQ
tyDa/HO8GQryXFurUCTVCFnnQUWqeMQqWTcMvStHLiipz5R4Yui7cbE5qMrUMjwZ
kemL0vKdKcMmht31aJ9z+wZmi4hZOHjeQOyMln1OQuP4y7WP5ORb1REEP98L6DAB
jpLetfFkLFAE5voCwc5s5cMRxLeLZs1rEGof5tKkutg/nfH2wkp5tpblCBSxEu4x
tjCnZ+HCcw4CSbcI/O09hMkxg8OIMwsrdo47jcwflzm8Lp2duKJt6zqNuDM6BRGj
5SvVEJe2EBAsufvf47lDHpAOhbP4et1WAb+LKtz0ie7Nd3f65zfcCPXcn81W2Dvf
CyToc1MKFP+p9a6XOc6R0Ve2hQsnWf13Tf9jvGHmAfmuvAsgp4BnMjo0Ju8kuQ2q
HW18JplSi6IEsbDScg9frq0OyINaW3eIROf6YU+2g5vwvGEm2F8o9PATNymm8Rmt
ZF9p2grhe8JBFuSM4960AH2F/+oqKEASVKORr8XGX4v9EAtchANVjQxjvwuNvbtg
44vfRcJ0VUHW6SsarR9FEsgD+B2jPLCXdN5Veot9clTPId6zfJS9I+1v5hHRQnJr
+R51Fr2cyaULjvtvB9aNmYPfUn1O32SFtFgjMKOVv75lZ28u9dq62Xi6ZvXINPzK
BrAiXdl4mjHImIxIuqvp089pip7kfPCvqTt6lmK/wL0x4DscRs6DmdoYMSyTLJkB
0MHGy8cgD2M0cwknRwl/uVu/u4W6XBWufvnRLRbCK3WrZrwcrr0Jl6Vk5cz2EZBj
KIEqRmPkdUArjTgmhIvMqH5650/EwAd+G+EJsS/VGxNlHPwwSLakc52ybwleuyXp
w4QV6NzEeGgS6xYm/rcW9Ar1nNgqwEXoHBZL0GpDX+0u5+G5PfCWOAtDYXNFLsHy
axsBynuxDSBNSsBm1bL0630RF83Qxcu9KtijIPG8Ci4nt8rgv1VEOfDaUr4zoCYu
jLAZIy5IOBRsNcRKFZyMtiDfY3IqNpypKwGCSvOcI+r29HqYBZWRl0ZOtK6JJk6I
Demf9wLL6mGvqvv4nyeBO1xUHx8D4/HHuzXnk3yrVwTHZyCsfZutty5icsYgXtWT
YsPwgpKjYmV45FoNer1MUfGjXIge8OkdGLnluLpixzB4l2nN1j2Zo5dqWmyoVjV+
pGbTvsJdpV7m9AVeEV4JSkQ5s/FOZvzrRYFozFO+vl2OQ0z9ZmtEnQVD3yDrwzyX
XP5IN/QjnRz6GUphdJrGV3Od/LA2GdNIccPY3E1ZbXLdK75NQcGZJOc/7h6txor2
GDFVQ8dciAG53EQbHIVamsgV2m2wpwfKc5zlYv3i1pN1o7io6aQyEJAiVHfvtgdK
+qlX7kF51lF2bFI24ILYONou0saMejjCodDHJbVtRvnTA1BCbPg1ryN9U7nguoV3
pSazaiFvRjs9RVlxhX6D8S4k83lH9/HTPzXGI5ICzza5aXH87s4R7f4BUd2pBlZw
Du7UQXFKzo/SAtiO05WnAdL9i6YtRiRgGRj8c4TwojNbsPpg72VQay3xM4rC0L88
F7Kp2q/sQ689pwikIafYHycM38lHrKraA0UQkZGnyjSh3sz3dONC7N0jBenmND6B
aOGyTX5yTlIv03cXiaiSl0orl0C7AFpaL4pkadudDM/AYdlgivOhIhcG9iyhRE1x
JlBMHNh8mnrYLgf4cMOsGAld+vGlGjACP4oUPGj7uPYUVo2hGxaXPWHY8AfqG6s8
Fy7w4/hfK/KXbC9a9qtDNeYHfQfA0QcZGti2fnooLNMkXRtbyixzjLQkxZhnv8JH
kL50vs6KH673Bh7mM1bjqskoxrqjiRmd9YJM5IgwWlF7784/eZVeuIhMt+QfkMmf
0blrOZwFLAJ4vvcLDicKdNQA+kwf6CTMM5RLxyYuqAyMDSLZ3SSVZ835R6BADPLP
WJcTBvpPCyzN6rDAg7mNhHLch2cjetGbTkNlikBFILg2BLsHeEFMFSg+CXkZ8PpG
cj0g00BN4m8FOOHxCXOji1G3fesrLgrQs+q8IwF8mEJC5OZGTMGasfAzfE/Tr7N4
QSwak91NroAgFxdCs0iH6ZN2MjLBXqa/MZLrekxKZen6+UcM114DCtZEGTn2pMC+
pf/Sd48a/YmjsVGz9IyYE6QLTtaXloOYtpBpQmyRiTsRWpMZQ0cbDujzZDrWom53
Zln31NBxQpTFp48tYOsmcW9UQ8J1DWsgcSG9cJeaT7si04yEuf/XYdOcnL5B8UiT
jOpZs8XMBlwO1A3AfZdADKUyRSU+AwFmluVS1h1SJZ4II0UkRPpEGzaThfSK9587
De3ad1SU6DfWkCsVMQjqLxvrG0BNusgmqmnZjxK3vbgkfMr2ResLnI2T52UZsN52
wboIYMeRR1LwdOdg4TWqxuoyjVnx8X719KinBnrRO5GS0zbB7I4uCLdcCOKMHpgw
Y2UtQigVFattsTAqZuOPhtfEeqLB2dCeaRe7RDeBnlpb8/FfPpzJqrhyJJ/KcKbY
xsT+nvRkqMp5utMODCeWcThhVbcpLiib3Xa7XQ+b56PcoA8r7M8pUsur/qchFX65
VTjvsBVXN10sdngu9/KDYr2TXl2D5al8bUbLHN8uGUaMNVYt6qBBlvMgmPQbcxjz
HUO6Vhav2BiPrspEB9EvfTahhMI8qT1xB26yenFWeHR4bl/yPE661DDlTuPOznTR
zadVANR6Y+CWQ7lkH8DBcjt5Q+LTAK9Pw3OLePoFpgT/DfrsR3/7V4IfvJCI/cM4
MwRVlKrQ4DtY8zN1rK95dTlxecSXdHwEG+tFCpME+YbELRc8YiuSNqCI+9IKq6QV
yE6ILblk4oN9TCNfBe54uabmyoIe9Dw1MzAGP8nSTgm1vtujQjhLaGiZD6+Aasxr
u5RgOX+XHjFP/OglPG6dhI8SmSNqyPZCEYcIiGsIpgbToZRuiUtISK34xiocKhVq
4D1BI/jG/yyhUJkei08qS+k1Wzz30yU0ZMT0SDxtWKhwMmLF9E+PgVPJG1RyJLtB
YZ5nWPj6MwPby3XKA1P5gFxRNquuQcinPPwjE33+e2GPKIYLXLvULwCWIr1fC4kF
3dCtJO4cy46AUa9D6cqeSQ/pj+9LF1+cLyNyZsHxSN1G4H/sJSuBQQNfmfjI/J39
CWfrGbotgb2sZ0eRGqRcn6WvCx61Gwzr3GcyxmibslVyNgAxnc3tZ2YodJNtHnUM
11m7HgVld0olNGwYfzvuXZ0U+GwLlZVmXufbMhf0Gn2s6ftC3gOJsXswPRhXeo3L
zSbs8DlLg2IY74iPLu39p2bfK56xUJ5Fazm+D6BVeHrj0sQ3ONkwYq+t3YRiMwZb
iR13A299NozKo/RcIhmvB0cDp38CXyQRfJqmfbp9f4jgr7R41w9DogfDAMv+6pHf
IVNohbKxs+Kgev27IISHaKND1v6qVh5xV0lXti8ez7qQ5Qkn8ATK82/JNE1pJExp
vGllvGp9gX9qqyrpO3f8CFXvIXICkTO2+OJcffnFo0ktL+N6eWje7y0s+ACll0LE
MQ68gd/wq5u7AhMAX+5PB8QEVoTHzR0cICwj3Bu6ZUcDdmFRjd4cLaSfkjBle0OA
VJ6KBrgy+POB9CkJrUzTJuuy5OELGJUV+5Jpuzk2fnAwv3YV5DUf1/3snxyUlFTW
f+Dv2FVECpPaM5TDXTBkqvWouTC/3n2tlu21s99g5fQSUutyP+OOGs9MbHgpqhL9
DE9horFDNAIzFozp56NKR1LCBHib9z5CHvp8Jwn4Mhwq4ydRt1PXC24Mcdcnx89v
3NdAWjLwtv/wjrm8IfFr2Yv27hSaB0OI56u80eAcZ9vcfua/0Ioy0P97erGAKaLZ
ViqUdBPlNRSLPLIfQmC5Pph/rQ8OPps3BBw3zUIMJYTKqLKzsSC4h33SqTwI3MK/
5rJnm4bt4ucrVWmjl5SLGq5usMgFtgnVi+alWA2M8X1zrbBc/B4OvSOSCz7ivUgO
sXSmH9VEvK9hkzPdoXPsZo/ZyZfPMq8jvM5lTw7cHrXa6fhCzuFg8qPG2eePY+z/
3iG/XzZhS+dFfb0MSh+yNlZbVeo+LpfYC0g8TFrq4eS6BlnxRsF6+xEo4q+Rx3Uu
va+jVYIRQomVeIx4iVoXyFSXmxvYtr7B8+uh2Jh8rQtItE1/L269LaxsaE1GIy/x
WwTTAr7ZgWhKcQlHG1cOEddlTM9xzfj3P9a5c260Sec+di45LEzOVMsB5L1tAJsR
zhlHpM/3Z4EE5Ko6S73jmfN1aIhTyeIb7au+nHjewyrQTYMgDufo8z1xOVnTOfo1
EPuroxWNzJkT2R/Z5+jyJn/xNI9GndYdT9oDR6pSULwxXYqEgbUFNsQNiOMabaug
1/lb59I/wcjYdo/yYVosIbMGWuXPeYA+TRVYz4nP1VqdKcjnK1ZEQNr9glUR1tKs
zfaVgl+WT5zYDdV5LSeB9QnQJPUBV1pJa9MhUw4BP7RT60nSKqpesY2s2mcm+UFe
rjAMBS8cDvoDHca00+bx8XUJVrIsCIJgij+w2kRuDwH2mKkLwYdVPbM7y+E9zUQO
Y8kbM0QGBRQluu45j/MSPmCxcrcmjm+Zsi+z/Fpvb6upIznw4zE76IpqX7oqaPPB
sX7Yz3r5RHKBRSX/h8TrzNdXGd8s0zl19ZguCF4DKwA8ZBxaSIBcSoC08tv/MVUQ
qqRvWwXssvznYnX9nAiAruk/Xs+GaMOXzN+xZ97tO2rK8Sc+2tkpdXsK+iZaQUgt
8Hjwk9tmnDrzZiz1K/gXQ1oHUTvBPyE8eppyI0KSkNCKpLqfS6b2H5rgCSOUEh51
bYRrP/Jb6tYrU94THjUJiNMkXvM1tQpBnJgsM+lrOZPm7bEc9UtJ20DbCdpbIAM0
MEY01tE8g5f1eyM0BFYDTpD9Hj/hsK2axhEgMnb/XkKLA6fOYR1idaWB2RUofDlf
5dYzctrlG9qbQQuHMAgcnWjxZg2bRNfNq4jeMXtVDZ6yoZUwkj68MJkVoOEC1/Nn
JcfwiS+PpNWS6FEkF9EknTYp3r/htZ7PKPA7czVXtlO/bejgE0oMi/rpezww8r6J
+rji7IvdfHSm5se+efJipIcgMtsFYXlboCHtUzxtLEAD3GsnRvwX5LsbkA9UgWV8
ZO7jgdZdF9EWg0R5fk4R/QibYqHkDyFUHu7GbcMteiQrrNzDaUB/6U8Z2C+ic7z2
ZArVfQ9pcWtwnGpmpAZrRoBRe3oH4OMyteDDBG+MfVT4HT4I7jMTxX1ZKufHe2hb
/keKE/vpVTyfUk52QUS9R+tvlC8kUrH5RpJV4mDnxv3H0Xkh2vzwpdS3cMcolB68
gCsj2pUwSYTWfdaePzYzwZ2kcLsMs/wE0grHgC924YsnaoUj0U3Q4KJo024Fabs+
DXaCHftibr75LaDEkOKej0ppKAQBU03AechvL3CjrNskjrIZx+mtx0SgqOAatMQS
t5wAbfiUj7nn8k1lebxZEsdjuCMQZ7jhM5p9MzSy9E/ozu/Tqb24nRGNipVXE4KA
Toi4wtoQgF6q/52ZWMJlaZXq88zY0o/5HwjBmc4WgH0+13hx2CFZl2AERWGokknH
4sbFMdE94Dkc5Qs4zl+4uGhbwZy23Y48HglCZjxEDIVqH8HHbEYO+PDoWKSVktsO
PlLjr/EX/cc6oC2rrpYFOpNF8RQS/7hHadmbqYkYIqo8MEuDxsjePqfqL4BqIgsa
xpjIYNYd9/lofYCwWERS/deA/ZjltBY7tn0mpPCr8PvGCnt8Ave7pSHTl6UCiy0X
7Wj3N6cXKGMyPmawMxA8Tj2kW/aj2TN6j+Y2bEW0akmZpYqWiDwdG72SgSodFQCk
1HRFoJLJdaFnXT1aZ6DeFIwN4bcvwcEBBxi1pvgujTRu05aQEDk5hFYksxOanFb/
yS87pfIvzRAJt4Srzi/1DUG7XDlZA7rGbSB+9EAOya1JO9Dd7ykE2FdC8Jx7zZK2
S2DMRDu3iAZ09FrfGMM1bq4+1Fe6Qk86+GyQecW3vQ0SXsXwI+L8l/StQ8moEadz
GrVj9WC2NQkWCsEKI3xLzd3uLMVneEPR+pHI/1evTzYF6Bk/EZMgSuCrl9iAZUzT
oSDjYrpfcVrP+oQPZ7u2GVLduMRtH09a9sOL4DEQgxUFIAQLgQfsXsoUjDDEu8pX
DRJWprjMQQRcj39wLXMUijKH9vGIKFM3Djn7kA6NMKtyeZ5otygIPSHgp5XPuSqV
L5LQ7m5TXMZH8rVULr80af57TEIMvMxnTWLDeW5I0xZJF7aq01Fv9yhyomS4fuSL
Dh61pUd+heptihx2fIQBA6piwZ38JLgwBhTIrM5ne1wyIyLIldHyvuUH6g9nTYam
YpWxGGqorEGid6BWXnWQ9Md0yCejZ6RtzyklV+nDD/wm8lAXz4mi4a4Nbzbv1+q4
YIkxrhwczyU9qsrqZTRi0BW9I9tz0wqwCvfYT307wUM2AQCOWZYYjnvSDiFRo6vV
t8lGa812eLmlWjkJqf0YivzVwFrsEVtGfJUEB2xcTrCXrRNdL3Ffu3yvRTETZa8n
wRnxQaEh6RAYfRsem43wsfubQnCMYhI0MuoITDo/GtwH3DbsUTQZzv95gdM+1/H1
WyFA8DEz0Sh/qovyu8t5Nh1eSPysBgObaenlUkfcyZGnXZFjArP+mBPvY7YodEKZ
Zv0oQXuu+qnVOsIVPLpKswK6k9e8M7oJNbkhfBPj4RUnGiTIMqD2VQGkgF4UUMvA
CknULa+OH8dha/7hcKnuUIXBZn60gwQ+d6qNMRhMvbMWs1x9ZJB+R83ztPR5RzY/
WP40ekqvXuZ5Mcsin7WXVTlNhRRqvBmoL84Pwb9X2TwesQA5KjdwYRaSpSXrvR7s
Ky97GMEBcMAF46ETwNIL/DnPn6C0KrFchUUaEJ+aew7ded8iYkxm416n9JqxLnyZ
uGGAFnlPzG6L061h1Q9CcfOpq1JnE9wdYhN26AEAaXkIaQ8vW3+0pVKOhEKO3s6a
vIG/zvoj7UF+MKjmzmukkTVFUaNi4awND9gFcJoqvMAJX6f8qlu/75kXhnjlwTcr
aUzn5L9+aGlBxmAcgeBiS5+DMP/Z1n1ASDYzZrj6qeGBVlz1WCrI/AyMtuYo/EtK
z35cWn0uWbWAwEDafoUXNXZCQgEVH42dd3255IHlbcCYDqLTm4hnRfEEB8fkrq6R
hA+bWg8K+AVEEM8CFZbFmWK3r7qYY2txJuS8n2/ok1tnkjxln2pp8qroeDpeUKxK
1wnpI30pAkH9dFsivMOU1YN+nd2GXKGNGdOPAQORlh9cxRWY2W02AnVhOuN90NuE
Ee5gc3TExWvl10CsU8mNXdbXOhv2iLRVcgIKQC9+wExhUcAgF0CS2Yk5q5Ay4T6S
DvjYTe9cOexupajeGsaj60DqaTsF3Jvd/GhAcIpSDaey3U3bPtdkHSRmXh7Fbp4N
dg6Dpllik+n62keV9Jtl5jtdZNdOZY3eJdcwxy4TCezDEgnt7RHILV5+niZUsx4d
/hd/h1DTHRWiOZzpZLMjYrVrgRJPrTKCfUy6X/aTiIiZUrNT9wm3tZ6l5zQVl0Qn
SWhWbYIsMpz3C2f7+4RHJP3TEtkwonBDyA9945HRri0EM3bo8NYWUTLH0p/e1qyu
ugaqAAZCZUyizDnxPBc7/i6yBMamAPuz5SaqGvvvNd3gwSrJ+o49cLkEGaPLpcT9
dP3HrfOiHSXvCnts+H2oJu+PzzDEwUK5h4KnQ/Bg8eUR5EugHEe7g/GIjbMi5l6J
3xyrxEztzwSWWYZ3ljzjKMkfb7t85SWuHndfQoqa2qDKR32BEeE7sd1B6/r52kcE
I8g/0XNOjx8bZsusgYOJZxj/y+AcN3MBWhNK3vf2nDNgXaBqQUm+N7CAhduKkoc2
8/Z/jyvrylXjgiqX6DuKyvNNFQ7og+Eva1LVrpBIMjHVhd3RV8NnQ8z7GyppFdEv
NbickfVFKmZ5YcYJsrJIADCqTH2uI9Jytksuida3sNdjvQHhnYAl5726GvydD2FJ
RPN9JQJRBNcw3ipQwVsHyfcpiNiI+0NUlG/RPM6SmqFYHemi3vK5NFOR9CYSTXrf
Lg9g5uaWGu5x8W2k7l2/VWsOYl/S/LibjcoB5gNe1a0iHv0v+8wwJv9qJ6EPDnZc
H4LWic5x9d/FtnBQ4Equb7xaAV7lHrXXZunkw175lMlb81LoOKj3KrctLAVsQTvz
1z0pfI8SQnE2SAFAWr7i34bnX5oLw46InwbU8RriS9dn2T90BZklbxqs8ATIwHVR
3cnTKwbQ+uIO6m8LVCWWUqxqwPwA13VkWHLUXaHKzL2YLerTuuvh3bkWV8ambFyM
DtJRzftLIpq60gA8K7LCwajZtaQijyLfJ++otM/302K1qIOfWRvzb9cM599+vBuw
ElLjlR6ndFR2rAHtsj8UPyhZ1BOibpJ+5LS0Cz2pUSLxxjHTkqLFtrIp4COds+lC
FErSoV2iQLk+iONfvlPfDzWyTBezKhoWynI2l8XjQ5YHFkgGXykzdstzLUo42D13
e0NbnipOUjwxBDx0gs+5uFtSn7B894HPkwAcS31SHjYvpJ4ZCSCpH8s4gS4/p+w1
ntjp+drZ0eQJsBzh0BSU/g2SR1D/oa/BEK06TkCop+KuzGD9zJw6DCYUq0ROzlXV
JsOySb1ySWcDb0Ni8jv5eNy5hEmR/l+V0IjknyxDJcS0Fy6Yv4gcQUJidvWxYEhi
leBNaQHGLKDm7RorGgnrYWB0bj0I8A3VzIWo8jeJdOqnLzsxNVhDu63mX01ZpIJC
rTGFsJ+SwbKwvQeE5XO/z1IH2VXDRLK31/eTsxfL9AJezR2WfFbZk9IH+FsKygrs
sW9W8iLD52aza6ls7REfvLJNQTPbAoTJdN8B+wTKXF2sgmcWnIfbg1y3wfc1eKQR
RFMs4RDO5jMD9C9b5TJIti3PJXpFOqDgQ/wqt/sDBU8UrAD9HH60pdsyClraMLei
yhjRSd99nMt3psDEWec61ejJejTQ3QtJHV9eVIydVySl0naizF+rwpOINePJNcTG
VyKtv6MxrAUOJeqIjlpGppOclJkc1lnB5M1FExAzB/WxJ84zUkcpRHFECLelJOMM
6w67bqhS0w3Xq0g65JKGZKdsZK+jmokm4O4AAsrvV7+3Cpcm4HrxrzfddtlI52Qp
Ui8DSZvnTfzcpkRiyotKVIO+lY6mlDbNkkImr8/THLhCRT3/5nYtRGpoVipaMf2b
gMXukdwRNEceneIT1rZmxPLqtSGu/R35lKjuFsf8NFoZergxOTqlwflg/Vxp/3Tu
BJXdH3Tn47V+3sfl3S6X/3JeAkCq2WIoM7s624wqxxp6VmWJaCT9/YpZGFZZdUzj
ttmJHcEF60UjTzxYf+D/wsrNDSegVaLSlpoMPxEohT5l9F3Ast1vByLKhqa/FLM6
HcosV8PKhEoDvLCBItCaO5bcmMO1MBF2gAplSbpFrTKMtNTzF1awHUlZ+tXOwgm1
Tk4W+5tGO799HMHdFQp9bbJfhXByJATFW3yQ+wH3HZQQfeGGNB9i02WNdHrQV37x
KpLMoaTXJ27MvWccrXvNMUJy36I3rKQWw/CwztQsHjMHh6U/1FL+woWKNT2Y5pJj
nMY2lGZw2oAJX0DmxF9qO/mloMmaZ1C/0nFWPH2vx+/Uq/o1iDAmBSgJyE6sZhC3
wvt9dHnK6lgAn7/DvoQljMzIgjdfFjQ7mZ8U+Elgi/XfPUWzH4pd59VgttflIndB
27CrS+XIIJjmLQcFLNyHLbW3tTblIcWNDOJasOZL7jRLpF+zjavAm6J6LqKE+mq7
jxQHGeOkqaX5FLXPF76CwBsh1oTjEcHBYc9jAdmaPoSprQBhNEEnlsQ/ILohcKIP
WbjPlL1r/Kg0SbnjSTPCw1pn+E3L8bO2BV3HloUWv2pJ+b4WXZrCNNJK74pr3o24
8Og8M9iLzRgG1rW/O9JMVdTnp40L7YcOrV9zQ/ZmorjjGBPfJj6eDgngiU+HWsAe
oONqGPiFML43TgqztipkcTV6e3ROVSSrJ86/i8JaWluwrmdHei2H9NHvHzrluHJi
LtOrP/Tvcye0Yo8ljY42mR1/I2rrwCUEUBldyJ4mNmv/TGl+KuaaMVQc9NnTnJ7b
vZBjYHYNtYKSy2t1Mn9Q2iZpMnIZdxA6b8x8WIb8s5cukZil5HrdNdaSsbRzePm+
9atxbiB0TuKtkuCjR7S105iIH0L4b2QNx8OmFIK8jpI/6UrmwJOUE9MpXxtninoL
3PUG0wMCUG5EjRT2zM1imYT76xcBVieMMzwFanDhFoUsqAkN69Fi4bICl4ahErWV
UDtM6b2ZEUDrJBlEemDzYI3a3i11tzLFdID3PXdCgE/zrHJNM0WU2I7Sz9CB6319
G7z5tA+XOEZABETS+s7/EmtUYoR0jpJiTIPDablxXfhDkYaM8taCA7q72rdbRzRm
5G8lQefaEdHfeSwcF7DwD9l/YDsupQX1eXJw3K6Y/IxVMTTj9RoiDOPAxTMo0A0k
qLagsvm5042OMHUxYIbovOoxiSJf2DVUSoG1nyv1+UHFBWcriVs8MqEDbX2/xfSx
40bDibV4/XN3Lfrbb5jqbjlrGwJrCfFHsXprQrMaIbnDtvLdJ4gQpIKmfhCliZO2
k0woRC0zXUpt0BzODoQ/0v01zZTBL39vK9L08D7rS3wXH6Z+es+wZxFzmwIWGkd5
uEMZ8KO9bxZbqrOodqCUI6ZdyAXLv7JQrI7tQwskYq3q1zsHR+XevQt07yWV21hl
BJ0MIdjNetlyGw5H5EQE8DeaBeNd6bkoD7/a+8QD2b9MCkg1zhAmu6xCr3VfWR11
AyvB7rS7iQ2JgKb/5z4rZnWwkSTNAITSV7LHjFuq1Se0t6u5RFo0UAqGtZzN4aR3
gFffuWfe3uaeRcoz5llO9rMcweVD/S5DgBRVNS3exnXoPi4K1qoBzWUbVix4m8f6
1vabHJDoUWz1IlQvXnG1Y7ntHGjM5+mfemyz23dWdj3elRjGQpfvU8H44D4w2m46
9SOfLV+QwI6TIGwuPD7998yjisY8m5/FvDty8sowzoOze7Pd3LA6UvOGj8t5aubO
r3U14IB9gdnxmMWKbhUoDPhVTOUv32ou3IjdNCs/2wM3HJI9Samn9TC5orl3Jpla
7u+9Bg1VySF5ylB9MrXDZI2A0xfJulwRqtob+4iHBivZ/1xe/Jo30A3+tFN2Pp2h
NbFCDGfNwX5Ws+1RmNWnFmf8iwnPWaR8zqXZ9uNR4ZA6p9DGQuaLDMkJ3944TygE
K645/GSHcMrJ7pFltlDqWLnAGDyEdYqgks2ssuqtLCsbIp//U9hudBWqzi6xaEZv
5x9uoB1CtbdG6WZK3SaCloau2x+O+NmD0K0yQKH/opeEFG8rHHrrDsHJkzGmxZu+
vmwaRmDu7/csWC+7/thqjIUDocsLJ21pMJWviLMPqc6r2qfDqQW1vbculIHda93b
BMTGz7Ofb3acj+d5TT17Q98wjNnnoz7xYCLMPQ8AEiW4HmoXIr2cxAsgrJ2eXHO2
zsdWeHwrC766BDMHrO8sr0aghGFL8HRu9jdBI0pntvU1tglkTg8mN8WQ07diMYLj
Xujb5yA0lRX8wGKk1vop6nttstlzE/D1fbVd9pbgM0UUSbG+17CGQtTFRGWtxEVc
hc7eehg3iWB8JnSklsl9Wj9NAd1OfbMo47EUK7pMwdEnhnDximLD0R9kwcbNvILy
0tUNu17JkfkSgDDfsUdF7+iuz5imYzFMag5FH5deDHtSa0QW8fqzDcETVAUGX8Ev
s1s6A+KhIZYvRsNC3JpIq6EVX4+Wm+2tUnEldBLxtunyIRwahln5n3jgrHpvnqrb
RF2hRr1t/do65ZmE7+Ua6zFXJYoaKwmkrq1dmaYimaH9iFvY1D5U7Q21RdzMpfar
W8P/0o9m+BGMu5oJRxc5wcdI57cn5ldRDdDkpdRm+ahILzPdW4Ek8/wP3trXXGrM
zuJ88xpFqJgJeEE51YDBo+X8iMW/gnRIx1LyrdWOGfPG5Iy7dWVqLSHmT1+FbGKb
cQbvMsDpL0Z7YUHa6ZlwIXelGkEbFiKvALnt9wXx56SBY8vCsdDbg6WNMU7IgrRX
Zrlr9hmTPzmnpt3ErtKCZ9SicpYD093noa04pMrdz/f0DtTeW3oLkW4aH+G0gFth
A5ucxbGsKb3w5q0jZA+H6Is80t1oPKv/NN+O2GRLhj7e2SjpaPbCh7SKNhNeTov5
oRYs1H/dtlPC7T2N8hNcOV8shsDZub5QAfwLA+6AbVJJpGW3RbDj0cHFdxQeG3Qx
T3T4Q5urNd9SGP1F2sh4erMrd++zGycWOynQp5nC8x6CvpfnzAtJ/XF5YS8PkdyJ
p7uqEMHTUpJ21a5cVSRzA3fL80ORw0lBx181G5ZJ8ozoDr2gJ9kFIafZoA5fCq7P
eG+OO/04EMQfdrQSvLLaxQgeICeoB+72A5PZIXWvrczkdq7+uOWqJaV7ZNGPsJGj
tULdp7E8WhRn5ihlkWvZF6+DFn+z/sJLEFpL4efXFHr97l9dCVyiWbPh1F07ZiRD
GPPyX3/EvoGip2Qm1Bw5m1XWX/1oToDh3uAyZ+sxDIIOziWFiqj1sqCgX/H65UP4
8dQLxl+wZqWYvKbWt1U+z2vb1YM2GT6lzeDvixH+cKuwOK3mAagO7XFyNqJtWzEA
iboHtto1oyaWz0F0CZsQokJj9kTOfIKtq6kk5rxqmboMsTmwPkdhdyNsUe3K66kq
VUTmpPJsXRD3MQq9n5udl7mpWguzDGH+NbPs7UAtVz04nbaTF1sU6uGhhqtRj7+P
Ourt0PdC51/Pp9ujLhI6SPEcaKwsWoMR/dFLxDEPrDS0D8sZh+DDLfRx4ZUJy7de
fXNcWXh4dD/Tb9ggJxUm6tw8RVk/eZm4NBdEx+zC2xKTkT2yFcuG9zWuGLGbGwqL
aFegWdSgZPOR6iMjU+3UD+if17imo6H0GFau2WXp1L/MWRUUZUecxwTb7dg55joi
tAWCgp8pndccjsmeZZKt0ZOYFruZwpFnBdB6j53vGm/c9uuFhPiwE2+pcUcuHcjY
aZh5HXaV0orGb9xmC5ps2lhrWgHVqd+VqGOJ1FEVYj635wkW4jd2NU9vfBviS/4+
WabAIxxPDqzoY7ghVbJ3pwyqzh04yVUdw2x8I6pon81K/svVQmNbEZv/u1iiKRSJ
Uoyp8giQUuXVPzShG6gtMrxJ79IkkfIsJXAnTZUSJMFE2kCKZrsSD4rZaZW/FY4M
S4rkJy46IjttN2Qx8MYejMjDp4Y4y2Lo2HvLax75HJMiHTT5VmORvvEddDwLBVo5
ouMmxbK7GZehBm0Uqga3J0j2xEq3fuqB5nljU75Bl0YWP+IFRJT7iFGiiFI6TD+F
0wesjbwpnat+QHwaHYNu85eocRWannLkeBoT/ZXhIY2hilAKJ8SqyQs3S4kDc46V
F1bv04hX7MO+7Nfn128xmaFSvhtS8nionw2xWQdpVWlLDd7PXqSJkHDat1xzQZC4
BYRA/VnRxsasDSU3yYU6J3HG/Pn7wNwP9omiiQgDm1yVm6+L2J5YZa+Vf2NXEEZ3
oTkYabpKE57mz2RxdOM2Yum1xHkcpMGKa8Bxj0MsHszMXWbnWRsJimHWGyhCVs/7
UHhHdTPbHqPtgZish0MmONXbHZdomACpYwA+MNrtYlI9M0asAGLYrSdOV10p4lw5
icGULdSp9Rk5Q5+TE+0wcR2ZdCCRu/J6+ju7+Z0RBO60fwbGeXH3VInWGbmGumIL
Q80ZKyugLcLpjas8SgXXWY8OEWQLIzGXYLcngNVLunuXX65Coe9Yult17EMZI9eB
i3ikcHpxlVM8ELtesYp0F1F5k++HMwsDl3QMXHmG0S7CSMpY5pr40nwcAi1R/YAc
qVouwtXVKzZZv1FLVYg+bX2/F29YGkQGAjnhk3CIijAuDQIoEd+TbhM8z3L5lzNf
TN+8TsjNmSzRtOWA/pKIJCpss63Ms8TwrbwdDFt44oqBH1cm3PGa05D6sl35e618
V6QMtQzczcoqnVA+KZ+cR87g70V48Sc0TkX+F+FkckkL3cJjqbDzI6cwLTzCgs4t
piBAXK1A6zIhPDNxr67SRPovZjw0BcJrwsS3ru+NMZt6kXyEppUGZmF/Z4QBHfjM
/9zoHoPWMXaDy5vjOilREDG935whNnnnOITrCTmiVegYF4GZfldpUCkbi2wo9jxy
L9g0GpPoBl+jMi5cVZA634VPAy+ILpRXLeH54EQsh85YR9phzmXvF8aDmfW5GZZt
H+xG+qXeWPhLbF8lYDKnLLqO5ODDMfGudBsgKWTeS4NPgUtJbNG8ipgZAtvlBpuU
CXUTqD3Gd4vJVyOkFHdfSSFM7pHRc02sXBTLn3gH/Jq+N0KClTYU27r1DrflEUSq
zCAQ4R4S1vcZqUhmVbfnAaKwmGgSNSbtlGBKlB5Rbn1pE7UqCOJP7U9Ifeyph0Rx
8+SqzR+u7kJRwFF5XXv7WL8CZLT+MGa704s2pxqnmDidsdAnP7KadCrWVLT4cTtJ
GB/5SY+TdAH2rWsZPuhMHx/BZJWTsVv+zdL4KPcw0r65ElNAYB5g+J9ctFkKN9so
raeaBcLkA9MoQcYlQCqw2ar7BFPOKKLB3OTcHqsD7tAWdJ2ZgjbD36rBy8HE29lM
AM7YLD8uk5KhXuY5WjExl/saeMFJP/nL+hJXZRwxByrJ6zN1qyStqOEe+RBvcnEf
36rx8bKXdSVbegkrohUcfn+88SE1Ksvc6Sv054FUEQ/haa+3aNXvqNGFV8yaIsDG
Wvc4JW6qIXvSWX9wZRhltTffnJfuYVpDmdGt3cBQOftcytq2mIF7NW2v7rc2jA9d
CtM41TVGbkZsvVe4lspbxt5CTq/SX+C+vzpNZ0h5DJF3L1KMMriWL/xTcm0AokYx
2KuHz7sy/CZv3Af1Typbd8tU1loDQb44yGUkTU1KaQiMTPd8tvD+3+FHfFuNajIP
+nd1/23umXPWYn1IGMYxiGQ9KTULkMLcCuy2U+ibrVxn6oKIxQCupFVmXp4T3ycg
jNagywHWjAwzHae594l6G8E+9KL71k6KGE60ZOTDx9n3aMsaL0os1aFzj4yHT9Dr
0dzTRXWclz5z20doyWUZzKu6tJ0e/gOM4nrQo8ubENLajob14O7cYKPF5ek9CQT9
Xa3GkqbgStVxufoIr8S3TLOfNTq+PugjWYCvEsjlAVTQ0a7upbDGbrOk9H10mCU1
MCrS5Ay0a/Wnz3ebB3frm3NqCym48bZ+s3P/odI8lDkQVr/DByjiq4QRBOlYYOiw
Wbx1kgkOefYzhIZz6JLoyJ2hJ2RAxKVE8v4kp98KVSphs7TWXiXQJqNLOfWIwT9n
hFvwGZYBiMflmPM5NG0eHf7PCGUaIq0mPnMpSSZbeh9VNmrqG25Xc94rwo09CAr3
qR3ugPoC+8dy28nCTStigXkhKcKJF8BuDGTeSI+x/ekCuBuEt0RFO/U7Y8f8nI6M
eqovpiDfiQAwEulahO2BrH68gOgnlZL1lBODMaJg5SXS2mYUdFZ4l+uO/OzFnHhr
gK4SKAOdhE5APGsRw6N9gsL4Rc6Bzey2naywmC2rooOtB6yzViv2z6/mSUjE+pkE
N/d39+P+zZwzlUM+WatzF3NGtYiBzrWeslih0qXnXh9ggr418aAB1byPEls0QhRN
pA5mjL8mAvvEMU6q5EbSsEXQJrc7DzJ1MbhDaHB8p47FeRdotE/eVmxvvlH8h8sI
CBm/QWSfMBuZUhM0/2dU+yWYN1GjNKo62PRID334dQxbLOlL3Y3p4hyDHbL7t8RI
3aTvmeIQAPPR6GLgYszoLdr8f5ZHEOMN433req9IrGQR2K84Bd88cX9neVysWsQj
u3XR8bUSGeptdT2SiXi0FbnltfC4Y+j4LKFe4N2J4z1DjtVINJW8/0FRJrniBTgt
b3Z/mawo1qKlDCuoO/owFpqjTUIRKAPSdXr5P4SjHpQWLlEDR95oZV/GL43sIZZw
QcLIWKX0hXgdxGZpAGRonAzcLTAChoDgL43RL2hi/GzAJ6chESxz/31LmYInS1iL
bl57fQPgiyYQCJWsd9rs4FzYji5w8appJuh0M5yceNGWrKBUtjsBzdXjrobXw+sB
vRAIDbGH3nUDIE9ymh4M4+pGvilS/rzKK7yOBY+MNYaEoKm3Rjdm/9MFkhKQMQ24
rLuUaHG8MKBtj26c9JVRa+QZypETO5P4XTg7eteUOpoC6h22hlQ4/6HOpqLjeWol
WvzDuVN6kESrtm+XHvC6N42hTNGZWfq8Pw3MV5CxFl6Lxn94hEuhXdrtV7rGl3k5
NLbn/hHxn36NCNoqWVjjSqvuvnxvCm+H8Z7MKuNX6VbUBV3sLbEZ6Ad6gsbCZf0k
MYKyb1S5AVMEQcL66anXAHIcy1zVsjiCfpgpQcw72+fcVU7IHcz7/J0CkD2r9M99
BTSFzYISAS7aJaVeIsukxnh27OrnH9NpgAA3Tmv+a82j85plf7zEEP9fZ8TmGu4i
2u1h3mV+mgF6mikqQhAmT2txc5/+hEkjWmE+yyx9wsA1+q3q2PjaCLurFSiEbOtV
ZBODGewmjLjwmQ9+eHIVtBaHvoPa8hvAJnuVaCiRaJnd+bzu3C66nZu5TaOVHbYf
EcLAPxUvKdgnU14+zUMp+P6hAKR0VedVaLR/dhDtP7Sj2y1WHH7AHU3WdzS6tRXT
jsTJhqfxmb3MDsvDyP1xZYNwBzFQ2uupVW+p18S8zZG/apItLbHEdzxfsTnluod+
Df7zfZo8SNKghQ0YrfxE1iAUhQG7/PFQeGlT8UWHOL0sOhL438av3BRmBRwtiRb5
Q23BXvO2QD8vS8T8WOGHMdPQav7qsEZrbEg4nMM6q9+2jD8kNJZEYdDzSIWWNw01
kw8dua+EJYvDBrgb1hpq/KlvM0JfJlFPezZKxkCP89caD87c57Ww4vvgQEscHK0V
R9VEPCSCaMWF19y/U3I00xgPrEUafMYCeG0WFbE9iH1MNisFjMCifb9Uhqgbn4ZT
cZzhw9X0GNZoJQH6EQeCJlU7p4uqqp0xyee2wXFMpG1Ha4k6oi5RpIwWS34/H67e
8SL5vCxd6FNFVCek79hTwWjkaG9LU50rKz/tV4geOH/NvmfjAfc3og5+8HOtrVYf
ZgDQyOxMq+5VXlot+RGQt4rDfHbyOsN6FC+yx+lI9MyZRDEmmDYL4Z7w2CL4NNE1
ddzF9Cj1oimwB7BXptCKUYBu3RRMRspeALJFJwJkxfO2onmCNmcrVM/Y2Y9ZUIkP
uHaUoZemq4k7CtTNxM0Ulu4OSBdwSi0Tf85Uy/O7QDAF7frWk+IF+46Eprvn2B10
LXom2sU28QEBBEzflShGQiqR84z79Q1T6DWHTUh3E9+xBYTR9jFDH6E5mahEvwpz
kcf8hjy9FbtYenBVrzv7jQBHaH8xco50pQqUuofVJ8QtHDdpZdsTSFf9u8xFL7GG
cm5lv0oe9MkwS8aUE9VwEy6bJmwYhM7Ki0FVgi/tpePC6ZSBPezJM0rPn2POPvOY
WuviWNBXl/NePKrf2CtyIMEQ97KahUehT7+uLB6eaNGqI+qp2XeSi1q/QGt3/pC6
lOffj+UH82YYp3SNdoKitNHGU4r0ywxQgrCjw/YS0SCeUlaC7DNrDOXy9+rsVvAX
hruhGui73WZ7RpZW5moc6ZE9mOL8C4hg9kzygSIVlPVHPmX70A6+U47BPBCuQUNA
tN6N1CPLB+k3dZCyz9jyto2uPs5Br+rrmrjUEkL9GtkoKGb1h1XFGQgT2WNGwPTm
T+76L3E+bcyvHdnSEpILzEXG+YRcjUWgnLDQdkyXqOzqdLGjJiVT4kfSTqA/QQCN
Jvg1k22+RVq0rz0u+JcfTlTcAPBaIy5NLnZWx6+o840Xm/Fq4JC7rJYd7LdH7wTf
a78MKjTn1+IsjujO9Q2zlX/KQq0zHDhjP5eUjf9K4ix0M49iBXFph7tf2wAupqtD
6iBGXfwq8KNtsF2+OFUkeU1mUnjXuPeb+vYSu/j35zvVCc8LnM5z/ZAM3fA+bys0
W5FTUNWVAXz5gRF9OyVttDWpjsnglNJ/ymf8ujsm5MfRaGPhgGHB8Z5z6XLbkJyI
uT2j3DABq9WmtK7+PBzXZAZUH4qmimbuxFJYRwVr5dj4PHACzWsHGS/WHOe6IuA8
k/SVO0M6l0j2WXlGv4rXHuCXBrGXbQUIYw3xE2q5yNCKc3F8ca0UscSRaSpoFTR/
CeTNalCMkE0V/wgBOhPrBAVn0J/yutRrr9/AqfvHYzYgkQCiqRyNTeLWuTIFHH56
ZQhtVIuw+A51Z7p5HKgEmJlkJRR9MM7taf0Qax4BRqGg24o+SCVhM323tGByft2X
/G3JvpamFynEOFBOg4jL4lC5Z/X2uD5veG54XqoFLCOZ9CR3SsNp615DRHAYdPd6
+xqf0E5VRFYgTH1trdKSEgEI5ouJDlBdT12qH/ah7i9m+GnybJG2WFOpyHItmlLm
8PvQcrQeH+N7yNo7B3ka+C+SgZ0zlrvuhQBsVZpZ/iXVmlOvRMamQdByDhv2f5YZ
giQqx7t1pS7TRBJ3yXBO3xZPInVweTqMDIGYmc9Hf6ek2t8z2Z6fAg+MBLfpf7B6
8tlFrvQsygYC7obMdBhn9n/Vs94/evyuPUbXxteffNARmaJftBpAPO0wrXYKTB3y
ecigGam1r5OOBx/8dCQrjYPmlpCTthuyBR29vkBJ+bRMq/IxFwWba17WBOgKqoJS
h9i2xDzljeeLZzONMPwr2sc8Qj7B1RWGB1aLg4iV2PKWfJPKm9jDA1LfRBpNqSun
n2prvWGis2CPxVz5oGXkz/opOXKrTGA0sRa4P5p7STwzrn8k8Y99/0XlM6BLiaZ/
S05C7SVlqUGIx1HUxYcP1ZBd0g60Fk5uWGjgl5gytkyuTYCTqWtVO/gcWd2zxnn9
SJFztrATHkA8LAFgVNpKiJAnk9T1DBSqbPv6nmbgudlZbWjIMa6WMW3MBsGk8Q3f
mxnBFbJF8W0ERxDaYY62DgWZ91jeH1LH8k28UPgTbpe73P8UIyIVhn6l5w3Ckb6l
fZISdlWhxiRvl+3Zpcxa6wEiCqRxt6nyEBiwUvonBNop7uM4yVlapbA7sTG8J3HZ
Rz5qIhvpX+7d/D826XqVDBA8pyPcd361MAF5iX2EEsfU03Ti6dTKzNYwv08Q0Zf1
AV0XK95S43pJeUeyeYl/edueLmJWEvKj/w1Ih45K8XVKTFU+wL9OsLUID/nbT4ab
gdbI4UCMFpNPcZ/dVBMfk7mL69MMc2KPvmzOqb3hEHIB0dOa4YP+JY35ObSlnlSU
u5k65qXZ+zoY8K+RkZNMU/YQKPsMxHt9WBWlIs6bZNu706+TrsAWL58oEK2xGDJ/
Ge3hNjPLPbsSc9xOR/RrjUNKMeThU+XTfEKeNI4dJowMLoOgiGqHVxArwVQ9J5vl
2dZGR+ll+XPHOgvL1bhLpMuhmP2/L6+01tc0EU2nB7DU8ZvZoBwfma2uVTu6SLBm
4/sHU0nEW4E2qgSBJaZBB3d6hIaHkvbdiNRRJ5bYLAAgcSOBHR9v9FsFHztHrnxm
aoF+HeEnvXjfjiVHarcY/nTjdy7kjyGsmI1luwsTFCHpaOv+5ndAjT1c5F9BwefR
b7QzHgSRA8L+c3O9Of+obflJMB/zc32Ram4dJYUXzani//RsD+ioOgpYUldFnX87
jeHGwHw26Gw0odSfRjpq2pm0iLCXcIeQ+rHRE82meOKU0a5iX7/DHY9N2tX6561U
iblSmXci9/fW16kAtqYelOCr4rCGdKk8QzdG2er89iC9yKG0l70BzEuxL8UX7bDt
hSxenKoaNzFVP5Gm5exjl5tLu5tXOtwHX0cnq3jjBh4lFaio9a6VqMp6iF7k5iQC
zDLrPGwmewgAGWXI2aQA2sxm/y77SHpdvxosvsjH77X44yYNV81nL0ZhRYhkcDK5
KDb8ZUITW4S53w5xitCYgk4ZG6q/JQ+TdOYkJ6kwUpbKL5xsLjjNtg0ykkoIdZKu
+ckLALWMfHzGxa9iPW5Sip1Mp2QuTcltuNUb5eonXXV8d6UNjpjyZKQcQ8fKj0LJ
sd8Z6cHF1rHCFxopzkx5xvikuiofDYYr4T6VnsuQcJN22XCJsTNqr8YjIDbvV9b4
jxVTpqVko1HSu/BYXL3N4TxpGN4OdMyD9E2gPFZHopAmn/Wli+H/ohpAMJFmU/77
ipZAFI1yfZV3pd0sL8rcFNemsiccgshMIx2gB+pGkEUPF3NSe6D1GDnrX3m8evId
zIRNbkLg++UJAZftBUntJ5jsrxKKVZlNoO3aA6KMuCbmtaQHoSZv0yMNHgaaeniE
Wka74vVHF3uBuboz0yGZu76As9jZ5MgnUevrEoa25MVtIyIF+ziEXAZre+XfareE
ygQFltou8wtnV+Ymy1VhYmJtFi3LNBaYb36wDY/wLziNZ3ZPr3diMqnvKx8RQ1Sv
BhvdSWFmiKHHIbalCNHSJ97eWLZXIjMLuMIS3z2RgLTg2tzJEPrn1YkuZHoEG4ui
0K5Y/2rlVwFN65suGQIF8iO3TjGGrrtUy0qQorA+ZkpWx3Kacm8GyOMgZ2IQQuSI
S8zXKHVfhPnggSs5AXP4MuNJx7aO3ep4aqfBfkrfOExvvvV1W83bkhXY2IPeCy8B
98AbT8xYhIv+snphyAWvAH2pDSIHybH/wMK5x8jtrksNlWrhPKLe8W1uA3pTK3lI
VU1EV4VIJZmBkuY1v63mrFJMLUDPENBiX2K7fSQvCIMQmwGXZjPVVLqA0hjyJ49q
ukEKXc+va6bGKIqZdjyE20+2Hbay7bvvgm5kEizNgVc3GKZxKcoIp2uDtgsx4r5s
Dxb3uaLO1LgQkAxrp6knGoZmC2pW5+g8D95DD1jHgqE7Vw5prSdcysouhORftO9p
SSuOTusDMCMFh/S9zALXmeKfdoyrfVVI8YwfPk6e239vmrrn/IaPirS61ru2Icnu
rjrKTqIzx6rRPJilYvftBidB/T+l8lStW6NR7YGMRs/A2ArpMDPLMIS7qIgJQwkn
0d4TZe1Id0fZK1aNwj5wiQ1a26o2LP+E9Co/daXh0oNBv6gmQMYXn3+Rbed9foM9
sHSLn9etuBwRzGb1oPcm9jG1gs3NHqr5ra4jgvb24hKjCNdN9XJo4VVdyTm8PBlo
MN4sLBncqPq0buXYJ+oj6ZVt4Sy/EVvVruwIH80HTOSKzEA4G7oso8Ff7OO25LMz
iRejffcIbqwJ3K5qKP5krdOavlHBXIrVAXUQLXq639+afd+7qo611Nqr4hTdso9G
Ji1XbqhbtK+/y/fSlJmf9atmmKON0KhY8bl1Gx2DOjEiaySKBd4MnhfY5ZsGaRzC
U29i3bhgR1kE/xFKeXrOGdqvFIBra550paJ91lsPdM1nU/A/rcIT9BP6U+esfszF
JN+YZDxzup7V7kii2WZ09sNKtFMsGrrLER0N21ETzYwH1xpIrbKhToqbrog+1C06
8XI9BEV3CgCmrntS/bduY5ZIdFTdN1Fsm8eMjFzstORTbyf/26hVg/1rBGz18B/f
JxaPxtc7M92wykIObZH20bemXLpEAXxsb6BE2H3Fulv0tgW9gaPN/Y3i6kL0skme
9FqRt2dPUiknFfXkbj9/2fxLFEfRbA8VLCb7NOvCtWtgD8IOgSLUKOEZJ/bTJbK2
0BmcdZ27ynPlgHKMbT6yCUc7UZyWOKxinPDaO2QvYy6D7owl9mWapvoLIV43l8vW
d/7eznwcJL4I1cD6Cas3XN3YfTiNUvxzPo4o4d7WM5QA58NPnf3RsPHiufaO3IYS
Ugoybat6ykwG7WqpIZY1NuHi1McNvqZ3DQ80OOOEp6nl2czqonR1cTT7AMd8zGJ/
wYsz3pZ7U8hwkazDEtVvzibMWw5Ju+h5oXp+QKA1k/IJGmwkaWdsobLe4BrS26ZH
WkJLDeuTdN0fHhtqY8A4AQgGcWhWsSoyfEy/nrQFpwsLk9JztYUXkHBY1oUlT6yx
zsOe8Vz/PSxQokvUBTv1sVIPUBDy2RDjy4F13kfZ0NHzQ/UmD13dFR+FS4UICfVq
kIFhyPhJ0r+OZ93gcDSrYQuAaOenVhp7sXcFcNvYkHRUAC7O9HnsO2ddGphB6ZW4
pBJa6dWocmRDlQ3W5OXySdwRtSXKlwkypE+L7wnES1Xa9aZqWNOOYb7emzAIGFGh
O5qG+rRFVRze3/CSUXJPWiRt5myiy6tJEdyTPBHIUXHcD/VRn1R/k1CRgKRly3Mz
5grzBNhzpM2WOSeuqPn37xMr7o8vW2+HwqkaUoSwZNvoArry092pSyruGuLpaxrQ
FVgyAXSCnkWUUQxkmNNGSciAAEHvDyNMqxXpbuDHan1gcv9HzftEkoZlrigT74ay
ZFt9YURxrwKrah/E/Tb0ilvvA++sQUkVEb7uL2oAiJOhoppDKh2Up/8Q2zEy6dB1
kHjeFF8CGlcT1YgI9jX8FWs+Rj+J/zF8fcI1ilHfAEN+rM2GMSSAHGd+xlgbH9CX
cYpI87TQ7zk5FzYrM3IARoihW/sT+PccZaVuWDG7mSeK8Jz2mEsd+dd7ZAbrcQyV
TrC654CAbNV6LTvN/RD5k0TUj3xTdXQm3us3U8K1qWTg7ylLgQLJUpqb47UzcBKj
wt6Yr67kynZXghb4DWvZ5fqbU3JLw3gDmrnToBYvz+2lSDg6DZVpJHxVngZjE7mq
16NzDd+jcEGrqUFS+uoM/iOhsr5j7ZPrCauwxJnrUpA9blqzaODn3gsFxmOKQov6
5A3d2uRuPR1N/gM3R+xkLSoBlbZyHHnftInYQUq93SxS90bs/lhMnW70jw/2BfJm
d32lB1IYXS6VG2eBGo6Mg8er5Mmt0zdJF7RjijVSiHJcaLSxjQYXlGYitb2tGZub
bLa7kHV13DB2cK7cP/U0gcaATWUhSt5lCXskZvi9tsu2cF9PDkICxA+eIbu7Qoty
vVYqVxr4JXzpkLv8NQ3RLKXZH42NQiydznZ2WK2WjGplBq9hmJE2gufthc/YEfcd
AEnhpFn0xn9C4ONw04CKkdIHemnjGeKJm8QO2N7cnokr+v387izUlvBUMORkw45a
ETQ8QbvmnRdlq/3QzZUDxfZL3+PSm0pei3OnN5yXDC2GOZMSgu7/4uuWez0W6/ws
KzAu/dqeeYby7kYlnBwrIF0NOVGFENuoru+b0z6ohNEec6W+JtoIxZ0kPBCF3WKu
YCpW/K/g5FJrruEgw7oNiaslveq/Sjsq7drH0gYB+G3sJXVY7D9BV9F2vA/4krKL
gGSpmAWb/eyOLQp56f2vedPjnYX1FO2c9JuvLLAD6LZTZ1+5+NGsdfm4T1oFx1hy
71lV/ghdP+AFVZfaG0QkBbK8mtSIu1LXWXDJxNxN761uoNMyNaxemSGHjBU4SPkk
53YzBQE0ZQVdmOtbBL9J0zyFgi2XYz4KCaG53tg8uOA9ibtNzIM96YtXMKcTPWoo
P9X/Cq95CRbE/Rj2RP13a5mnQ02i4lWAsDY/v8cUdqWJfAOfVt3AgmKczmgp6GNL
QccFUw3apJjHS1dkhFwBTyTMn2XR2CL/TtDANg4+/BVe4ubXClSVcjG7WoIQq0nj
nfEIxkKF+TL6OLc1TmC9WdukxZ7f7K3FYQH5DFHoGX24J0nbL3j9IIC5zmzN6AvW
rxGlATJJFAoj/i8PULrOYtNsYOsHzFxCvqGINNpCp+rd0xBzD4viBf/7VK5wgHnH
XmW1NYouODCBqGo8rc7uQFH1wed9ekJU5/2gEI6xRx9vqVBCfZb8cyMMhEjmeTei
DhcvL7zl3iv8re62TQpGw/qr+ZGrwSOppn+o19HDtE2qougsFhVI6E4C2iGtgqq3
UPXFGCj39ETm1IdA0GLVCzKTO+DHjZZHewUqRGIfr8018KnI5DitR+UxxmY5zc94
Bnfp+rvzib53KhSp37tzlC4HhJ7YxDNgvXFY/U3cvbQoBz6gUkm18RBm8p3+5okH
ybD8vmndwhb6Y8o78z/EBkGg8VXoIei7a38eNyu9iEwStd7xdtMCw4+q0NbbPCC/
AtBHKL7bl8xAaApKpoCj3HqAjDKoZi4AQA6z0uFGqoS11g04Eb30gdGTuT2jRq81
x7yMT5xxpPFHMmG2bMvuFy1PE0V+CFAKwY6l1mfTGvIqLV/9V5tBZGBGlLZtg49+
sAEYjw6cC2DHghmj2LL/aezN/HXR27IMF6J5kbysIWG9QA9IifnX+p1N1HhalvXY
cJY+PwRQwwjVN/N+QEgu4gBrPKjzURcsyZ6CBvUetKWhNEtAEwjJHIb+BYOFc8B2
BgLC0bIoEjqxxuYKJ+AzjR7O97bOqAN7T+jf3F+L/G2txdkNBkqxKvhQ0/EHhZBE
Q9TBmhJjBESKwWpwlJpDg49T0p76uTqiNvr5iKsvxh/ggZfXyEDeJsq//16VhpNc
L5gnbeeQ+nCCa0njggmyc5KsUTRKYRdzHQcrcOVkAsD+o1rBmVNYSIWoYyJJeKo4
YZFuWXpmlut3+fiuvsjn0TXXfOljsG51ZN0Avy1p7Gx667gj4RuO8cfQffBRmOit
UAOMEA86CGeZI4ltgP1taYLMyXfMTqvz398kkOKGW9SHH/6aXexWwuoOD1CwQgc6
zokggTDIr9YWVIsPPSBgBqYcnjD4RVVO7YZnTE7IqXnJk3R9Uihr8dKERSByyNVs
5IWxHwsmUfKtUHVkRPvPy4P6ArBSbXvw2XciOFwO9vqiM/I4isllxXrxxj3GgPpT
TzoZQf6EaSLnLI2m6JafP1dVBVToHwxkMYvrkDLBkHeNaGinoj/yjD6YAM9hBTIj
btDL5G+hTwiTMFsoF25Bhik9CcQPuPMiEa25HcTVgnL5GGNOXPnFUh+cK7LP43sY
9Y4D8MYmKj9UjTRuQXhaX8L/lNIf6c4fnOyDhF89moimMGpYfraD6N+xZ0RuQVr2
uO+W97AOszvqM/yN//yhkMdT9U9vQOyDsq1caPFispRyGOk+b6uFpFCqPJLj6Ca9
XF6pceYxBcK5qeQF4JtzMpwSlhypNQ6vNKWzwlb8DAYS/qeCjNZ5rm4q1aETWqna
OhT+NeW5mKQREDjmO4GKg959B5unDRuNRNGVNLzUZVnHmjjzxVVLU9vDNCwFCOpg
VSyPO40X+oVE0BmVY48gczF+LjGsuCa8xxWrAw6IXNKkL78Y/tTmsXhjcXkBDUjx
WozBkCizZiiEImKZxJoKgdzYU9lwqoxy5hzTw2WdL4kG5ZCq7J3/rEtdUi8ofUFr
xsXGbBb0muZM/qSj3ATke+2T0pyh7U+dVLsVq0+8TCRhoELK5YHtvBmNjVjbgTcH
R089INLZ4uiGYIAxtO71k6h/vrGOpVg0qUna5diWXZswNlLJ3bJ7qAwUP8RYRfdz
C0D6KBnjThOTpygS/LiFTlfloAAbB8tLT9TFbsowjtU2kSU+Xc3CKz3ky0V4NXeU
dzGWtmqnRdC/QYN+DD7z0LUcGNck4AGykiI9PdZjsWSCvYrJnfXo3BvdkgS77SPd
tE3UnPIyxaD13rLttH+71fNpGlNg7ynAWgpXAnmIgJi0lrLjhqW4JRov8vLXxOHI
wO6nfG/z27EA8TA6MsaZAqodQ2acWK4i2Wyz6K+4m1fMLHV14D03/mEWs9oqsd5v
Qrj/z8YWeTrGGCIdfl4tLa28eWi0yxWyz2Wq8y2aoJxDFZci30v77pBNaSJ19hQs
hqil//ZB8rsaLW4YaH5SMxcoVM5vJCDap3UcfV9TYzGo40GM2UJwRipufB7gzjRJ
GD2tRi2NpEAYOmQZw6U9avAbB9GWYvt52Ddt6rpj/IeRYhI+4PvSK7Xa9B4Prxpx
jHLMAKEbfOahAvB3vSecWQX3K4pmpiBLlBmV2ZkruA1d8JOOCXY3Cu1DQgSsgbJ9
prNmSFWXqQPpS5aokuc9QFcGk2GBTBGeJlmkBHTdJUreLN1qsNdM9I9eXb9jiROL
HXm9LtAjddKuq/rmgB/lgUxn0f2PwpHEDHqg6U3/jsrcvJ+MY/2yhfTqV3GWAHhd
tD17SD2LQ0qCFFoDRxUJEL8SbBLkkQSw2e/58JzttDG8TM/0HLhBL3+Hswy/Ve7A
fi2I86JyHMUoRSI20Z9BvbyWuvTnEa3H0VZ+9jie7aKs0xlgS2omRpnOXikGvWC9
69njieaDAGbGZvXEeveU26/YmT6h6SBI6INerUUYg5qIIagCgV1LjObhyohv5iKE
J49nJgDETTkK9aUAsjodLzmexqKUCotkEhqvHZ64zQJk1HCEIv250JWQGnVfnPTS
+VJWPODKoDDRsNOsoZSmUKpJVvM7PyitcQG1bkvpMxtOL5luO0PXQ1bm1HMwJIF+
Q7QUEJ/P+V8lS5o2I5IyVuhGefCGv4lpEFK0zkw5oxFkb/5OvvtXptVV9d8IMegO
F5IYrmUPRGIdQYm+GoGzAdxnRm8uKeOg7XBP1d4oZTG5x2OKpsindncwt2kcMpmS
cEsVyST+7d1IovBzUFU3Owm6LXqjHUH+yOzlO3V5+bcuyCbBlBQtBbzpWcBVcqjw
6IW3PsnIKQfwdqG87MeARy8a7C2tZcfGqmpfU2FqXVmVx9GWIB73me+BVtVa88Nl
XRsQIYNRghbk1GhW8Wk9ueqwizB27KaElqB6ZQL4rPS9ecTu3FM8MBU4hqf0phPz
m6EAEunqH6GyjhQVcB+9Xzwlnkq8IVscIuzvyaXmH/bREooiiMNPR2cgJH8i3+YW
cLVS1r0c/6m7lbfuUiZnrqtRJ2FcCl1x9gqIfgkcSR1p4KwLayJNxeTcaSvnH9xq
89dvB272qiLx16sNDI5LOaS5xwYmKLgE7roR6nN3g2MZDiY0gFotkF6LEjze7g50
3c7AEQE+p+1hXNSE0N8/M8yF/ATd+Fu3jjCkas4aXVAG2TaVX1gN+Y208uV9O8SX
BPmdICteiT2DtUsJtGGTaCUVkm3SI/LH37Bsu7u5Z8RNySw++xZy9tDg23IZvqTh
1ePum/+GhS6yceLw4VepkkESFT1jAjhq4G8G/TegfbCbsH/FWp06Xnz5bXm0R4je
0sa+ISaCtYHQGx4ktUO9qB8SiFm/J2JUQLqK7tQIMHlwItw2c1CVyt4VL7EwT293
/FggCC28G+RhioHBZWt0IGtlwC2Idcg3I+uTb+S+2CoW2KMvQVlo7pe8NHUXPvw9
1JyJFTIYOM2Ucp5FmyUEw+gxb5oyHFroQvNTKQB66uryMxaVN9K37W0iSaNajDgi
unP7THXFBtZTujt7Ca0fx8uElk8oW1b2WX07Mc5nz7hQt83h/4haI6bjd/kFY6nO
ptq/6ZeVkI0TpJkh8BT6LS0gOr0hYVpLqR42BZVmckNuz4ugFN/iSleom5Y3ia+Q
/DM2lsYNJHDwUJcuqJaMl68SqXgl2bGvfRAnKGyoRdaeFDe8y3R59RE8sY0eeq95
Ais+O/VJceGPO8VdMTIxVG7B62OrM/CkNUFn7trX9oRkkTyvugmFJU4etRW+93QY
jr1B6fIA5QWsO25h+BDMDiaqfWvM1P+Fy03N76Jkb9yly/uqOJMEemXYzo3WfIVZ
FfJhDC3ELk3mS7s5g2QOzr6TSCWSkLeuU6SuQQSnWS5EyaUoRQ5GAOdrglT1ZSDB
R7ONkDli5WAW4IyYVVpo1WpBSrkGLQxcWn+J2/b5xGH7dpeyY2A9uNEdCpSFJNG0
U7NemLzZQqY0DCG1P/JvGA5f+Zs2OXv4uiHvPzFA/qdc80KXf3NjTFIaLAmwjm1p
liaqg7b4QWdZER1gb2MfaJdYHSPvlLaHhBc9YuPKpkXqpejV+Bu3Jzpot+/ifa0T
G9uXZkpODX98HBVFhgTkyNP5eNv3W7PzP26xulTy0PH4wq8jcqN+OU1/sysQjWie
AMNm1/2FBsC3Sji7PnswSJ65w8Y9dnjMkc0WwAQOYpjXA2wfzFJxesmHQQ48rQe3
UyLn0R4eEpzKNd0pjkr8D33ciyZFNyUGGf8j8LxJTTNGc5WxpUdEI6K01n5u/psw
fgCBA0RyBTw993EVWXx2OieDFFACVY4Apm8vBZq9/wQC8tExHjpiD4ipLAxcTZCI
qooPKfZN2+3ssVHe1I2lwq9vhskHvruAmUsmPh/zTjZwgrMz7YJW6Bba5Ek/iQiW
8f3KZSq1K6RLPlnXa/J0WOcivYaREu2D5aoodmUisiXgrruAuO/hIBESXJKMWC28
nn4nbwNu1SHlixHOueycNTEXwQc400SfiFcDiKmk6R5hZwDJLs7yyBGGWUnPEzbk
E66cftywgcs4/V2KTqVD4EvzCOoxgMQwyz251ugv4vXJWS0ylQICub3dBKmSQ9pj
7248KeNXz1IcNKrW82ia9r7fqAjxDf5WIx2LZDjrx8vGEPUP4j1k0DVfRw65P9Ya
rUo7Ufj8oVX5McVF5WQde1qbOVbrAHQoCeWfiqDHRXZBqdBAud2f/j9iurLP/VWt
5TKBGjTekE040suHe5q+C/YvaIk7xRjMHjV8NwjZ9GifVhXttJnHflYOvwHe7POG
B0RYgEALkrXKyK2WqCoMSkJRw+aBi2/ngvUMe/Ay/XeIIgLsG32o4wg4t8mXp4Bk
N5u3zfraLQMutU71A92EfYwJwOSXvasiAZwLWcpAsHfTkE/jUDo+cTk3c+wyj8Em
N5HQQxfi4GOcYX83q0RDo80qJg6ddQzsY6MYFPs4ke3FNGRHX8ZH/ybd3Ue5ye99
SxnnyoOyxI+qEb900J8aq3AP0CluGvZRLlAt4sjLW29hhIERCzkiZi49sFOmjfj1
EGdMuxbN4MwCMcfhrNYyqoNtUwnD0O8ERC7pBs9abTfzAz20bpuSbQAgd2+AjrfV
B98HCFZvi0WX3bXnGAW2plvsnQy28cjMvpmFhtp+hZUQgyBJyoFXcgHTogxGmmcP
DYx6PK41rPW5ia4xze9i/AdAbGXXWwEFXuJIyMdiLZTuOK4/MW2RO0FKI12EaiRG
tm20igvqN4LWHkcLpt4lB3Sduu6SKjR3Es/PDee4EooRAOMO85PSDVQso49ecnd3
wBTN0KDn/vRXdvFCBTbEN8vJ7Vw5AA41d5aEDX9+A3JumxJDTLZY1wv2S+6zfU0w
ppYj1HTX9SnuNUqup7W2NASQZLGKQ7t9g3q9DTZ3CqswkA5D+5DRYQPdQVwINPO8
KXakM+43qzf9IHxPApzJ4EovCc1fPpbZfKcF0hvyW9HPvONWwWCP/KsrXTZ/+1Eb
ZIRq+SMOH36eYkEoNSPpktuXIx8QwcJvQ7wmMRqkA8meZjlumaTuduMqUX4jXD1q
MFS7jXqXPMdcbqPUlaN/8YHH8wChiNWMyvzNCr48vsdmrE2vGt/nYGNVvMULtYct
NHiwejzldeSqZXLlg+PLXiI+0mrpmWsj+yjr/kqgXHJa1q5Q8QAQ6ob9C7go9Oqw
mlXH4dnImCj2DeWrQUrLcOxlw+iih07dd0CPHGEZIevI2CPBgiOKwEF9VVbRhXU9
ILlQ2cq6QS5MLSrC3uhQtnv/hW+1QwEtKaLhc1w1kBAQTmngzmi2OccwEckHDs13
oEnA06SLp8mPxex0wCeEDpWCJqx7+5+Q36dJvZaG3N1uPBSwfb66jKhPi/xldyfx
DsNtW3Lj/Y6TXQ6Kj1axd55TEE87G+NwP6LE3kZK94YPuXB/k4iu+kZ2i+PTRDUr
fK/NcMs8aNDY4Qj++0xNzMyq9lL/3++38zjwsGqQ7ZTdOZq5x3P8pB91aLu1puGe
WF2Ir/Vmp047zrKadlQI5uQ/mfJqnSAusg4JYAnaM+KuROEqkd0UqgvZqUR66zuh
ssWJxSchELELoQy/on1hMcpgFNk4KZahpYHzy5J7OZ4iSfDoqlSrLupfSuSLvIeX
FFSVJx2+nXMI0RZIm03bQhXlTGpwrJIJaACzEWrPcPyGXu7vg8a1dE06azgHhmXJ
9Fmz675I+GKnVkLn8AVBOP4nJjS0fDSSVMxXcHhBx1C3ZEa2s/xmXgJmMpA0wpAf
SS6f5cMT1Ny3LA86A/8eTqk7vpcvfItpJeiqMM26udkVBm3QWieoIa+JC1CiQR9y
JLdwrvfyT2et43L7weN5dKYx/hbGyW1q06qkAm95GWXgP7vAkIYJyI5aFcwZ8c9k
p5zOPG+feWIoVcMcC70mRChkhpfnvahOOLJbFZLCUpIeSyFb5L2lOw33LUwqLxKe
N+HJiEYFBS+kqImkYbGxDJLfnVHsJEG/GaQ1yBdwkpsaR4knGZ4ZTNCpo+RvZLV6
GnccYnIM7RWprXbuwiOnjM7EqQD/2d5FrFeul5kByAG8Y1Lrtzn3D1Rk0sAt+DVg
EmTLcqmXaS6sVY5+//Elt7oJpiprUIKAymNHiudqUfGMOk7TQFCqVuDFEf6RXJjq
sSEVQmwGvPHYq9FSH4gOS08JJ/JNRt2PHRbVs3PAQxrKnGc6T9dLm0mIN/ZVmWop
Yq2oaRNVfn06H/+BuOoGDrHLjRMiI9ZoUvFCDk6qetOL1Da9fG+VPmGiGjyK1jww
qWOEKzXpHNLGhKr1dAs/PW8Sc6TvYs11nzfynKgsI2+SNX832zdESgsAiUQAqOgp
6oCraQ2kjknmnSCy1K7vWQlG16+vXPWwrWG3nK/ukd35/AbVi834/UwmNujD6v5i
TJaBg3epyxiOr3Lqzn/Yqr9ECVv4MxverpCEyRsgZ7dMppE2lK5TXQPQ/WmcJLxS
GPUCcrm7MHU7WZjllSu0kFDqT1bcuxbFZhBcCmSayiM9i0FcQDkoGdrT5huHlgXZ
abLtgXdxt2pprkA8+TBtCHJrwaRNs6WUr8ZjlDWcbZIK+MKTcoyLBTRA7D+vXBOY
muDveuK8ofDbAmpXlftblizPh18c6LnbBSta17hnp398h2BBTJ86F4vh7Hkt6d3C
6/F88qf80bhPjkCM8/QX2bunihBmMNU2nWFpM6q3MCDhRIt806pkGwwAKDR5RM90
mbcPMwLTvjViFtXPTwZxnXGy2n49VeDpRAREt9fUTR+d3cXL5c14M8oqgOGvu05y
Pza7qaiuDbCNqapvKuWQ0dBdhEajOo2EDLeAx6qmbG0Vbu61yBtpoA5EMrWw8Nil
Qe81IRZnZgfQaMxKHfR5hpLU2C7CTIgTypGlmfC26Ukb/52aK8TF20SY7LlE7lIc
ouhEh2e99sgK0lfuGtvnk/3IazXpiEyYf3PL1hnaj7W2/gOyzpg43jO0WETvm/Cl
oU1IilkRuzcjGMdBhdNtiqP3uZ7o/gHHKzLKhIaY2lX+z/EcyQNW1L0J2hk6LXDU
69mI6URwofUaziMZZmfNhCUx7bMyLxarAYXvRFuQHKdt0gwglkAMV6RJZspd8mAF
JvU1BEG8g920QYL9XsRjeV6DciW2QcR+L4fWhrZ4ruN3+gZc/vF4MdxFGMbtcvqi
9klCmd4w0k0wa6f/MhwknzD1WME73lMi89UUbiRnNARfa7XWYRDG/4blQuRf/3t5
6vHG75zP2hth5rL4Jl02zhR/o7DET2xNovEOnkgnatK1kh0sST/d8TkLTGsCrz6b
sOn/TfuWrT0bTkwiA3lelFSD8sAD3XfANsB8OpoA2PONtw8iH6K2Ay7FEr89tYah
5UVyhsexkTapTppYZizFSuXK3WOzgAfbMDdU8QKt/PEkqnpvJj/PfdDmCvFb+cjR
FxmIw1Jfg5XoD0+HmXEv91CXlEZbSpEqg/DMSJbfAdPYP/t22PJ7yTueGNQpTChf
yLM2e7kfEznixm5GfSNilLO5ckVZWcNKY/22EzLL5nDs9TvscT0lsJdZG08477n/
wBpxLONUl2H0846PsyW34TEImvEnmgRnWLeMH+eJVYt+XX3GYuCxsp6wtCWLwUSh
H2e7WQrEJLHNoHWERiDsMUob4ckvOjMuqLLV2GfVUlLCORP67SAhw40kOzYJTI1R
YIH15xYyH2uDZQljG/Xa/364/H28VQxpm37VxH12pDY/nMNSB1W9S+KbUrmXbMuh
Otzr2gu2b4TyOzxM/3td+qHwzIEHT5+hS7G58NbGaWd8ymye0lWnyRP9ewKwBxp5
JCqAtv3kRqDxYSbJsK6Bc5I2PvwvWWmEDR5dU1Brvboc+tGdrGLEUFQjfTEbJ79B
MRYJX9aKbxF0E7XOz0kbwocB3Tpz0HnNl/HsOpp+eJM4kU8qkJ5BunTzXALZ1g1D
AoOq7NAsSUNg4hQWmmoHxp+xwroUSEoVDcxFFMEoHiL2FBm5CD2lh2JpqrgovbVo
0mXMAEe0WvGy9IT7E/M51/lmVMNO6A0ODg7SmEA064vWpLqPiVE19WOJoxB7mdPh
cBm1z32/h/sCktoqnD2JMg2oMNAEXCkuussPrH6kfurUOB5/F03+4zhNVwqGJBvr
VZexMY0kA1Lonr1ta5sBqDB8/t9HpdFLnchGSmvmENgUGfQxOrLfH8Wrq0LifMRT
JmDtkbur1PtKXXAtYP7QAiWRQsEuhOBuM/FNctvThbJJkRNzz+qOEOBjkkTxs2sx
7Rkrq7BKFXMSRu/mRbAVcxo0zmkM/4aM1TLfdgOa8QUpLamPwslrd+bkHxjRZ9gV
Tho08CYtk6LoGeoV1G507E3i+hukkkf9l2NCnE60qXOkl6Ln7p/Qn7BbXyG+OUWn
2J8bdDRCRDoY8OxuV9HO++FUiTZDovKsche4ly8h8MlIfWMduROFeO8vvfcEF5ex
9+8az/Ae5geEBTMsvdJ7E9mnxNE8DeFm86qR8wBHSU9OhXcu/ZYTFkta21+0vmFN
7GVtmzGBA+I0ISW5t9xKkKLi1EwngGGEEbGR5szo+gLnmrFzDIzw6eH1I37va5XB
vy9j9ucGTpK91pzSS4XA4aJCpXf3jPF3usFwkVcnQkhRN2dtKVak/Sc9NDxPfBex
ZUyUAho91jF7bNDqBS019E7NuweJlTfqgjGwR+l41QuOxdCIgY4kSVyhtCisQ1xl
66giY3OsmANEG8WngQNNF3kLuhqHT3xb44WPB9hNCxH401NEP0EqTH/Zjzk45COI
m6m6CooPYLkeNRMQ4a6CUiEN8+TQJZkqS+JGdqRKgdvQbyph0Rue8DA3Iter9BG5
3uO+G7TaJjCA7YYvTEkOExGIo/Qu4JJTbPzWN4LH4SLIeyygBstZYWihNERGoQnb
w1lcacejhORVMBGUdnuFMlJnnSQreBS6BoZsumOyUJhsJCbrXUzPp166KUQVTLUQ
rrJ84z+HrpJB/ceQgJ69ufbrKwPwRe8IX0pEITzx/dhEZ8GsY3IKksQALve/tZif
bMsGlOLslLEauhXmvOBNEGtbiRu4bTP4Ra8Na57RrnURnnt9Fb/fh2MfOfaO7/DA
WLOuHmlEoXB8CUWhoau9uXSKZ9glbq7/cYB3g3MCBI3qDvi6nVdN48O96wm8iNU9
LpwHsbbGIlNPsn3RVxOQEtmBymsPXsq9Wz2jRT/E2kJQ+0Pdmb+8/zkUWn4ZRhf8
gFFjrlKCdMP8NbmeoxMnMfJLOJN2pLwF34QkfkJydbbxklEx4LFEP45f7vd9g7VO
OEF6HR0GfRz2Vw5tT2JUoE/rTfCyJnRD/nq1DrGmVAqkymYuuGVi7W1N7kn1VYh2
kKMGD6s4Ycu2lE4aVBPpvd/Oe798U799Q5JcYd2zY1z1s+rB0ZsbJF9mAUJz4gPf
+A14on1fm5Uxox+DKOlZeO+fSxE1ea4kKGhYqP+fwqY+uabuEmKGKbuQ086BBI0a
L9sPRbipsIevGh+R0I7CB22W0VQ+SCSJ95gaM3AcRFM3YELDh6aoMR/M7rQerS/7
UtciZdGFZ0W0R/8pEwN/RaS7XlU17+ZRfXKS/wOS5lV1RAz5Bkaz9A8q0sWcl7aK
1jYOgq52U5yQmMpWO1uzli4mEJFy01stXgbfTR0ESCn2k6OxphvU4uvAFT73lqJ2
V9Rv77DCWzXawEzJbz4yrxVme845nefq92cYMFcxFfz+7HAe3EswGRfdMa2FpaXl
xYQ9eX9XuS+3JI9rSDU2ReTrOCiRMiXMkjqRwzg7jfNj6kMzWepraBbSThmbLMy1
SKNZxvoMluUSzLkdD5n4ySFcAFYsql45AeuQYF9bx6bLoYHlM2cwqqx3W4JKz928
1+cJQ6NYYe0WoFLdUQ5K9+K29vc8iU9KZoCak9coVN568hl1aD57tFNJqhv4PI/p
Sep47Aqnfr3hyFWeUtf82BuHeOy6pfstKvFgNB+oPGimm2DmKlaoicgFirXwrKO+
C+h56CgX3W8tnh0dSTngH+xewXfl6DHTbofhfI2gdqTjMpdNu5T5kcY1xCufwfd2
bMb8UOxZyCWwnV5W1DvgxCoHqrBAr5dFgE+cHgXw8A2UPg2b5o7VMdQsZfiz2/Sy
qJcfVelwnB7Idu5dksEWCyyqF2LGsjEbnG8PSGYHTPUsiWh3qNK9YgBGN8jTgUOD
5GPFdrOIEvG4jWpnRo01RYknMuxvKZBH0JQx0vRmZDAwKpiOggGwxOd0i/Na1rP2
PJU5UmbT9td20A6L2ctHuH8YYTGDQq8JpxuQyB41ljB7zpjwtmiTRZ5jH4RPgoUF
kgUFDvd3JYNHz1y0nKuY6BVpMV7QNB15XwH4/vjlXBXONLFdjqyEu3U8kP2d9rLQ
T/qVT99i2mKg6/M1Fh6gvEb4Gg1dGiuff6RaUhtHqoV9+I0wrN2ldYAhI/UoWDOv
W18144AB380R6O6rzkqiPByRFl7+W+/C7uuOVUZrr0vB/f9ErKXldtzqhotTEtYR
pd7J4DiQ2QtCDs3J0qmfCqm3Bib4WoKXkIFkEUeJ3ZJ5U6PWCdCplougTAWpoJSV
Sn4/IasqUEZITcfDaaKVN8LWXtMOD5OnVNiLDAFmI0mMs1Y7r5YTKe1dx5Wj+MQz
EdxH5TO69zisZV6dWlXKGaEIei5zYcOMY8KyGz+nrc+EPVCkpgMOs3+zLlOBoa1n
fAKaA8f+rA956/jMmN0V+KRWMYxYjqe/ywepllVL+a2DwdSlvbAWOaPLrekTZA30
WDidj4iuI1jEl2D3nsY94KCcMh3/4m72zjQiww1U4PeyCwBMRNfPIi0jYff9EirR
bdVUSUOJrQg58rlbiFSqe5yse37YmtI6wnZ27jx660SKF8uHAGehosKd7QBFsRVl
u4+E8oeIDy9xAK5SzDu4fe+/52DQpAMnqGaMkSG7ERER645Q7Qducz4kC0Ge0zcz
igTMk/PtMDtVwKIxQmFsmMNfToVeq5T7IN1h4v7tHqZ2h3W51t+FAZRyy4EIUofX
OFtAMT7lSDu3fPgo/EnfACyapSc5E/HwJcrwlSgf9lxGMmZu5QKP5AcyG0uZ47qm
4MM6L/lzQckg5DudZ/U1GvVBtLZYJy0miMox/3EXKTFFF+ehDEU0clHJXDJGabGL
iSu1YNEn214qWBzh5N64/kL4XZ86tb52dT/69w1HBfDzisqu3+0qAQcVymC2ab//
Bzr6P1l13A+DGupJ8TTMLYGCDndm+lAm+DkDIbZS9J3BEHeScKczvcDZX9zMWXbD
zzBAr7gJ06Q8lAJS4g5vBkoE9ySwrM5q8lPAZkMad7X4ct0R4bYJKO4/TNLahHia
mOkzln8NaU/ODHvjv2gqBZlQlJ3xgTmPrKSA1MmmtL8llbT4M5uL4dfhCZzMqNGe
7W8dwIGF27TPRKm4kK5kWqBqlOLoukth69vqYCa+yqxufc60uPwlBXQxcaa+E733
PSLHERIUNruAbBUk/C9EfEgExS2QJ9DBpqspdSiNQE6zbAXhOxrmYOG3jnqvzbtr
ISg//TgCnBa/Atg6v3tLocy6irpQARzhtPDbi7DpeurBFF4CGkGaK1+BfyIh9RFt
gddeSrO2BV+TfY+0QhqhHVRUpYma0dHw1ykWZ22kbNH8ch61GdvOsEkI9WNbwvyn
KZJ/mGrpXgPzM25ae8F0KdaHogPSoWks4QY8Q2GW/VcmqVUKuJu6iYs6f+C+dsTB
Ez+qz+ccm42cVx307xXCKNbujrXPlpv09tmA2jh4nOZbRODHq1zNq7CS0iMClVxJ
Nli/Z/YXDTIm/TBRKbXp/X8uBSwk2rmmuNmmrfKhN27W8xJ5cFQQEVBirDXahl0O
fZNaTNkiZt2Jatx0jqtZsMh84Td7q10/3Wi0fhkvg5F4xMPYu2bQ40s+nox5tggO
7zeLRZMWoa47BnTGMsgzcXPDcxb9o7KoWZt1Wcr7uJZMLiWHGHyt3/kMupT3UXDq
8ZL6PfHnwiKMPSImVHDlteWn89zQiCUhOG2GK7g4BPjqXOw7MTB8YXNIq7LGSb6o
qcR8TWD6et3ncXNZdyvKX7lL3msi1AGIz2ZtPvizmij1Hyvu07L2WewjYDjn7IOA
mNZoMF40oCKivE4x6wvMQ9FocgABcBnlYkgaaZqafsMVPgFlKICjeaffXDRUSnyB
TmYzz0SvixKUoRxAIUPhVrqxxcnFFwVF/83c8m/U5uHKjuA3IZulPaPsWI5zfGX+
sOjBKNzoezVEk15xWNVryKxzIdQQtCg2b9zoHYBCNHFo/WcOxKl+6XwH4Os5K79N
5eRRZ4XEJeYLMK9b6ywmJO7LfBSW8mdGSkKEOCnh57191Ld3t4f++wOrd3iOXDfb
vMfzsr7q9thwbogIINCuLVzXJXTrgTpDHlx04RYqqy83Pxlhag4TDjVF8jnoFO+E
JqPYo5B3/Z8+CdvhxZgfjKKtCXEVUldkbVQfneslj064YjHTgA0uvAM2LbfwvN9v
LJtXbr+uxCBBHwy9107kpGs3yW+syuAjb2xsRYPifnKF+6iVuyThN6YedK8g2DD7
JRY0ZelmVEvBf4O+RjZBW5ZzQ1cAMujHc3xOk9iibqilgKe1oRYnYWgM9CMlqrJV
4kTTH7MeZXiFLAoYRUvGrAGUyDJcQtmXzyXLXIo5KkEcdwzkezeARJIIVOe9s07J
EwUofflvxRQa4Xy3IvxRCvu6rMvT+596WXHsY3yOlyJu7u6RFmlu33ApNMNA7dWA
d8JTFOt2h/6KcmjEV0CzGMaUmtjodpM2sfBo+GBtijxoxb2v9LxrDUsdi5ysp7/r
aBDhVSWOCRG8BMr3GV6tKjoKMV7DuQ53DOELAQ8OS8jTfeITtTWUBrdSInHcA/0F
kdxqNPYTqjJSdyEkVnHQBhcY/QTqiX65NZBqhcIorFAxGAgWibrvgXBnQ13T5yIo
5G7gZz0vdtBCBxJsZkM/HLXoBQ7mhPC8RJ4mlqmguGoHI1nxaEBIfYg6Rfkhhx59
ydHf00m/ihfAQHuR5KwtdYGvRKEw9LhQ0y5wrI8L0bLq6KXMiJlKQrp29aunH5AY
6UgTxWAABzFshZZf/6/WoWgepCPNbqAM11TWXRJS+JCCjiVcx5RexvG0HfyG3NJc
LRav3BfxAW/VHfN3qFC8U5Thq/alKWlIN6QpQ3UssDwviri88kLc/KnEUWXuwONI
2dvpcjSVJynLQSTvv/UYg6/cgwCZ7cnoesmc/ViisB9c2FhAgY/qv5RH1bbM8svY
WE8rFeqQ2NzusL3jHo7u8tBNUZW+o/XOFv94i4D4h9FIOXc8qL8MEq9wwTucs2As
apzO8XwBNym5jDzQjAffH36dDTH921ixLr4Ny950UKK6RF1c83PNYg7n+CosCwOQ
fMpaTIehvfx1U+E+1WcBu42DUn3/g0r4lubyxHK5lJsE+mF/p6qIYztAechiuA6w
fEOO3XPdCvw/Azfb/JL8UuS2YE7dV01+jkqH0V3aXngsiuXgQgchpRPIFJZhXrVN
7H+OOs2GHe8WHNLnlRiEy3H7/d6KWoTPNJbmnlIug/hTVLs8iKUNF9dbEjSC0IR4
smuvMN5Q8D6FZBhpUV3PdJCELNnCmnC5rY6CaYtv0SU/YJKKBvOBt9WwiBuHlbf7
SEKrfkaD4XKeM/wVzq1r9bGkWvf+jyfJtwsbWAn6ZcOPEDLzVe8tpWJiChIxzEJJ
BSr5ecchOoe7qS8motKSCyjS+iUfnF9AK9/MkXB/X8ZAINdbWQVUNIELEwMSU2er
35YqsOmbRH/eYbSUTuGIa2GL2kxn4rzPgcQOSoBGeDsEB7EMLz9q4xXyihIYfG2N
RptobCGKPu8fjQAiJxkFrbsWyOCo8ymhsQwclTMTU6kHRhFm3GBu5ZafoOykKrya
C2ub9NkSGO7f2cFOil0k8IQGiazNMEUEFGJ+gsfPOx0oyJbpP3+55I6gMgEyHNse
PZ5cagw2FoDZF5+THpFk3Y/jxavVLi+UQwYs36AC75zmK+UCJNqKBs3W61oCRRfH
36MWbSnFUA6ZPCeTRmdc0zDfc3x4HETpgzZ3OQWfCB6vx6yRWNXISnwFCWoR+Wch
PNdYlkzUmPiaWxUU9VrmpZpkFiy0xU/1pn036lHsp6c66KvOa5VVIvv90KwkdKzC
DJKwm74EsCtZhqT5lmR7GMC9ROdCZII7iDXk+hRNjysXCfY4pX1H2kFVM8BeCb/C
MBzmUP/2yr4HJbVPH2GELEZjGzqql3ZhMtC9gRYbqpjnm5CvbPzv7gyDQ1vgGRi0
b+TeCLQ6iD3/yKYvi/+Vbgb0Y8f34apeJMCtnbohb6QFtkEkiAoGzGY1Op/9sXSW
+7iqfqxYl+iGuggxhlX3viebqd5AX3BhLhikpuxF2WfiZWBstgxmFQBT/lORiuD6
1XU9tRfLvzl9P3jXPgzt62DiCBdAiuB37tR4H9F2gCVvsJwiUlGxFbrxMQ0nTb9/
BVeuNQ9NvSuKz5KRXUNFQs4yvTqX6ppaOx6R0jii/+6GI1o0ZvFt6bh0p2eqMpZl
vCyV9NqqxyYN6yd8R7k6O6EqBzskesBChIsB+og7cZMfiVvbJdttR088bUL4ECsO
FqLEL2eZh54DIqBfIKO8f2Tet79IMZv9yJF6ZmffaB8G3QG418iNSTcVEvqYZMAj
SNxS/B0fSDTkPYGKapsHvPCKqTMFRDzCrMtsN9RgtLwMTcuLtEDacyAhPDd2dx4H
yOx80OlcOK3UaNsOXLFNxD1u+a2o6v7NqlEsY7LxksGA5ERhmK5poVduPXy/9i8N
v7ESODA5JGjmFAlerLi4J8p3k1aLMbMAme4U8hqoms/p1y+A3ALAmmq0pDPPq9fm
d7Q6HiekTGtwVZH1YFCgdVCnP9i52anezLX2JM4LrjFyJitNG7JJmWDLhZlicb7e
H3J3rTbrX4oeIGtSu/Xy+mKaGhmFPMXyZj4Me5DMtvFApZEWc0RuOjpstoErpGGf
UjofMo8VhNKiEOo5j2fNUebyBoAL0rM5SG3sz+tf/CjUua2sr/SdTkdeilwvNDdS
enbwB2Rfyjmj3tzq8u2gkqVDpHMZNTCo53WjEtmz0JSx5BOZyvwLHEDVqhijBfFw
c+An4EX4LqRRPpp08z0HwenxD70wxR3QZV2yy9qVrxbh5oH88IeVwGJUhA9izHN5
Qv93fSNhzscYEwTb/u9qXMBCm4FpT+PGxAxnpkHB9CfxLTFs975TMC8yx48ssRR8
Tc1ZxL3ghevfUEQXRn0todPHyAtSu1O/qS9Wgd6cWW9WM6GhppQNs10hTlhEpqc1
/hINnQhTP/OvoTkUXh7kZRYhtTyZ81u6lknyj54B8ZciK2/P88uemMGB6N4mjfrP
h6PSISWevtpLWvsue/kHS0UYcu5UW3zhTJdYHNsdwN5aaZWbMt5Kh40/IrNav5xb
drGnTruT0backze3ZESfpAYY4g01k+KJ0bDMg9c8WdEk8RcoP1rwKpq2h9lGaySx
AsUPeLcxGg22tRWKkzlmvtG5TyUj4bul+G8ZkwEQZWcpMaxvQHpjFMOchtGdrIsz
BGUXgLtK7SXzymeugLMQlapMeKVB5KOnGCW0Uv2ttSjooKROsDk68g3z12V4cauw
dSAD6ZUEWRhoIKNF8sZbaBOL0If6F62JWKa9ewQDsateVwMBldW7VxrSVI8ps/lW
BkvOuJemyQPOvGNADWNiQ6rHsoESQJgI74jRItdP8YTKhJfVxrioK7LvzwkR5WSB
KC11INzXjOzhVc5YvHLDP0MF6J3CnePmfp92aC4ZihBZbgBIIlpv7VpmQtdpXYUl
yN8btHGbz7Pjxy0HUoF5/6eeeaV1mMaLj3E5azgefke8uut0dvcljWetbWG6zIWj
ivf6FUx0GqlGilvkJS93Fd7C65tboxT+yAXdrDViIhLlt8tOFhcvJAIpodVFoIZu
R6tFD8vCqsSI/t2TE+AwuOtFqMyt5pVClO7Yoi9Q9/DOxuPFUuwYEVyoqpNaTdrH
YafN8RfcXrAkGWZhN27/1bNW+0TziBcezgJodWWVV6B3XN7bW5yN+x0ieyPD/rkS
GxuJA9dT0SGa8e9P+dKVYWP566cL/VE5t2ncRsJrXjgqMYzzJ66EehXjP9hiSoD2
vWKMTk8ZlV5nCTtJIQm37bcRdbi1dUS+AJPLEYk9V28DJHhBCZYByV2cNo2+zBLv
k2Pvi7O1ZYLLNa6Th9RTtRvCVJD+kEjUqt3zShKWOQ0L735i4FICjpDBKdgP+kAH
6ueQtbO+0yTzAVy7C83FUsXs1wM/kgg8sAh7tcl9Iilaq+NOCyfdj+edXAN8emiY
YN/DA7GR32Uxk5mVm61g0FpZyD3gNktUttrarOpgRr3MIU8gOPo2oTGTjIoIZevq
VU7n8tgVnM0v+4GfeJzkZi74pjPoOq0dSA+BSu7MpwlkgE6apcx2ni14CiuZHpZd
OVMYro2EWz3HJ8X6KlQGy7a+jbMAIQHrE1lwScoSGDrHErQbvXKAqqfTKtiSn5DH
/vVJanETp7w+bI5/aYUsRioDK5I1dkqhyqIjhnO7Nfb1bkOk5rMaHq/fZyGd1/Ql
kS4IfJiGMERps2FFGkiS4wgjzSnMhsPNUZo0NHmXmLq3ch9Rw58tuHxgHmQOUoq9
qqxM8HNUfe+7kvb//OWOh3hmDei5KNu9EeQ7K0geYRzSkpPbNgSgSLsdyYQhQrZB
ivTxS7eGQiOur5mCXFVGM98WaMBJRoggMoUBihTkE7qxIfidgrrfIJXWeGJrU33z
DFSpA8f/n7CecTw1Z7LjCqI4xyxrBfkZEgc2KSb1tnUfWFkd3FwGu3SM2eUiFs1z
F83EDpMe4V5RRYx5/PH1bYUmqlFMS2RUBVhx+VZCCfjf2IKV/Cb4O/Dw0nP0ZJMk
H1mdiuNcdyLzIWW7qdEjZ3Wh13tontGJVSuB3Y0PAqearAj+KHenMNTlPefGbRDv
AGvgyu7JTjnJB5IEM5ZbtMipWDvIW3/h+/b+jChY8ZMP8fkmVhbYa2mI0W+VlCOv
CpKmbQ+c9XEcr8iDszcVWB+X2b4J0oKLwv+PYFl/g6Jl4NcmJVwRE856pVB5HylV
JQo7AxQX9vYt+4MfjHq6PcP6ChUYxsZQKOCZ2O5L4UT8FUdfarXfe7lwv6jSTTiC
xN4vglNhYl8TfGWyVXJQy4bNDRI0XyYphKM4OLa2bwPGifqflJpXrYNAY6q9cAH+
RpJoIAcQxgZvw/QwI0Rqfu3mEen6LdGb1R0ITC1Fv4bn/JV3ujQM4wT08OCt1qLE
DVU0kuzRo+KD4RRHzWF2zcoZfI+jNyVPdjUvo0HWe8yFsbWMn2zZ/fS4VV06AMDu
VtdmvYAxYOrpBlX3s0sVs4q5YcWgHTl5j9aYoT/3QrF/4TDLKF4zgtFrlDKFx7fI
sgYMr1owXZ+uzuf+OerUY4t9nogEy8yk5VbiAYOr14AEeSZZgvQOj3Iv/VGCf4+o
s7GNMO4iHVuj6Az3aEnCYcuEgzNLGBwVAF/dEYcRXjzpkZv4ZqUm+o5ibQmwtfhs
wBBal15X4k8Woi1P7/EXYshbZ/PGwbhfdzMyDD+ndR2XV33pEpei0bqA+QCu3D4b
G4e39JWe7RWo70HrbVvqljltAcu3qeHZrWujexlkUPLgjIIP/pY/A/+KGViWD+En
0owttDTq3PZlP2QX6342vmsHlgXnHGKz/4ly+P4F+dFu3ISX7wsRtUNC9Ub42Wut
7H5lqnrTpuc9RgNE5L0rahPkkn2oR7BqZJXjARemnWym+D60nyevYgFUwUkeoqEk
xMweChPS8Pbmu2Cn3E30PD7qNqs9yPi8FqqtMLooNQI5scegDfv93pM41su04h7J
2YzjyZBoDPJbSsmit20yCb2DOeWvOxtVMNgwd0VksZlNqfoTcdLsJPKygvAgmap7
jR7Cm8k6ZnQuSEBlkCAlX9lppXPLkRaP/vYHdePU4FCPK0MX7scdQzcWLfh2tRPd
q1dadG9e0eLzg7hyYZ9T4iSgkocGYiAM/P+cCEzZ6CplfCzte527qpBQU/Y0NttD
5yVadrKlQiU5uuWOh/9RcVr8n6ZskQ3PRvvcqe48ykOH/aG3CKeSlpKYItwhWgLj
rOIqGspYo7R7rpQCgK77dGGph5/BZYb0hgXqjQSRis3f8Ubi+TLuvR6aqO6saJjQ
77sQDWmcxryS4Ngm5lywMvmRa3BtverdVSFJMhAXlftXycyU8WWexBLoy83gzlPT
19CF0lh8RnyDnusB16a/IJjglIB9FavVh4bsFgRfWfwis3IZXoKH/890vUBAaJOA
zgSO3SotntedvBkxG3bYCxXBt546fIbjmJBJ3Sr/7aOv+Eu5dozbDCMdnE/MHP4u
92xpYUPGUi0ba6Hix7Xb+lI+Tcmj2aOSBKbq6qfErXyKQl8wuNd9yXr1GAKtAE6a
ftEA1cIThzoySzXyHu+7NOqxZwMFFcbznSbWv2Aqz7fuX5XrvpAIuTGhkQHmJOWJ
GTZGMs3EAfnQSCTh2HcmJ4ZTj2AM/wmJGMK2XE4r/rxPP9sv6rx7ZJR/h/ngg+S8
SkjDubTA4PkSBUZAv7ZQBuTg0BYSdkfBql6MR/42GITtgSvDonhUsWxuY4/KEsJG
Esdv4nM8nIjkyMfOjf4ZiIsa5Zy7TY3s4lddCwX7vErmouiFf1/1QiYCAmAMYyJG
PBZAQRA9PpFqGPSjrRS5f3ZfmMEozqcA3odMhzUGq7OG27hLZAWIEXJE+fY+tjrM
KS0BHo4ztfU8Vgtm1stohSgqFWHpDruX38UWz5DKxFXyW6hYtDoDdIqp37OgMiXq
eS4U3H0uFSUNyKEdHWu/C7NWEek65ETNUBq1q1iAlKPJYKpgm2FQsX8f5DhYjPh1
rEapUZuOIfQsVt9wk3/gCD61/PqxGa5kw/vHmpRUPDf7qiixp1+XVDcBkzHdhWP0
KEq95ohlqtf6xr8WR8xdK42taGXx2Q66QwmYMEAShLfTilusNaAN8LGI+VTNq3oj
kt7v16tdaxTez1cCJWBt8gmF1Bt0F/7/GKyqaLNgBFbOvkdAQlYS047pa7ahrPzS
BZlSlA68ZK8IcBrlDKhcmSLjhPBjDrDmoZ4YlmdAvKr7VDcnF2cM6tEnhv1dtIDr
J4vBvWW/bqphX6XgsgKW2wo4GWAkCXRCa2CyJRbxL0qxBZwmBgw2D3LCnLltVkBH
1d127MJXy5EDXgMdLI0y3t0ka0G+4IMvIOvHei7mtgAyoE2iLfvqnKVD+8u0bhtA
xWA9SDLKf3FmkzWbxzp/MQ8rLxZl3EMRX5baAPY9qcxoKF8VjFldKieCGYqoRwrA
c6F1g4LsAhgKPfaDKgBZZPrt2UXlH8LmAET1TMjuGGaZDvuwJZLqwx8Py+4mDVzV
9SPGlDpUCO6oJyGxd6JF52ynMlI1OKdCsnTJnrrAFG2Ko9tVm/XhWOA73G+SfoBe
TeBGLGQAY1/yBRNQ2HKfkH/RKN31+PrA2Od9GDlOgWAWGHSP5tTFpNGI6+gvvPNj
OzccQd7VnBRP5kbVbkLUxHR5Cy+JXcUvcRkU1dntl75lBc2eX/GQmADddcYTG7TF
qvujqu/Vdd+MVDvGIQPMaAWrg5zaAimk+ls0knAZtlSiNgI0jWYNGh/tIwWKniwp
92rwRJ8juUf5UY+m4zNpIdlccG7s2tdqX+MlNqtibEuQQ7sC5NNKQwQ/RJLRUoUO
UECHs8NBU1VXGKEz6Qt40+/97oJ4LPBbzbfMXNKNdNbo+DXWbDt6vPe4anQ+lhxU
+bstfYLo38LA5sSe6okvyYcMgDpFvVyzsZOdtUhwS8rGwdbMrrv7U8Gs+oiIcg5S
+vfwVQ3bs1mYBAwx4YayTUqPSKhguyxHC6MKmtClJ4LNhnhq231nsd8CVIKFXH5k
7X/GeDH2/Gni6C3JhhnjQEzvjgcstkxAteEv+FR8gi0w1cRyzZjDiWasW06B04eJ
Gn8lqZdJMP19PDoktgaHMtQk6GwO8BdepJErQkJXNgEg3LrkIOTomF95//KehcA6
EZS+FHRj+olJ3L2cPY+jHIakvclthDCXWCRxPNy7f3HKVPWcbQv4LrwlnvkA4yuv
GTgHPpih0K51Kl3Yvt6jZv2FYl5MrOAlS6FBJWUNuFLqW0uvh5GRCZaPfrlZtGVO
RIYg5G8ZuCk4gdWgpaYDZlgW0kRuA2zlU4ygsQy9kl0gsRW5ygf5qAnmSocYBdne
5mGDzFiNjIoZwcC3acwPrzzs0vJluZS3MAZgnR2CZtFQtNSrpOqSDioHBOXhYG9b
22B4jo0C5GSdn3uiSj28Uxs+9zOLXQrI37S0KUTABAXCkoZTETMT2sd+alMCQCL2
YBnOBZwHb3jupP07zxfQjyV/toYfhc9+0eo++cVt+OCOUAyvUnMF8FxC5R6V8+1h
etoJl55ae1Z9APTd0sgib5FfqhC7y9Om1CvETx5KIG/UuwAfAvZK7zWqqGQYVeQW
d5Fxf+kcaNVUB/Uz3L1+wzMt+actC6MYGCIQKQnFW4Bjvx4UhvAGcTxApdw5JLAL
+eS0+8qTVpIk4DFsypJlshnKfMr/mG2nM/D5XGhFBKhYmmgkgCNb3XZeuMqCLvwW
/woQ/VhGOvpFIJD0fWIAib5vZFXNIqsLnKl6un6xyQ6Ctw3sovqT+E0x0e+P3/4c
dv77VYntrwi01ueRHS4jOMW1+bVAX8KeKwHIuoysLr08bDOgFUPk/bby3RS9m2MD
i8PFePdpuhewTu15Mhj+zEfVImkKMNvu87XdXZNkvG24iZXwQnoAIf0JBT5w0QC3
/JRSaj7ZxW3P4PbflpVkeiMxWsLhYLvXYdVzCvSlCj3x5bShMHG1NvjqPmdpBU6/
nuuFr6IxgvLoNpzcsMto2w81M+Hpv/tuhzr+E6BhY3lD3oUwyr+9c895LdLcaLo7
HVkgin6bPUg1D2ScV80rQg7H4OlcWOOCRAqF+UctOGSxilqpj0BuBNflrrmSVIHo
6M6v7+0HlSmwz33co/4+Jk8k+9D12lkGcGs9xuTTEwoDbSiKBodTRgUNVPEnGGea
5Lo8MBUZRdImGrrlKAYU6tYX7ot1uc4BBf4z3t5FENsTe1RigkIALXPwncNLy6Wq
ZHAU9+qQAw6pGJ57b1EqH5y5HxIqyhtBFS2ArIt3wkdkhCIh3+tQsQVYP+bSUlnN
ggIPFghopw/PZRii87HVKTEoea8QSAjidEMqPCCB4Ytd2yFeIuhmB0brUbpSHfpc
ifVk9JsgFpIM+sK2HbRB21mFoClleCuKxpmt5iLsUGt1pKabEbYpmRDwkdY1ikR0
57dFMFXPUrVleQWln351+Ezb3NRUbWPIQ4ZyB84pk11HiCOIpNAbJnHwPGWxXCnT
qryjSyCmsZ5ieUhR+farvlqbdLkgReIIUq8U2GH+b2Fj8I+YpLXyIoi4mRnR69vo
jfrlR4zrx5+e8QYH6aKK9KTJARgxD62JRqJboBXpxWRqPGtHivR2x1vnUBPG2y7y
AA7Ss9mMGveYGeo2NgNl0/XLblLQAWapcWJE7VSU9kMvUDz9R2MQTpRdPvPW9VnL
Hs9bIe3a7GimfFSuhe0UpcT+XvTZGulssrfL/a7usqnu17DxCGgw143jcRYq3qjc
QwXfAIHnAupQHtjXFkkbAM+LqIPSEjjpvYfRNUOomPcrrwn/WmWYy5wzoVcDf6Th
tNiIOLzKDPodRCdCO06iEZJGaL0/39U078MVFVxKssPYrUmkxxnEwCzLlE276nh6
d2p5UMMz2JjeP+VP165tS9RBDa46r82P3p4NuOzg/lVbUEI/ljf9AGtyvbPExIpA
+SpsVJWqKhOTF2jKbwu2kScXce3qtHjKl+MIAPgb6wO46lTpA417JD1gfmIZECCx
X2igjTbBwy55oHtPIfNSB46XQjbJVLMwCjLvXVGHxsC9LgFpf0fVfc0D4yamo1aR
R6wMIonTgmQ2Wy2yFnBmOMSTrQkayCHrVyZzINyboK7FlX9bQaBjHpAcZr4E+DrF
BNPL3EVhh4StnVoCa3Bn+zNzjGA/QY6BbNp+NXurW8YCPW6h65cboM/IFeZpccxK
QVhBOhF+BQffohwn4/YeNrZ3vmUN2U1bF+JjUH0fip0AqnZlZVGb4rLye9zpq8q2
zkEe9VSeW0kz7OFeTiB3z/Fl4iqugbeFiPmRbzJEuoiHObpwIuXKbxhoSjigp8Mj
YJCXtstftK/O7DTS51WLEiQKwhd0PET6VrReYiO8CUy0fQPFwesyq6vVBLz048Ey
uUMEyEgzUO0jGYYZxCryraF8omO1wJWTcKt7LcEr5cnTp5xWyLOtACTGk/IPELmf
exnCBGU/ogHX7QRMc6yQHDNxpi3uWuD3xwYV9oVQ49MmtXVi+kHPVkDJIZXdYRdc
eonATSr6fqhiOFfnoqwBqBxV6j+uma1Vgbr4bcpATSz4n0a0d4QZDAbV0Vhdipl3
vVnuh1J1GBYVFk/N+3weLS50mRSw9iCdOoJ3qt+DULC4iphGq31EL3CeFzXuTkeK
lIKBMG0LRHl4k1fpFLMwYyiVsnIJz8B3+1cu/5dxjhziNVwwvkx4XuUPhVHbEiR/
qLUbMHs50dP3g0EynJ0TxrhHZjyaP47Cr2cl1BGERLggmQjgQNZc8/5tZ02p5fPK
G1xBaDrXDMdnztsdszR54M8pSca7f9Pzo2cGjkj9eGatVST6ce64NKvtB2Z9VZ5Z
N2dR2d7CMJmF2/NHD66kiNKPnB42Wq6gnSGfJbIZfInaEB8XMblM8KS95nK/719q
rFiJsyBjG2g4jyaFjv9ECDL3bpYNCWaLzDVyOLILrDE1amHhdah4x162I7/+Ib5B
8eu0+DV/CfG83C8mabRoGawxFua4GAZAsUZ0rsmqJU0FgV/bUJNov1GO7Nxg27LL
GTEY8Vcj8TDNn/OF5u9JBEbrjeMXcKxG3ZvksvGVCyE2gKWQJgw5XPkXD8tQnHDN
xnyIMGj3VRokE3dVfq1WB3rRBBbYO/d3FlQS9scGkDZHAT3M7on2GI19RUSvVGGs
0Fv4Yg/h0dPt5DrssIaNOMGy7QvJUiZbhGfoVSr2MjKwnESDXKEQKghWb+6zzxtS
OjozqH8wcCVTRnAyvsTygjEy5qAut+81AOhmaOuTo8wffZFtsf+8VlL7g5J/PW0G
9CqjJcoRVHxjlaEqBnqqEVzvaigoldPMO4OkfBpmH2K1owdTQ7BztB2ZMbAenDr6
DnMgHpViHs36Q26P9VFho/w3268gieAqZge2rQADfev4YrlsOX6rC9UaOiBHfAEY
vJa5rn9HgFbHrhRbVxeb96sSnNZKEdZ2uTJ51CLIUsuhcDgEemNF/IbqYAyltyma
Fjad77N8nxNCSGFYYY7KOtx780skHejZJIlTTawDk0Q5LdM28fz4/fxFsd7kP9y7
z6XRydhmgfcRp9IQp/+XXWYduztcURdNJDSZmZT48YldkuGn+aHtFsihcWKEOJFs
HkaOIMk3GvmAB1gzANm00La8fHSj7eNKddZ1pczluHi1TUvll3+XrOeFKUGwHVDj
Aa4aItb9K2WWLMcZfgoxfQeOeQkXperC/xpEKOTWIpu1qpz3FSaYdZNbBfW7bAaK
QJ5pvecp3NvHyoH3AY0C2HKHrXnS9AT/l5FK9jHZ9JGj23hSAAhPZaKo8WvJtbaw
wBVzes8eJi1iIAW8DzLDZzn2/zrHC8gJC0nFW/ZwERuLTo0RFSw71Xp9Jhegswtb
aBfilgh4UbMyBhZ03ZsBcoXA3NtTckfDzQ0sIy3d6sD3TDCV3HQ1DKFs8Vv65S3O
yS3leHMYMmMtK0HOq4he4BK04E+Eo7k61hpHhc0+2yHTX6gE1yL8F7lVAoZoBlCe
TmCHfUBiWoITCfM5kaSqXPcL3OO9QhKGz1+TVkXoKCZ6yrkyqFDdAtU3hYwKVh+K
AmeWCI/HjunDWqw+pioGDiCQvgwXQopa+EF/maRgflS/Ox53SFdD0V57DXdXUUbe
pR6xAR6Ovqd+6mGxLcdUiUBAFggmmCiy0cxHTGUyAmz5BU8mwZ+4LeEgII0WgqbL
qyCFZHpoolxMkBx1lYRSBsVT7DnIoP5aCpGKlqQ+qNUSnd3BT5/D+5ulr+OByXNB
GSgU7Zmn2fNldYtzDLXPYlIuyIgQd86sGhBL9r2KlCpHKp/hNGOHQ1DN9WP9r+oq
fOolDSKX97d//ouvJ0Yt+Ua12QylX82Undz1xVOtO7hmPlguqMAgOTQSf2cP9jlf
b/qioJYGSZdJMIsnFPgSdS/KSPQQCUjtXHw5FwakKwXutk+krEgXoHQ3qi9nPrNT
BO1Sr0FdmHRfOf0OdGOO1WLOlx57tontzezsR51dGglaryAXXLDzBKhwu9eJMNwS
WylwLd5Vqj7jrg25pixCSQOjKGjJxrsKh4T19cr8wfj0alqY/WyuFvvlhzCcNs7f
w2vmJm1iNvXmy/opmz50nZdv6PXAcQOHWO59P17WOQL5bvG79JulA3u8o+K/juom
pstgCSpKMmzOasDETkonn707Ys/6XWT/4uzv6Be7oyQhEJ5z4yo6nnTB5PYunrsC
X/1tMFkmwvntnAtv90IrdNintAUW/hp9lpRQUriusxU9wgiScLrmdww9x1rj77J5
4J44nXIu35oBOajxYFstR9ACxs3gcclxbasF/Vi1eWbKmW9ykC7JZiRBnJCskWFV
CFPlcsOqijtsPQc4aBqc/adjCEUM7YccDFuvV4zeMR6b5ZztDI1NYam6ah/Z+6Sz
2Vm1lxezRKAlCmxfkUwUaw/1w+z5cC4NJuONXR90Li9Po1AmX+XXTOYdy0e/62D7
qTYKF3ba+jyotydTwV95R4frFbXb6a2cZFSMXQUnA9ks4a2F3cWe4Ao2s0rQArKe
5MfR0dCKT1j/aoewQfmmECbgjsVvaoDgzyaaaMl8+ixu057cCJn/+PVsQlHHxxY7
jpDSMqavBAXvXcuo8l4QJ3UngPWuWxj/72hBYQvAQPjxxiPtPZeiXvAlWpAiHaPS
3Tf+g1sJdYWUSrSrCwgj3xQmq56l5Hi41bMcxhtdfWUYU2l36CNMCJU/UVQQeKdL
MW7oDA8dp8GnHnjbrfoL3wJTcyZGONDHoeiNlewcA8VGZP1mLQMUxMJIxSU0ALC4
Pguig9Ox3FpdNyAev+9X5Elhoxlvmd35AVuZOamwikllDgNqMyBvfNZnTFClUGXH
rg1FkC6SOApmVkJdDTPdnicYyRXeasIYDgG62LC7hfVV0ozZ8cW7czOhsO2l/9Y+
YfswyUyhY8y7VNoySjAxbI1WJ5kpy/NUrU/fjYMWwWF4gg2cYrurH3qeZznODKiM
OIHc6BCC9SHlaaVBjOXMCk003N/UKvi5BgSh5SluL1DbKZxupGgj6hAtIepCnNxk
yCbSJv11DwUS9eHUJXR8J8ROnlK4F87AjZJnLrYf5UCxeR//ilFKqrZ9eyynVEjh
tXoBhGuH2Zud5ISfPIsw1eA11k7Skk0ZaoVc19NA17aXn2z9NfRvJx1eH8/9oxQb
FmbEUFHkAVWGLcNBdTz9bcnP04nnu2rHQXEYzmxnKryWnOBD75EJKrI/u9/NOXqK
0zpOvyJ0YUlUYtJkgl59l0bz37D+ltE7sQcVt1zqCuNPGDIOMqJKjmhV27KchrIv
sWnbo28aMw47xcDYr3Ry0cBhSemXddbAtUTEMHVl+7bk8gHPtONH5JW6G/yloH69
woGL0LUXwMQumH9PzXOYKFvFEEzNs49XVz0TtnFNeKorYIEAVGtsEz2wHZ1QACGO
ihx/bgy+d2Butldu7OBONTkvMylerrWMNOnbY/U6jrOSLiD0s+4j7SSObR7zisq9
IaCz0SMWvVA2ORNILh1eQEPQogAR4GNCtSwTxLMUE3EsJ59RM0k4rYiUlwumi5pk
5Mfp6sPW99EkyRNL7PtvX4CBF2mTYzDaG5rpvCQ8ndEDH0cQhDV4EQR1BtsVx91P
jrxCtYs2soltIrFrIJiv9IohFUe/LIVesr2luFog+0klYa23zZc8AgdLJ6/xbs+q
tO9x5xQHdvdcmUvFhDpNHDa7LObXRnZtJOtIwK7AODW4dJAoQ7GRyqjnFkIrYK0j
FzGTavjf9cvc8WO2fpSnC2T+8uTK9+13pmk/a19z84RXxOfIcd/BtlT477MJVJNa
MWgJp8XEjHbOEmmYhOm28fwVkghdkaFbeyP0EQgJfElcQKe3klI+dWum+RD0sBxl
ZOT7U9owvyZCL3ZBllqMktj5vbKigWhpD4bqlA/WDFLufVktqhjloLHApq/jH0Tc
I7fHa7VlRXZvmpdDNfCdVrOL5EJj+/IyRZ8sHTPfVAT2ioawtFEdnSclly96+42u
D+5ZhH6KgZGwM2+J9W6PO6KwBNwILk2aWzB4st7Qw1OUX5K17Da3rpg4l/qMQV3z
L+moqo9xzDBcg9/eFb8EdzzZ2KzX5Nvz/NPDYXc+y4AKkoJD1YYOKx0mF3UxRTPW
m7lgma1mpTdcW/AJC7zLQRFEDKTzMX3MqHA/jDbCuz/cIIjflimgOLsYjplIvp5D
lKRPT4zEVm8RtdXkEkTYjxuVcRRXdAD1NNAg3/+4zm/UYeaTDRlziOIq5zkwS4SS
av3hykpmGLRuAV0pOO24CAzAcYdfwuhf/9YtA9/2TUglyu/Pi5W730EaSG0P1HGY
jyDVfN+WC/qMidBVe3IF00q39JDsD15StD1AsS0ttfQEnPgPfFgHlQWwAx047lb9
X4xczgs2lXGtv57IlIfmorxX/8/cPYHaQ+7LqUyjsoaU7c69U0ShixoixZgpeg5R
6E+XQ5DL4Cvy6Ob8UNl+RX+/ZMR40GLeFeBpD8lMadXMIZIt6J1W3fSE+mmQW4bT
snzOKb56ZGMaK0iJXckhr5kD2dT9NVfNgQiEHUAAbHMsiEVPBs2kMokJboPSpYbK
kffOUWCOjsakgl7VJRwJfljCRlj1leIt/b57/U7mz1pklxf8B6PHOZLWFDDWSgnB
AAoJLqGXK9kVsYO4q5GDZPmTdEtOK7HGfsvlbg3AE1EVG2LUQOReRGab18Fg76f0
gJKhGOpjHUId5XWf+/oPlJgC2jtLtpRWe/cIJxn9kW59WyfFORIDFqsVZY0WjcFU
0iTfz5uiMq0BWqAoT/PG1G/QO38PsD1vpcDaBdrwOaPQARO9ZGWbqoCNaEKA+Mwg
Lsc9tPU8dxvb3YIoQuQdVK9fKUv29gS3+lkpHK0Xag3PVmBndTuvS4hxPguiSWqg
dA7P3W9fy+nfoPnbPZ2gPWu7JeXZBmKkE1erhmbksvsmkeYvhF96zoe0c+QkjWx7
jZMIHDg2VeO4/nmlnjmsjQz5z5bX+GN9LfnWXxHsm1ag6I3CKML3dFzpsj+ZWm5q
hnBPlim5OdsmRqF4kFNUXwa+LmYHW5z+2Aa3N8Gg/oiye4c819H2fpVp2YQTLh3O
rL/6aKviKM+TMBBdPMGGPvkO9KL+1HnVJQgxvEl1ofPyRsQ2f1eMg3Aze5d8UP9s
7RuwtoS4DY9tvy/LzOBgIgnOamP+D+PIXt/sP87A2HrblmPvjXzuX0hN0VnEfob+
FfC6b/iVQ6dFrkFVFZk7uKLdVcKPCy8OdC3XImuhJ0pIRo830CbkuUT9aXWFktw0
ONC6PxIkKPDBp7aOf1POFzmEJrulKFXTd1eX7gxVufYpNBP6/Txh6e+wxSSG8wAa
EluqpupdkpJ5AZdCnIbDqZ+/C3t24fvxk6hARjeGHfN0Pi6NU8D8E8iLLbQFI6OC
vsYc3N3e151ph+jqqGgHrNSijh/EX3DtJ6e/3CRBEhISXbRaMq9HpnnTh/HjD/XY
OT7z7pwQeaIPlMaxULpkWT20RSG54OW2uTpU7fIdmhHUaIa4XfFXzTI/bKfT5GOF
Ne+Ts4AHYKW5fCaTeGVBUy311qKx+9RctgcaDtaD100txj8dDW4XtPvCxYxaBae1
i2+7it0qiIpEeYHPn5Q5IjPa4iEMn02AnbLS42d6JoL+N6gB3D/pppBYalgbYGxH
uiARcYIktFLHgXi2KNtR2YRWdH/WiGbVMx3wfcfsQpObqe99d9F+1UtZw1PO9geQ
kVvpfAfzltbWqrcRw77XwNXtY5PHpF7u5AzbNTQ9Y7wskd9VsaYiviKHrCxkMWzJ
1Pt46J0Mko8QnOiJYldPdwoYgmpYCaD4GgDMYOhUqhrl/55gMIYI97lvoRcgzYYG
rfFai2oArA1d2y5BlwBeAWMr5yFDobMNX1wS+7kSe8GJowaxrzy8JaHJ/2Tapt7N
BreFwaFmNo1cKV+lg1V28tEqaAuybe33OMXhTt9z7orzNodfDTevR7+XAQJdbdaL
2QQL3luWNEImrKT5yFh7Gfd0CjkqhRqhzkO+bs+cNZvPtjXXo1CuzY1lL3fepFYI
YEEnd/ORCMrfgo+ZdUHG/H5I1fnoTaezX9dw1HOtWv08/kVKL2FhvEyjA/JK+aIZ
UEiqy9Laju36YXjyRjLWeOk8n72a1bHIAHX085Gq8Y5gjdsF2/geZCKk/+qierIr
hOhlbKtT+qOIURq/erh8mTJ0mLtRry1ad2sfjlZorBKEZPDYzDscKXZ8bDTJAP3f
PF3/IiKKiPIbzgpm9zhtvrpRBNmITyaxn2ghsqm5Sze9qSQyCizkENUh+8Ba9/m8
GLKwt4dbJ4U3tmBNy3NWbwP/qlbrNs4m9mMW8otfYzOccEEnbCHZwE8YVZFtmTdz
wx17+nm2k0NUXY61gGMKfRvOw+ELFFyQ+HSQK8uGOeyh8ibcW/vbvT03h095VGH6
MXtz+chvp0QTD32zqMFpLazzx+pog7yu/mkkloqwNMSjX29SrrVCmbzyw6HT6UIV
cKe0cYFBvOdp/8knHgSy8/2kGgjRGP1ZDMam/s6TtJMi0ReFaD/FpGCGRlWlCL78
jXZ4pjqLr1DkddsW0A7avBXlvRGMwao4x0CjQcoTvGAExWLu+glrd77ZoPovyFp6
DrGILh+mN2BqirmRAZijN2OtK8mleNAx13pJxJhd5oO8Him5X2rDrLkxaG1Fvkzu
11hT5KaWy8O86Q1yWLWuHlbZ9VngfWcJvSpyKA9GE3wVn1USNni2Zm/b664jb+5j
+FzYOvcbuE6MliJdLsSVPFf09p/1EhjD0VaDNIkfv6bub1NSifcisjprRGJH3jZM
Fuv4XvHGIDzUpv9Jio5AymEedeBUESuI0tBKXH6y9W/IuTZrjD+Nezup9zvUBmiX
brbJHP4geE90hiiOuCDVJtYQA3pdorMPDM/XB+OhTfsFOzUH6FGV0pKw4HeAZv2d
uF5NtA6qTtTPsydhbT9JWcpMeQSYkh4DJyHOl9Mym8bz62MauavnHr/9T56kG/aY
tJDhEHHEva/taTcoWFXrpvcqnufzVJTHhlwwTmhBMWbNU+l6c9QSCbUFR5nXxj1o
jxODovl/1krArmZwoM0LgfqwA6VRxIvD4i/ZqVFU4HamhnAaV6G6/oGjbtTtWzrV
EQsg8Dl+hX2gQXvHRTywqrsomejY9Yk8s1vlh2cKyDRuc2xipEH/i/iI+H5d941y
Ya/3maUu1CDkxOGGqzDdeobfFIP4630zwk7rFmgC6r8fHquQuOB292557FJhpbGs
sCjTN94+2YADlTpXsYTYWWWLuxeVbjBqFx+IP8iuFmr//STqtuJiDyLs8eUTYKi4
8jpuV3jld2hM6iqckgzFhT+KweF+6E4c/ZXtqkAijSDrd9wfmHUalht4ttdMva8z
QtxP/tW9OQyib2DFinWORiXJCcAbu1eq7+t6aAOV619LCBZPtBwJprM3lpDZZ7e+
k3i5C34g3PbJxo7TgdgQgpxlWbKJVBJtFWbFfsnsBbSOnyyTzVS0V/YvTStv5cUk
76ZQITx58eRXTchi8DZCMI2jnxPkIO6HpXgexfFokwG680ugQ6LoJU2PCdsNQMpx
BzekApv2uN+99GYQYopFS09+2EzbxaYsFB85tXc0GzO1mX3VZApw+qJpseBOMk4c
gx3VWzvEKPqYGeGquZO96sWqUyrs3sOpwihBGzPwoTCmPU2rIshyyFxbfSrSyfy7
R0gTfvAdAElQmumVAaGryLC9PXlxnZDNWRSEZSVZ5+xMDxrXtSIC2kH7sfM8bDPm
CAvaiYPzm7FyMJpKlSnEbKEO9WqwLbj4Pq7D0m41FrBNjtgfODMbhVxFw3TkktQE
m0aHFzt89t9UltmiD1r8lgP60KYCj+Ya81VAXwbbZDsQSErWQtrKT+6yO+cv+FeF
CPEg0EtsiI+9EKowAkQLqNqGqt9+BdLhjANy4dsxHGPjwCJpoeBhMIwXqfz8jW8o
OavPsO3f4T9b88EUroAZGbru/A4KnI92e7VaSjX59cdTKhAb9RDTdYZ7ymhwoCiV
0vk5bLU6Esy4UrV7Nd+AJqHgkpRqtev+bRitM5Jbi03jQ9Vy8bB/HasgCgoCtNZd
nSijjyAqZBcZ/5pGQTTm+DSo6KOrF1iEoibZBMe4b0YIb9TcrgKvFoDlchaNSAYD
Xob51qBsQ/Lj0djgG5/+01X3bVU5+mCDMjCsIHYK7aiZ452FHk1+zEDGxgyjUO3H
qi0s+aW4oVuSQgZ1VI1LPZqrwcL4MAWu5hzlclcL/QbIDjwcybldQVjvGuVGQ2BQ
3TmqC9S6m/d73CX/bXaLqnDShKN6I8Up/b7h130frVT9aR9iZpdVVOEa07Hd9n5W
N92OINNFEwH1ifd1Sr/pHVJVuuumZ8xakPKmGG5UDVbe65K97r/PKK8nLBI9vBk+
Ac6hjurqBslBaHY3+vIhbU4h5DnByCHKvgWTYiKP4l25+02ylOhce22CF8L8apMk
vn6grqmGKgGEXK9PQlajLkppTkK0Cz9MxZOXJVLdowinKPES6hFnfOuD/hN1V855
RsoagVRR2by0fi6UAUse1eD+MYpbPEe9Ct0TYk4pmJ+dmSF4pd6t1RCN4DNHC2q/
RdD+7JItl7RsHoN0RSdoyToYmw00xZynoj7p2DrFJeWutDQFVPRfU8AKZZG2bWwp
wexwOGNYGE9X4sHm+ohuy6LA+gxonqIu3DOcskUqG47oGFvUAEqalIuZpwWMveN1
hejnMVOZmfU+yaL1xDcdZ+4UUQeF5hB/x6hBXnrpAinSerYVNvqSWx0l9xO3YkrN
rU99xurNRxRREIcqp5umpx42SRJHbz9E/3mWxHK/ssJUmT7wyLymdMmtOm985GSI
5Q4w4nfFCBQRbZVJqu2RUT98CDE233E1BvIQEs5+W77+Bgla2e6nBrJICzQVAQMf
r6bY8CGPbGtWKVnZzl1x01blQeaYl7kCfI1sGl556jT/XKGlp3IpP5wnvqwf77o/
bwNAAcVvrSESkEJyanRb1PBYEoeZNGaiS3j0GQ6Q2pgixJm7SiouZQYfUNuOreDk
j780PwBVGIQ1x97wqWmYQStm5HOn/AVa+6KAl00VRzx2tl9ZlNArTq7UUIprhSWL
fuIkIfAVTeNT9MXG85g6YkgbUy6LRkX7GRUa3VB/GZYAXfRdZyQ6oxDvaEwlaTYK
0JHNKyLhk4/m+QMXIo3eSDPAU6fWta61oQTqwCvsor1CyfbiYbN0eQmnvKSTbaVr
GpDdVaPBLZISR6pp2OR+MMKavjTjWeIVHzswyXeX+omYaNMvwphypdC5if7KruoG
0vNHW8wopFyCnMitA6mkfDw5+rnAQytepjZKeqtW0FbZ+AuYmUzUeuZBBok6pkvW
y/SrLFQt6I06q7Ow40nH5j+/4nV6nFDBbYptMcgBlm8KFkUx4vTYjrCF95XX/amE
dd9lPCG54a3Cw0HFwYrR+vFT9fpZ9DpAg+Xrf4gS6bMCPweZNIqv9YxI00VllDZI
msJtxiP2xP3aI3C4UvGCAI5la4JepFk8aAZGIFS4Xkl4ebBjoEaUdmEZFq7vGjc6
OtHaR/xRP9bR+JV6p49E5GyoI4dG+P/JtO305sGseQS8ezF/z31+EyzLVQmPO/Qd
ScTGlqUpOnhwSZJXeLpFHqrMMHGkoPe3Ab8MURW4HYJ6XGUCsbgkJKamJHxDBgWA
bCaQQPAninLOqBzXB6EnLNzjfKWcQzWE+6louNeoz1q4l0TRZNsWyGTQ9b32rfkw
PNAzz2jSlGfYAeDZYSG4gLXETHrrLaQrqcs7cEFIkhj74QFdLHmv3MH7DMJZCoip
KkB+Tm21wkiz+pjdOzRW8tlCQTDaxH+vCRb/GtXnZ8bphu6P/f3erVNhS7ymff3Y
mIAejXeJYx+Rl6W/lOyLwu5dBglVlbMuER290CR9iwnG30oZEwhJX95y7m69i0jS
gHRRK/V4LDYrRE48vsKrrRim/i9rhmkRMX3bVm8rGKmz2qcbh8LVQwQITQ5mqY3V
cWRw7iX3lHsJfbaTucBa7/qbDTbGaxaU5sLT8hyVZ15HKU27lXD03dfGaEF8rssN
Brh9s6an7OA5sgu/XNzZitfuB69ab9A6OYAP0IIILOMm60MoLzfh4m7/E1y8AcM5
T4eDSH2ZauTGS+0MM7Jt+IKoZti5yl9fipgtmmJoTSwMvWcd59ibCDFJfow40oQd
Nh9b1YFc3Z116pnkpM1NjSyqWcf4iUotnkAPtFNBn/xX10Y+b7LtbzNRPEmu82tS
rAceJrapBMFchR7lNf0EhLr79HUtVQBkqYDU1E1G/VVHznSLJvz5D+KRTfTVXWsy
n8JZP+SSC6WiDxpB4R5A/S75JG8UmvFN6Xqh9gNdX8nsyeBlEW1vutm5efIoxl0j
jhAou7XaY1XxVVhVMMd8yoSZLqi8Nrr5vLIj97ueP9xuHIZOonKtTIrr2ljzlYhM
jztpT0c+3prRTNsg3z7zmiMem0C1KL+njkQo9LRfj3gHbmaiJAfZ9Vtk4macKewp
4u+skKiiPkf7j/uU/ePzYuKtpisL0WW4bpymFrW+OhS4csSWB217JJ5A4MGOEIsB
Xrv8B5gBBTDnJwHDZsJ1LO5fLqD4Ngrj27UkrcTS5gzS1CBKougtUapm0wS2FIUi
iPqJ08SaO96dB0/cqh0FxZUUMyWgL4qcjgSEQQnqzJIYa9CgDH0JfRnuVi8EtPWa
TPiO0yVgw7KGaJ9DzL0tM404IcmikJQoGtcz7vL7Ywleuwf/rmfKi9wOJLURcH9K
3pwnX/YzvW/1p8eCHY5B/XOia970v76udqrgUgpqbbjYNIleVZ3gzqOHFthKTUVo
ZDpBtCK8GAUftoPEGZR+L6jrT/ahLwViDnpW5fGPS+z6+toQHJ+MXfsQFldnnAwx
/bPO17OrG7I4K2k4yuYiwvBx/he34aBEQ1rXBiVr02XWrxu7LPyA9/bZ7s6dLSt0
N/sKJ49s/B5GoXuMKPIENmWBALb1DPoKZAiE8NwnmiQ+SQ+JgnQesam+U/me74lx
f9gqu+aT4tO19XYVwtx1vwkWKgFeqzpLeUfD0r9JTwREmEXs5bHVNAFg3yT+Pwnr
atineLosdqVDoPnhykLSsDSAkT8P0RliNv3sN6LCJaBnRqA/UeJVvyPfIH5pYVai
UfhQaTyXL3Bbnmitxf0Zzb6YOVqXPeY4TcBnjXhumKSgAvamLgSww4TthYMv+ulq
bsYloxAlIH49lyOS4U2LKc0YlJHxH0UNQyxrOb1tePI0Bg9DEsuI5kymZUlRdQ4b
0NcRL0Jy6G7dwmA5pnNEdMBcKErPCntTglqFOh9XUK4WbB0Q6l8Rxe6JsnxTwrQ2
sXshXfrAwVMwHfu1+UXBMW8u/6OvsdpUKbvI1G2CpDGPAWbXL/zMHKK2szbeDoz+
ULDGS5qtCEWOaOujfJh57jql0IefvtOp2KOfBCwRwrLB2f8eifTVLupD0BPz12E2
HSLQ0GT8S9lQphL/uCmdDI+I+E6jNoVLaoiashZ2RlDr5QvCIrZx8OqA+oV1hGyE
e8d+IPj85+XWPj6wLST0VWsw7pj+kL3E6Kq2jlhN+aWkiQ/+Fu5cL4JnqLgsUXPn
EHfTqP0PIYQ5hX6GQrHGII70kkLcVd/iT95Dl8Uj5fhvOK3FzIIsqkqHzi11jrNa
+vosmvs6ogHKFjFa16ipp4meQdIeYQYeR/cawS6GV/3FCVWNax84uif/MZ4GZQka
tFpNBYBhwItxfvTQkCVhe5DV/Wq9gYFsqZPlT3MRb1SrSndLdOHezKlnOu6EQCfb
m3SnC5pWm3mnfYA176gmFrQ70ZtW1PhNypIhYIA0fUUfgFjKNYGiScYWr9hoNFeY
axvQ50xjy3z4hlqLXVnrC0B5MvCVg0XSsedIevfHF06FLWVh8T3tqT8CUVDLnjoV
8J2YI1QuR0hkZ6MzuNUUX7nrjuuY5MxYgC67A+SXnvMc1qW87tn/wO2yuevHPfVI
ZizkeAVWkSUEyoaMUuV7CQI9p836GI1TFiILtpVnn/KPGzPjYnsofRoSp/a8MaTM
MD08gmYSdZDs5AUEuuG5Z0OR/94O4d6z7T2AUhET2SvpIaRsHeqxOhI7sR2rEy41
SBBWLSPusjfz/FfMHv/wT06LXlTeGAvOaan3Js2bP1CS5pPSHM7CwmXGzPSIcKAM
nVKNwEv35w7+dgJWM1SeJiQIOV5MUD5IJfEZdDH9sy9bEkaTAT88urBEpssgjkm2
7C9k0rnsug4mKq4QS27yPLS6GtTWD7/5AR07T14cBEk0P/xOEu1oQ2z7dKGdPMH0
QwlZkNfLHJRnW8Y6ITFQFu8g+cCJ5ExeamZ/mOFaEJZwUAxCukSLMFQMpzVbr48z
VAH1peH3fWW3LPazuizN2Wgf5oUYJccbp2BKENg9e8m64Z3qpRN8yDMfNajh7q2L
ObE4g+yuxV9bBBP7E58xTIBEPQ13Yqj8qOg469dyklKCOleEWSClnWlSB5M2yPVh
4SLRAwksqI7CDo4Pznd2hscJ0TgxSKVQlX/aovk1MZRvJTrvUGMOZvPyAW8U97Fg
UhjlQZNaLm+dbj2/x9ofjLkcFLKduOnpTcJtgVfYskA5YF7oYo0LLo+/wj4DKS9h
+43REP9bAzFawrNcwG51+3XMkavTrDMr96APdsQk6+ZoWZvu61uG/zP7ezfXkZop
1WX39TZ5PxIFUXVTDD1wERcGUw2cw5Dr+Q4DgFxuPTGJpqfAuzBEDA+BvnsNrZyT
yrtZEMMFuoeawDPqcYAprq581FwLLijjKSyusDK/M5EGiVvg2UIzs1GXzlCWQhQM
owY79z2bzluFInvTLSURpU1+KEgjWxMKZ2hw2fW2TgpfrZGoovrbti3qYRYyDGH3
5udTaOvChBXXjSwmflBVnqEAeVwKgBANeQaUSqF4zTHcvViyzmSCqmuherM5v6dP
mvJfdO2wEi0/zy5fAEbNWg0xQSmYxFVygpedoM2u5jYvHU5WSY+L7RI5EV7ovFWs
7z4gjYrITQRnIgec7s0QvWDXtLbTDHOubbaPhGZYFA//nN0qTwtPt9Nbi0CIPEhD
XwXBTZTWfSB7fvczmJP1vLxxUKEkZt3ue+v8hc5zqEoGrPidHFkGn+VntNiJ3rab
AB1NWiJC/oe/BAjGGGOLXvHq1O+IUNfWwa8x2rI+QleEfdJIKWC/ogDe/QGpvfRj
HVVX9vZ/kaKwQDzhhi7KQ07aT+RaAOFGA9/TTG5WDI1KXO6p+3GeFEYuLL8yRp0f
06/hfGKLfGAvEcjkQO2WEFhqMsZA47+KYWcjX6eVZK6ePOZgzYQ2pORpQvzjVzM7
60yn0A/VQUrTxhjt7vgee2GFkO8tfXc8O7qKtih+A9LQrwiunlRf/qQMCXQsNCeg
8iWGd1UZ5z5WW87GBcruUA5cuxpZdnEfwyS25P8x4HvWVGIPTgLwOX4cS/oq93o7
0uK7G5c0qrLIsUTRDYUptfxcF2mUYtH55A4XSpIaFIcpjZs4/u9WXavR1aDkYAHr
jjQP/pAnk6ASa1A/LgeagSug0TJXBOLnJakTwawo5+SQ97q4rY1mJIf8hWdT7ibn
KQALUPCJkmnRoi1o3z3/uJVLthpeBt586s1KAXl4wIPgaPWwhft2B8aoPJH/M+g+
qk80mbK+/lvDXoXjnIYexw==
`pragma protect end_protected
