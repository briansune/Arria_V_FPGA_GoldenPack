// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:22:24 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JQzMcDOpr7fY1e/ffJdiY2Mbf5UQHjZztbN98pfwVzHj2zMQ6Fsk6cCpSMjNdx/v
m4BMQMHrpv3FkDvPXGQP+RdH8ajTMd8H00lV7aNcVt9ksdtSgtPbHflyN7h+FQCM
R+J+U9z/Gh/cFKDmbl6Yoe/k8bravLKdGGb+kM406RE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 93888)
eJY01PDguCGJkBAcohK+TMhTFRkvK40zsB8zxrRfrDHTs3G5/I/JjFrgHUeLofT3
zVKJmy1q7aDsKVZIYbkMPOHhZvPDb5QeKkxWhlBCJEvtVi9Kk0c3b1fajp21RACO
5axRq1RPwT5NdHgqvsNTGwtoZFaJWp+r/1WjhTEZL1xOg5v0RKVHdjG/L7BUC0d3
FIU+EaBTzgIpc8t4cYqbNipvsXDf0JxXTVHBdB6bW07BJPjszMAHz0F+Asfau6EM
mEW+doaP0P3oBJprpWS4IlKf67JuEzt6KaYRGLp6kpjU1ELzqLkTFHuanJc6yXN2
d9S1XlqFAy+3r9KBz0Q2T/2rQvcUitWWQoltT+Z7vkmlTXXnVifm2BSdLYGVjrpK
nItI8ToRcKB28B8tey4ourGn4zRiM3vlXEMpQ2FxezbFIvq9SkjQ5W/Xyeh5FQh5
PmIlE04nTB66FJaNx7ijivrOYlzX1wGLHvg7os+Uwxeax/iQ+ZEV6bjJYiYVH8vT
FbK87PHWkCSxV6NA4IKH1JurqfyDQ6sgFDWQ3S7/DXQW+mDCa7ewqtfn88RKauhN
E9WBKRXzMUWtUzADQFFpNaHQ3Aq3yoIpflZvufOlV+Cx7O/PyQkhgFOnT4oNvS1a
uSnkcWg3+lrQrA+PVdRsCx2bead9DpRb9jEBkjeJrI2JZWVQeUh+kSXF67jSJoRR
bOy92echUd8yA3jUNtVxtzTIOFuhf7J28gjRYbi68Mq2UDljhlffJmzyUM6BFWn/
IKnBA3audUrMEh8/GFLvRXcVHvcE+Sizaxxp4h1X1gLw52nuqo5PiJLuSAVPnxQt
cTvYqSX/1KPS8H/hAJjA+085W4Oq+6Om+zbq4RJVNrjDxSxyt8VrAIjrR7yByg/Y
jpNWS/QNWTv1kwyopEJ07CnMUzUi9MDOKr6edXqJolihK7CFjKfDMO3fEWa5fhbQ
sjxH/AuUfgf1Y9Z1AEONwAIdsdvA/wZW17yc5C9r3dMTN/bt/C0Llc913uK3DHlB
fMXZVIt3PpgF9UIz7uYe6m4F5epBYbOeP0q7AnONT1KBM1Y9EeelYE5B9Z1LSJ0E
kyWI7UQh5jT3ziZnY4ce58z4bV1NQTFletD4CHh9Ryd7jpd3mCcF4AYPBZ5UlrpO
+eRtUfbPHww16/hizxizihB75p90hA9Y+TRtVcoH0iFZ86pR2urct+cRIoox2C/b
lfXSnAAp6qY2mZLux8A/mxpkfN9drIPdO9dnMDNtraLInxOStdqVxJym7nzdbUOr
M99CTD3th1SmvB4rYBQhsosM3uBHI8+BeAQF1eDF4/crkfn2ixtavIXi0ZXzshUI
78n/30oywABdwQN16Bga3astWB3+m2dBqPnwA4wqNVpLVaCeAbsNDDXx2Oknz5mc
aL9qUcf6OAjPjxEfnDABBSiasrYIlpsHfz4JsFAoe/CzVYC0uzy60c/H1BeSqxYy
aeSHFnBq+EqkWbFcB5wfqrPfjKvVMvktYpVomr0Mtsl/lEbdLUj2Dl5+OXr0rhVv
UzoF8HBi/k6nXVUJnfrQnJ+qRQVlYTQR5RHUpelmu3Wylj3vNeLFXGXfLvWZ67lE
1q41T5KUYkZCizTeM8u7cCRthDyw5atPP/Np7d8//WRCq8SdK22irK/3/y/V4Rk/
yHpU5pQ7MfdEe8n2g9z3sCGSZOM9CDqSWt+YPe2xt4hCymZMDEacDcA+q7arrD2P
qVjJWRvv80m8NCRcKGTRF5tuD4aXHrm2mrwaZFhTz8AtJZf7rwg6VcxmwV/jzu6+
2Lt8E04ufea3H6e/X9cjgbfigCboIf8NdGIf16txUEJI/KY7JdV20fB/E7tPfLFj
TSrlJyunZmA1O+0AInbj1pube8xOAv9lrbRF2+46zuZpyuRsKTh99Tco1iULfcU7
5UiCd0SFGFv7unsaiw9CC5C2nobA9WjDjPVHHgaFatkAij9TFsBg9JR/OVZ5H6U+
r/uPLtvi8Sl0zFFjzaL4+l6QstIYw78MuUrDJZ1VWgPqm64GysZpCrxo4Y86NTjU
IqocLAx5AAT97SvvvVphddPSihBrMM//T0OjLX6B9wf66RmB1/89xa/KIFp6av/K
z1XZfonF5J4Chg6pgK+sHXx3tgJIi2meOur7Q6qN/fPPs9n/3IhzKjUxKj9bReUq
s8gG1k0M+7aZfdTJStLB9ljiLZ6H9G87BLXtn60cqQlW2/QE0GqkEabDq8Jl071I
VwUF7Sp11xN+nFMFfM+ebLAGW8IPeslA3TOic49xUHiPsp9yGGAsHCB87h5J54Wy
9sQy8adOr8FLfs9nxOH45tW0nhr+84ZV+dNgRDs3qKpa1U5jIY4s7hw8LQwhKinx
hHOAf47ss6e+rVphL1jolDP72wbRJw8YFvd1u4OS0VXBwiqb8FjlONKvwGjUOZul
csIbi/44x+5ZiFEptMYZaZkNNjXJAby0/hw0P/7E5aO/HypobohQXYcMvvy9jMFl
PLwf88D8K7Xna3UlWnWqj2kIiFbGlf+31mZuRg9gsMLYhouQTiT1uBbBQ3ZE0VLm
L/5SR8axvr3l+h0Vb9hHihPI/V90WeocECi8K5hwDRtwjUoJy5vQbZyx1gNrWlIo
s/zKcCWzeecI6zjdZTHQXN7PJ9gZRevW0k7vYK7ijpeMGz0ru0d6X6UmEY63RmEM
Ria9ribGXky2Web3BZ3yD98yVrh1JfH4yLWTPJzYmx/CVEXDqbUEHOooS0U7n6x0
V7pQseXhV+GVULMZn2J6kQRb8pQqjXVfEAGZvwIgXcUShZIUEaJxH4Wb/VxVhy4q
AlYL/olclUlTgZlgIRCuIWQlCtUgiR0lLe4+rgae3VW7DcBODLpegEAYlq6G6+a6
AuL6a3Kw1yPvCEiVoj0qdIaVsZ1WYuvHbgcE5whjLvWP2SxmE1QJVEJdkW8NBYM9
XM4pdaKsPFBITVYaeu853trc28zRFTAFV4uldpuqcR3hOCjlEH3v4PPCK2NyNHf1
qMSP3xUG/3HrG+pWIPLgPEq3b2t4DxRWNrvRY+UdaJtzLgwkBpVPYCd1QcIwCYtM
pZ6fqIIwD6YwTgGKM5ypShqNkP3pQsNozEL/Em5LlFWA0Q5YRGbiqjb8SwZeYvus
hAuaeAZaSPIy1UfJ2dfcP1pAeGSkGc44/bfmGjpivVcCO8C5IhMoRHvsfCwL+xDe
D+2HKc5lmRXrPtqQabB2Ij0+9fs2HH8ZO31+3nMeLPHFGFmOLBttNyhvwH5KRhvh
6fLcpuBIfOI6euoXaZB6FjMMJk19kQSQEzAyZqjvG3AVAgGj8j6qExPkBzjphJ1F
A/YtWZQIG7qkiyO+kF/G13XyA1g1XLD0ocUZEk+Kr2VVHGzhx1UjI3TtR/QrRR2L
siQsAbWU0i7D2hrOktghC6GbK7vM91ztn6Ly+PVg4Jhmh//0jqF1OZWXr4c1G8xO
Ry1EzMkIKuZBr+LJAFFVdM2unL/YLa0FS1PxlWA+lr++QsxSeMFq5uGUzm093UA3
Yzky51m9jUVGOs4fAZJu5lTfvbdhF5C2fO0MSai3Sg6P0iWoQupBVWuy2YhkWamn
H+L43EL+c+qsN1fafKSlcx6yYNNXK12n7uwL8iW+ml90bYY2mWDQamQ7jclaeFZz
a5oLlj67Icq4VA4OJoMadxUaxcecCTum6tXAFxxE3vEufZbMjDnqrkSW+n0W+wXJ
ZdCBfPY6MNTo77qHpcCKIyEu/seytxgDjZhY2l2+kpPXcr0QvEnJw9f4N18Ir+id
CS7jeNXW2b+P+n66mWSN9NfcZqvF7UbM+hGX9QnhOj52nlewmmbRXjrr4AxBOzri
9gx5JUxsVdprkDl91O/yr8nBZ8ElY8tNP8J3hezIGSGC3CfiYPgGMfYeHdSKMgek
2pZivSpNEBKlhJh+ns7FRihz8jdgenXBhXNwSq/Jqd9cxt3xOsZCJjDvXTgJi+od
ByCEpAZ+cRWf1R+zVPmLtbeEsjP1tl4jnPD0Tpc0JPNxCKidU0f8yaVLTzKOAfzp
PPWfsiV7kvpjT+FDbKgIqcHF+2eC4NZATxTH3xcxwZbFKebNH1IYDr3rWXQRywyn
X7G3Bt0XhV87EMMmuIwgPlZoQ4cpHWdUG8/9XdNjySUq238/H1bRfM1wXEkadED7
pCrV1MSsCRNYX3NoqxgTnqBW4g2QnK7UMS+CJdWqc23Jm16472xqX50U1jbP/BFR
ECX551UpHcm+Zk0qTkXlObgqNPsCQSfYyiCso+cf6jkc4JfRkZBGjNRXzLRLB2PL
1I6I7/nHGD0Qz1u0NxsX2uLSkC7JsH0CdOAnANr7QQDAFzEOmboFDBx4myMg6fIh
Md+9SUw5rIX26kWzcohRKpV5CscB0Q3Z1drciEujkDtGlRKJCe3ejtWxi2RQJlgJ
8A+6XTwuOLorzWM34668b73brI5QVvnxN/mix2zNyf2WV7u7HkryJsXn9dW2iVz6
p7UjkcqvsmO4fUGv3e6o/BFexGYo3I2nAQZXr51nrxq4XXHyOuPs2drIOv4S8cbn
77css01uodd41xMXVMf87uKh8QkcRTXIW7cjeyMluUrwEFJb8Zi9XVEloYsD8XVC
y+M3T4+D1ShwcXupEDFnX3rVyXiBkGAyjsfZ/ea1tR/X6mnK0a538WSJGhgnbq3O
Z3+WSAkVimAbLWYTlVhWfRBHT0RtPRpcf/RGM1wj4JJ29vkQtVduZc1AUnB/ddQY
QabBnf3OOjZuDIDr25uvvy/d2PPNYkL7GqXKFhQ5xVZqgQT1AsoSbRacOQveIFba
4ta7HokHq/MLGWu8Gv2eDxIN17hUo1vgcfp/Eb3a5IVeug4B8lv+ktX6C+sR1Sc7
OXtrcmUINH/WG2gviR8hxaBw4qj/sB73T29vLK1MoZZ++M4h01TZAOmpcgqwrDmy
q8LyFbz45/xurnhOKuPAyTQLVXKs4BF38A6qmwZfFumUYr0NxOxOZ5m926m7yJzZ
e/OPuH2g/LbAU1AaMmC+0kcQV3KEX7AJ9r3BJBxLh65DErNiCnCPE8pPIFl3Xc6C
TooiIwHcc/B5QC+Z9a8VfN/1MzEW8B/228ux6lH3p+FjS3VTKnojP8BoNEJa2HDK
YyhWYwxolBzP9uBM5njVBRoEYkQ1bDdZaG+p/je/Wi4brQxWjxmjBlS3vitW4gVW
nFFUv3QB58x/11EEyzhBCbHCEsGHUof00eptRYdFsEEquXWTchIJojvIM/V5S3bw
VR167gbZCgOOGUUGEWU7h3oTgOZNprh09h0TEc8E4hQT5G5fem4cCW9TjvnyGTrv
MCdKpH7cIlGSelbTkFRR2bjnjTRFsBqF8MxXAlGNavCpyqwJvTZRAygbakZlZUT+
2eLmPRGl7x6n6cz4SuNkrc0jslxdOtSkd6N9PkNbRMA7HLGDY610vlveHaYm7xKL
o761USZWrpadQlSv4Fih7aKoXxZm+zZCJTc9E6R3h+pcHg4Vh6qlR05ddSFVRiaq
WrT4HGJBlQID9avHgElTyrYVNd2CNOnOJjtDzn+GdisRt3JM6jduIK3c6RYFzy6O
GsrU26ktdum1QnjYvuI2dvVluWRDffydf3z2wCEEx+xyvWpC28DOIaK+LLpdRN35
e8oqCFvi7GNoDhoPWk2Sbibqm10cf2aR2m04emoXd8pSiRYFN043A+X6WEf6sWCK
CWZ2TBSw70MzjORBhu6RoB2ZlhY/d9NT/MlnXQoUiVALTsSD8Tpn8uofLV2DH3hY
jWFvk7r0lZ3ramnbwHKeX2bzr3NJfwiCpRtDh3X+PLPHTZa5kwcwzXthyvw7pAOs
fDSDGqumXkGkadpFS+Ia2WY0mN65OKCduOfT4/J/gg4qW0ta0OEksAvxrK3XuzN+
X7ZehZ9ZM3J+gF2kYZQPHT+DiXIxtHAXdXi9+K5AW3NXPQ5V1ionmh7I2X8m6BVj
0kqLZBXXvS4Nm8+rfgn+PnWoRl74zdYt53mPcKKAP2f2kWa5hcoiDqAbA1OJ+Uhg
+vysib/WsJ1X9sAWDxi6lnZZI769nNafTq34LDq2DoFQz9pOrwltINGSwGzZi9iK
5TpYauDB9B1pAzf26oapQScAbo+6oB2X5R7WKz5KnBJc0Ws74dmIrIfh3GZNa3T0
mPgNZMYZ+sRb0DqSvPaByLELEHEk3/UDAyQJoCHRUtKznBfKTHv0ygpmCUsjth56
ufr3gp6txBoyoJuVykNYhAoMGk8g2z1UYqCDIgZLec9AWKYnX/VNf+45VIIVd15w
LhjdT7yqha/2JrgguDoMW5svmfYhounrMWPEFjSIANigNbVK+aXo/plkOoMAZtJc
Bnki2WfquFk03sd4YXw62rfPyiqMBW8Cv08/3bDmBjjVrAmClRIQddtel/WrO99/
6DoS3rlobhjRWVEnbi7siYWgOJfBaEkIDJu9NWaZPpFhhyxnSHsjR0GnYx+1LYQY
YFcZbB5/3DAwds3b+ov9AY7QiOIKLILU7vci8bU48v5izz+qMHjv/+mnDDv324xG
eff2Mcld8cjb85n+clhaBi3GVM5OTlbtw52JM5Vnl5khRIy6WTVC7vW+ueo2ywTU
YeR1NnB1TmZSSSxYpOysAUyj7ipM/oCaVa9xV4s7WTERWciuUWJ160p+drD9MlJ9
eQbWzSkJ96UWOPIv3EwG/1OR3KzJq7OvT+UaHQW72ge5MvBCiwZuAiIwoeqUmQNP
yMJVKEfP4zNKpMWtpxUx0TfPT3AeHRb/jkRaVprHjjyHDHXfMihwIlfsz1c0lyLs
vgpoQtEEvfkRZ681JnxCQUBDX+tZQ/YcDgzReiEMUNLiqKViB+FyYJc9aPjkv0IM
b95vxTVvALlTCNh/oo2ulRr4w7Nwk1cUgjwkVoI5KU7KokIqB4G7Cbdhndaj4Fdm
g0pB1nQA81ufYmiwda5ARKy/VPnHOfqfhqK3pRTia6gEPJ+UoDy+nSQC/WcxtWcJ
9dkcUFL5r09xt1eddQhcrFb7XXBJwYgIFAAXKxwKpayrgXCrWpC1UU1I0gKMoamk
5G70GTTo+5+mRulCO6hsBQ8yd4Ie1dO9M7jkvSt9RDm0RPyAOFw7P+HFQfj8oQOe
BQLZuYWUKt0CvAten0tFA/xEDSMzy0rpSGbplSCZwqOS1Re6KAgFJGXz2pV6d7X7
5cOns2I6uc39qQRQBRK/AyfgfdwhrodB+Rjlz+edggm6DLIekTEYAdB+HtSbtIS/
eg9HJtIXn0q/r+nvydUz3T4xYm1eyzuRD14/27fj4gAcMkE6A+/jbACZScPI7iOe
UZvOSiZKLkQy/y+NgVbdw362wbv+LLggudEroi+P7+Sbu4EVKjaa0CH7CETD7frS
H/NmCyZvxiiC3d6xV7bRjC2DEzKFeYbCR2c/dAlhJ2ZDGfOYizxFpAVfG5EL/TQi
aquw2LRd7RsIG0jEpzRg1g/rvDeNP+Kn5UWsovyoNEuZ/P/8Y51nt5nXHkAoazmI
id1CA0E9MYskmOAuATQLAIFCV5sD6wtXXlSKgBYuvVgV73LPg056MSZAUpAh0w71
5JvFaC75p6oysC/9wUW/rTUvPWrcarURoOcV7V19v7Be46FZKd/TpO4W0pZSkzQ4
gGZ4UwLyH8sibSfZG+fxqxCiQgRIhbhQWhraEHuXHoMJpH3oA50ToJlAFJkho1Y/
TV0dJZxJPec0Cc+0JXs766rHKwWmis6quTulNPR/LQAwvcqShQD+OQlfU2xE6PyB
6Sg6fm5k/dKwnipdR6cjvSqdhDTbF0A6yr25xYdnYeVU/CdlK2mWELHAmb3cVfBu
MmFAGRtksLXSTxyfzOJEOZZUxjF10Us1Kde1r3xUkqjfy1sgOnEmJsKwxrIGCVEI
/D1cjqW4alcKeWmEyCUg5WzTfQq1MPe8bL0hkrsxc37TDz5pj6g5iVv2ju5aHjWw
hTd52p/CFnhjkJYPTRu2UzMbVEXGmOQDQkA5m6nNkBDDjtF/wYRd2ASDHm4uEWG+
i34TV4kO6GwvF9joqjeJszCCCjJRvVA+VqGZyCnvQw/JLkhYX58OkIdDS0UIZxmI
nlO6Gg3rb9XA4p6jt+mzH7SDIEAl6nhqG7FIT0Hj62J5jBIQG49e/NChC0E8Ed9Q
C+7z2ZYSJpQ3+yEz+N0ihICkYLvGc3zOS40EpIejjRagkUKQGuUetN0LOOe9oijh
QxNEgfdktf95KuYSskrgtLAQe0MvMCD1YtlBXj9S3j38zaorp54vd/2IktXgoJLb
GsQgk9xB0zuHYVH2nI5/rIkHGnp9kMqAUiwSyuZ47I1F2k2KjVV425cDd4EwL7GI
Emlajc00aQ8WZc3SaEmluM9FlvMleS9XtYHI72BopGbt7TVsREof2koUD6Chiiq8
R13JZJIVF9hPWhK7GLcYPpe/wsQelfGmJG3l+DLmNKS77/eJHOPOTUXb/yBLP1HA
3In3HQ6d9sp3/tzmfQGO7PdaA56j3U17HplsW4FmXghNfs0PS3M7KD1PGiE83LQ2
xT+NI3jcrd8brGkAAf7sNbgLVize3reYQIuuYBgdiIM9CGjYqk2O8EBEhfFi+Nmk
0qJIKQhdGZZLDBbllG6fxMsgb0o5Y8qu7eJSaNjO7Y61k64LtRJpDhH0CJkzR0Xz
+9XIfEBiRylGJI7wYij3rmUf1lgSD16Iydk7AsATErIR9CIrzFY3FkxIE2o++8lb
l+N/sIIaShx1bkL2ZLBZirmNkxz6dunvWD6BfNkOVqT41fp2pap9UUgOGCBsFBLs
H0a/lXBSBtqnw6n8AJ05Mwgvaen+g9cDhw/n+MwWIwgqXpuLMwUmE8NfARejmT4v
yO5ja/+Ny9sKKXYEAFi77z/xMU0pd0d/UDSp9bYOLzuqGjWRrBgtwe+DK2Q2M8m8
0o2QbLlAQUDs8/vucRp/iVFaaj9SpguzXO9aBmTxrFRyryKFYGMORuuc0uXVu8YX
XZcHuqkx4KQSpafIJdmz61Bsn8uvm/C2UIdFTaBLRJlXcVUtcXuWkEt7HvKWQR+x
YoWygWhJAvbz2JASozSiprqkFmmboBLwh7reB8RgtL6MvFCr/Z74Zc9QnoxNcXu5
MDkcgC+TChE9A4TitGjG7tZoJdIMDfd5X2T8Drb02mJJDIBjykB7c3bKFEhJIM6K
Rq+n/IT9/iy2xcK9V9cfI7OWDveX61xndTxx9O6A0es8U5qEWN2lujB7MSllOKE9
RjpJKGrsSsgwqitoBQw3PY3raAMaYrwBDKruhL6+bVEIf3ekqCq/abfQnRn52cCG
F0PFKG9AXmYamvhiqherxjvcEyVVIYn4JvodYh4bQEvrGwbyNEpnMXb8N+AXZ0pq
UfBn/ySuBbA1XOAwZvP5vOEAiS0vasuYpxe+hEJnAnPXNwzwjQuLiU951hHLakxz
nF11HoJC0Ikt/VqYGkhEvc66FPnwEYw7pIYiARgC7rTvv2Rh5N/q9j9qL6mLLC9B
AP9WSvmz261LrFsV2dlLvEvL9vXnquPvgXKRBJ6HLq3HzJRdmYQngDvJPjm+gP6P
YlaaV1TqxHpCdUrY7CuJwAEldsdZY4+UIrJzmHQfwVttH3ooq9H4Zdwp89PC43yu
oqzrPOu+CrWei1y8I1WsAQyY57frBZD59IcYBG/qKtKKmdP9WavvrS8ZdYZfoI0n
vq+oUhzMEUczTP+z4cKPH5XXGz8R0mRCGvkN9gzO9vnHIBIaxuyPd1cB4JaZFUNt
dm2TwkpXh1gero/YC0C94NsoE0zLoKMmnPjJTUJ4de9Dov9NapQuBi91UGAWhAkS
+KGS0KUCKiAEmEK/ueNFzoHTIjWbU+NoUqvzoN/hGxjtDHQ3+aXkgButTEaTS/v0
hBL3nk57EIK/I+IaI71Ws2pCa+5aj4lprNtxIyBhvovCDwTUS2etmsGXcwyT0WQ+
1RX6TUC6OVH4xNIU9MOi9t7uNxI2MAhp24YfrD5xliKo+aZtlsnCK3IBgOkWioJa
mUitzIrx5j3+t6EdBGxf7uygSRSnMCO+WK63c+RXDDHJO/rWO+EpC1bk5St5N7vj
fcQ8CnpUdHPo2gv/Scr/uGicmdlcc71ByII14LqFLRNezwjYx0xM3V7c9OgSR0+h
6U0S+8e66W71vDQMjoGWVH38hUZEJPj7Jjd0Y3RcF2dB1IH/XnjuphrMfS1rDWIc
fHDw9HM7oCrPpdO+FL/1Wxqta7I0jw2hGFJC0J2s5RSb0UA3tOqlbKIfGEzqRYWf
xnietlOyJBiDdQV3bpuTidzteicsLUAgiIKTDLX8nNT1SVieBcutdzf3c80lPNkZ
gLJXyVTjuMMdqVvCGAHLojZ5FWAxOOzgx3qHFOeyc9u7BzCBtRotCI6gUd7pZp5E
dcyYtZIloGoE5g/J4l/MdCSpAyd2nWyBtaAwVMr9f30Hy7nCsn2/xrZfoHbtOqAR
kAaBoThWnJyEMKYqbLBnflc2+ANBoEdWVSvnZSsteN3WIThfWgB59GAR6wbTBCm+
nVdSdORMvFIVDs4ec9nydlhcyFdFp7rRGPVfsBqp+s3o7198iILBBugQFhUCK+F9
HipUJbNFcsGXzWPFVYrPbctED3qhzf2o41QN+ykGxpGysOOLymEzuFyNoS9SHq8S
wTBilS3itKbD8pSNvdY79OaxcQTS/rPFu4Y8i21/BZZeXyv0Fa87Hn+pOYv2zTf5
SGlbYuYtoQxpPuT1IsPLL4C6c3l6F06BjU7SlStS2s7KKrUGJM0FCZh+FNLY0saa
ru1ILQQulJQIZ0alvZEDniaGvANOLY9Na0qfkL4dsnJzy8Q2eeXJfAZmtvl8Kjbr
dUNFRFZvYyh5tFTekM8kkIU+OhHuSL9h2wTxydmgOwmyL2UMRQYPoZ/xI+bTt4Y0
SPK2DutdfOyHXUgR/xZAI8jqx9AafMteBTZjUt4JStT/Snah5DqWFFliLgjoTNBJ
6YS2HiiwD4Dm5bbiYcPRwHTli92xm4nBvym3CgfR+DXrnMnsIsGAwgz9pL8WaEUd
Jm55eCtKeTTxts6wPlNpJk2TSYwWYWwjbcPNPVCu9TqohIm91EJKucSmAGcGSA8D
xiPQQ7b2bCb2eicxzrNhQZSneHX8RId8kPauh1pY9YM2qYgu7NtudoOAGlbaCoJa
+k9J4ETP6Tn6TgHxhMbs672ybNg7ngD9bv2SfI/N2Fv5I5GlAGaPHytBKSqGlBcF
hZ/ZFgn9vnLMHPXEMzp9Xep4scQ+yTWVq6+242GmQwxXHOV3i+G4SIZ0NWCrroz5
dyewyIV5U01Vh0Ux5o6A1eW8qTsytmypfjPpN/B1l0bjZm8WucUpwbFkJz37x3hK
pnwytiWGmiSC1wX0G3cTPvdiv8Pigi2Nij9R6Lzg/sbiJI1+06m3pqMcOJfO+MK3
CwVvXUHv5R7wd3zTZOPMNRNXCTRJh8by5yfyMosdFhh5KGvFPXpxjsQQhfBxqA/G
H16r6H1yEs+sqVSOVFWyuqEh6vXNTweudh0Rb4BofxzTY92Hmpyp1HqcAIP5oGix
DbKmRfDn73VVuA2N5/SYSt7zi/26N+cooOLe7GmRgyjEqwZo+9QHZMwzTwQLYeDA
zg5Sz0fPwPAAyCcgIxHl8OY3a5U4XdECElQxXtU8/bdOdaaFHUd9rkeCuy79c3ur
vDkemuERQJAx08R9HgD2w7CeFVnCHzMxBtrb5H12h2yaOxKFIvDYn/xueRsoIs9q
T0azkG7/SAWg5N1Pf12Bm+hlsqmnclnmFJDGEBQBkQVh3lZM1j+jvR4M3ej7X+jY
KT/P29Y/1AFb2ydtHjhD7CRMVYnVvKga5ovA9NNNwd3f93yx4xXn2IeCIHGHMiPe
wgEeeGH4X4oES7Dq6PwlJdRwyfz1rHXNVB64PkXeCUXWi+pSJKo5ubuhgjLew1tA
cL6Z8JDh9r2/fqEtd8cVSirAgYl5FhGi9Ll1wwK7HPSNs+KpiixTCyApdFYXUbDi
D6oYdldXgV384Jjbyb8amAGQ6tHX2IOiNA/AWKK/4ZO9yr0Q7I0q/R4cuI3AkLGg
BnB8zB8tVJhzq11qI9av0oRJvnIl5vTCv1TzUXY6sC4nMAzu8A8HN3Yy/SMGn9qX
12nv1+M8IEoVeVxog4rDDnyQQEL4ro+eQctljtsqRPfnDxCfXQ/MqsO0wz2xL14N
D5wR2GaAMqtPzPCtxnDY/Jrx8pGrnDcMn2Vcsq+lw1npb1aRAodyuTNmkA2fNySZ
vKp6blZi4t6Q9s6cBgeIYS2/R7L7BGJ78AtJpod2YP9fwbOekBM4YYbPFqprYr5H
OBjjhVg5NsItTwkuFyvgMFvsMcSVvpdtNi5wrQp8Jq9gA+1KuyuhU4CSoh+wPUK2
jcCUkdiQ0w+P4BAaDSPisR3UJV8SSoPEMg+Q0dxVd79IGKGzqElZBRdipnRN1cjS
WP2Ft3GMFcOUeBxjIwH2jkKWBucBkV/EiJRdyFrBtQnO5/nRQzMJO6nuOjg8Abn6
7Dasdh6rmIaT9B89tsEzll6/uEemZGkh1BHtj4i+goRBlgrBfiGRS2gJYpv1EXc1
Y4IwvEgj7qPcftAx+v4rvTlG7OKGgwEd4byifEoTFkfLHDu10LcKAB0ZHZ0HkGCK
U8mwJ9JH3K/LacGa+h/bE8kDhn195W0ZDK8Q2eVrO/O2R+B+GPCmLT6nnj3qH4Vd
l+9D5vqX/q3C2/MdzFtBUemH3kmQ1gfvxUeHQoTLDoHX4Atr3fuL5Ei/t1Shi9tb
8JrAEaGr4TF2QRu99bqKBvhT3P5xll0S03qoGNOQN2MUegLcdk1ELLwvE2OZWOTs
VvdxC/IqbzpZqATTLR5BIhxLJQPOQENJKnWl3kHW1VvT1+5lHudXEdP9jOjT0mRI
Zc8Dd+x4R2JDfVLr8elKd5gHqCjbLzixmjhrmqHoUvSXHjT6nI3Q3i45iGueCnqC
/U4yLNx8pELneEsqQLXtKx6JZNVJgag9/k58ie9vxmRuzQ2QlpJE4StvfSGI3DTA
/U34oLcYOT5qnWJJj/psYtPzE9z1tatTR/oOqZMijud0M9LoRQi3A82HLi08hcwY
fLfxpbR3YYQG2BKJoHtRhcOzcs/QsUjic4fSGC6QvzPgKRjB8E0/XtuTmnTfuZbb
O5rVak0+epmISAcqvA7JhE0p/fSvfl2ZKqZVZICSEy3bcwe9YTxMP/GrB+mZ9Yr8
moLob67PqB07PWVJ3MNjuUW/K015UPwcr0a1/ZgBkmgcpPrU9XD32mMfdXr+EcUs
pUs4LG8bvACCVeeFSvROpQNVnZCUPiWgI+l5zhTrdSDK/ZhOuB5e82+EjtIasB/m
NVp1KJHZgegfzlEK7p6e8LFe4bwYHpcSk50P7itRkSKns503Gp+ZUAq2n0kr9QI/
XKl3kDZQwA3kpFxZ9awxgpEMipwUSq7r9uwa9SC/zEsuAm9Q43oirM72f/e31HEe
pR2qK0dX3VqLjqNYIVWVpmRmvDrKlVRbW0m8jVuHi96/4d4YGTYEztQ3LKciZOFT
zMZS3hbEFhtTvLKrNJaP58W3UBJP1ql3sM2uY4nNpXsRvgdBk3MD3C66kxE6TqRy
IYzKwX0VHANcEHqMRy5Sjnjl77YmBu/Ny0i2gd5C32zuqnZgTdu5lnLfbpoAbG90
VhhtT1MDCyUyOoF6zA1di7DrfZ2hMoF3w3OGUL8lq/I1VN6Rk14CGDhMU7gw9qxc
NlLk+yoMHGFOji46FnUr06OMhrahSTw/SGgH7gUXVoxkfbo9/1eBzslw7p4at9Sr
bQ8vHYkOoIVuued8EQSg5vXlu3Vn2qrwkLp/08z4+nytsHEG0b7sB188gRgpuNCQ
SEFyxNiZ0Ansbjv0noSREtsZNAam/tkQvn4UT4iRi+N39NjlHnGIA3JM2EVWeqPS
tSHd6cYhuIOSbNJvwyfgv/0Alm5505Zdql8LmCbpMQ16KK+Yjfbg7f6X+A3UybeE
CIuUszfU5XyUIr8g5rVnBj/3p9ov41MHTh2bJ3rFxYjzHnMekeO5vbCRaNTDTRdN
4rbH+RNfmYWZAwbC7mxEyYFxXhWOaE/NQB5z93XC2kP/+ZZXqRcju5q0arB18vmo
sr9MEO9b9Nqpt8PeyEbX8aS74xidX5WhEpTpxHPmefhq+NB0hERSIUIJ2RDEC4lD
BWxNxaWWr8eCnxbmu+JV50BGyEAESVWwbMzKL3cgN3V4U4JUicrBa/FAtz87squH
sFu21pFE2oK1TFat6oG9FLEIHMlM1Lq6fA9wjS7E1H9eFOgPYsMedOqU3TedvGwS
LbCYztU6UI5Fz8Su+emg5F/PRF/1MOFZMlLeISOqNASex9Fl/lfqZK0VK5Gl/WFc
yc/axfdZ0oOB2Yq66nTS8SvLIURNC2wdwzqBRxVVMqzbu564lmbtKOANgNw9WKfm
iE8wXDves+2gklBvewAtb7O+R01/jV3U+w/zCOMnQnMuXYzYPF0Aw82aTSz4uDso
QPTd9eGmiSNr8yG4XvAb62NIZQiGKNT5IYnxyoxdNU4m+7JTZwIcQgZuTXXWUcnv
B0x1vTJqIGlSd1T5yEPstZEJZ/KcXD9Zr43DCGNgEGnNBag+W3D6JoDw81+hZfzJ
lG9i+uhscNq78DqaXgNewJgGDhLq1Uw6GX9t9ZELxW2GSkE5P8fXcaGCnD70o9og
/ZqSn75bvMyehZoceW0XGtlnd9DYGx/LcS2bHVoWjj9R7d8bQO7CkN7013ahWHrK
0NgGLTz0EtVl7N12gxrFKQlit3dQNVLfdjRdRdyn1hEcHm3WTZudnliDht+CX4Af
CJDCniJIOHZ12A/v/unsvsAZtVWkmGA8Pmg3+T7GeiBmMWPHROef8ppSMOAimTur
/Z+hQkLa9lvWOw+io6nxo4uqqRz/mthN3OdQ7ljlo6ZUZ7vRlvv0BXwEhwshUxhw
DguUlkIT3ly7UVixy0vrKBcM6FTESQB7lo2jQpvJdJtyYCWIDt0h0RaMwXnn3Yhm
G3vUidgl9G/G0gHVLg+wWVGhuFlr8brw7WdM9L4GJ/nXDFdHDE+RiYXE6Ng2Xy2U
fqbr/7z9aPPrGpyWyMkDI0wCo6kYrv9Q76XbfeKD9cafA+2LWyp3K4rv1IRvOj0i
dxQiH2lEIv2/GrbqwY9oafnmdICyWIpKe+kyrjLf8cxUahnLcVXZoMSg7295qEOX
gyg7ywb0gBa8S0t7Es4dEC1ITw45AVTyAHLbf6arCIiuG1V7MzAsthOSBWEu3dcT
0IK+B0/YGDTaMekoSNk5uKpJdbfbpT6d/oTf8FFgUZQOuA+jhcg9Q4UC+YRqhtHx
7uVNtwlT8WLz43rgTH/C2DCIYmasjGmkq0Qpsz/7esUgnkhxDoU/G6I0FkIp4dMK
Zk5euiXCguhCEkNV19V8pr+Jd0eSAmDs/dpMTqbkPXqhnoBQ81KoYeYxj44rmJ9R
e1Mgo2ANXf51Oz6katwcLUuufvHrjoOIAZgjkMPlULd9TdW08B+unvbkXK43vG4R
wpzCtbvtI1kxrZCIMeXvQh3fmUEO7aUqY+rzaLQhV7JISpTsz3q0YFfgRptSdOKq
1f0L3UVhpQ+PiL0lyMPauEcrVIt6iJHoYJOSRy/ikRtpF1O+AjeUXYlG5v1sOWmV
Cp20wjr577JdfvsbxKlThrMjZR/H2kISNG393Ve4jtTQX6oeU0ZM7xCjUSOXtPs4
S/tE3IBJ+F5ehqNLSG6UKopZG5/Qz05xPkVaAo7GEoHrM4/MWmbrN/8J1SrVrlL5
QsUZ1g3YVW+FBS1akcEQ8knBsarjgYGWlbTkfaYNm++KBHWvhFdzQe5MoUDOoCvF
u9yj2wnis1J1w5qxo5mBNS4nba5eLzx0+UrqY4sbqj6RpY+SAVnqELPRNnunFwFc
VZ5SU94D/4dO5nLvpobijJ8kPm6ueg/I+grbnVUsXk8DIKhFVgQ0fJpIsKUJHe6K
+fC7Sm3ByhPceeyZD02mz4+KRDzFo56owwZY1/R6RtrI5/fBJuOzugLmqX8DCcqy
XwewGmW7tGVR7ggvCNnEv+03bBW4sZkTguoStuJir6Efx4cXgETt/SWWTEH38Phu
6WOCvRd1PlvtrIFsMLNtAdwA/UW+FdX7aaghbBKVVxKBgkeguXTGelMjWwHvrtV4
JqTfvpqd3Y1OCFIIY8md82ffZGwFX528mqxn/6SS/uigUzBd5J+jiHaxMaYQwGYm
HDrYlDjzJSXMngkkb5knym9S0/4bA16phEV/a4MZUkKV6MjOxGmD9NY690wjECvL
p4Ad8PDFY/JDkTrxmuiYjM821vJjaEUN2ZKnAMbL7IWLxFWY/i93gvfMpMwpkYoG
ApQCP1sZf1xEbxtlXSADPmsNb7zWM+WsWP1zub2rcCawxyEwEr6kDFzJ3JIQ4I6T
hfNLHI5LCUkhmzSMCcZVvuLZXv5fq1QLN8dp5KYZ3tDYd4ugvmB+ExxtDW4eNxgx
gZpQJWVxWDDHgmR/6ixjtuf3IO6oEZnkHP9aGryq9I2ZR5V+zthGKeAb6W2MHNJM
jtE3IoyuC70nHyILAj1irQrUKkJB8BbTf7mGB02L5DlHYm6YNVrNMBkTfAzzHnx+
6e4EdTDhadk6klqOX/rJL9JK3K/CuyY5Ers5xk/CciwpMiv05R3JH1pewf4f9Bv7
slT1cgoxaRCIONtEbaLWMoldYJENRIiMhA1zaVpe5UShuFv8w/rP2vA6ipBYMpKF
vOFIdmDBeSlVTLxJJcbOIi2PnjDQI9m6CghZ6j3ulBsmnZ+aukMXcD1dMnZfCPvP
vp3vM5AMoimedcYwAMg73KSmG61xd+LHKJC/eTcVO+tod3srC3/V0R8LWbKbKRsD
/VPvTnfep4mjYKeQbTGtmFmWyC4TSSOGkhEmZCt2shyOhiQSPAS8IUcSY4ptGZ2w
OCcYUATXBw4XnNvSdcVuv4kHjAKJ59/0/S3bHRv2sK4hifpKMLfLGHFYXKW5hnBp
UnNTGwk/mDzqeDmD8uBQAti0kX4LdalG9XnLbOP6Q74dFv56jAoizysNsNOAAlRT
WqBXh/Ak+GyttNYVePCf8f5kHAVxuXtyryKrbz4y+a703kBuitjd+kFCC3kFy0D4
IypOhSA6uOOJK2D7AAdnD3xBgpM25Fk0BCvHuOpsoaA/Ef3UyoLQcPOSg9hQyNCD
WCftL0lGwEjIdmkHX4HRS+LpBCzrPNuFMMYMj/ra/TSFdAwfRA/58iTbKp4M0Fn9
yjPu0YA5bN8F7l1036Bd09XOKkabZHSB1fZLfnuiQwjOMIW3BdneZeqsE4SYXueY
pC1Itk84smt84EFh/i+Ocw+f4zJq1ydRtzqsMiBavs8sHZQF3jsv5T1OkG8RzSSu
ZA16xv6XsaSWTN7FwNa3GAPHcCqugyhkrUD+XFctLAIV59PObSscf8NkR+Ruyy2v
tu2z7zUHV8oI0sQ1+VdZ8PmXmDLNKU6zhE/4+lI9uAcOup0QuTZpAW354OhMe2W7
rykfo7x5GEVxvsa5qXqXVSjC5K8YtOiDtuEc7OWVRoOECmepmfIvAYIa2GkIg98/
CjsJsJ17/jqdorEEttwCD14tSaFSC83ZI79fKa7DfqR5E7gZ0nvkMqwBpjK8yCFT
ccx3YruzzGERTU4qYCTA9FOX74kRO8ytWW6x6g+oHdy1PBqfKZeV8Wini3WesCsc
TFLZ/nQtkXbZ2PZdO8T1JUw2nxIbl1Gcj+gzFKf6bf4pciwkf8I5+/Ds/BVsIIJz
pBYeZLPilq2Wy+AsRuwETZormFCD5+Npzev1bQMl2yvMgQwLbR3FPht1vrdpwKrO
yP5GP3k1dVGVUt0aqu4KqTcfFnZ69zefeZsj/VfQ8PgTpGxFG8PPO8jtKR3Sp/N9
jSGBSKXDmJV2/fc6asXRpDqXbP5TjUI0IqbcYoR+0hE5jaVODomU6xo6BDXace6o
yc7qYC5Zqz2GwjgUNhJc05eQyuAC6yu4Lm/ZCVHdlRH5fZC96ycTYNgmRQDqt3Ec
hsZ1lXcXk1TQA9GafdO7a3Q964GZCT8EDdYGuUIvpkaIXQ1npa/fOa2BabHY8jZF
wJJlk14NrrIGvVsnL78nt85T90XFUM/uLhqrg0xUNohsndRCsNyFoOgfKYIDRVpq
paF4a/y+wa1McrtJIgH01Bt/VkfXsUiGKlTzrtoGnRljv4x2m0bJ8aYPJ9cIDUQc
0ghHMkOPupI6XEEdh/nWGNRz2Tiw0prKlESZKQc24ayNL24RcRUr8tsIFTxys11E
FMsVQ1KCqfkcAMMzPi/bbVHkJ57ATVonqAPb6yrTFM08bAnTsWzFHgIxg2uWzXxg
e8InIUBvOQ8s3si4/1QN7MdD5cq/7uNfAyNpbd5q2IuLUg1StpTIdkcJdx8AkOjq
T10j8gzUFaiSYR9+5deB214I9U0dR9QKHx0Ma6OmAmTlSh4+gCKGmnYmUkHvzAJ3
d6jKQE9ul6TQobwHOpzzrh37IhoN+6EMVKr/6bk1vgFDozCszgkC3yY/ClIezIOQ
Mmdb6c00t/sIpD4Ik2MyAqakVujqfLw8eQo+LfuSrOWPzEHIuUezc7aBFHF5g8Ou
WhzaG4Hv4Se2/6rWXLBiJ0NsFi0lRK2J9qrxIdvm5OMPEoLeJM7PmN8ipKj+z4K3
QpWn/nQ94zsCIUQDh37ps/hBjkYVGUMWJ8U01v6wI2fvqsbJIUL2T0sWCUxdcFv0
hfdoZapnXi0rXeV9xygou5SMxT47a0zTmwd6pDDKzIZ5OuB8QiWLUQzXYc00TYxa
+SPlCmtJX1P9L+CMHrq8m75UGhdGMqDlaJGsYIf8l8m+b499qH1LufyZ198sH5h2
3qakFjO1ngnNd8uJzbZt2z4Ckinf2h8SfQ2KTzVjj+H9pnSJv0QhCgmGuoITLVtV
jSkZBOpzUs1cKYyHWLLC0uDndPs/ed/q1txThIjHhse705lpqRdK1VUTZZgqcYqu
x8GrRpRFHeeveIm2nl5bcwHjcgYB0H11buScFqfoLXS1nwJHu5bdbpRtxhXIgOg4
KX8t3/Om2Rc/bGOuzZ7x7tRS+oAGF5R/CxHvrBJA5zq/Fyty3az4Ch6HJm3lsUif
MXOyS/RL8H46TSp7VzTKib1MxPmQEDsb/ijz6pv/GQPGyE7WnBMwXNcT2/063rSZ
nVZbRyrUsKQX/M/Qu4SOSZJyoN0A9dgD1+6ne0KhuwoXTNSQrr9EvvvmB9HGHSPZ
n/ErQuNbYSVUB8zZLCO0FlGpw0FW5yyrliQiT+8DPe4cFIRUJHSDAeASJ6fk6jBv
xL6SNynOY9zNRUy7hu1iyIeA+ZsDUUA1uTDxAWwPAtoBMCQgVNvfmeJHpGNteDyf
InM7spj1tYA+kfyVUQJK8XL7SuKZJvcGa2sGZfYRGm63umS+/xZWS1AtFQnItN/j
ryFiEgoqIgjsahz1R5DFkRAzF3ospXtRs4D64XWu1ylG8YPYQouXrnaMhCYGkXrc
LVBmbXCRM+BPqANW7sP2jogNlayMAIzGt5FGqck9lkz7FyVhonnmOJpHE4+29JJ3
U07/j3Coau0q9IrTIDFWS4DlbgWpTAOrbAEXDy+ifHknDfkro7V8VJFoh2Y3tW0p
6ZLZwfjld85swj/wyogTRFsSaSFcnh+YlKztvjlpLY8K0lmegsvjamahhEaobd9I
nJ0wCILY9dpWMxc8IUof4hYueyU6Xa6LaCIDyW0AD35+nfeI/0urcf3BaSk5FsRN
CQFO93RHNYhNouh92RiMIhq6QRo52b7wSBeRublY1LMUfLrG2GLwNyNBfslwwDnD
aBpS+Konq/o9qdUAO/PzXZ1O07vY6RuWUZtK164Rqu1Aw2l/U+fr97V1dHgpT4k1
P0AwfyFQcvuLex3kmnelMdBiBFxA8YYLUnEBeejy6uFzFOfj+1nwfISbq8Nwn6RZ
dTOkm3ouOuZkCFMINzax5/Lx2SXPEWkzsLUUvTBC8B7AOmj2Cb0CcnJb0jB15jwN
z/sEFlDa36OJD0AXXdL0zFkuyZ279pCHKGaPU6es3QmVYzRjPLW5sJOFvSnraee+
lgYRfr9I5huyNwcVlGHiFBx919RxfAVBjQVFKWCUPnODC8mYunzpG2RfrIciIy1+
zOxUk7aiUdIrHzVPMw+/JrXToYcF96IxDDiqTc3ygl6+eF0yv0T6P1D8CdSG+g2l
9DRWDJDEGrxOaELijYZA7Q5+/2pgw7AXBtCc8tGfWs8ZMTb9oSAi4fyk8h1VTC3F
rTGuYLl7v8pHEo4lty7yJLYcCRgLq1qTpS1rQ1gg2915kmbRUn4yWWrPOpSsLRL1
z9PfD0fgQzkd1loN6QPGUeujpIbgeLRVxK4vsVwnhsD8c5hdRE1GagUZLJtgCkCe
AAm/o8rBUT7+0dfgRrBZOl79SZgbCrT3LycF93rVmJ9asCqRxDK1y9chD7p8lmt9
JIVPfzXXTqh96Pw39KcGVcwVIuZSGRiXWU2iG7fy9ShZeMFITLDVBaJ5MeMpSI3F
Exi4zt6p1lxPVu5g3p1xI1PyFeQ38mBuBWWdBHkWOglWQN7pjZTrmZFOQn9wmEXb
hxwOaDsf4cKUgOs9cRn+DPP0YLxuNfTTYdGpDB3WCckPVqXddT7yB92KJGPu4lsu
bkDGLcWq3UI+ns4QfkVIXUh2yusgxIWroWvan0ATx1iIjXW156yfe4kBorHVQunP
99akUE/4Ey1W7DEMrueOnIBlZObkNtkHwo/ti9XlYB+I+QeNHTBFmYe3eB6pA89D
fimwVkXC5b6/D81kjJbzMfbthCf+VkdaNs9wy8fw9f6H/Y85ASD34kViNhxZjBop
6G+bUcj8DG5quvIZSAYiZoZOPpSrmWB2z2ISTs1fEi1V5IIMoQWorF72VXNBJzrC
FX/kvtAMyBspyUwhgA4yzB6Y6U5swaklmMUkRh+hGDGwaXvicp7kQMnDNJjNydXm
EBkkEearg1YN46HGBKQ80gfZWHvVKJF2wCr1VYm86RLuf7HzyAxG+wNLj5y0zLP6
3n0v2E6MiuZ1tPvf3AE89xEx9bG3FF4pasb7wdAyFLUueelQg6R44ovMuH9phmyO
0BLVcRQ6huE8EPckw+ooap0Y2aplezSeuu6US9HJ39rYLl5fz3g08eEUolBGcgr7
+o09omNaHmJEYrrnZS7dcFgoyd0y9S9dSo7jq2r0jGIZioPhMMKV49Ynjy16T5AT
JyJ//ETojs+W/D/JqDTFzghJL2kDtJu2YY/Z2GWa0H/bRD3lvRBR22jG+P3mWfWX
TCzfPcg9Gp7Lqcuf/QK08EGRoS5WkoPECrzmncfYIwDETW7ErmVLCD50LhvuGvBr
IUSRKRhTySNYaPWAeV9dC+h9JLgpJvqUnpPu7Ttaf6siCBB0CohvfS/tiHyk+G0M
xzCYORRQswFJSQEXGvOnAg5Equ1oBCSl+EYmPNSS83hq1CZJY5gaURVQ9kqgYOMy
JJPrHWxsL6lXTrTr2w6piL+9k0nljt1yHfRI8dVfNvudKI3wVXNE190tJZQr/u13
FsVNnnD1+JYaaLPm7+L9YC4LLfYBvBk+Lon6Ik/K8r+jXELhNTmRMbnULl5jm6us
ElujuQ2NwfRcOx0YyMtrsTIGTjftbMncDG3AZjQziid/JCSMVh19UpEMyzqBpbpp
fSjU7nFDaRywpMmbSbFJbt9QOUGQoZBkf8YduNImK0Z5JPyo64VLRPtxQ5UvMrYw
T0AIM7Q2h0V5D5aR6rI7Q83gCeLfoMMBWwDAc4joG2HgXDfNQk1027Wwqfl+WFGe
t8Tz44d+BN7Jq9UntKOPIYCkt03YNLPyp1TTKmq0hS0ZtBaxn7m/oadH0YXVSrEz
ukPVVFgq0SDQwZqWKos8knIoc2hCe9fPYV8s1NQp20HYwg1+wfijDtKfWKldxQ85
28C1ND1yMLqcJeyI2d4aJmneSpl82x6QMcpxgaQkolp6tnm9euHqRz3qiOHHJ0pK
SMI/eMYEvU4nTf4+zdkmpMx6TN/AdUt8MDV+NJRlA1h5rGNRss5Hj6fUgPHt2C8D
6Pbf9OMW6NiY45W5QwY09XbJn/ynykUZ54gt/kW0CdlIbivWgCWAnoVTsG+Q7rew
yhzSw1hxZ+h6y1aXN8Fpp4DsJQcspbzMMI0v/g34nXPmb9vrAa7aL5wDvqcTrJf6
jIxnqTxuTGawgyIuINioEHWvPBRGOBh3qgzwaL5CbUwzeO+i7Z+f6MTQ/hdmB/D3
9t7nwORAmfdv4rG0vMqebu+As1kqYIJR4NYzbB+S2Hhp7aGm3vJvzroXRo6MCjgQ
cy3+Iu1Wq3Ot314qoekL6FdFrIhYK5bAxX8w/dfjNOvkMCb+2gNaKx/vzv0nDCL0
z9UgFyUZJCd7dqRMKWQh2hwiG0AM//mG9TMZw6JO3hs1N6vUtRPLeJV+Z0D1W+IQ
1Mc3Ib0Ps12MmYKlTe5uDWLMe4CMvUIeg+jCKZHgFKeY9Mkjuw1yO2TifukEoOZU
YFor70A7006DH87/oOEwKBM5cPmWIalSNCSYXlUtY1UEKvX3v1MZ7UmhpV8K8+ld
0o+HBJQjEOyiuKGCx3wY/9gVFa5CAqg6tV5S+l9GbO5O3xNKZb5mOGuiglQwXWMO
yJ0flkkCNxWJ3bMHbHwXYucxyyuKsbu8RMtYvA/B+mvfulXeH0cr3mnrH4FZQzbb
A0NYQ5CBH9P0q6wSdRFd5KFAeMT/B8v5yrUewl8HbmkyKihuJESGl2R4JWlo0SN8
r0s7OKEiOnWI29yfeXJ7YdW0VrZwFgjgp0SIyCet6hSQ/mt2rXc72ncJuLnpwKdf
DVtkOwJnwz/Y9w0jEcFAjE+VGp0CozGl+PxIu4RswTOjwkCmlvlLARkHCsEpBSAn
DXy32e0pYPSNGw6lUdaDdKUSUq+CziXruNOrq0euivO6poB5tkMHYE+0C/pcgPmn
4pWwR9WntplYsla/m2eobemPHDL4QniXVgY7f0sdnmHI8rU6S7CMzMPoNXjXIPk3
0Yifd29Dqx0K2CRAALJEt5ky0wHgZZHL8B34ejScJq8tkf84RIUMKglEuL1liKm8
ZhPLUjTIy5kWlk0jorqhMTChUPvfqnJzT1zsWe9Nq7fwiwCkGL/BoD65ANOSy1OI
7TnZR1WI+rPxbxkPSECOjBkH8HE1EvZzPQpWCZloJBWtiAJ4Edd8Ffs81vXSOAOk
mWHBY6Wep6HOdFqjH3jpPWhFOfjGYq2ecUGanCBJvWFmXq9+WFI0sKtuMc4e4CnH
8ANN58Lr7An8WTW3BPBskPn/BO8n4ZNeS0qJ+njUaNoSEe3rFwNf9BzBvJT9HblJ
XlSiizWMWTrjQZPfoULimeg0h01/d+k2oaPItEmcUnVv+zcfsXhQUUpzbWqtdjdK
mQhUZmM5VB03vRRVS5idIP/R/g07F2kTHI+7iQkRan8XrOOErvH1gjhhBPe3sx5U
4F3MYvXeX/sdkgEzzVUF1zdOtY/reOWFfiyXmhUmGKhdCtAmGG85s9isCKGUTsBz
iKaxUcnATGzQp9Kaak4DCa5W1cCuCzUjRgi8UD/xfKa2KDTXcIQvYvE0WGJfhoc1
7nxSH9cqB4TDZXyJWw1zFKWNpk8GznaGM3Mx34w690z/736dH2TUYddkhquWLTye
XShRYLZFMZf7uquJiEnANIZGBQOKDQnGrKfE1uc+kTRgc6uoKzcdEY7sGonA/G/R
DQLdVi2aNeLJEqotfUQUqWistl3lJavq1Ws89qMafKNOOq2QJ+NeNhn+UIw8N8Kk
MITXXeEkzNMJ5WToD8awHpB/Ji14WDuDMxNoMICvBYbvz9kOnCQgYkwJ0XtZEHDk
llhTVJ/g1vs9znOUlPhECWUOB7b4S1340eQu5RilCJBNE4ttFlNsr7uKBiiFNdaQ
qCNXrfKgcAvquxyIx7b9QXlXZj1x1sTloTbb39Pk5i8wg/OHjB9jj5BHh80UzXW5
3M9v5mEoXCMNUwoaEAFvwVII2s5ovNzdCzHksRtxZr04Yf4b7TsZpVRMuoBu2Tu+
ldY3xlUAc93qBDlP91VNk4WtJSGU9jE+64syB76POMTJp2vz7+tKmCwmNRzio/Nd
ilLDhAaZlfIowK5FihFITjx0gd7A2BjBNhbbXMqu7P8kREEZk68t5b1ZKDXhleq5
nS5OFXomWljrtS54eav9bNOAnwzs4qYncFjgaMQYEcS4RrMi9+IUH13GXThfgF0y
3L2p3YAk6ym8+f6kZAwZ1ARMFRypcHyWqcEcwzzVW7/V5cr5SzWQwnGsHCMUbHrD
xUp4uLkXZYMlqZKAG6KeFlFjgCxII9F7d9gsgXojGGDWYDWEGQZNaMqG/GtSY1vz
fUR0CSX6hF9bZOsfN3pbqEr1r8KBrP74EusXfOqnwnqZEx0IkiFQoTV6I0ZCK83K
CfyW4lO8HtPbS+v7K1+JcogCjn3HAsvScpp2vtrVK2bSJdmQzFnnYtSZ0PvXk68V
vb0PADENE90p219F6h+KHgKkiBPrXYHLZ4pijyW754RTVi2ZziDLdSOU03g/ih1A
uN+eiRV1R8Vq2EHtZZ5hNEnBu0RaJlDeDzENQOGiqIgU9VMKj02jJETzg+Qphqzk
Kw9YT10gGx3LdniPfdsF2MuHSUL9STPEJSV3mmCrjxWi+ZtR/IY8xDrUgX469ucW
B6wbiOR1weHtfOqQpDU/d/ykkxzEjlQ/SvpbLmyiHtuXBUX87ozAFilgz9ycOED5
00lyW6hS9ym4Ec7P9MCmEf8HKH3DpJPWCcNcm8nfDot7baii5ifFB5SGbIckrHZz
Z5g5HXRLDR9csSjhWvXDV7N6eZWBdTo5imcNSetWpol/vGnVRZ/IhxKyq3XXRYeg
qLlIn8kTCDXeFzznNkl6Ja3Wl74zOJ7yQlu3U7Fsuo1cilH71mgFBzAqlH0gGZIx
H1+lgjKsYh+7jpTQ+8DbXMBEDUv4/v6GiPeKBkwSgr00opu1Jo+II/fbsaV3PG68
na6MtN4LEyXbLQ0zNsI64tS6BjQt6GKqpZC4ygBvAPbU0TDxGGhYwE6tHvrbQ7i5
lheh03qTsJRpNPES4NdazzEqfKXX4qjrJTyOAi4K4ougElENolSPppmD1WRxHXJP
5Uc4fVdfkQHuW5CwGhOL7/Ec+dHsIwKWttGyxy/yiQWuhkGCVeJWaWKHXhcfCKoE
qMT46fU3Pu7hVsepPRKGPpuYWoYM4/HxFaDt4gIFWcVMNC3yN02gAFKlFMF8xUO1
Z6/xXW4MZFiC+LFu2A05O/jdSF+b8lnQDyXXq+hK5pUxb+kSDaUYjQeEDw0kjE0B
yyIgso//KYY5K4I6vmQNJWbl60FgVGb/NnRG9LxrAaoa5jILImADM3Dw9kaj00iZ
n+CF0w4b+kF0pPJQWXRbCBsbHnKali3tQRTQl/G8sXENLuc51ha+EOwh1Y9/Ag3t
k2NfG6Dkuy0aXzcVzj2ucrR31/SjxUTl7l5qMV4sKNcIRg82mfOStQSoEOccaKsh
iE3s+JMkZ3naeog93BkNaI7UUZa8JlpIx0YkcyyWyKwt771MVhVSB4lCXksp09aw
ZOn+3JqEiyc+xpz/OzTRDVWM0qsY27yUfVzF1f97INyzTQVGYDEKAtfEGnSO6MDB
uOldJ2WyY9XmkTYvoaer7lBzh3z0z4ELMKMdZcjo11vm4wLCT4nMq7a193yvWwnL
WbKRYRRgW38XTfCutg/jxR21jjNeGFagJq1jd5Mb5dQrqw7aVQccZ5t3EBDlNX+A
REDuTzoYYCoHDN/BP1rMy8UF/9ijZQH+koIG3y7eKAMc+gSWsjRk8CAbrqaa9U6b
/K9aGnvDAoR1h4Pf7fX+nJgaHYMl1BNROIUbPB3RsI331gsicDAIZ4GdBpNgI1BE
wHlaNTGa5ZON/Eu0W4BRA6zhivEI8cvrqcg+pxNW//5fP5CT5/NuE2MrCy9w0GkC
4t6RBB20hlF7EH77bxFdjQZIKGhI56wdyYgqjVxSb3tyfQftntPclcFK0CC6a/Vs
RuIE+/gy6uXxAJHyQUsUE5FqNZZfeU6rRisBmVu07emgFQ1Vksek82qGe7iwOyqi
BMLRhHX4ingPC5wO3lpIWC04I/MhfqIcDQQusTGI9y0gcTcTi10NjlgWSImELznV
ciqU1X30oeHXtJlyhAz4mTEJr9HMujoZfsQ+eqB5lVXXx7OFL2LkrpVz2nlQAwwD
k1oYK9vlA3j3F9uYNbQLyU5COX4Fkoc43u+1HCe/AZYNsiLq1X1DRXYG6Z3Jltx4
LtWDbZWlEH1/VdzuJ6x+HTJOKpq1SN7QP5z78NDL9wBreYvuoF86R1GXIhHPsPDp
sEqiTkPHIv09J/ohFfnevL+487+bisukuaPTA9kNFVhGvsL6b+DFBIxjgNp8GtaL
KFzRP6bEGzBaET1sZulllTVNBZ6pEmUDmL1NpbtVHmGUdsZ7Yf/AliiNf+vCDQXb
yyqFAAl9kLmUM8aZyYUrwmMlPH/V9SglK6+s5XfL0/a7KfWqMzJOVEbO3vm7PrF4
bDg6eg3rDnv3J7J7Srtau+kP7+23L9x8gL7cW46VshGvuE9JR/6BcXmASk67kIOj
nin9SbTKZ+qqIsr5U4YtRYZ0MrrOfocbqbY1xX94YhvrLKrY64yFCl94X0s8lspP
GF37nNrXO7BZJXMa4N7VWmroJ0yd5q9tMon8vrrSDKsVrz4S9eXWtm8idA2ri7yL
YQoZExtagJjJLFmF54IINGw2LSTyJfKN4puZKvr/Pb77qZbjL6o+EA9gCKT2Dn2L
4W/p+YHrgiDxS47ev7AkPp1b3PBeQEr+QCoZPi307YCntk8Jb+g9EQA4yoqsJXUq
JlLs3No26uYbl1sZOFK7WFLODAkBp4WI1IVLMVvogoPUN9pm+4EpM8zkFRZr2JMG
+WZcFL+hSVn6GSM3i0EKGpkMPmHkXfKJLZu0vYGWpTu3sPMJyeac5cvojYT1TOWM
R2uVE2E5RxEJH9ezM/gEk8NSZqxBPzkZ3UusDsfLX/RU5+adyIuj+TLq2X9cSXRP
qZCo2G1c759H5olHIcklYpIeX7K9R0uQdh0yVJX73+7cRadsgzLyUOrbKytc9/Vt
7krvhIFzcHVjsCaIQuAc2NuQ5uOonTjyYihz1zEb2wEDF3QXITW4lGrKAJLaVzjY
UsV7AsO2gFMp/GrFxwnUduCsSCyh42I0wn2dUAmUJE6USsEoB9nPoIgBx1iP9WEv
6Xccn5XTkRDzGo5EjBb2Jwy1/yZWxRILQkg8o/yBw9ne65wDWXWs/P8vB5KSSm6G
vT2meSyKlFb6Fi0Vqa+4izJOWzTZtq6zKHFmOo4NiaGBOvDjpc8EWx3Gi0xfx8RA
qlHlPNwOTBskRQF7MSvpeMEYsYsgM3zniWZTPCPmkjgFvuXNbyqVdW8TN29eH3YH
u0iHjA3C6T6tsBux1fMVs6NC1cn568BFN6iZfo8ySSKhcmmkAZlTdY3szj9oiQKW
iTHEylooe7V4vHN9dCrmvOaNJ5nyLAuwBSpwrCDtvE5gjwNhbrofrA82Oa9DzES9
tuQ/f3WX9aGgeOW1LgoxCqkAVoxW3fNWCirJvoOiL7IDsd+YSw2FtbloMaAJNIOJ
9RXKSJHO951owqIffAu17uC9DjlgxsJQA8LMJYetXNbKFLVsnS/vJX2OB+ya5Jxg
fzyRywK9w4CLbHfTZdJBniKAAKTRZxuBVckz9TEXtUO+5kXGaiW+Atx/1etLtNKe
rYVhTg71jEXkwrEbno4nqmInBoNWx6fT3pLkzck/7QjXV1RppZ3C073ahYtNinqw
QEW7XAzzvr6qL+pGtqH4lxiQiDPDlLlAdDzPfhNU6AoAOjFIRHL3oAnjizRjdVyC
8i6mmM31ed4M7HL9VN9qQHbok0KBL6ZENrqEbTitBcnAa9KKetA7A+/KnZqfYr1t
O5ApmplARLIk7mBQ+7m1DsuyjL8QIdB/veDhIgijVukUv1ukO6Nd7DC76KiUokCB
YtvKGzBQGTIbu6VjVVpLEq77Ge3ULFRMF5AUOrwvjWyJTemisZfL3qBksoEjYO1T
9qluQSXolPlyo4sAmA6ZYIyWlUF8TacZmVNQXREBticdREvq9FiyoPA9rMLG6n0M
nZuP5St6e8Q3yOfFdje1F/ejGgPFi+6+K4oP6/QSYN3RwdN+TOXxw6EKHJCpKwuM
t3OzSqY+/I5bhuRCvpQlmEX3gPW3b/qpzIP2E4DpTS3s77cG6gwc2KkXbFqSxEjF
VhiABXv7VQgxJ/J/h19rE/Hq7kFs12+XhnVV1ZO6wEmWz8QnKAjM5TZ8K12K4lDq
Bfn+GJg5tqhSLKVMrU33USvf7WLmHdg1/be9XbqAli8e4yM6GYlGuQu00S7gTbM0
fjnazCBc6/Tfl1EJ7y6owuZWSHuuOzNU+We10uB7WoY6FbTvGOTN9Jouz4k9UNkh
7NB6HRcyAdBBO/3bjobkDohRKSmlVzyF9RJpo/cWWkBGXCgMNNB4sOhJJr5wPXN6
1L8EaCW8b4SIlbRMKzr62NYtiTqs7FzPybU4LRrGea+LKrzdh20z78/qTL9lnKS4
rukXeI5+oUymOx3Vt7Z47MHTh2J3nHglxe6soYa+VRz1zIjti2qxzlc0XymjEo6+
QQsIaxuYT5FQT1S2RGOH6N16Niii35C1obpHO8CiMf197f3WCiB+sWKeSJ8B1xw4
krjzqXhFASdV3O9xvk1P6oaqK2j7uqrTTuUpmbRobgK0BoVyQhOdEWAYsDWyykqu
iT02xrWL9epL94lDD3rFYVVHl9yVSM4z8LLrmFYsnhkJrhO27RiFZtFWzYkNWb/u
kP2V5+TXPUXGULYORucCxFPqzKt504hx6sC7zEMCMOG9gW53BLkJzRFO49tloJT5
K3IlCbX5lN/v5vRhsnriiRt3wgiBt4JQKf+bWdonzvY+Z6UDNjMjUE3MNAqLb8HJ
ii0I1lSDI38wpG6svN0e7mALzhm+yceNFLutZYX3rcuTZoPsHURNXJPSzODBw+Q+
5zfw/wV6ErZe/Sq4V6RfHcYuTAsA/HgpiCWdV6lrWYea+OYOvFw+1E/wroTBT1CT
aiiWvm76p8qVM4CXATWwibg5B19sCQVheW0VcrCOkJX6nllFr4nM1cPg57h8+AxX
G0N2IfCc8aQtGco44osqhMgQm+PtmifqO/zWT3jtOsy9U6lYXOvLmFGtwlL0vRZt
M/TmZtLE8lIbMPwqjgZSnOblCbUomN4PeVv6nUarMGoIFcVJNCbJaXFUoTaQ7rSg
dA62hs84Rh6RPCCfriyuFWapyEGq360cdPiEKwmG/nMw8YBRoM441LUQRXlm/qrW
3XD90VkChON6vHgVhIp/6kY5R7jYeUgOoXOPib9srbJLQZ1+0yIpqtQZvV7eClEt
P3dXnnG8xGY4q9CXn+hG/XyXCXjygIW32hhpVhxpydMHrhKlPW+m/29n/JKiB8j1
z/YVbsXj0yhasFJi6tXAbyNH7q+oPCk443SQFRZW9e1hqVkAQhH3f1X7SBAfjnHz
5Zpg63Jxpdon82LWaHIy0VenU8y7w5twes97Y/D+QVj/5qFapzDXvMwhrJlyyPZa
0Rsl0uoCIzRou7SAvXz74IA6Bu9dLD5vJfY+g+hyFq175HfVKHQ95zwg7SFqTiX3
SP4iABteNhszwRaYs/blVHnlxK1R0R38WW9aYYht0VuyUparkNZUyKH8aRwHiIEw
gPi683vXvt4ATA7WRZVCS0+XuEqfThQM1RsBQ+brfvqiDOtG4tOVepNsVKcyHfiD
Z/mT33TzvtQtzf8MT8O8PwtIkEqKEAHlRqXXdF0Opu7dU+NGeJtv6Uhd/BCG78no
d5hcHNgrT7uszfgE3WcaHxeevlYEdB8oMAAlkLoKPJqECAFQOdmoPhzgxKgYvbn/
/LEZ9hrMKXZz1NaaIzUOClGxBmVvzh9UbVK4J8cMOjEW4R1bJ4FBaO/PQXnQ7iA7
YeZ+Xic+NSLTUNOCaE1qOKNVYy8BwfbNKzlhus6TEJWhGXKDqpbtsZhjnYGlF7Z1
N4vDhMs4vQ11smos15GkH2xyYhLRa8HJRYGdD4LDSM8CTVpvB3/6VB+f7aZqbSF9
QaU9kPOi7Wc09HvVd3a00FZCqTff9xLErt/ZFUrFSTRICXFjoeDw8zbv6wW+1ATr
dWrJQn4cH3Liq84DcI4VJlh9qcNbUcUBbY8V9Zjv9lJz453AFOQr9BkVS9LWFCj7
H2w6HoUJMdKwKHsbGF0drz5sXlk4z3E+jWMSyMkXhQf5KRj4Rl+QH4vIAQv1iN62
9x2lUjXuGdRwE7t+V9ijBGtXR5Sl50yG3AmI1AMKBUmjI3MhF0LQFnVBERDR6PKK
mVfgD7xrpYdUK5QF5FNGgj6CsZ+qXH7mu09pUeRoLL3cz6kpKTrQFKRkB0bVmHrM
Pp+kuZU6fESTt/mcjX17QyGdWq3ZhMTkqCMZmzr8Q3iQ8c0olwBAfd9Yk1R58e3B
lhgY7gNnT9OLYtexq04cHHraix9HSHm5A5Woat5EUE/AY5IzTH+w7rH8A7Vug9Do
d+QJqsxX80LDOKmmlURH1/aIxiEKfkWZWvKxFWAI/uTvXoyVyPdRL0O31J4hrNGy
l/UgU/4Idnp9kJX3idbujP1ZflfCU3vS4quxEuWXH8I9F2XDKdOT9BCyI9QBS8//
hTmk/P69cv2Ufpl7rf0WsaIH6BlWTe8pUQ9vuUo7ITybsuWq+ma3sSh1ObtO/mO+
0jrHfjpLW0rF4Azjkqfmk3kVtXza5Quy1OenFMbNbQundzFpx9AzMQ9oasPc7iyL
avxe/EbZYJjO1OI/kgCVIeMrurbAzWpOAq71BQE5L4Q+AhzA1ILjD2CMrvT8So8h
pZeHvwucRyg/F7M9i5fEs9DVLYFIRe+PDRL16ddqexZTZyWlCdwjuUn0SpHX3QlM
xUJ59c3UkejMn2jyfOEHYO/0wxt/Nn0fuFX5x1KpL+YahxVjzgUAb1BDScmBeTuo
1esQsvJAtS416OgE9eSpqcwzxp658lVTv+7/zLGa9QasjwOnP3AgdhbQ9r4wQABn
nW9Y2Um6wzFr5jQAEmDDjP9urHwm0xqbSDISI0tlqqg2S1r/F4ZRHQdJ7TYRVlRL
mRbZ5ogGVLmHQhOI/TDtvex0qHzQ9lafaTtAwe7yeazYwfzypg6eA0Ke6NswjWl8
vmZxUxAOiQZiKGmxqA2/MSkukdUNK3w4J2wfX1SRHVL+FMYGiiiR/qZI4AoukiY1
hvd7EeKy2SgiAWi9fyATzh/Ciu6ie/Eb3p9ugHHNcMAyB+KaUHbTHU61memBt9Uw
V+FMnPJtMAr6N2dQf1uBCDzBs2ydXolJd7lDlYYxiJ/YKX0AQXHdocFAW15ZlP5F
9jhW56+121rKe5gtkL9EygoN6BdRlwOzvxnMjOO6Gr2KJ61vjtNWcWESTEz0D7W7
jAppPsGwFTqXf3a/JV0xUkr5k/wZbGbGKfbfB/934Frn0akSdJfZQvPOf/AOOXfd
1S37LHGK6QJWh2NOQSdolW2+Uoxf4z/F1xSNSjwEIag51kqQmphEXTJfAPjyaSKo
hLkZ4A0IqFd0j6eK/v+QtFrOwIKHkgfi2qmeZHpk8Ch2iOZVgrSrHOT6QNWNZcjb
QrGJ9ABPlp7Y4pbKxcYDbFVntKuQP7PAZ8moCOMpuz/EF//JiklR7UXqhXNSFjbt
RZoCCPmwH+112rVJwRWnc1dpYsOD565d+Yti5TbF1ArjEowBvyiyRXzJ5YJ5+bnR
Any9HKBMn1Qbaa4bn2NdtF63poEbVFzrzdMA2BlkZFCr+slmrnqgLLyn0X0cTTG5
nMIC+piskwuoGRtLUTIO2/sZBvPnE3e4/7l2Jkm57CKr46ymblw+kQoCqN0M809m
4DmPwhp3PR9GZhsYV9QiS1eBkmgCQVaMnmCQeuT4UWwkiQblPFbBUrF81vF4C7Am
i10b+2hE96XJDQbGRCHYV8k/2a6C7AuHQJzgfVaEVYND6AnD1kJktnoGE89NdDvp
0TfaMizR3/YMH4UaRMoJqqT85DRTyCXvM64Rnqfh6KYsD1H2YHbrCeXkU8Aa+3g/
+ayEH9gdm3zUW13tMJlU90Sw2QRD+WcNsuYh/llvufwdyD2ajPCXeTS7uBkMsvlq
zK8dLZU6welPzo63cm3Y/hxKOs7sZyp2ud9Uky3C5ZH27MeVmzM+HbitK5C14XPN
oaU6A9rJbLGqzH8+b+OF3g6CxNrKd9NYe/j1RKowORlHJvqHQRl9c5gbtH+FMp5W
t5KR/NO0YaTqtrDgG4f2IEuu7O1IY2c1pxCwFT/mLwQ6mxBgckR8AXAWhSi1RlIP
/fhgf+DT7UV98k75O6VlOl0TElh8occwQROfsF1YFH9VY0K3hzC35PhKu4IsmfQ3
236p8JxqdsrtdBXvFg0s3lHB9C7noc9izcD8wKEExFKzNeZJVoVQLDIPQXc4+xyp
ZsFiItRiclbZex/2FDhq0dDQvitVP+vNCzLxCd+WsWSJzHYY//NOg1mUQm3DJHeg
67Rem3pwCNJ1cXOo/3xnNBzPQZM1hScnhZzJFeZns5IMJFxfZa0pNbrjDbNEF/tQ
/F4sjYCHIRaITSsMoMK5b0Ye5fzhnOcMukg75QjbOd3oDEzWl6jxRZAMgfo8/tii
5I9G8zFQVMMS939r7KXadh1x+uh4XumnrNB46qDB6LMF9/PVMIXQU5NXWNF0gbxz
GpNlGODHlGBJvrH0OsGoYMmE9bLX9Mzu4IKJP841wjXKLVVTjmZg214a0wq5Q5Yf
4L56DqKxr1cz40R3aT004BF59NBhh87HnNWKtJcrDb+BuasymLa6Ba5L+6nI2VyX
kZmY+gQ+HI6klKXlL07hVvrLR/d2ZNhEn3jLjo4QgnFyRiAITu1ZIf2LSjTsrxlN
OjHsN13RkWm3aIa7OvnVQBKPib7FQKdNqRsDUlOJWj8HvPPWBYS4765fQYaPNrF6
zdEVsxc/fB3l57ieVRfI9vw2GLLP1dV9qshhE4ShKa0trL1aGsjnd6LtNzP/XnVB
lvvVZ4K8DiW4OQhWE2BWjlDTrskz57NxaUv8FvF6AZCsktSVc7bLAKtZhRyt3V7d
FObFbIzJ9jdE8S/XjDUBbcD/JgcOKVwD64GfDVFutiU//7ClJFAk1sK7xtlSrWTj
ncJp85oFJIsfyBY4r+qx5ogpXInOqDYb3qQT+AMAGKh2KsLxb/HRZXUtrAw5gyMN
3JWV0jji4MRZ8UBwOJpKfEu5mpsPfzXwsNTFp5rHPytRbxT02xbubQeLvnWvhGeQ
FDEgyj0CjWuYZHyXzc4k+qMsqXDTUKk2z3z5cuS8bm/WCnGu5TDkB8EcKZTSrOqm
5WhE1RUqRNnTcOUbKFRc5MUbOrx88RFvvuud99p8q2l7dnYiHobNHXhysbGVb9q6
XLeJOjbq/BnVLu43JB2Bg1IFkj4gXdSfnMUsElSf16QvonQepxdVl1USXZRW2OoB
ECjcmdO5NU5Ds4yks4wTRUMIS4WRkDAO0/Kz+OY7jU0PgxO0RS3yV4700spLxk7Y
Wk8OLnFIKvDnImXT/aWEiHMEWSBETt1PJ/iyMJbu0PVUx6AESzRyc5V9jOFx95d+
7NlCnT+90oYWpzrCSsf0pKeBE4z80hSqccg3ykYWVib7/UDSR/Pd8fBK4+dyDkI2
CPuk60icy7h7uLJb3HTAwrPyBtNtDlt8lpugM98OPGAEYScSCRuNQgN6vQWSIDqE
nY5YCJuXoYY52OtwyGzqsme22/GPjzGG94ggAcxZ0Pd9jym/p00XCePlHp8gwf75
Ai8DJTWiMCREZRErgMAidwBmfDzIK5lKNH8ez99284tuPAp5unj6hyInSU31Oyr6
cy8rMJErUO64cvdHB/2A2vpZtWQyhte3zloDTrdzSz6J8J7Ravv/kMZHQ/jZc4om
iACsIgXrHsEXpfmIb/42fR+CIoTGgoBCNthkOGmKXB28G2AHQORxj0h9OZq6otA0
WbSa2HI898Pt06w5mjydq+zAi5C5ErN219qoUrCoUGMs7Wd7/9Jfjw7uds4WBM5l
IgQ30ELSiVeIw3IzbubNnYZFkYncF9BD0FOg+W5Kd7LVjG/jID6ygraUpQ1lQMXr
mHydMzqQ9TSkDMJag0EZzQ+naGoVLQomqh0qZSeJ1ZQjWvmAgzd3FyFiTkrUH7dC
5Oc+UJC1gKZDmPN/Lpx+61BeGe7DMO6fxVLjdT7O5UqR480dJQqflWOyC1LvfSM2
tNUx7V12qwswGNn4t+SLs1b+NfhAtXAdFlp1cXkutknpxfnrFMwmFf0e05xbOC0G
SHZArkXOLqAmJo0VGxFEMiNUJQvTxoyWRf7mlyr6HmUwlNo+9sijJZcdPi1utGzE
r0wExT7j2p+QZAlRPIJ+5+z/gr1F6PPyET8zqq6SLfL2VNdIPNxYoDDlK12aIEus
9FlnnuypIsjrokQmDCbiTiQ0Xm3Ge4Jb8zLCqLqomadut+xHTmXByf/QQg9oROWq
LVZYQZNBSLfBJuQsJ+JnebKMjraQ10TFpXxniiB3t3JNa8j1EVMCw1wzKAZ63QUN
zrG4wK1e/JkLZgEI/A75zfqWbfPhqAiQMDsj9wgp1NIBoFg5h9lV7CKGtSrGfRUo
HtNyPK038hA9h2lQ1bZF5LstYKQPD0aad/xYe3MOnVJXl1mrQ/TxKCICGS0EWTAc
/jvokghF2ZRcj+9qkTMRXk4d3/VYm/zADXXwDYUEKo468/ypShTYkpzmL7QEnL08
u+b/ZwE9WrSmerjcb7y5KfuGA/KjcPCCD3hHL6re1V7kM3rVz67RhtM8h9vJvLSg
uB3JdJr7+o6vl4GEpQ8T7M9qoSivnTy+R0SIWakhTUAmDo2PaNtotL3tztZVIIs0
qsEOXphuoU9ZM2NnKqzqJUkf+zyU3MVb4FQ3CfDz2Ul2HqluOG5S92vpKG6I+IPj
I+DnbHzjmjJqNhSxHD9FO/Ez+JIY5mMlHyFTn8M7se9P9AlELKxVhZxtTVj4A7Vf
Y/FewuDzI/dhwVtRDODQ8XFy+TUQYflQ2nUHoO/o3zy8QqnHtuBrotT1tZXDPbwI
3IOfxOz9f+BudtBcqpBwk5+2zb7cNkm8C5WPS3ebY32omyd/5Nb1SbK5sdNesqZL
v0RvfZyQ6cA0E9tPwEaf8pSKw8wv64PKhEbMRCyazmUGZTmb4OYvYl1jPOkQ65S6
IRO5uK/PqUX3u+XlleBrGZIFMu20Q7hbUndxTpTVvHmXqktrgYoGs7hrT1p3AHRT
qBLUeuQH4YvrynaPCuhdwPomLL3ChGIYTpGNIrZ+O/iTViD8CVqnsV3ELWgT4FOy
Ga20K26SUO5NicCQmyMjYiqUsUMWedoAIbz5c8Wj9hCVR/PxquqA4C9kUZmGtd9E
vcKsSsn+M8i3Dev/gxm0JxegRE77A+uQ6MPi5KuyIhxaTYwcn5hXAzByflxfuRDH
SJrdu4Oc+y7gk8nKKNwZTTez7CebHWJEmwbJYPd0K7zorLWmb9b5Qc6vPcvYIvtF
FrmXi8Lgj73lNEEV9VBm4oGBW56amfFY8ox8RMa+DXU/XGtnlcD4d5kML86En34Z
esyoZhiivPkSBl/Fcng7N2z+qqcIUrpmp14xSz2IWADWgZ32RfK3XRguly7GNt7p
fCqf/luQrYbDJfduM8SpnB7+jAJG5WzWWUROeaLE48b20Z6+ODhHUi31CxfBySdx
AlXOyIAnpPMmzOLO+F34/4gIG7AKr6BJGijxg38nJm88oYhQOqzZJEf0G15ddbsp
29NaBbH1rVW0IDGsryzpH71i7dwjetA8gRiSxASa5TH9+wgPhq7f9AhaR/PFmIDf
hK8UwHJl/hBpk+xK0Nif5ROvRaG0/mBJHhKiZ5CP+wLhpw6z47t2M1DJDzE7n0QX
mZRxTcJawmn7COul7/TPckSWtPzsYjKTy5KREUEo19ho2cuPfBNbKdcc1CQMdcNJ
fM5IpULihlcmHO2S7jnZBnLOnBW9IZTowik8MOIzZTpiBAYDEivtHU3JO94HRxwD
ZJrbVfn1rYxYWC5ymL3f7T/MjwY35eDW5HSU30RR3kgcuockMbiKhyLwPO89Ykgm
3srlTJZiBMgELji5yeCkreVQ14rcgqtZmxxDDe1MMUBfb+r+16KXNqiOuoBGnUTl
Pk9uY1zwsounPydmAoJ3iU9G722z3aM8MqHpQCDwGpSK8OjAJNZ0Yx6eTN39qc/S
rB57+5xcf/1qtslGk7dH3x5j6GjIocH75eTKsHirkYTwwXLHZ/qHNxihxjAzzFgb
ablwT5LGsCGs0rpcVyD+uZopNMEgCIwvkBr9n+aStxPJoApnta5UChEnNxQOuqfy
C+4LpaldZRwfZNP9An/ZlRSOd1E8Y1VSnNNdUrHIjrvOywxi0Yo1Sj4khSxU1pKo
6kyks0yfRNKYnDaFR3vN9AMZmoXahtbBdwIQbJMABBZCEiIBKaGUkuJRegfrlObU
IvZsFBpUTqw4saFikODs7Wrk34B7gV0VtRcXGkZrnsMvYtyWNwMscBnYrhSCZv4f
QXquVTgyDFvFwNk1/K0kL2X80IqE690PgWj/FvWva9GOa95/ERgWnhccSjVxJntL
DDl1fnVjQlWMbN1LcBdt22Uq3qJCtSp8Qf1ZfYk9UnDlxSDVn/J96d/v+gn971oX
6ADOQck6mZMZ4CYGN4rFCNh0yBsB+9KPnX8NSxWrhjnupt5UxN3BtpCQLmO4v3rI
gRd4o67EeFHQl3RECbphca2EkkGmOOFGQA+wZseN2UQxk0IJix5C3csU23L585Gb
3rFmzaVwjz5L2B4ayOdknfE01ORCjzxovJa88rEy92sMrXitLUMtO2NvPcgROKG6
6NIuchMApMJ4i3ZReXGk0lU416zuMQAM74YlqUO+Q03FAHO2d4F/AwMSlZH+yLkG
oJ7RaBbb+Ls4teS1Exc86QAXD+SPJGtsOnQ6sL1cepa9bBkjfTYgSuH1VChkV5jt
K2VKmGpjw+S3wgHBxJaRCS5pxzDMfknnNzMG0G1lh7KaoJFhfEOXBgm0kbia867W
gVPDK6CqBfjCWxzyHJJZw9smR2UGYpitV9PnBkKZDyjuj64wVNupUSJ17OLGYT/r
f89RNkoGW1tdkLYM1TcRo8mddyRRhytZ2nVHHeNOCZdiu43ykWInMTOssnBLa4/g
6EiKIzYAqdsZuqYXDTsHOmVbk1nQykl1q2illzaSZ1jIqUqsS4Q1NEODdC9fiiSy
vKekMQCT3nO1NsxOzuUDVk460brLQYr1iefAtjcHST2EvjMESu5wHY9F97ic9swe
UMHfJh4v82HVuCrSsuC6CxpR4IycAfZU0wXKQk6BIfG4dqCGYJcXu7dhaFeb4Fb3
FKACAgs5jMFqWkT3GxKkRuDGE6LRLqWQd7R1nGIEbR1H+uaZAUUo5CR31IZ1/Tit
02YNB5Qj+w79q1rEU/umhkszoBdFzn6VSWtO9LTId5N+CRTcNL38ZQmLp8A/HzVy
RJeXiKoh5ZrVtbjelZZFdV4PvAtF8WbKMaukDqj/hm0EbrgFreoQfLVJ5s3Pyz3g
XzrZ7rI3XkZTsCYqnPk8UkdCyaItv+mX3NdCEPOpxRqBGxgIm/4bzlg+/59yucJ2
YyxMOSZsSZUBjX/hkGadwPdvV5XXnnH+zBUIQ9gf14urN5Q6bv205djEYw2nEF6z
3da/1GXDS6aF3kO+Xrkc/26jx7MOR2+QSaLXsTTIBlznmx+Ws+TfcV12JVoEbO15
yvnwIKvhV1fxCwOFojB1TbRZD7T63S/rsU/h9SQuMTaQcUsuG8I0XOZ1sfocf7m6
ECu4c88l2nbeu9tfGXc+ZjKfvJAf63tWv+A+rEz/VsElbUkPZQNmxo/WJfNmxkW5
j5+BZ4tAdirn6eL90g1fY4g20wG7eUHQOTf96Arqeyn0W/K+7Xiot5KQwMHMtj9X
SE+UqLTFKUBgkQqSa1OOpF7Z0yVaR/Bfr/K5upSUNQTHYQzBCyXpk596Ju1Guhbi
9C9bygOyC7Pk69P+YAliZKUeRbUpeoXqL9PnQpi8hxxn3OZNzl3Ms0aFFK6xpYBu
x3+Q8ajWLNRKmIcF02qJKhOQOb4lbSQ/NEx7qDqXl2U5n6Ik/Y3r/ljmSFJwSNi+
Wehl8eSuix63rWKmpflS7ou+wHSj1zs009QzcREbRWjgmBJfBz16CTgoiy+NV9Vl
J8bgGOPwoRDQSObCeRatehQr48dMBh52J3QIOnwcArXdsw48p00122pQZvtliEFU
2OuR8h8sYIk6J2/DmxwQ9bypTSKWnO/3MvfAIZg7cHCsLJ/oFH/sdhyyuArAQvm6
sAGnzkebUIaQqB7i+Vx8d6tbxQ5KOYDNSMLkTBmcD6Um3jpgnnF6JeQXwYsLEHrV
4B/+ahaRNVtCN4VSNJEh3gpZara/8DPm9d+29nF+JuE/dSetxvHvxPluOkqzCyF4
uDpiRbIyJ+kv+D4gBzMKMeyobCXjUx55siRIDG7eG7oRlyThuN4M22gyWY+gXX8U
jyQxhuUvtUIZGtEI2Cpin66QL/ip8qCZ6HH62hq8oPrt4BQhkiZ1EITq37K+/6yp
OMGI3P5Y6h7vxFlidqs+n4Z1OX8XDFwnSr8j5/JmXDYFZE6yrwzRCjeUi1Dzs9bH
BrywKEN+co6ZsX6Z7H6Gw0jdFT1SNTipi1Yq19Uw7bvMtSj/IMCg1UYgHbkRaFK2
YLJxqVAsjJ6zvCn0T9IlZvjz5cAiyrfjZzidxtlOnAQd5Dg7NJ+4LPzH1+E7GiBa
MGNM3EQxEw1NxrcSJHEDLKMFGMWltuA4KjbIC2LYbEXEwhxuJUkJll9FgFhbOMKV
Xw2AzuC/rDBVxV1gALMwz1HNKKh41ZQhadOPqF0LU++VugnpodTjoEfBQ60oETUD
/l0RfrnOv2AxMcBdDujFFGuHC1DGwMrE8WWy5dTOD/l4dh8ORQyJRqdHl6GBCGPC
oCQjWRo7xcR0wel9KzKkHlz9lzTsw7HxPjI4Bj1R6uTVCH7buU0060WG9kTeE+SG
IiOYdpyC91+7O/j/UnvSFK9MDULywLRNWXeXdXPJA7Zsv9X5BZCVDWcw2df+1dYZ
YmdsBzPiF8Usdh3/dGtg1SKkivlsbhJizm+BLrm2Vqs8YZUUmhW8WVDbsdv88+x3
9bvrlbgGyC7Dx47nFeFsQvs/DCQYMTbIJ/lS9Jh/SYMR559hUByOjrI50pIZw/UM
MOvaUd1d62iwa6tvbjwQgjH4IbKSDj5WgfJ1lyOSHVgbDwuz7Z6XkeUsrbfB5Aqw
OM6FGr93fshCUoRtItNUJ97a8h8D0luIRumrLshR/Lu+YdZZnRcYewPHFiyO5ZF9
1U1ynFiiKkuIT12eIuQRFPLouDYD6AUwxyNfxUNDZVUKNE97WsJmhi3Rr1hEo8DU
KoDYiIPC7cwMavg2ACymKY2LWPpOy7oF80TmO75NUhri/8MEb/e/HqnBe2qxjPtS
nflehDu7kFittB5Qc57/7TKRjoAhAQ1RELKhN4cGyq+EoFDyzFoJwcxfFVw5GBGb
rhxfitbDKC6YeUzDQeaAKowOm+laBhYE4+sKnqnWd/bgfEZBoa1+0jIqBSBotje6
C5BvsSevt38y81ynlHuMhN4UAY/5mZEdVPD9ad0XEyK2DM2Xv5JEo1IYg06d1i8K
eICTfpSeuV4791mnWA4fNOZBKaS8b7McrFuaFj3jP2eBqPDx0aS546CutsBH0Jih
8M//OfZgn76bYGD4R4jfYLHavNkD9Y8OQqrUwgs7BEgfWaiHnYonAfpBxYzqoER0
b/fQ69SrZ9tbLWhJwgdmfcc0+WZsp8/vxHJ/JELKmLQO8IMGZncgpv+LYR2AKBES
LjBiCLvdI2clM0ox8fq2SArX8COtQ4ssqNvaliUEvX48JR1ezN3CtoMel8ExrwZd
ii1rjb6E6WLl3bdAeSNizv4eC9BGD3rslDvfJHHOS/riRdUsVyhitXQo8nDKnvuH
l6K1Wxfxsmu1WfCEviqM0m/v3yF0Uc1pmvMm9hgCE81S+paCrKxP3TqeIYVQA+z9
k7df+ahevZ511jdh5D6cSKGdEzHBpEIsJAiTpyH9JACRbqdSUAddpWspKRwYrmhm
ZrGYI0X08bVX2NXuX3tSDkRP0Rki1GZgU1Lj1xw/pC1URgHfx1d4UaFt//tfOQ3p
CjJht4BzlEAeF3EngUJRntqEFcCVgu2Mq4E56nQr8wRd/zKxVb+bddn+1YnGsXrv
rpJF7boU715/HJJbgCO66XfAE3hnyJL0BwHXuHUAgyjxm8Es/R/DB9aybeaRQoFC
RqO1dmPE+WzQrTuxUa3XmBs+RhO+oSp+ibm+T+n07fu5auzK+CGDfDLfOnFncmV+
qgOGYC9/ssNuwjpoP1MZCyp4fYQWYp210c2p7yiDv4Fz4yn3/6ZeqHinoiYsQLc2
yfSldyTeFLhUmOCuXWzolRAWO5n/+Bjqx3qgSXj4L1+PVm8EoyncRrR6U78hFdhw
6zmJcbVvB7N78hwrSUF0UB2Vu9rj2PgEcPC16vdP+HpZZQg1psozVmW8SQAxVxfF
HqLFpxXQtxGntBjL/zh4zqc1o6WoyPuki0HlWp0KRRLTsCG/cWGrWyCAOCsrvrL5
OA23HrIkJYsGcDqkDwPYCpzDgNt4pedrtQyKrOBmcofilhhvdXDH4vCaQuSSInaC
d0lg2W5dDRuNijxn3gWsCqn+MlAffyOR4kPC1iPPVPvxTUzfQk+MBzxgJ4NAbJiO
GrrHT2JTZenVH6xnrML9T2/gpdyTwUNylf9gPdim8oktdxdJQpqW1UOV3HrlWj49
3NqCTgvJ9xvuJ8x6pCDdDto6CbMvdIQuOXGXhpQmxmYINBKc5O+yegriKyNT2O9X
srwYeWTqhwcrFmU6Achy+55HItDwVK09D8NGDsbKKv/hz0Pe2jX3ueX1s1qDJzo0
pvkRPewYK0BtpErJv3Jl4ZHefJzJ76YexmvXL0yLpvSr4J4PHQku8aH7X0sEEHor
osK4zM/c2wyMqSKmsoIVW/dfIkPi4D/VfZ726q0s9MRl1yCgwzixqZrLKzsrbCc9
UhCdrnVhJxomMYjS7LyG8yeLRmADSuMadkHo7eknr94YAQaTMFnmGA+Dqeou8PwC
mMz3Tz4boFdLbat0uVVI6A1p0ZChKCP688jeBnV2Ds7iMk0yTNltWSo9Vw7mMKJ5
EFdW4b/gYw4WCRFqOqkJsMe7IvTb9nx6CfVuonBaK6jjGFq8h76q4qC9b8PDrvEV
YJOujId+eAMndfKJR0R1UeFLgFfr6PiLXJod2NDqflpMqsNY5Pb6kur4nDA/QJGX
gGsQEgMfNP0cjeEglHIvCBbzyipNHeufG3RbbmYKsAnPfkIYiRIWvAQgar7VVOgX
vRcsPMD3nn9pHtmXXwjZDWwcFZPa5O5LxaO4WG6Rux83wkWYRhh1phgNz12THt5q
++qZXmsuPxfhCNBTf7POig/W3Kjeq0GfIeqSj9oMvXAuH8+VOQLWG72BeXaKwrNj
syUueiDMkCr35HruN6Uu51AOnVkAkya+NxM71ZyoQPdEbp5jELggBNW0X9WuXtt7
b3gpU7pARaXzJYnnNKLpdxXj5Mx2IjpwCHH+NSe2KjWSulgd7Dy+LVlUke/L/jdu
p4PYMP6bJHlOZ2zPzjn8MkH/4m1YyTpBh9XpipVmsaYW8Mf4WdPw5/Qh4QrgNVnm
bvcbcyjM/8G2bQlCIGA3Lj3qvs3g36ackba10/fLWDxBB4a4y2uIbETY8f+g9Q+5
SbZHEzNAK7JmudUSPnEC3hjHz+Qond00SNvZpXdhsQSHpCioOsPBsyjiYhFbpkYP
82h28MIJED+XcF6YLCPaWaF/yt8NJBY+TYkSfD270Z4YW7oVz8KXhDclvkctZ4eT
/spT4NIfh+hoNCCqK1KeUK5p5A1CB77qVhuNUSgcT2VhW1rE8t6OnDFpT9XSUycj
vjcsf2PEz7qxJilUszMqMhcQrIWA3lIIpRcwWXX29eoEmCcHP8Xoh8AOm5ZqP2SL
8k3CSDUG3rqm9dMSNFXfhg0hVAEBSIpZgOe5Wy6fIMd3gcusMU6cs2+Ik0xBhrpC
JJu4IdCvLNYJqeCJpG8rx3yL80YnmvcmucSgNILIZV1ij+oDvWNbfJTmYPO/XKxT
WO7RdSHJTOxkhFqE6HdekMRphISO2Laqa0saz3RpIja9E6/907KW8h0AUcfCAImN
djbnxhGiQYZBSIpE5AcCy3uQncdd/S18A9lMy1rVJvWSw8iIlXM3cCpj/fF64dou
+0rNqpNjtqNulIALYJN4y66WluYtALf0EyGPhhqMK8WL6t1ka2uQwVQK5SFT3WzC
fhC7pMc8WXgnXYT/e1GXgc3zQ6KGNyYEmpPqHH7N/lhcwofRb/amjcDFlgzd98Vn
SrwB0WUL9kowxQrb4kQJqbWgrkvpt+iL4v8mWxyY43aAgMKasehHa8xOo4V2Mdz3
hMrtUvMXxP7ZojbvoSd//nNDps52xhGlCTNxNZuxvHoevLPkZsUIvPTd/SSK2o0r
N3YDpwEa8nEWy587f7JZOH2cJjavS33RKuGeLwsVh7QoV+ps1E4M9sUllNr7Q5Ya
6Iu2aRj/xkQ+qsCptfRRBf/dLzNxOdgWC3ewN1qVnALuiGLU5Oy61qz6Tn/Q1sYL
Mve4Ssald+DdpgcARyNFJOIR2tDaCHBgvT8NvAHqD9CcEh+uvL8MAbKOQwGv3lq/
5RIZFNiwzYb5lJEI9sVcEthd6M6mE0LATTR0NNrAYNDsLAS9yxsRVLD/RcX12OVo
EfkVHkbJH9rFyazxF4a6R0AjRVOEzIRPk1jGnYz7XhswORMXM6/GHjRek172SttU
2yNzAleTAPo05Uv8RXe9jjrtKKzldOBm5Z1rl4nAGW6ddyMXafyhKPiI3Bwq+jg+
nV4gYk5Yq8cn6fZ5xgHt7KNQIqS061hT5wjhGLWO3tEqpzKCJXS0i9ZeFCaCVabc
RAxtJtQtWs3QUxMb3bd3xg4oROiS/ax0TbNLQ4+WhhBsMoGyucvdYQ70O18Sxjel
68/Ts3ztwMxzjyP+sPGZVIjhSp0IL3J751DFvPqVRUvxOgXbKzBcXbNasdAtrauH
ph9bln8CP8PxOrDaASRUkUa/qS0GPjJa63fMUfDrx1v/Ch/aIYtr5k7RUwLidH21
H6lEvP6u7c30aTRxypyMLyJuXWn+x+33w/qtS4+PEVGlIUbbY167U6WbvOQCtiOr
CUGdq6qDAvith8eTMeI79hdn+iKOqL1UMkfZV4lEvcLYttxzuMXK5CmssY9P1A3a
Ltx5YhcYKd9oCYnxWErzfVT+bLuTX9unCWapIUAjeLOy8GUZLa1JVPvnbs1oLxnQ
MJGt86i87yAb6yFEWmDbGMBhDCODXH7LoN/ltwD59kk/NK5VABVzoPfi2p9Sd9LC
nvWS7YfTyBlxsyuy140Po1siUKlmU1L+eQZ2PSkUxXroLYOH3O+UrbBEB18ET+7s
ENCEF9AyI1lUKRC/JY6r7Sy2CbOyXzZv5tpb6xmvVNbHRRvx7YYWByQNDH6Z224Y
Nv7XzyxiWi6Ap+oejf5kSO3Hh7L2d/Sz7FK3Fsmsu5CC+QpgXjA8Clo0SecnMwQa
9DNYx3bYItHXbJDUQdoTi6mXx2b+8RLEz60inTCMfRzRX+Nx2kft7NEgqDC+BUR5
oaC6CCizuAPUzDQ0G6nOB3YP2s7ZxgeYopSAxBZWg/4CugqX0Dj2vATRhVtdaM5y
2DQbhpWFsSk0gC/is6umbrLQKxEi2tvb05EcGi4cj8bxIWUB5FJipsinYsTjx7BI
84Hnjk/4U3DLABbLUbZjjdRsXggMncjWW+ldJsrylwp/Ih0QXqy6gi4xMcHcq77d
lhxqOS/hnQFMC7ScIQT74NzUH5z16hCq3QTXEk+03Znv2ZPHOF2Vpv4Um/MJuBeD
weDbqXw5QIPAxfnpTz0quI+H0vjQRzoLXIvpfc17qO6ZMLbV+ym5mR3PZwBrAtuT
q3hLNDWeXmLUo3b8psyQ/4hSEPe/5CdrjNKonFCtboTpGd/OXRDCdy9aBD+MZ9Dj
rKE2Hfjljne9fRNPL6nmgf127hQR+R5FvzmgRa4Gq3H4TQ3uE9zPXgxw+qLBRejJ
GPJB58jsYgiAExaUIgPbfnWgAOIM85wKCuav9xZcYj/YzqDWE+8RSrPocG2UcFlx
dBikwvYxOltaYgjW/7Qxgb4Qm6gM6vXi0KUkvD1y8NDK0uBqSssp7O6DOUWbhCZ4
StwlMjiHfVXQ+2rmkZeSq/rJVwtbkrqTdm9tBzTe/rRhCmTEhTkV6zHdOEie1SbP
yDn40yFnMVyEjTt9OD/KUaoT6D92q7EBgTuJrowUftBxPnhsfO16OJsZN/9SgmS5
7HQc9xL7LVcMCHUTREFKtKfKLSX3BEPy98r1pydYH2uBSPw8+jdtn3TXRi1Q/Ux7
+ksTvcYf269vQ24zf8VftVKpoIHyNdqpv/jfWX+ybg/JBZQgTRWt/SCEH7f7JolG
D01KbA78Z9+utIEcatSGXBQuz0jjkvf+Uv5nlboahylw7aLK9JTj/hwjWXl7D5Jz
+28nfVqnl6Z0B2ea6tQ1s+P6d7RVzZii/8xLHROg9hpJ26UJgrInbvkJ7ZkvFnpQ
gxYT3g40d1fKrr1cM/ioTwFcPut/z5pHsv+ohXBmUROlc0Y9t8/4zc4qLqcoUaGv
7s9Tm75Hxxo/snvsc6Zw+FFDTmyevRnwGoQbCvPKKFBkp0oYBzVTIM0Qhh3b9Hbi
+BIWMxm+ae8mxySFvKobLtdrfGwLjNAszI9DCEgBZ2vpPrB1kVj+4IuZqXqSj+RZ
g4tovPq1UitgmT8zNSE3S9ns+RMPyJKN9rgH7J7+JULYXeFEdMx1kuJpEeh/mxC2
DQZnfVXZ3PKa51TZgcCZYCaxu7S5qKN2Nr+Ua7XSn4ltC7gwOKchA8L0DKzjsInC
EEY/t2sJDrc90lpntZuHsg108Ij1C9RxEqY8t+hKZijyV7drmOnwH/UhpepZybnV
9c7OHodsm0C5cEc8T3o0seJMKf8VuGuC3NQUpNsHm0rnJWTFM8J1IPGxl0t5g0tH
XlmlVYTu9/2KbTi6qjX0w4dGiVerIPq/eQOC+BpaSp9cwFj7himHMSNoaow2Gka2
u88dYWGJ85JFJKgptyYq68xqXSPOPTOeVAeSf13RZfkAC49T+TxW2O1xCHGPwgh1
Lxj2SbO8jX8PUAuUtnUD2UclSAGDnyfKgsgQnLfQd4xlJ2pr4xnymu6wFy0jK7IH
uMnXiYqi+hj5tHRbm5wjvMzihFmNGonxkXoo/sbQIVlECYAuvplGWaG/qnHTWVEl
Lt/9KymKOJm62irvsEhJxqrkudAoNE+ONB8ZAgbGX3L0l/ZmATudKD0IXH56w3Na
bX5DxVvGtVO5Ub3HXpJwjZub/XkyjYBq+EbG7KOlbPYAVHRK/KoWip2h/SOSnCtx
ku4GX3tOUl3+KuXyeTAJFPh8elaFeR+VMtXEPnRTiBKtM8gCmR5665pVnqR6RVKZ
bNwhRGXnfs789c/Dij6cTch5NXO0x9n/AefiBqLqwTIeldqZMsfht+nwgLqT1d9C
0eaueIC9+7Gns1Hc+DAsDLAQYYHUKF1I4erQU9GdsYf0qZxqlx0eCxuTTXbp3T6T
+xrYGqLPYPUX9YIbKx7zcTYsxnzJ0yQN6OzKn7/wAb13LZ/M2cF7XVtSQCkjs7mk
sCjoIQ61svkz2dZ6i7Y8BajlioCfEYS6MZ9rBDQ7TMwKoiLCi/UKr24EnHxBvRuk
/3kOWutcGG61cHeNcANiipmZZhJKQtYs5gSlCXOs0F4PsnLiUN5oNGfYF2IoTeZe
H+hvv+5rRxRxju8d6iUPOyrnaism1FzYKm9MdBLXAskL3yYRBD0ErgoXcvpB0vYg
A9QsXQzjdabeSom4fCHSJcUHD4Uvwrv0kmfORue6whUMD4l/SNETWrvDKB1Crxx3
lh3rrDygvoPPfYAYoG8sEeXT2Gp5MqZ/QgGSmZywnUjTWYsZGUfg/hucnLu9LL11
N9xEtAHd764G0GWGfuf+HilY8jaONOEr3Ni/XffA3QKRFDUdGI5QXgguLgpJp6o+
I9PV98P9EBYUtWwD/hMX8gBQRbyCrKROmREYUixdtsfYw7rZ0H9mJLlV3I+btwfW
1CF5DPa2DaAlt4dmt5EU+Jl5x61SHIZpyRjVXKSQfYVEKFO/4oDlK67g0YQ+zpZo
YZya/m28hrro/EmNovPsrQiEvE6EcqUY6T1jgCGpLwK5gpMepQ8gGx/o7VUAHc4I
FPyS3WBl/QDDM/aG3Oo1G3AdIO+xf8ltfjSbZDe1iMTwD1IdcUS/YcxwddrlJZz0
BwDmLarBcwOJ/26bzoE8lAvcL5xZMzpJ9Ewf0QxkKx+2vGV92+mUCpzaF4dbh7gV
8oQ1HJbG5FzHNTQUcPzSrbJQjXQrbWQz5zzttKrkRxLocLINmFLrdmiW1fOWxniq
g+CZoyQAssoD6ab9VLiGnBX9jzHB9hxKLUMCb1+wIvN6VNn9cm972BSAE+NMWhxg
APQ5zTtyZUf32zYueWtExd/jA5C0LFKeJ0ckYulmuh0NgKmQxKM+1d4W+BUDsvJh
QwlJ1mxwF6dK+sOuefaIR5/srv3h6Euyx2kDBTynTmz0jQPGpdmjUuzIUEC5+VUa
qcTCVFPCkRUr8T2I0Yn4rXqrNadZ+VwxdmEM8dV+z8ecjUBxyEAEoefD54XYZmDe
aNS4sScQD3NnTfKDSrtgk/cqesaOmqgc7T4/JrDOulU52FU1TqHbuF2JYzwLnLFv
fI/C3yjQeHjYfGUvnlHVOhiT1K4jFnwiTYx9AQev7n0owPoDj2xE5xH2M3lmpLXN
AT626tSWZn35jEvsnROunuhdvR2AWxLtae8HhawiYJ9gEnaJiTJofth5gYDTVbiA
TXIViraMd48o4s5CNzqnh9VSRxUpzSFW78BkNhElChvoXZv7XwluAaLLBOaA73Qr
MDFdJ84LJqepe7FcaqyDcfStPHAVcNzOJ8vS+W5+spFBqTcUn8TtV9jqwxanIpP3
ci7u8k2igvsbsA6o5F1J9vRVrkeTxLJfcjAcgCEoLu/hqBKV4PI1SYG14iTEc7vT
n0W6v/z5rNQMyMvl6+irflZhLysXKszsKIYctPOo9U9cFFVwL/XHl4S9suHyDfR8
tA/2ktDs6IFBdYiDVdL2Y1vBUqTAMwLtllHYxB7lMNsz7+gLBFtPJxGSnJq7wvR0
c0lEDCNHUyYUIaEG6NPTT/VtYX+C9ZDpOSOW3hpWxEDTTKcDmuycMxya+kZhrAyU
lrLzTWzrvOq/vnTotaX1kL2Ooc5gXfLZ+JVX19qm+TxrefU4IP2YkdiDptKEkvHE
Jtll0ofNTbtxJ3/pW7t1Q0XNdhHI6RoHDDafn4TbloDFHsq0JIlvMz9AsF/EWQMV
qxOUAiMgjJ7AQGOu6Hzeyy1t3kWXBxNUN6+4ZPqCnbX+EsS5rmPdQOx75SbgPfKl
uiuqSJ3xo/M0jKwkvSdOlmHuKB266jL1RjK3bca/nEn5al7BIkeSjU89d3qBqE4h
uTYZV0wxaMZUsdlTBue+HJb9l02nBJIondOLAp4XM+jJZxsBkNT7MF8cNtmqzp8O
DAxN/oGsAKi3wZnG3bmn87wuHqrvqPrbDKEptzQlbDHfSpUd5ygN3tPmy+YRz2AC
oyI5O19Z7B8UINX/jNIr8mE1GJQ/lxpeQDPf3PxHTUOK4oc6aKwkrpE3hav9tel9
1NcJwJoFNFdOndUqD4Mz/JwGeIXGMJWu/CG7+m7L7BsbFrHduUg4tiT5BGC41UgT
+jYCY7Uec50RZhFZpxhf9Wk9FepobfilPZwZ0NeqX06aIxSd8IxONREZmgcXUTXg
5NzLC1Hak7O7fdmZIM4ay39Lin75w9iSMVO/l/eVRqzaAwCn2e5wIpuMA0h0M8md
w48fTD7huekYhEQIoi4C1GHGFMRbL7BOsq4gF4D+zJ/GsgKbrbk5axqwKETmG/X2
K9mRPhWk1Ev/4OnTZJE/w4W5Ci14dpb9vh6hg9G8bOtPrn61J+TWEXDjxWeONxZT
kDZHh6AniohS+7F/6TvlpWWcxdqdjhH0SAZb9zHb2MsaRQY6N9JYl86gr3I+nmyr
vIjazy+tesaIcflwICdUmfgEkeVPUgjx3+OT8lQrc1Ngh1FB+AmInXs3/QAp+Dll
mUYAqx5NkPgK6weq0TCtICJSeEPrtPRAAdWy52wddHePv03glI/hrWkbKHqTg+Tj
YpLllOSjfujxJuS2ETG/ccOVzDLgpoR/UoR3SPuuStwMxqXghcJAqypX8Xv8DYhd
6YLTr1i7k8moHH/7GflVecTa/94bhTeigTdXiD3STw9ofPujJGkbQdFdwtGsEA2n
2YGTzO267R+axMDE7CgXZyhMDsWCpC9CSquL4R445OWc9PNU3sCMI/2Wg6pSi3w1
tQdY230TN7u/aNQ/LsO9YtG2IwV6G69j9Vcj3aMYMWE+NNmEPdjI9x8ZfKzP4O01
0aP6dDt9CRikULDhPmee16SxvUlzhlpb3VVLAElo6m+u1Q7IRHa8PD38vtTTZtzL
wJ5VGiEU9aqcZCtFARc72ZAzCTq39OPF5YRk8rfP4MaqesNSDAp/6FTXny63nuN/
OfEeDEsYaxd//bAfPumrpl/IkU1JF9TnGVFpRa0LBxS82EAeCpuN7dGpXPjTTg+p
/FTYfFq/wV2RXZQFma3ouFTORfNsFzZT177v+xX7i7txpuvX9xGWEzr1tve7lBQO
OCYW6gfygrNwR2r+8VnoWLYG4MyqUlwtOg60oufDpG9h2S4n8RFu+UQ2h9byfW5V
aOq6jhplwOicAg+MkvlQ4z4k/Mr5ZgpzFJ0O7W5XDJgWmqfw+SoOGmGTbNSL0lcN
JzDK9r6ysESYI5VTSjFeOTQyc2uSQF2AebZtBiAadaLXY3sZBDFXuHedgDgf2kvL
beUMPApUoeKlNf73Vzwg3ScMAwyUELFLkSDSAKMwAqzKM9XJz66g0lPc341FEheT
EA5l/VyVTf6K5YegcciU//W9AsWbpGGY8Yvby2YSyrq3eu/WAFT+c3y1gC9nsoLV
OoirJkLUNGHqHj7PLNxkR2qwUYxDtOrd52WG8MZdfd0FAwmzkjFSVr+9iPmCEySI
oYVgjpqL/YJCctoW7NDC8qlL3eVjtDnFClfbbYv9/h1QwFl7+sdpZIMDfzaKx96W
ttjkioBLBm0uvQgsr/F4uOzZkkCOmVcNKFTVLS7k5oxeNxsLNZptYOhQ7IlrwibP
UFPPBhJ+SzrWRcwmSfHLFgWupqvpXsYUu7/v7xox42ZDRF9t5xs6cPc6txTNoX1O
oLE97ve1OCfl/VtfdZOD9jFfhL3sNquspxTwtIWduN39pSK4boHNQeHQeIFX183O
0TBKSS5/prEzt9hSzrKCwhYjDQTDpPW18LHrv1+1SSYZINOOvaKP+Jj9mnrRxxok
RnGbEm2WjB5kqe/MVnkDMFs5dXXY71kImVpIaxBxLUlbLtn1LrWw7VKtTMecAV4W
A6PMJe4H1D1rH7I159llQg6ryEp8T5GA7AAQ7BveHCQyNIVYiRoEWlawMv345Y+I
V64FTs/G9+PZPyuzCaS1pz6pA5fWwLKr8n8s+d2vZhVqX9Au6wo/ipe2gjVpIsOX
nuCMDhFoADZULBdYQjzDOyYUujuQrz0HR/XHKkJ8p25lxM2kDlXDFPEjiJZxH2zM
+XJ3Mnf7Gj4V6Px/hHIY+zhDBBEs8DeavkWMQTcB9312nOVGT4eY9Q2iJ2KMVkzD
FDgl3Tmy3O6Mc5LoXw9c5deeedYQHSp9et4kwBmn4TIBRh6n0JD9pi36ZTk8U+Wh
1FnlKFawxFufxa0B3ZPCsw7RMdnA5GP11mNoJBHwLj9OdltvnCxytihXuAxwY83A
S9XtmKxstNXXzl7CJPl/VELNpzspuQDn6HG9G12PS6LFQWP4mFPGJqHDWrkQ2A1Y
iBlKvFwnAGsdbgN6C99jaeAD710nVzYbx4cxasQPkcSI4pE3h8dSTVH2woeE0o/0
DDllV39Cr+zhZX68T7J67lp3n/vDbvp0/WNDIM4LP9zkenABGTSPLxNnolHPWdii
ybm1zzgzBCzWd52qQTr+368+kpC2qBZVdd+x6h7LDjEHAkcJS1d+5w2y3Mlpx41T
W9EJMD4QIzgIP3T/NfI6LWy6jEu0LFRybUxOObVi09LINVEOfp3yd3TfWNSysfvj
9WiE7NTMqhj8is83hAEabaZi3kY6zrYb54ElY14sCvydZKT+dBiLRlMpEnNR+Hpu
bvKW1/DW1YenuNHTSf6BZ+OmmyGQ5k9Pm9oOCAa1xAjmRyU6if8gRHjmzBCOoIfB
bV7k4e1spO1ge+yu/jdwgWHnJnlt6ZZ1M3RK2pNjkg+ltJwhdbvUh2eNIf9hN/1o
VmaEt6bLtuhTWcRYzBXb8SLTOh/i2fK2zq9M9sKyROmrz6op/QsxgJ0aDZw7aVxV
GB+RNVVnVpmFLyqbB7jm2BwHyVFGdag40OS5nE7u3DzGTBIbtNa11kuMJPVyo9CS
qHua8sP6FoPF57oT/KC1VSIESIIjUeQQaHl5paxFYAod6Q2v63VuI6U6AtXtnmSx
1fpITzNZTPtxZJbJzkr8pYtpctIHn7lfQh+uHDYdreOEQMQUJNSO/xWlrIWwg8nQ
QKEiR9YmCtf8Kb/pBCD4+Znw5NeFeJgXeAAiUvI1WTDa+o1hBInb9tN7V047xIwL
wC2bFYPxTe77QDhMWyiM+aTChovjYf40qn7QUgj/wRXaaJl3kkt7A3b2vs8Ez8/V
xqPLPMIsfw6+P8fdyFdmqTFUxGMZNOT0nPK+lHOo+Xq51v0LX4wqXoGVgUvK17NK
JoOCY3bcmTk26lmg5+TI6rDO5EYKzOp5yPTFTgQhtQrZu7HE9lTQBfYJncX8DcgL
Yco5vCqtnN5ReEmcVm5cgoFvGjOS8d2DO/Tpr+PrM+ND/d2fHe70eFBVFm5Qi/yw
jIfLlhDbTC/M7cwRIOADfaU8PxRArlvE0dY2oWt6XfIRULr4agyl7XGg8I6LPPsz
eg6TFqqeNPhjkkeLmFiJwn9nFMAIynNjczqplUXsKQ2mNwPzKHDtJx9v4U6SA4JO
56/p4vDU6D+8IHDJe686fDvzygO9XvK33Xl+5PWY23CHLM+CzuXdIFmV1JNozjpD
wN5N7A6FpAQNDHy0c+PP+zjFMqEozd1eOL2bmjhgL82alI4PhrXom8k/1LidySFl
7Ner55aarWngPDjbw+Ujjq+GRSZ0NwCBBonD4Y5Yhthaacoi3iwb/cs1FJtqcYLt
MW+Lu0jEjerq+sAbj1RnxQMW2xfa4sQMgued0rFI3yVCUB1jotAyJfcqhMGFtYqA
hc2ckwOrxkdHaiMTlb1lAI5w0ylafgjHPHvi1HQpngZ8C2pnCTEGiePaZ180vyEu
ZshZi0kXwkYIRZNNI9uDUeVgg+tBl8/ej95jMnydSXZiAG1W9pRktWbw8qln42sX
A3lja3rvNFG6pK2vIeqYKGZagboVoFhU+XIwn6hEyk9U+BiVApfBilI7EZLwP65n
oUHruDOeeLbN9bQNxCD7P4RIPqSzx4XB+N5aNRXt5Ttr1A+PQILXqD0g+hug+CK4
v6UjMVp/8yUE4SWMKa9F7MF5FbZK79vo6Lba3crs2Zr3Qrvif2E0UMJxr0CM/gMl
x6/XxFXdy0uVABRnO4jGRJUSnqa+2YWLsvhAQxkIOm478YpfuDJPS9J3QYdD3lDG
0+icvXg/Z/GfkH1Tn9WfA/sjHzjGo4NeyieKO2XtaiEVPk5wPGXNJOgJVZjLc9HC
ToEWHGF/p2i0DfszroDAn4Mqud2fl3/fle3LTfwNxhMpNa9XYmFanS7a5USGeY27
ub2C9Ig2tarJfwgBYVZWq9loi2l9Ny8Dg5emEwrVCJc6JHAnz/MdDCC7ki9lK8Dc
/lp66Vi1oh2jhSCqIM3YKaUtgGi7RWoKkuAw6dmtNCjahXXCOuEsNmcxgcrvxZ0h
2QwVkg3z7uS8rqY/++pdtF9wahOB8ngWbAFpzkS/ZatkMxhLhnD1goOHa2ETrY0q
fmPjs0etlrQ7JT0whL1BYz/PdAmuH02ut8HZ+D8ACzds6taqtwI96YRVobEeUcYF
zMdKEluyOttoCHKncJdkDSVMl25VtBkrv3O5K40NcEvy+TRRpoSfVph2tYrg97SR
Qau64uVr5HLpMimWdokrmtOdrdybofcMpE9Z+Au1sB2m3JcZbcCeJw6DxiO9tK/5
6z5IoQx4QzmBdiQZlRpgrtbIvjkLDco2wmfpiaF0kO146t3vW3VaF8h6648t4GbJ
0x4te/NLWzl8HpNrHf4WUqHPmXUBxQbTjowI7kap+VWPmGnpRKLdQFd2AmMdcmbf
DuFuaWenJh/PoC+MJuBrW5QsjhuGIwfZR2jY0xQRb9k4BgEBtY/Ys60DPBhWFXMI
U+nVkucz01rEu5hSGY8VJspg22o3vb0GnE0CX22yh+G6rOJZfjmtLqEzv41tGgkC
DmTQuzQer1hdMoH19gn65h6d9hfJIb7EcjX2VbHUfDQUo5bN8RPWamTwaY7CeXON
MLkgiL75PEpvQT+quhiicgTcHm9SMG9FVVrE4qSAFpnfBLsytUhV0mi9SLnmdMaS
OiItR3PeyzOBaJgfokKY+VTetF7T2dQFHpCdzpeEhsazp97lfIjD9CeVR4Jz15HT
rRmTqUzVaLFVYwCfdXEZ84Dy6uWJRdSSs8jh+EYmn8vN5md3RuyD0oxICFONhS+7
UryxkkbZgeVd2IIr11di5L9VVhzgyf1U/pEDp8YBYK4wghHbz6AE5SD0zPbG0Xs7
KvAoYa8m3Sf5NBavx5KYWhg2xOZZyugYrx2/F7IIE4sGyUguLFNjiEfH/0R1yhdx
2vt1uJGjIVioP/96x5moO7PALDxgmlP+4EkEVJAd26ZcM4yZ6SZRxkgAHeWfnZ6H
PS6r7Qh1Pe3feop/qVV8fk8r2R5qW7V6LmifMWcLp+/q/wf9mHLSYuRpLyYveKxW
XooSGudLraTpPlMHIsP3gDtrnbYloJs+xpdGDo2B93zvUj0QSFyWOBFgUa6WIoqo
HEqgPHdCaQdxyg5pkyB2iHBGXopfzgYwHR+ipWEcDWQ+YDTaWEmNB+8aAbrC7j37
g/MnhbBx9cQ1P4uB60i9gVHpNTJ2YAnOdnuMzCjHBkZWUse2Nze47Qk7F8iQNpt0
XodduZAE/xwHtePiZcLb0uGHyEk8iBRe4WL2av/qur+H3D/kvYL3qsn4plLCh9GV
r8vng56LHYscdkc4DqTOSnJg2f0vz57xFLmE5dY61X6Ilf6x67Uhyn2TF+iAo+a9
nj6NaKv5zVNB7k4T8/ZoCSSxq8DZ+3fTqmw3M+gz9FQBjcWqgeKWzEvPR3/hzaxW
SkyUOqXE2IvSNt3qvm06GHEj5v5YPf86T9RYhCOJKNk6S6aDiXaErwSx8FK0gos7
325Bmxjlrfj8t0KTfKXYLbZWCvbPxRaYH958pzPuI8XFmeNlp6Yu/36iCYrx+tBO
XUVRXYiL165kCWXLy+kKnXH4aLUGFXtM17YWxjGk2SpAXppaRBDhnIgmwLcH0tvt
y5AYgm5XtAE655HTWmpo+okUcaRUP+qa6pJNbCqkbW9AvF88Tzdyh0ZcLWUhcNS1
YBQ2gqsJwmVR2bAK7xjK84O0WSa60NSf0Pw12MU4YXS8oqxaTgRnDBXc/KYxv+Bu
1AleifShf0mUujt6+LePn+Zekf+lOBWf2snlqSVOPHFac5BSHKiHXqOcQxLEjO2z
OCrA5ttT7aqwGfkjHO/S30GYW3yYuzU6ENvv7LrqNdCsG6GErq+BEhK4ez60ADZW
9hTp3sa5SCPlYUYF2b8IGJxRY+Gde7cECHMcnMsHlELRb+9Jg1lk7e5G3ADkk/s+
ryakQjTL2koF3j+Kmp5RxqmG3Y3tmxm0NtkAVa3mYUUgTNiYl+XerGKcvvVxHica
EGwlKncjx57kZ4YrloO6N/JR55HXlyNY+AT++SE/eJfwdKtO0TDPncERyI1D8Xt1
OC/4/FCKw8/kaK/7+ySVuCwmMRR717M4YUAj0pK8wOVR23MlymYWfgiE7BsGpC0Z
XsTYTjS9UkmovVTkHivkLN2PvP4M6vmqyKHHVOEkafhrVFioVg7xDLS5cf9lTLqB
Wh3cq9lPWm0byJKvVqM2c9eY3rrQcPbjAJjNt8MVGJGfO+CXwdUiFQ0BFKDFoYXa
IVzz7VO8p6vCpsY33eIHGaBsgIN1lR9PQ+RMZZa8K6BJ3mHAMDKU8yXZGtn4nDay
PSVE72+lSe4K6XSinbmttq4ZhwzmZ1E4xwXYBynpkxI/xsdcD/T3LVCvb7WlqVPk
gag/S7jtoNyhgxJfiIOJWPqHZ8B84dOtOWvdBteEPsfe4xOJ/kxwKDbcypRV6aUb
KKaMV9V5Fdz/Y+DAUXzUDKySK/dRCmgHelu7TSBYRHIyAxZI8grz7//MvvVkXNFp
om49kY1hrrPcFy2fGO/nhqZeoNFkRQIP/ZGGH9ZSGTvlJLb1ejyOMz2RvDHP0n63
mYLCHkGjRAOxb1Qbj5424QTW0ZQhbwHquzBm68TuDzN7qxLePawyyA+3rTRMKJBW
1KMOCll7Xqb2OxdNQ1hMlBoMmqrqHVJBv5YcypNqbrXqIc99LELS3tgvEFIubd8y
o1lLfyvIf5ecYr2JtOWdLDwM/5VEQ8y5efvDNPrVT5JDpRiejHtovjxQWEj+0e0C
b87rNHJ2yI1INq8DrYSDwGdmbUXBNtO1u8yuOhayJKnUBqnut/RsrToYla1rnrqi
qX9MFHMd4V4FsiZ27DwyXvB7yAR2HoPZ8Ggul5mr2WDl/LIHtiO7SlqCQyB/fvK/
K1UOftB6y6ARAS/+wZnUEEIQDQyzH5aKncm+GnSC10yBwF/Fzu9wl/KeqhA4C6jM
xdTy6xAeInQYkLJ+yeGAxLqivqsDOFSfcgVsOOdD0eywcOOhgyiebP2YUudwp0RZ
lYJDFWKQaGoqtQxamsfHxws06UPBv9v/lgOTZlaUCOHzox7MlFfsE9ouwUVN7/Fg
dQQw+LtYUMGrxO9NODlKT3uwFQH79CxdhNDFVCrdaDIOkRyuDuh1AduRP8u+kZ06
O1kPRRQQs5oPLndcM6juSo0YWW7zIFxqX+AvcoCreyJZiYgwwHSaW5/OKC9ejsbO
GxChUTABaFebtIu7xsuJl88pnQPwq1tiYSuL8MgCVyxmb4yWa0ZYYrbkamPY0RKS
393MU7r8rAizzlp3FN7UN8ezrRU+m3EEPdKlHF5qnk8Pv18TX0wgMyxu+gDPq0qk
OMD2IMEc9aDRpdA4QteUyreoqonL3oSssW4U+fEDYGfwVmitwORbYW+NVYjbm0zk
f0gTj7sXbVJzL9SrtVULbMJPKCukZ3Aolj27RLys4ugjNYNd2Ohx9aCkFvkLeTgO
UrdYqKeQLCGJid/GnpiFM5KeAyheHRZp1Uy9qKuiQK9kCfznWErLLult9yOv9KRN
RySo3XaI1GWNGM2Ch/lsReUwUruwrAPUK8ha1BYfnlGsREwHDPooj/8j6zQsqhkI
FBfZaiG9qIzeRy9gAz4upV/oRRRQts3BpMlzt/j2qvSxa4i4anOJHgSDnbMC/hU1
SzS1XKXFACfxzBrULFq2nlVf4f8lBYBg6vgSDSyU19WJa/d4QNGhvag46oWTJq5g
yUtPSZ4/5LJDYNMdNouKvIwqGL0Ln0pZBTPFtLIZQgUNFb4h2RW9Q6P0RNBGfp83
fsXN/CzPzyJQ0pSDhlVuyp7awVjiYb1Hys/9llVmqVzrB6X7caMaBtFbwUiYgMW2
2PruEZqz8sAmgIs0q3Uve4NCn/qH9RJn1JrPZiLVW9l/ETmxBTWUDt2JXeZVxWrf
LzR2c6qX5iYb43w4+4RRrvAh75FI8N6qVUTt2pdnPbq4uzfE/wruT3MehkCm9wjh
KraJw70W0fv8zDrvtLbDW/zL64afpPJOccbWf1QCPzIaGUfbiObgpZBLzPAISfis
cF9lUYZYXL7U8DXoRwl1kN1/SSa9W7XLp1DO+VAPFNrGzVhSdc8yDLL6RhBSDIcN
xo58CjC68NBiwTjy4cR04V3WANLMyYofPO5EAX6s3SmT72gKsVcnIoR3xt5ZMEGl
qiTalLbWDsxB+anVVm+JyriBpa82ihA4wSvSARh9uAIeEechFndDUlCRy52+C5cL
ICFy3eLXmKU3D2j6eDgv/xhFx6ZZlJFk9w7yKpbwTeAatrcWE5ZuoNlaU6icxYc5
yp3PdYWHRu2TcROcM2sU1Yo+1RCzAKnMEx/B/vy9xBkXvANz8YajXyz3P3knWi1b
kk+AvIoyyIZ8wfG/XC0SNOWoCaISCHqtDPlMcRd3/OREiY0LTa8fg2eTp4GV6uAh
56i0QqFrZx2m/cRkDzp2gHYwFbQMuTsAXqmWjVw7CuwcSQjvVmxfAVyuafxYPjiu
3QYKB3T8k/XWlEWBafqhoYyvP8/JGUGQykefupZYHovkUQCjX2XZqvTzzVWHV7rO
xePlMYzhoUQk73opcCLPQyC2xzMBsxJxzLmwY4AgpyeKBiSVgE/NY2WY3gPy6KHU
byeaI7mvsVZqHF+DH/EzqHyy8pikYqudA74JMEav0PpCMbaR70cigDMxgYGn7TLu
6xPn4f2pUOFEUvAnkG2wk3reV0ZwhN5WqcwqlnEQfu/+0eyv5AK0xwB3Sq2+4dq1
x0wmEPbhXlxSOtwLaKtYuXPFO5TCrDMkCGPDCvfCojj7w8qY9fJwACPuTJktSbHr
ymLMkiQc0ESd424HEYwMtIB2z+ipDS7D9SAuIh1z/lB3PAjfR9tSbW+E3VLWCdyY
CFilHkLkoe+NZgL47Sw+3rmxIZrTKgfkSmN30UvlNt+q/xZVEb9qWyhDsfHW9TY5
cBOcndUxicqIEX2/YP/clKULbYDtPibwFOHyBH8/VjTnBKORxz57VBv60+cOuePZ
LpKvlIHA4Dsry7fVTF9urQ0nvrGDOvFtUBM4R0ZRU2ahaJBQhOB/DxvPeONeqR3R
HmukJXoJB60u4GKtWJKxSG3UcJL3LAaZjoX+w0VhUFNV1KlBygtpf+yxBUhwftEQ
lSBZYjbizk3FDMXmkvRdxOHie/rmi8KJeRCbfGKy4zJFzh63eCkVw0TxXdKuZB07
I7SGrNzkMbqaOFY2cY0AbBIeZaismFO9l4SxsFXpQuFr1mXpmA1ScAaEw5szy9tD
szBFCgSp8zkzf4C8AEMpzdy7/ESRQZXFvGfOh+UQzjpUmpHETN7Rlp7CZ55REK78
VTH8w6GXP8o0tqqs00Thzq33ZO3gCpPev6/041i/8n6oHRdE4WGczw1aZzF+EJ95
S6C/W9n1vg+xtXta4haZthU0igJMOFw3rmxwapdaBk+ObSiJlr5QHj9tAFTEX7hj
9i0bIWDGsWPdonlOGw7sxb8yim9yHGBrJRReEmviMXEn3aRyDDCDd2EYi7Zdsi3O
CH8ZAvVmHdGjuoOEm1NP/83Yr2hLlgVsAo6LK22Gzyr/YVrrU3cbJqHjyFmpmBiq
10P2sXjV0brnrRfXN05n+zrsYhvsC0eUv0a49N7SSC0hVdt08JTf0dywTH+7fGG3
szk9TfhjqDBWf4hHIzZwtlFzDT4m18NlB6B2i+EHOre2LYXCqwtUaoNk72l0RvsJ
CPREXaiFWGmmSyVRX+NkhDXwjrCtIXu9g6jCDwBSabweymYemOoxa2oFGthFfegt
G7s2KHLvqYaeSU86VZdTgnuG0WAXO924UjMp2W86ODqweEfCz0SBRM/+GO91Q089
z9YonKpRQMtWPnKoB+WeeQI3OCYk2YRUKS8jcY9OsZCUll113cHk+jcQm4IUTtNk
k32+FaFkuheEPuSD3YZ3kqEsi7LqNvZA3rJB1JQKfZeJ98PbOf53LVkAkFBw6DP3
ujr79m/pdrnBipGwiJI+/MQP5d+IO5L24Q386Z+w28Tb6n2X0RfSwgdykWl5mGLA
v04zvW61NuAYl7AWcN9YA8R2nCC8ATD7DkU/aQUBp/8nEndiLxtZXyrWAsgWjXz0
vKM15EjvCibSVqviYch00LyXu6HvwZan9BSOfvoi9Wq0nNKxX5viKWcplk17+f6K
O8LdSTR/z0ZcVkYrPB7JbtTaDAQ8uhmHLKbUnlfth897Eef/niYo7SzyqboDMqnc
ofe1SJU4Uestkb+wy3JhT0VJX8Jv8/aRuQ8SS3ijnjSeZiiF+TlHGipw/nvXb9wN
VUUeo/PfaygqA10cKr/UCNHQYfOhAf8ikVKkTo5EdUO7eYhsVETtGK72JX6rZlCX
480gabIAx+w9OE2Prm6E73WbVUVvStIvxbE9fvy3UUH7vKNSvqnItTDbKlRh6YI7
2po0RkFrfpuJLK5eFXGDJfCt5K84UAALUXV5hCqR0jfoNbDu1QaWN+KDpSdcJ9q7
ol4g08rOGocZv4UMl5zdpeXe7JxS4mDpUVFajbSCRTxMMX7vIVFYc022+vc5ms+x
mHS3EaDN75m8unURZT/O0K/twGeQlaInfq+AHiyGHZkaSYTmGd+mjoV7SlkiZExy
1KkVk5lo+BAq4XTRTboSiPOeE/HzdPG/NrTi0FMCSQnp41b6V3FAIph73JF0HRYH
idg+PPMOIyEnI9JYU1QZ/OkgJ+Ea+kEMMKjsr+tYURjQnuO5daOGMsFnZgUpGTgs
Z6oUuCXMTveh1ogruxxoYYfk66S4xI/xWs8Z2+xncWhZLyS/TH3gL6325w9MdMQr
IofUlyCDIm/yAbA+eVw3u3PRyb5eT6vXkuKurs36rHgErXlLCEh/dxZHqTSmupPU
cIY1hgHapPRPIbt14LlM7aDBTwb2K3SlJc1z3E7K1DweSuaZQneaq8pOKH+xlLD5
ev6ZvSo+jrWOORv/24IDjgUScP4FpL/3/ziDu1JO6Sgzf0tRjS0EmnHwHUnuGu2A
9awsl3enpA1FS0VtXNaSaP8ZaxcIRnBex6mx5T8lavWYU8r1He+UjtIP3d6iJWw1
Nhge9bXwg7gn6gPbYsi11MiqqCFr+eULFqxKQPP+p3PkAvuqQUmJ8ATiyL/eKUxd
eMnuiofAo1paPf7MGqHt/lfYJnMu6+CbZdtoCf8wqATuUBrmMjiW/3aph/QACk9X
L3GjGGppI5Lc04j+bqw1I4dfeiES0J39ExzrmAmuDlwqU/JO5W6Eupf+s7oda685
/yA5/24wXSw4ijrTFpsVT4UZZWdWa7cJ+Zw/DRXGvwBIM6DHA0+g7siWBcQRVAPN
pzn2UGmYWtfA+qKeZ3zEkUENnmHvBSZQ78V1Qjr/GPUb4cIMOHK6YyH5uaazGoBy
wALjrwh79/VAIdoxXmbxL4dTzrFkpjvu8D5+h617OPJYjhc3XVHB+OShJkfOQq2x
ViOttSVUERa/4RYXEnacVYPIvD7EzpQpnOxLoykLdmxx8uF6T8l4d1q+5qNbgySC
x9Jsw5yAXFEPpmn4E05uTLBm76Rg2W/VqDj4NhPhkNiHnQx/5ZPvmhQ4NBT0IGw4
xxOS8qEtm96pcA36Rs2YPt5otyynQzEEYf8f+wJHGlSlOPYaZbGpfgb8Fyj3viHZ
HLB5TfIvcYzfCFQ/MgsR6xynxOQt4pyc00ZcOdKynmSvkSnIQTIcRTOnDJAfh4dY
B+CXdl+upXQjJAWqEg9utu4XYm3EJNW2busPlaO932GmfZiJOIMtY424CZ03tXCg
Erep+Cq6NGYEdMgiN/vvX2WWFmkj8q+4LQJCwOgRRFRfU78dy9Ryz6ApRTVKJrQd
nVAKbwQzDd1s11gtyXiSeXt+NxgzqdUCGndU2Y7eFn5YANmQze8SFPwy0rYBqR8R
QsXkpPQUYimIOZZh3qI3fWNovTKzjpsWp8BP0pgMCcG274VX1+RS3brI+220q/IQ
l8yq+z4m/eFhDXKzDOdf5n8kILPISz9YsuPobLYmfIKXpXmFcVs3/1B167Pg+1PU
qrgikMxkg1QTjhW41Uvl8NbI6yEjihNyodxBBmAvcb5TgBOGmb98D5J/MWBkO4ub
QvO9fC3TKZ+WXXp96zfmbz48UDr4XjMASlrnwKZhMCIEu9hC0m7GmLtnL0fAlVbb
X55YetEsjVbXy8UYe4skWcXofkOAF5JoKBN34RGgotNyhtFvdQQL+fz7lVfAN1Ks
71NyH0+ksAkE/VXQpRzeh+aimgji6GPxw2jCG+HUMffXpbPfe8OX0VkRIxs8Im/i
T+LfAaPEtK6qQc7qjQ6nMcvxNnNhB+ZJubfsj5ajFE5dLDlVhbGP/f3SvjjecMMj
Yc84nB9XPFYHcwQcnnDsiNw6qFgLfxx7VIHssXokRWJEBRvgmF1HgWbY9h6dxu5N
Cf6gU/gdIscudzyvzFVyUIvbYj1Yh7qu2cb0VPZOdWz8jh7EPhxSCPb+4d6JEwmH
CKbQNCycb+hcgQMSlhhKJCgW3prRrG47nRj6K/72oAPzbH5QKgof3QkxJpnoQz7h
+ex6RmClRmgYZgzYNvbB7RwSZCq7kFGRXI+iMNxEQrCq0AyMItGIANUAIeZ731KQ
UDK6K+7GuOeLXGvqJa+r/Wbdbkw/re8j8R15QeFg9zEZPrKouC3xEPRZtDbU/MVM
zfLUpwBACNxwbWvMjms65EjRhwKMezfAKFJGOQ3I98q2ayjZMSCQdguduwiUlf9j
e928Vo1F9Ik9PjfMSBrS/jqTppa278oGnW07QkGhzdIwaOJU881aRtsINU8AALao
zlHj/tOMkpDaOUtVNkGd9RyM2OiuS9m1U5CZlvu33I06BDRkqZCRkdjOBwGNIFXx
9Oit7m8ZGz/YvU+4gI+Gt1On61v1qmqvJ6hHkWOS5Gh2iSvgvrgAiEcBes/YzHde
NFfzt+vhZz/wQ1GK4d6YBxPTxDFRZt6aM7zKH9gs2dkzOrjqswksLBKSPMH5lanq
LC/fdXS98PpxCnM3McRTMJ8SpShJG54THDDbso7r0TdlHLwXC3/nkZcF0K/s+kLh
sQlWayCevRCzRLCUJ7qb4q1rdnAe4oQbRfQ/dJ7yQPHnVXWv+EaebCHqNgol1frq
U9vGp/7m4szCERFju3d9uTLB9pksldFwZ1XH6zpfSfX/qmU16tmwpgkhn6YOQr/f
TD7F59ybZXim37Lt318kxb3IHTbbhseXiVIeGxRRH3ZaCu4gfHay0NXSezMOYswb
AmkQatLVkrzYVxIllFcQNkIPcpv7pAoMMITmTEcP7bL9qyeOOz3pb56WPFMw9xyW
AT1FrxSwo42kV2Io8DbbqHNJ6fEIlfHdtAc5FusR37y13difT47yZ85XoXsUI1LX
Y41PTfjehtfQuJqwDu3GkQabxQgImbzfThp53GJdeUrjT+PDHfcHDNYouBO1BUSK
RiG4vYoOznCFoUus0PVtwqh07lmxOR6y329+5MZsFzxoQP5IPXYBpj1FSPQdzTAt
p8hSMq0qDHMeehSXzF+kKSLpcLhUR3qw/l5Tuwyjk6fzIEtGjrQOO+hVZ1Tdqhvu
HFQnVzSb0sS1kUD7sHpYYr8HxEcMv7bPd2DkPAmJpDmyOslsduo/5RD4/x14VLcA
6HUhoGckeIFv7ENSkydaj7cKCNBlWt1Dqs8yglSMEMW3apMfGYje9vnHOW3lzSSS
W/Z3ayrsipN2i84kgVrYtYfIAYoPKAgDPjGPMn7C97AUkRgB7tJWQO3kQLXqZPVG
SVEGy/NKKOoQTXfAokd3TfP6PJ5mhfVgvt+LCxfPf/2V7tqxzjTCoU3/1ubt31IU
7rOaoCiLx9AVfAOlVazjsdxgfJXQBajTeRC+kt1ChkbgBAFv7ZU2a2PeYWtj1o2J
g2VsbWS+t7H/y9GRbfSoOOwNx1IG2zhYzG6U7yoPxtoOMwk+7Tpc3lc5/2H35Fiz
PyFjpM0GYS62HO9IcfcIypNvOsfrnMfD9kiV6UYFvi1bXOnBAiEgpCGIe5Zv9C5R
E3KunzEd4vhDFeRZe8wGi2ci3I/bIvDjZ55deJHFYuGRNVx6NrURvwFjBAjMn+FB
nyo1EaMvDJdH8erl49CEvz+OkaGL88Xc0/4b54lenWCNo0n50sdH+e9m82soOAKK
2fcF7HacV3CUwsweL6QW1H5tbir2GNLaOdfx7hsBPQA2QbmW4Gpn1d4oatIH1ERx
CUdFGsBc5Esnex9qfGy56G62ZJSxPcwI2UEB8mlq25UtU7cZ4z7A/tngfziCOQRq
BtzsMVLT4tpBBs+lriqbAvwT7Ir/NIyVyjTf598DnHQBitcQ2wIbozCmoGYqlMww
GlR2R4F2L05XMtp3BZ71oM4lLC+Bmx7xoTMc+j1u0xGRP6mVa843fRJqwnwKGUc2
5BSzh01N5O+7VWR/YfEzY5EEOreCG4oFB/hGtFIyf2smAD8GA/n2er9AzTTfMIh9
3AWXmfNDBPa/Hz+9fJ1p0ZqXpvW1RP0IbveE8OVge5K5LUWjI04MxjFSa3yc1Tim
gQimZUAZf3TKjXRIqo30OLwgriNrUOtPFKbfVITxyuKAvaCPa6To+3dNcZDpM69D
vBEMXOJSN/L3DdPPNCRwm0BQD0qhu5MXeo7wDDrVnn6kHUq/h53LpfFvnR/o/T09
1Dn+kpjNfZZwuolpBeJOSOfFVywsbVZTse3rwaNUbddyk/HZY3H5UZMe29MAYs2w
ZR7bKL/JLzobynxb9GovY+sjefi3idssQOW3v3MEzLifK1adlSXn1fclJzIORpMJ
l0ptF+n2n0xas4P4QdWo4o3uVHuDAAQK6ez/jWIeAeQO/4t0lnC43JrVKS9AaTjB
DVywDQ8ft5n30nIi0G6ICQqp1hTTWH5c08zvR1QrgQpCBK9h/O+BdUIrbXSOGzP3
WUrqZv3fWzOsMQ89H3p0lf5eETSJW5n8qFWJxGVEWStL0FZ4U45YTOkpyd6oe+2U
0ObGkrH+6tSJhyLjeMv+tTPZl8m/k5h/VpCTpemb51X1W/FwKyUQBg9pKj/Q9aV7
u1OhLOzkaG0V8cCqOTuXU6BMHme7A4w0QQ4nawFXW+4bd7TiXh8MDFhWzirJ67pO
TCJx2pq6SBKg3rLabNuo4CfiOFpTHB8A0caPcOAEo6oVMW5Q5QdKIi3dunpeuuLP
NVYi3AN77L1js0InZd6ZF7lGR1ae1xDbIWAq58zT15LOfCAnvp92DdoPmhQxd0eQ
M7ghPLnraWjHCKbw6HyLqH6shm0P0V8UslmhTccpK/fDkibiuDOldewa4NH8NgrX
zCPvcHXC/qEUX0ohyQnoA+OGzBOSBbJjFmCe2da3ZTa7wL2BnjHnE2tWlPqW65/6
fGIp2eTVoukOZKBr0tyb9Qb9UJBQzDlHJGaWlTtFjHOLqjF0l3clSuevHRX4EJUv
029gifJG0f88Y9plPHVVDlewobfa0ySO2dZIfpawvRCZLiKlANWJDcyDJ3zbk/3M
lnU+PhH3e5DIq0k9ilyPeocEEBkZKuBvfxdSijkdqYuA5cytM6Tcv77OoTBYyVwQ
OnDnUH7YWX4Cc16AWk58uy6AIWiFrEzLvrg/7C0kIDUvn4Rntg+i4DxRhyfx+h5d
if9IzHgsNDUV2zoxlaVX6oEGfzF7bsgPWfjEuMJu6+wXla6+NVO8pAZfupwfduJn
OuS52GJFSWr7JoF8qm2XWVweBBaW/NSjC2inTxAJsoBRZoXTdIm1ZEvJyeQ7pfgk
oj5FrUSr7azcDKGDFROz228FgFuORhqLhE0gbzHJmVkOdBMAczuySySAen9FvHwN
O5s/CMTSpQfIhLYmMCRLh6LzbIt2kQuq43eTcIDVVxtBATmujyl8m6xWs+YKTzdP
ujsa5lYghUArcnJUXXtPlaxXtCn98AcjisjQ+bW2ezk1qW1c9QcanuIlq0mMTPpt
5IIxQKwLxj/XLHMPPyejZS78IdfdT0pMybDv+q7Xr8D2UEhTnq4qQl/UbAx2AmrE
xs3lnaoac3+QUq7Ie+0CH6NCujZozCEWPJwAtL/uACFxDt64EpL+59gb7PwhVjI+
j7WS1s6d9X/nRcL0HYEhkAYW9qIlqx/76yS+tNZi5/QOa7v8YTxWil9hti6Rn4Ho
2NyMYPMwod8YkEp+Mj/lPJ+3DI2e9JIgrw/IqM8Gw5LkeQ3nC8rn/WU7kWA9tXoY
U/fSYIcuaFZ2h+DmVH4tlMgmC/UQqv2t8FD4G88T+CpRoQJGhwea6p+b9bjG9pc7
Jmn6ZEGZaE6BCHNbf1zUi5sNcOaxHEFdCqfaOZq10HTLRSrTwKJYsiFmEXPkMiIh
LotWKFiE1ZIDdrhCDn1rAJLazVxZryrASKOh9MRigOMESAyroOVyExi5O6WSYlaa
Bjr3EKqoaHQvQWgdfPTj/a2oj3WeyIwkhE3wKQ/iNef7JztuVk1pJwD52xY8EWu+
7uQsb0tyDwh5T97gym2L75a3iJ7ft2oiJOU46yWj7gfkcy4fwDlP8JvD64wRWpWV
HDuu13y3xJofimrfNZYfV4sP62lZboJ65jMyzXrF7s08M7ktNg7mHeE28GBxhQ/5
XsWD2I6DFzzS0cYaVN+qc5ue+wOOUtXslE1TIZD6Xfl8f9hDs62hGYxCvUep5fRn
sqXrHyJImrx3ILM+F3pLzNQXBBDN8Iy2zbAZZ1CF18bzwuJC2Gu8DsJTBRcq9OTf
jwG5hjrKLQ1GRDfFJ7hOvX7v9rgOL3690RHD8q7ck+DHajwWRelKCYoPegP2On+Q
CJLemW/6iyu+RhjEbbabtYWP1jvkVmw8VKyqOCOdd+Vc9Q7HcM+ElHtNcAWQWCFj
n0xL1mgpcaLEJVXj2w8/u5WtUH/tvv8+VgkN0glr5p8dT4H1Ddqeny/dDsS3dveR
GW98hfHy8je/35RnhBSA0lUqFaB7hHjYrIox8pHPksCc3s5G+43g0Q7vGTp2B4AW
GNSl3WEunuXXRlwhK6IN2vxmDcSDjhPPT16rjx3TnezbcE5VeBV6Wwp/K9GBMmOA
P/awe9r4Sj4Oy4ddh28PlBGUbeamKWMclN/GztDmJi11LWI4ZkjWXrcflF4LdRNm
IGQuqXPxSNb//uINcIee3OamJyVAfUmlqPijoZLOock/ptdK8WgTHs2+vAh1oAD+
/K9CIv2X+WWvrMwuAdkbAiPZHjAiansuOs5ZMafjXC+tfOCn7tPRNuR5JfygEDBh
QRCfg9RxFNFU7CuXvR7h4ulFjvwxLJDmxKrJ4/nfvesx/jJ2zPm1zh/4tR+2tr5z
j3VHrNB3wg6tzl81g1sHfc4qR26rpWFkvyAkB1GLvUI/4l2fMtwa5g7jDILn+RnM
f2ZdD/lGkeMWreU2GWZhrDm41uORwmy6yS2inO5ndIagAIpmVPMzT9fr0pKVsE90
Bbqjp4YtMtlbVCvubCd5F8iH8lZZm5KWJ/FfUiilzimEKVoxbkChynGahK8lSUQD
N0fAWMWqM8CxOt8+SeAoeiv9g1xGX1gjyHIFl+7zFQbW+t8atjOlrB7XeFk94Win
me9ahT3JLZznFUs3fKFBTBlBTn6ktgvTNm8ki6B2PSOwKC25JwKBuxLe6HAoJliV
4ZAQ98wSQJPwX2JbeLmPv3Rzg1D3PFo/G+z5yjPl6VeCQQXdQulN5/D5GfAYAliD
au5qFzjgz2npalo/RI4e6hsrZxrcItWMFPtDM8AYjbX4ELwbC8C5uGewbyQPWT6p
sXdmQx7ZWtwbLVOsj4HvQQe4FrBlrDNCfujgI4bQKPNG16DHyO+nbJumBsXPwJna
j3fsPzc2AEK7j3uHFMT+hNIXQuCMSB/jO8Yw+tTlBmcO3rw0sY+wljyQoLWhFO5b
vJKyzMM4cHUlKaI8/lU2mKuQ3ol1gDkVOrX6ZWP948FrDy96Tr606HL/M7xuxM/p
F4Q8G8AWsxkyLdVmx7RVvRIWJgxdAf16+dQGgErwA58GVizaeV6/AnVFbkHG1G6T
9uNK5gVSCc3V+z3zpxk3hCEDcOLSOvsien6dRcjNlrGuN2g6RBUrcl8CPOrz1AEa
U12/+rtToUNz8ur1SzBpp3FnaxiF+X2yCDvwTXzBGjuJGvlvzaaC3irAOGiVA1n5
fvzteJnRU0r/ASiZ6yzi6RhAao/1RkCAodpshjMS+dvTGnvIiWryRWUI0vrGs6vJ
tML09e+AaSgzOYFhVvWj8KCvNsHR8j5ywbJP8FkPhKxT9V8r2mnW5c9d/8IRNWG2
wPBPz9Rlc1a0ah/r8vc5a6QLJW1Z05Q6kqf7nBYm9eHhyF0Nz98EXXGFB3VNeqJ6
qfPj40sLXHml71tPg5XHnH73MqTrAmYgXYb+TpbTMWFCy1ftLYcWhjGkFrzHG8Qq
fkUPKiNXjLz8gFi295NFN8SpgX864rlf1memxzm4eEFHboEZBFAMNDXFqJO1k/8s
UylZbaVW5KokFVkeFi9KXO2NlZ9dCN9DHuoYp26K94IitV6vwaX6ABQScDYg7ABD
aRPPvut3NeSEqEJDgKgzSodE2j4AAxnGf+gACGvHAbpHbI+h6iTbmtcHTk2+0ClD
PuUpQha234xM8j0cxCjtyHaiVFgZT0sQi1rsKvXjdSrm1UYfkJfhnMZ5cw7EbSqS
iTNMOPhgJaxriUSLJyqxHLzfN5haorO37vmAeeB8B5fmyzq7VQI54SCF809BZZVv
SGxBMelfHuSeHKVCzpeC4Ijw0irfusp6lcfsDP4XDFkojQ4lp2A0ZmuwEDTwD3Y8
ebAxliG9NMoNveUATckd1naBhfQcR6HFnhb5/RDdO8DrL7Sw7LO1P/KxApbi9G0m
xcXKpsVzVCy9AFsOUmXPhObloVzvwicZkVS5NWT/OsuHXy5Cq3mmCkV8YDWYLTcf
mNGzHF4rcTRdEfRoze3Cjp+Wp/kkU1QYtODJtzCNMqT9rza1+ZELYT2FJofGqqgq
VrE3Rv900aic1/SeFNByNOaznGAabzEljN9DmvVRPUln8czp8mQqWNl1NljhKrDW
HHliVJ0qVsFg3ulrAEPFa2saghWWip21VWTGVJU0rhE7LcbeISv2Q40Q6IjyS+bZ
OnrA4kBxYYJdOZlWXhFX1ENBu5laqSx9TLDlh3mDvrumm2Rgg1jyAfh9INC4NzKH
AZDtJVhyzZJMdxWEwSy2sl0fPceFdLFrPnFxzyg0HWlTJysPd75Z4QXyvd9F7bcR
AmbYTpk8Abp7ZiTMMFAdryf3qQqHkXZyQ1SqW8qy6WAOA3yEqV8FUohbdK5mN+gG
H9X+9KI5rKM3SmvI0akAuv3xA1ExfgUZ3bIC6o5HoXyOvCWaqj/9GP2g8IjR2EpI
4RCMt1SeLkNJRQ/wR6+8rEeBlQuYSOX4JZAqp+CdvXDRplO6qou0riK61i33qYWb
Ib5U4GU27hgOWCAQJA7WRSTDkYrAMQqFE7lwtXrlPrmoARfEvEDn0828Xn9lYfr/
s8+s6nbtyNKW3Di69Ptg+BuolM2lnMxEPTb6UIMjgOcPMchp+AHdvYoUmCUCr59r
/paFdIupZ0gcGXXfx4Peq1fR39x3t6PIr1lo/yqFDhFZmQEn7p+AeznCChgb9Mso
S6EVPUiaUi/uhrcvBI4jtgqJpeoY+oIrvvxLBVQCRGswWfly+Jh64JD8nVaaLMNJ
s9SlGQhWmQ1/V2DDMxzCxg2ZDgd7DUuJBgNqiSsPjJ0GaQEM359eogW6NmjGQGd5
KFgw6VfbgwtCrrf8JLPHUzABFO7ak+bUtgtj/JpGlGa5+zWayH9kQvmIFfgd9g1q
yfVHCoSO2MqKG0QtYbiCR9yRCteGQQk0K6ZVQQQMoEQscfuGXKZhnYlCM69aVDGK
HP6397MSQ3NeXIpHuhSRrpE92TMW3PJHgx8n9RwCAiLW4OHHv3XmG2PNZQDorzL6
+ME+Uk5+FCMpnmOc0nnkEkcmQ8dpbgGVB/W2Tq+UtgqjlSETeZkBa9ot1tQbh1J+
q/IGoIa597NYJYTVWd219TWK/zKJ97MnH3uXFPXBukZ7sWmxDVLO0Ys/G7X6WhBG
YFT5VvF3INteYMQ1gJwLREyZ+lDYHqJ7FVIg+kbwMhMjmLhtn7MSn33HS6drwri0
CA6y+pC92CDXa/da5D7mQai6PPEtBH8WUw5S1z7VmOvfL96N2M6QMowSZGbbA5iY
NkIbKmu0qNAlRUHUAMT8xpvFShK0CRV7VNQBYkXYa997Ces6CCkb6vvhJAkwoX1H
9xbDglCV7JNsvoKKUHfoZ/aGUxrpumaR8CtWC6aY1KU75rJQ8foDCpW3DBI4Cpnm
YCE7ZQI4ckimzF9PFDQ3ECoq2fnDvZPA6PW0oJU+oZ8AcBqdFCWjOTUMvmrWWbqt
0EJw9gf8EReEd9RLAyQdzZt7qsJRxe/TNDX6+RBhsFL5TTmhkzs/iDp8EExPpsBe
dyZCxC1vkoO46WroL0sq5LXetzwog5uxF7OajrOvnENXXZcFe1puAqeCketB15cl
NHihPd8lOb5Op3VSik1cfGCYYJGvOz64bsfXDLvhdMUkz5fXEaSFkaB6q0fhQEF5
El/hvFUGCqFOoyWsrV7Y0SDQge4WscnENmTTvUErTA9HhymSOhN5IPnFQQT7z5b7
QWYfl0uGkx28TCE4pIZwDp6m/UPQijZEsvZTU4d8qp26UB1bH5K3xi1eSllQlmEn
ZXIQUFDSd5rgP1kcxWHYbSRki6YR9MWY/g3fXGPEe3CRbcjkUnPT5kyaCgmO407Z
YWgsBaESHuMb5g77l1jaILfB9GIKz9it256bENs5Das+dmZTftyGJ0iYUPJuZNk0
Tx1tdkQAL/5X6phxuRv++GZfMpKgJnBxZymvDRQzMYXDmRKPthXcRvpv4DsVD/Wu
lc2NMf+SZeJAqJzUer+qZht/fpDFMNB1fM8TCbZTTvb8aGubCxvwHFp3pvPE+oNE
MOjX3XhzoKNhxKAY/V0h1VIvTTRYu06Xp4powS77D7LgpnzliWtmjG1rqogC908V
/1h97iCIla+9z5fkw9Q34yHnhPL8mGWCGBk/FGFG4mXp4+9/0DHh1kncLr/qbXxG
2gkweaW865ITjEAr9Q3d/Cwze1fIS1Dm4g9UTZm9316O6X65coU9CDxWmQlved52
04YH+9/aa4jJkYN31WnTozzpJ86fWv9f/Kfph6+Tc/lv1zL9BuS62GT6ap9yFDQU
vMPrS9BqUr0kGqHYdBjOBoL3YAmk6KPChwNqGxSljlpCs4Infb6uTf/1s+6mLcy2
EaDgnABLiKMWGQ8xmZT6SYQCdPtql7aM7u4jNWOCt91x3Xkk8rfgI/R7uxKOFB0Q
Qf6BN+RXxpYRj18WdD30hE23L+oF+2ygi/M1cjSOhoQ2c3baqcZ3kw1D1hnll+Za
kefUO2Cf1ybNupysIuLm4EGv6rmgJm+LeKmxiwhvQeQY4T6XboGDvBu0zssVn+E2
sNZ0zRhVL1R35tTI1hAQcK2pbmFrARIGcim37pAHIbaIYmN47byXN729A19EJRZC
DaY8q4t+w5o6tt1gLkumORaIpSTe5hDBD6yNeaVt+G3Hi80P8KED7mPU3jfLjwKh
wS6/znUMYPxjjx43qWJO99d1NeVb6z9dwn6aQojpYCinzNQ2LKSlBl9LzgeWHS3h
qi/zy4LUPZ9ycgBExyC+soWjzT0vepv2fxEH7i2kuEXQJM+Exny8llJMvEzSXu5f
I9gQXXwtuXKy/qZ+VvmjOifwu07zSX9P1KRIQPMg5T6zcHZdb6RrpSnbau8nktR+
SwZXYIA/49LYn9jNwX14d3wmJmQimB+nK+N0gbJ8HSJsfy7o+E8x6k8Tkz2ik8MX
8+yYxPfgWyYXyV9T8lv+4DLeo9ioWtKQv5qdH4Qe9G4neNCWFnDPu0AIeAryCVcx
jm8K3HHIX1//THq3JYhmliLTT8V0zF1T0fcLN2TU61EWqEkfbFl2p10ky/TXiEAr
+Rc4HO4mH2WwQ86mX0+LwYvezE4lXETkG7f2cGa2hUQv+SdhXUYNM7CgGAmuZfhm
F8830FwrgZWrrumBU70v6eJw07ldtaRI8nmJv1sjhuFUYwqxb173MtyokfJcHPnS
P4XLRyqLtcjC2c17AyF1m2A/58dt3wPpfnijfMNRSOLwK7StJou7ZGQIQbH53yDg
Xm9fmUXqZwQzL2WMO064uAhdIC5IdaEFO1+Dr5jvUSWbgLE0MKBn1VCjupca4qww
OIec8s1bIYhcasm0VBz8L6vRfsRrmgwKu5XgjdVe2pnvOlVP50DP+/ju+qMBfSBZ
QsLH58jSBqnN074Io1hXRgtEsEWj8bl0cssAKKfRJqRwBu90oJINYiiKCd6Z0YJb
Z8hP/AYL/3/G+jdI1bhiH8LByP+VfJmrwYgJAPJNj3wRDr+aq6YLhA5jh71yARfz
G3M9lqNO1z82Dj5hmE6eoLr5IwioaKSJj2Km7471W38auwUkgdaPkXgTT7EANP2o
SLMIDDq21yA6f+b7ZJK0vNkeYzE3RO0QHixb8dbl+sQqukQAtTwW1Ca8AIj7Df0S
UmwxcvytOvBx8xfCnQ4a5TDCP0TYEl2DMAKMSz9tl+XSQkYq3TRq+Wy2bCn+fbos
K4jvHLf7fgFYiQ33A1PQnhk2+vgCujLi9w/5fz6a+UMTx6k36wE7d9+S8mDVBBKf
ddHfzrXe3/ifciHF7VPCDVlV/698BjwUp/aMOS+4I0ehFzfUUvWvKnRwd5JuEhS2
HNL5TCUMvBuhTp1i2ipNV+QzXe5XJqgKKl+zSC8BhA2/RcaRgT2XaDjjC9agrKoO
URocFPlMcYXiZrRWFa6Q2ToNCBJSpjnmYKUK4a7ayrWtgaKpUKKVVBuFDb7xaxGG
ke+hk7e/WwSYifOWSgUV61wWO6C33vESUvJ49iCeJrKWD5mLPMrybYU1kjfZBm1v
+Z+TcmdrkoFMABab8ouni72plNagSIfyAaKhQlxB1+dNExqZ6+dbCMu6SByL7owX
/S72kTcb1AAmq3dVpMSoNrEBzDYJTh2nqjMc+KZUjn0QYnDujb9B1YNE6gYe1LUG
aHeiumuccdGDq/JSS72pqQwhwIyigKPp42aiXYv4ceayHF4jDF+DqoHNUVOq9+8f
zG/+rtXvpDOvNu/5wx4i8h6mB4+PBFYwVb9HKNFgATLvAeAm78B2Al37rL0YwOYj
1y6PAfW37EyS6IOZeD7a8EOwt8t1v75n586tCMx7l4WeL+zGvAuDk3LbQVp9Mxeh
mV8/mHU/li/mDC8pkqS9zBFhebpbT5ZfQ7KRzhLSBh9P0VYLUlDTfCtzndjbVUsK
nQNoe320/VDTW/VwvhuvFw2wl7C0MKXd9o0AStAZi9tHqcYF1EjpzHNmgue7tgyd
58VnqXbLPsJyGX7ZsQWmXz2Q/iSXIUfZ0vFnHUYb2oIGc8H4Ehn+oWQyyiBZGFwU
kkwTiEFOE2mkZPAAovMEdzGl1A0MJFMoXNIPJixgj9pHrlhYJDDsNE7eFW9uIvYG
3ln72ZIrgLNK4oZk7zrDc8ku4Au5jFB08pDQpmADr7ZHk41NQJ161yeFbSuFzUof
ljehU+RbO8sATqbfioMhQWv/4hXFSuoHRSIyrMiXweGGXnU+zIXDKzV/LNuRKO8S
60vgBjkupNOlo28Oum1yqtXO4Ehf77RkBbIMBih7XzaWXKCpLyx/ikIstMkbqG9r
Rbu4/KgkvXy3o7J2wEPGu6mb6RKholcfQ4MKfB9faZHHw85V2iQ9oq5TLMV4eN4S
0j1Yjcis4h7vfvQsAResFBBOXeXpYiiJDRjSol5j6dpympw4KKigkVvmnT0WNlA0
Wy4Ajg9sZ0ynGFXqEMDBS0yVxsDQPB2U4Kjneu3v6ttclcOBAOk1lzR/8ZSDpOcV
4ISXezlhom+BaKYtarekQuWib1Z9cPmPeBRi86mkkHy/F+Ibd49+gOQ5IL1feGx+
6x872mwSP8BOL7iH/8B+lt6wJlwKIAcjxq+/HY2MsgafQPzNdh83jyZU3T4dO/a0
w0nSf6cAje9GeepdmhJbuKSu2SuWtz/1NGEecOT2Ew9rEn9rOX8p7iVHqj/lnUaH
WuWZf2K2HtlZvz5VzT2kODp9oY3GKTXvftnkqnzQXjkBZlOFf7305Xknuo2pxPjH
pjo/q07tCe7idb3lrTyTiabRkrJk3qSk5vvAJkkBpW8jrl9robksxvPboqb4GgxM
w1Mw9gGdVbmfsuV7bXGFksKCLOJ6d5vHLy9S1ZLATsycDaXS1yYa3qAHA8+aCTIZ
pQHXoUTWbAjekg6+Eakhh1jd/yaTMc7WAcw4F31jaR65T/R2EDCDlzi7ypGIVgbv
O0rJbKQyBfReXlvUIk52aCawuo4rfGSDDX0O/mij+VbKDIXxLMPXF80vWXJtB7/m
uYW3zlRtnHr7OmKVORp65oPMUf4Tk8iEEM72FhhBnJkEqX28NgVcfa8RkdfV4Ui5
8Ztp17FEJVe8iEUq3kLkYN1JtRDml6pbYKFSL0ENHsf58JU5Whifx2ELFyLSNMAo
fkeWja8B1mmNtCkEOMEjeIufT0EcuezWFeOB2kmnM0cEQSYsDlMzs3cotwiC4zVb
2jgda/Q86yZYphRItYR+f0Vzb+YVTBAsXiqw05l86Xr8GRn7m3HzGeZnSMqZSgOb
PLiD+ucfMjnIFg4FRRnfX118nio5r2dQ4nYsDlW/yZT1CFJ8h6JxkSr7dEzdvZIN
0J8jRYdbO/ScY919Jso7nGsc/aIFy4YJuh7/L6GzUOD94obukRWLJBk3q81h42AG
H1pXC90YdA76Vl29ZjwCamQux0ODxMTh6WwURdWJICIbHV8qNzWqHiRWPwWirUuM
wCGTcLX9kBDHkWVL1/bUvOmBLAr0dCyV0KqJt9EZumS/ZFtyY5KTjAsSMYDXeCur
bib/cqqoLfA0Mflkfqi6kJBTE1FP40Go2DD5/mgsTq2068sQwi160isA8tNTY8M3
sWwoySVBShhri+6DWsfsh7wXdxgGL+fxBGbO3tXFuRkvjK9dbrye0novnVwtzoHu
qHSt+7QfrWh71jpoxETMPqTnBoRtU/bQgi5CThxGLgfBCDPTJTIshWnNAAFosdpe
02m4NNhU42dynwJNWNMlKMJIHuHFMRYPR/GRanCvbtULeN0uRAaWyrfyja+YwStJ
T4OIl0pqe2w+FtXJaqlmFhKTdY7feDEyIPvY3gMWRI9SGn2w5473AeOVKgzjUMeZ
b7otOE4s9aFBnD7Rh0bxn2deBGjEkS1PGU44/AdQ9Wc0c1yYmy/enZK6+K6zGx8t
qD7xstJ5wYvubyZvoxGgCkzgLvPTWPy9HTkKJDrQFAf8ABCGRMEYdjgRknzqa5xN
hbsOLUixtZFvIEm1BUTcvhBGdQlO0DRG9dRnG+d2rF10sFYGP9y/mUZDx8mGaLAA
GUadE76MRV3bofNkGWQsINaUhxms05oB5i9hYCFEEQaJEXyNbYIR6G3zTEipt2TD
kx0VG+JDiccjarAG01iUG/QJqV13FCqerZho8U4cLGhAMl/sv9m7AfLWsXshDQwi
XksShYYYzH71KEW6A5tgm7+cpxAZK49o2AeCvMfQTYoU7mP3csyviKFtSH/3lMhC
HBpEMPaYTGmspg2ciPP6VxTamtogv5fI8Rn1h61/UH0K8faQq4Y8cBjgFnj07I8M
DKHGbC2yUMl6yMnJclr8SLq/3sx7kRggMkLWSPAlboffQ9W6LfdB2dOQd/eC6Uqx
5soGHMdVEpYcqasiGxXu34S5CLfbeoeI2CHhGXWUhb5FeMpylqGJSJBIwD9wsuEb
xjsiGPfk99nyVZ34mybUnvT3h+SxdUkRHpDq33Qhn2Yt+zK6C2up76D+p5l5+9h7
2LwZTQ9PExHORg30rQ0exgirBNkvrGvLM3tL2gFi0YZs9UFfd9fkjGClMJCaAwOT
iWc6YgeYEvswRNG1fczuoe0yAKo0IkJRJuXU7DBcCEChtNvLHzQ4x2q/IAdfDz4V
K23TRalY7Pm7M7dzb2KQtlWt8XoxEVzKF1mrTOlgtlXuZKcidHx9Cx0wG8nnB8Yi
MdjDdAZ/OsLHNJ0XElpiCUfhCLgTAyNNY52AXoRicaXYo7vl68N42gAa4bFrCW0z
pRyj6D3Hj45wDIcvlpXo9uxsS5CCbjuyE9LKd+oiHqVvCCjZnunXcL4I00qlKXBD
Se9aItyb7pHlEBmhaewk4ewKD3Y+6pJC6fcR28oSxf9aVDXobG7A29xCE5B2NNes
GD5ELsVePQ+8+Htf9423dHot06hGaDcLStTOy0nZoU/om6ghfg1Dg75yVwDzNpJf
oNY4a2SXqzN8fWCDE8RT2bj14gP4ZhDatCyjWzlJUIlIfF/36jztgbZXDtVQQSFz
bb+hy8V1egg21kszosdBWW/ntQQx3ALJ+kiDYUrMNzSMS13NOMrIuRJkPqcJdqWd
g5M7uQ8+vbJhotZthtpzDx7M+ArgjFFKyVfPQyk8agvb9ad4o0dPnWbUxgon3lox
WGlnnr6TfjPyLXL1sF+1Rq/McVy24YBcLP5dSgiqgWm540EWFi5aS3BsoWy9JZxF
QPe+JndNYpPoCLsLIdPzFUww0YM89BOyGL1XhO9aGs/6JISRJWgOdy4nA8Ty+xNp
3EcfPHVWK07qSDk+EhKVj8Uk1SB8tH4SLS8TFgA1oXrG1ZFJ982VM5LJS+/+i1ah
8vEnn8mAX2JCkpjsGGaMKbziZFtiBvvS2rnJm1N/u28twcOsqgCp8gxdXv+idtUh
cCspgU94D4/mtLzAPtDPe40N+1iZ7KS7O/rX3O7gK2D+bvema5ckzD9c6IiK5M3a
4sqLaByhq9Wh02TKX8AOC2nXycueURJYF7OErIITLrA4ESO2xRuuztIZiGxhwa4O
Ckk+viIFZ1FoDxnO5JuSeq6045C27siYwqLpoFFSNit4/hhXKG39wnn+AB2EVE/Y
IA/FykjUyiKT8wpdpQd6mHd2u0VuAZjnT91JF6iSpzcEgrsXxO+H5VGLGFGk8yuz
GvmfeDbRdlO2v8ZEox/9pedh33FMnysIIv9pG+v4AQU7/VYgfrg70Sh6qr+C7+qV
75BCFzEgtAonmHzUMD+lA89mljDoGuKrI2y0x3jJsQFEzOJ/2sjWYwyZDeDmWl1b
lSKM9UUMemLE+5J+3MVpn9I/IVIwwkTh6/nBnBk1+CjMlWgdq/lQsj3UZ23/qe02
+HshPea21/Re0ehIvPwqyd0m5YkJiowBECUjZHmAxpdBt1geW63SRuXuCDcZSr9B
KWMfmWTRHMvLsER/8XHVYfJdZpairqrIuqucH1dIyhBC2QQSgDRd4G6aDMieDvtm
cBMT5+qibu3tZqPkbbxk3hZAqE5uBZkHitxfs0t/0BhN13ZAqiAOr4VS5bS5DcTK
4pmT8JNMsSh3pIHuCIbZH/CvEIgwMKSmnK6XEHDmIHrVO+3tz7eIk9OzeDIbNPtb
/3LK4qvFPmuSmgC44kxCB/0xPG6jQZ4uZWB8bAORiT8pUgMxnv4CsmPTl2lIfE0y
OYDjobLtme16N8d9XahoaMeH6gDsXtBj4iV1i7CXiqcDbCL/N1oUNC0CUMY2jxG8
XFpplKMKlJwRLjBlWZzsRNWukA7LtpLDXEIGdkX+cnd8ATazYTbWASPE35vSTRu4
mVO/rrG4yxAaB5DkPRKwy9xYpUBrnlO+T3MeTWDUFX+OUARt9uhN1xalqguPim1W
h9NEkC3Bvys0R8zPNq0bgS1HHovQNkyRRb02m5ItwjeULNgoYdvhRGFVhTTZM7Jm
xkxU4q78uZfVI0PKpptwsPeO9NEyj+APFkWAyQJyy5pMMHjsK/fXeoA+gA+LAdu4
GnCpXAZUbQ6apT12GnPWrWWAl+Kf7pvyI2RouHzlgYtnl2K7WiBXBW2Mr6IGgd7K
P/qG/IEzuk+2uHtA3XW36TPkwU8NDECrGT7XnJXSGlRC/XgMekfKPcXS5KaYQWdb
Fk8X4Rpzwd+usgyZQxTd3V2MZvVTAd0+Jd5MG9y3zeK+/iphpZ25H1ELrWSyoyyE
V/B7b/skUq+RobSuEp35Ao8QMBSQOsv3l6bVwoyOHebtOF4Zvw+DW6+K/QjQOR0z
L1L+MCSd0gECMp+bEkag3hdHr6cm05k2ziUzWCnvrNow6FsVgaK83RmTpTLXIlkE
iAOX5Mhdqg+lP60CYGHos2ajO6tTYs7tjCGkMZJ9dl4KZxQOfevRoGFy5YwQs19N
PAMty2zSpcSRP8BTZ5tAqChLiVDDmqVeUNESckkAXQOelFY3viBsp0LRAHs/f7+K
ustaoDCbJf4zgDK9nYq6jcQAcAeumO98966b0HXEdwrwuLz0jsftTZFAIW90vHXj
x76nzj1/nrDD3vT5whUJfpL7h7+t2bU79wlLwFxKUJijHs/hMhRiNAn3fmQ6TJbB
X2VvvVM4ro+qVTL4SpvLVanWw91qYAXTBGvYNKB4nCsr9wxuPC4OXWAsHKKzYUxZ
2m0lBT+Pb7iIx/LMkXIQMINriPDgZljEFiGoqd1qHmb7CRGtO/DsK9j8d55PbgQA
BqCJyredPcrx2j0fGOi+XqHt9rZb4Pr79qvhhkMAsPr1Y69cJWYEj9kGIdlDvRFr
XBiRN1Up8Lwow1ANm/s/Fz462nYUbGPzs0HRk9uvYtqZ7HgSFt19Mxg0tehXVDv9
20OiOnzSeImEWa32ofuYLbVRWXonRDcUjGeqYCdygCznzeVvJoCF3i4qiT2rgGQO
Bur3XPKAmyBGJvi5zYdh980I5v1ERSlh5c5ge6riWs6gcBfNEo4yCHyXVZlsaKOJ
3IlNgeuB0NhTPNkaq5ta7hDYDosKRxpVU0LAcpzTbkVQEfZqjNd8wQUoxjQVXyqP
3D+/h5WsyRz8WKKFKf4kuIN0KNwNIk65rb0iflBgWl+6oX5z7TNuVcV7A8e5Ue1+
AmQiHQqJANl1VjgRJVqyIqRX25SIh4OyJ66kpKuMphWFoZhBW2VwPqOxCWdqfTss
IRRcTLTs9jxVz7/Tbb0lz/Yy+RzaNGHG/fh0yiEGBMM+Elufl0V1lbzmzmPvXozo
mymzAhT82Qx/PG7818P4qcF8A3+S9pbh1q9f0guj8d1bAgk8Ae3D20wjIeisgfzR
zm3sTn94BH2n/vfpcDQjFIMzdtkAtQp3iYEfO8NJCjlyRDZULCpB/mv6VT04d6+F
OfOfCfO22ek+nngy3mFcLcBMucRVE+O7gL1aoHC+vsQQ9EI/lFu+iKnJ/EpKmDmo
gQGgkCeC/o4huZh0rse2Y+94Q7ktq6DBOZrrGXzK5IDOiHE8ekG9AuR/gtF/VJzS
IFD4wVVJGJhS5b6Pzo7IRYb+C+B3c5LmTUJ8BFQR49FTiA9alPyPdnr8wzpxJXXD
xwSVKLT7vSRun20kbgNfD4zYqTaOh0m3XE/WuPu5BML0vg9ImJnHN1ST9+iRBRhP
5uFDUlUoaeK8nq7XrS2l+026G8+ZneHFOlbB1Hf+Kt1XZh3jzPUcnOirT4xnKfdb
9pxyy2xRAFp9jkxe7OtgFSpvnPkPoLm5NONFu14CklPw8+Ee0tf0S0I6nmxiigMQ
CdpvnGY/g6HJyp8F7KM4Lj0UM+g9T0OVJxTGyRsue4kaxGVUiD1z4UMcGDhNGuJ2
neht3gwjOXVe1VQ3TGO7UoSjWl/1unqZfK+FhNqMt4MXEpsQZ7aWZUPSalq5cWer
umULkiVCr3o9POQxbyAhd6V2Q9zy5bzFN9zz9QMUwvWAyIws9ZCwsGMMojTKweDb
lF2rXru3fNFdUYGkbah7DNCbKDSuoloFTAdbCxmn2+1jWn1xX6+K6duezr9tnOv0
3vLwexKofz9sXsFvtgByxmxGC3PMT7OTgpPJTq3PaJ/vmzboL104uni337TNnA6Y
qA+4wjulEZj2gVX7ZvOnqHTL1VuNQil9anzsMGww5bVKiUCAKpyQx161YIRvY2b7
R7Bx9v4nAB/i6r+ZDZoAUa4ukTgHwPWHZw3vckfMyGLjtitMUQkQOa898KKvFKVz
McrXNINmiRnThS6L7rxWR/WpyaE0N+BLDElWzcMGzFuCEvOnczlKDpX9sSVSgHob
1O6DdVrzr62ujkt8KRMNVh1tUGU/SMgoYiEs0+2e26rnCJaAjCsdufqHuGKLoY35
6QYJF9tDvwUc52fNVJybnmAvdAKSiO9IWjM6ClWK5qUIv5hlE2XeQalrzNWLJFUL
BQT/F7cWc9/82tJ44IuoBXSPBgBaQvxPnRnIGlsdUGZQnus69/7LJqQ3umt4E/hK
PU/D95rIPiYf8lAPdUKZzeGcoAAFnq+2k3+qxE6iuUtSAKUz9ixKOvvmVJ2rTw5w
4w4aZA5dBkT2ffCrSJ2PiDg4sydEcc4isKSieMVqOAe0hdisXob7CFFXBaBTuc1p
Dm1bGo+vMR13VgVuFYECjXCXjYWPgySPAh0oblJEvg3Ew3HlFqypKbDdXFeD6CZK
xuOxiv5lGubobbCOdNwK1sBSuoSFCodbx4SCeodHPYRC5WCVmFeFG3a2ykFgXFG3
u1OIkm5ypXBriBAUbEW67W2YqXfELSkFNnF27EPWfjZ87JWh/OhG3pjjRJy/IHdO
/K//J/S2D5vpyjIw/OQKrDZpLg8K4k1+NyfKRiwbyf05jS+ilXkQn2AZNrzkuJ0q
pojedkzJArQWZS1shbBXhKDqd1Iq2uDd7aDIkhz8DhdhQNr8J/YULj02/FmRyBw3
l/fCs6Qqu1uIp5piFEsjERoW8cexj1xMfvioqd1yTP7Jp+koJJm//Su45n2loLRo
2+8I9+saGvFhjPKQ9XRo/PLxO3EK1HYgaRvrctd6PD/lYdDT8Nmzu7ew9DfwRN5A
mpk/8uofANJRKKqJejy2TUaL+wEJORI1MXkwUNcf9jd3UGF4QoNNv9XODLZLmHl1
rqqRIuXmh84iyeDwnYbaVLNfS3mV5WORzGBBKtZ0EjazMBvuUXOaIM2y9dv0EDrT
FfI37vJx/tlqhyIVGTGAPrqSmY5vXk9uz/jv8c+lMkfajC0/nPe4nKkpSM/h5BQG
x7ltkOyKnyZPInSc2OTTxVpSX8+Jbp22xx7pNHMgrrqhYV25LiiFrrt5sU9pO6I6
bEk4/QFUZy05B7UIbd0QlcfAu+WCugO41SJ4e4X5RtMDa4MtuP78mGwpSwh7fCFa
JO/AoYPBQ1ZjC1VhVEurMx6mXXa+WQeV1izBW7QkUeVMt+B1e0xQij93UVR/E3tA
vf5t827SaPuKVyjh7uodr69RpBENu6X8z9rEYO0laW7+2scaPUPCEpZihu+R3WlF
+dyf9uEVh6rmsugDB4y4J9LIUxzuIQ1r0F+yRnIDEMukk4+V4mssrm+Eqix2ukpR
cquiimi6xfQvT3yRsxVAY4biIK6fXUFINCTqLwUyZNfeJftNtXwvvs4SduvpBfZf
OYo+8dguAKwpeupjPc77bAyqOEpJNjZrLF5GNDDjTXqwtCS/Hrec0RriR5z5tNJZ
hAna99fdWBvu6CSmptw3swbofiU1yPTJzWpkp90sdv3dsz0JxFjlcZr2PWyMO+rt
TBtyBMjs6CliGtcWoaWL3pe8hviGT/ga35gNyAA47Dfw393TbXFKJoDK+jApmj1v
dGL+Bz+ECHGLvuYeoGYuAkp/OOKEt5lIu5Drx0LegW7iiXCGP5RvBusBcqdHBpmK
SKeR1nNL/Q7XvhseGAFpja68d99hzrIVd1RbwhyY9hqySedde5u0CjV1WZEDm1zY
+AEH5W31uKVU1bqSbIgTa2/JD7vKAfVgCJWKir/zDDemNMsRuiimuhF4M9FD5ubI
Co7cQ0NlpZklLTUY4KYWoGVwc7iS7XV2CEGEfmPdbXyzfIQAe/jAOxcZXWGxjOTx
SmkYC/G3HrduVmkO9yxe2ZHmrFabweuJSAzbaS5Fh2Sb2D8Vk/hHWVthJ4EgrOam
NOUndFEjN2DcORg/a3xvute/Fg3Vnx1BzpRPxBrc0ePwreIqxJar7QRVHwuLC3f2
gh+DqWddH3v1ML2UW76wXs0uRTs5SVXyV9DNyVr/DSHUyEQfiIOgWpwdKhFjTyRU
BE9TAzZGJBxEL3iKbbhNqbNoNMqNX2FmuSyLzfPYUNlxtcNEcN5JHt3TanVz/7kr
CbR2vVaDAnuYeSOqzuWaMWItplVSAnOUkHvhKexst8PfG2NHhcXvyX79XiWX7lkA
lWVJBMVWFCeSehRJXWCLNfIjrZORjyigTEP/cuP4u5h7Zodhcla6OSHzb/RSad/n
UUgsF/DBUvSBkaBly0vGWZuPtx8lZc1aO3v+K7j1g5cN8N+bakLyjU+qlnPNmBVK
WSYo8JFqW7al24tAMoyocBpL1A/WCkbgj8POAqQHM2LErQ0xY25VlvhhXy9aK/OU
tOhQVxO1rtmi0BoutcnooxcCRRHDDnGZw6Kl8SbmRG2Y5bxARvPlPXcl3orJ0i/A
bYWWKmHpm7dYU/FTzcBY4iLK6rhW+pyBZ85X9bL3AhVfrPHQHLz/52Xa6/tuutnw
jgVcvc6Vga20tbqYLhY9mE/D3Mb2GbxL5cBs9iBtwUwS7YJrZiH3KTzhC9gtjtgL
B0dE6r0pQdIBGZu9aVVNBU2rSxp3VQPFljtoZon3g5KMQXNC8q+Kob8EZ9f+eWj4
M5LD4VLTH07hmbMnP2pf8R/GxR8ROMVG/skcxziCVgORYdLx8QuZdw8YmpQYt2LV
zw8WfwxcEXeZ+z32qIgnbQs0ze35d2nE4swlHp6UY4yNWvbM/Ov3oM5QGRxRclaE
pxqRStHd8PFvwqbSyTXV9393wyX4bdMolrZ6R/dSu6prqBDgardtCEhFxvSMP2lJ
m1BQMzXCKdujC5UB3hwLLhqJJLR9Ka3HO2eI8UlOafABos6fzkhvKF1yLBtcrHSR
AX6dI3wFf2lpVI36CE7kU7QjFl+bufWH1oMLskoYry1HRAVlyMyf6biGE7GtoTwi
XKsk7gIoVYsdw5UFJHX7iL+Y18oWBE4YQSp7tsTUjMM1ysNx9TL1L51GcU5vMkyi
MTtv1v5n/Zqay7i/7Xo7MCmv8Pf1MV3F2IkkNKmxBEhlasYhDzx0vmrhOfcSO4pM
u12DnzVN6fxCIbbgfRdBO86VVx7OYTiUp1JhxSKJ9UATZWJeK2Tsd5BUjgiwetcp
LiE1+fYwQQj1OHVqHli9Kg07NaMdbyqNgGLki8eLOuKz6vSDUzwZyeNtVhTM26XR
ei7A7j3zUoqrT29AHTXHHF8VWpIBi7V1tBs/iJuvmcYaTrBZP0lTA7hVZaQsmtnb
2VPGUGuROWhuv2fH5HeClJOBpr+3JJSnTRj7K+6cXhfjcgU9mpbTS+C3/PQU2a3d
0HPw9EssPQRKOLFYjFaO0DkWqyD9210CugE3zpJxFtxcqssJGQmvl9IQ2YjJOKTJ
1BmbQDnNrn1p5yGUfVirnrc3VW/fj0EEAtcIG352MdlmWZsqKLGeGYumrrW4o5rJ
IDwdXsFz5nsxs1JiR1q349gqWNPQrHyWQObDlcbKgZQXZpVebs3ZBMV5WS7BQ0go
IEn/iMkfWlBbc/gE+a1zszskiXW38Fxr9MQLOenGNfuOpvxouK3Nds2SrLB8czeX
xieopllKhmwUkvcp5n81XD46xbqZEU839q6+9fQsf1FsJlhuz+DpdaVNOQl9AbxJ
L0xpnePyCtXa861EX1kG0VsX2HyupZYPwsq138rwtAThy+HwN7qZWrtDk+9Hhdmq
foUlg78N1ohcobeGWiWTWIWqBje8c9JreVQaQv3KiF3ZTu+wws4u0tlBhjzl1B4e
w3fV1HPk3TGZyi7edre+MBUDbHtTrh14emdz3rw4R7ERMnMoxU5VTap3Yp7Z9Sld
xCQc/1lR14B8YA94nwBCgk/ojLg40PtXN77KUczaigGeLJVPB4v7w6F5Gezaro32
z8ko1RXrzrgjLL/gr3uj8nT7D3fzyK0T8WJwqMfs33cH/cn2LstauUToPTgqa8Pj
YZV0oVLDRSF/jyqByiAq6ZTpv+BiRibM8FewjM9Grdd1Dsfh8hKlphBoIVjP6eRb
Zxh+uweS9CnAuyA4LW+auHWe15gV7VsYKNJ7WD65WiiOAcXl596g2WKZUcN+8HFI
AzqMmV3oCOctV6zV39HescR+u9OnvLvBMBXC98X4NUnbQGdX0iasOOSwXrdh+FBd
nb1ZBEY+lTsskYDKQWkC0nPQp0XkifnT0Rxj8yQ8Rn2nMI35msj5/LRjZACWDSaL
EvcCdHd5X53sS2f80JHu0a7Orjt1VEVitVNMUIQlM6YND5xfVbiIdxOPpDFqV5IV
jJMzRa90Tuh4ddlQEwegXpyO/7IM7YeTgX4Op+sYwfXzEzhryY9s9QN8UNGQL4CM
8OgJzcK7N7/WKc2JjDsSKYnzP7wupglOxRQK9VcitWUkHDCcjlYOcWPqp6g8csQ3
HinunFMqjTEE0FW18BvKTGuYXzrJNNU4n8VDqZeO8JKhPkPe3pBvU5KjEx5s/mxH
ZWf5hBF/HHEEFiL0ys58xrih9GKjP598yro3yAe9z+g4jzcLPKl82SPWE04VsacF
ZzmlnQpOcb78JqcLnDom0zhIpvP5AuOSi0EraUMVOZ6p2Dhdfj3IcVWhk1lNpAJu
5qZyG5oeS+VUOtmO1faMtN2Lfdi8h+RPP7rX7dVwcD75WyoOdwjR6HdpZ3LfqSxu
LU00shLvIQ+gc4weZObXmYZ0pUwR0iH7CY7Le+bgWDHH32BtpZUjKCM4RWY2VFZv
eBa734aXwkoS/6yuWwurtsBmGO7LXtxE4YGW8hoNQHxcgybwaMsJ7mc7jNXwmfu2
w/PfRkP6X7s5B9j8f2lu6IDb5RXVYJIkjQBMRTN4Q7PomMIDjR9w31x8Qxis7JJd
5vjLfPh9tKcweJLlOVYPpc8yS+slSTKW1jocOJXlm7zHx6AS+qUrAZS+XoJWX1oh
2dXhNFFtrKLLpmMzwa1OswpZqNagzaJB56uaq5CB804/FxeLN5MrHQ2Abot6lUG8
N6hjjzYKWAAZBN16jDVVtPvfktJt9BbObTs3nYDJYr2LM2/0l/ZYa5px14QggiBM
5T05Gz8rX/dYEdqMscsre4RsP8Fhe+FLgvdxCENCotf+7A6XkfPggep1SwjjaNfL
kTyx3fUmM7L5Fxf3TWzguvsJL1Iw/iDcXpPzdcX6M6rjEV+qqSQ13fuJ7lpoSqoZ
+rhtOuPTneMoX2YPpkn0TTz6yFBNGKJCCK1MynZtsqbeYTGFz0n7Cdf2jylKbGLY
krD/6bZDwg/tMHGONh2su9g5rfm4keY9JaEHaBRO6ebSTje/0qXicbuWLLO4JCli
bGqoG1eiZwl8JeYFoO37DUoc8SsNuzjn00Pltv0pCtmHT0GUFa/Pzqf+ZQLF4ZAi
FE4GfjzaUr6QiMP0C03jf0GvEjgBuKSKZ9d2MBmpkF562nH9ArjSVg6wFQVQU2Hp
kQAHYKG9hY6NctARpyw/DB53KQUojQlynsr2hFtiuircTQLj/fEmpczN9ZBDZNp6
KiNy8DfIj+7z23cf4AbZEXIX5c+PHnD6/OrPtrNSWT7UcRb5mN6wypI+wJXhvU9a
pePy3brtTP9yeI+70YuOKAm4/ou6Sur75Nnq29Je9aXA3K2+CnDPlM5Tk6ER2lOK
iQEG/LbdV6Ohmh/XbpyJyLkIcPtlSlUyixwcBNEtrUtimKCmdXLTyGyS5bl4NTNR
KUlqV2d9QI6bGpTKlVBvdhlQPK54CrdqIexPM46gzh7WCF9J9z3+iyC22ZioJhSM
dsUp9430a830XRAtmHz2Fn34ZqQLx3a9tQcUA/spU7AUJylSLHpZ4l8MrhHHSK+Z
iwqituIWtp7q4qM7rUHrry0MIn6pbB0I7Nl19dwtxIbq45ixr5KlFzvvQCee05XI
8au9xfzEKsYiBSqTs2Cwwf3HxqE2hkraWMaK44z+DogW67fUh+oG1DcOd+QrrTyZ
mBe6td85lsnQXlFc+1Wqe+0iywBxSSs3k10Bzc6EYvdxx1b3WPpiJPn0ZTD6yABl
iw4vt8o3T8uTnTPo0U007ZsAcNgbuemLs2z1VdUSGLYolbOJPVZ8EfetaANCK05s
yLdHCQFiNs3c9rk1Ym3w8Hp4v75Uj8XUR6VPE7Okjeiar1IXY2KSEi/c7GKTyL2M
msjaTWTRlIsxrOtbKvDeiBg0UvqUtO1EdkprGEhtP11DYfqkegXHnWVQfPnmuDpE
s/1AvhojqR+tyVhpsaj641hXlgaF44tkVaq+HO805NiOrAwZB7+Hqr5fOh4/itOP
SPuVg9mBINaf7dbAw2GMW5DbUCF01sptH1obPzOAP7rXoPGgE1GAYHp1f7dEwTjU
IgRVNQdXoqtnQgFg2zQr3rjj7oRXRs9nocsx1hUVCqQnptYVBqFoDXIWVW4/IcmX
meyY9ExarymJfxnV+TRxc2ZoILqqjOkq34/KcsM5ikit2oDDYYNYA5rj8x1GRdqx
I3UCRbYCOXCweubLWmojpx9QcDLoIyvZ/z8mXjIc4PGvo8P8vOfkTpPRGZ1HRXJv
iwlLS4OmuFWSOdhEUCezDIYWpJvQ5QCL5aZi3LVvKzgRpLXeqEhtNJg2xanbo+4F
TgknP7zP+DqDAJy8i+iRc3EB9u0RJAk/myIQwnv8q2jZmdYCMPfNz/oA3Xp8Z5Ia
Q/eGDJaL+5YSweWYZVBjM7bJN9LcTADS8T35KOFPMDActnDyKruOCkY31ejUQFI5
Jqhb5bklM9SSaiyBhR5nCY3kWhvHYUgA3Dp+p6O5eKPqvPR1l6t+jAeOd9bSrOHF
Uf2o7tGCg+ZyiKM5uAP4sLHDfOA1rVg1yO24h6dxaxQOoKnedwfIBar1Rp2A4zw0
x07hAyVnzc2EpmdYQW4ZgoL75Z9bBlJgLA/eD4ceUyHn8KplGTooV9FKSNxxoTB5
zGCmnOSgI3Mlub+E0D24AQqKXmW8ostdlTkOeEOQ6wJ6NOzx2NouPXUIJO31oK/n
tNBX1rGTISWea4zBLImvw4mfstTSYS4sDyZdE7O47xOgRllsxNMHNkm7J7Yhk5+/
arlYX+rl1pSIdSKYQTq8PWJg7JKXrjYxC5w529Cqxn+yyx1iiH+yXUcntDzqc+FK
WgHTVyWnzUTXNStThmVMmLyNVCC3DxJejMmkhykocribcLv+SuLFuXTZJn/Yg1P0
h0tFyl67Y9iY3X0VpUNIletSqNChQ/ROh+XJG5gfWgVT7MiTs1XyoKfJySqs09dw
t14aeAQtn6TD1YWIUk9ik1Hm+b7hoEIyxhxovlbe4s1vKTHH8H5VP9p9c20caNuG
c6+GCuKlq4gpKuA0Te6wJrD4kRaaxuAQGAdlejom32PlTB4YGuz0M/El7zt84SJM
iCAvTSjIV/3CfIlsqQyiZaDmkIz5ZaKicKbePTqFFD5+NQYsGWsEzKPYAZLEuuO8
+qkWRvA54H1+P078bSxSbZdNi4/eIHy2L1sVcwhTzOWvnxcaE5OS6peR+RceqmRG
jVl9+BuaWx+G7ApTQwUEpzVUnXuLtijh2XgXhEHJLZijh4QO60xhlAPzj5ZUOYEc
64lOnoMpzFlw+splau6Szmkb6UurDB9y6tabeNzIPriZ/9b5Gyor/DwjVdsbmSLX
K9pGpNaVT9R6NtEbtJqfGCj9bSpn7EbDwoe3zmrywBJ8h1rzzf5IMVn8DP1AwqNv
Nvepomq/MkAjhEsFFf2Udd/aQvdNT+E0YfOGTRwklDjbG8GzUUOVCXR/A+YWxrsi
h6U4RdHS631L1heOCKsCaTcsUvH0olTBA59fLUXj1aN0iwPDfAXnE6KC4NhvvyIL
MtlpEzl1eKZxMQHD/11t6Zvf/FulSY9xaW408oomAoXYInTmHRCFuIfSAVgYjTHZ
RhZNf0O5tLcHU7c079WqlaZJxfgqDWhnF6Ro0ejCXa6Lj6C55CFefnkvL3/53DKa
GghF6Th2PVYj7+sAQMQkhSmtt3+kG4Lx/uGuswSVNUtmjoGoK4ixNRumOGHZv4e1
wf4uzDTYstrJdlnyfsEWPM2MK+dDvtTyoPOcXHNRnfaW+/5qedSCXNYCenfB4I6u
0GJJ5zz68ct403cGTMY5TvhaP+gvfUtgTaCQzMMWbAfZu3JIwBVk4Pg9EH+HxPAi
UPNMKp69+DCd2zuWz7VDtYP6GBupBydLGZ/iS3DEVzNn93tU/4203XRWVwgt8c3X
ckfKlWPYy7vPMSYyBYvYVfziOVfwP4VKRL/F+hzc+MRLJ0Q19OiXwL3Q5Lpg2uJf
e8hzpegEcoFy4T+JuDhg5H0iyRD2ilJRuVNvVOIu+IGcR7LH+SPiiUn1nUXOVine
jn/ZwBgUP/LoPwXdJFvpMgCoqH+WNGHsrngQSl18bf69T5YB5Maj28UxNo/Ag2ZI
x5h454hqW3YUPVH/exAOcuRS+d46TrMzfMlixDELBihf9Mr9ZEqRY4MQ+c/tXmsH
SK0AAVPrLQc9tuJnQ9Evel2Q3SmNd175NtUUNp9ro/4zMFz3igBxyCPBru+JanEQ
80YaYKou6rhknEwPqKpWPXgqJ2ga0tq1AUF710kFoZdeblrLh7seFKL3L0bEAvfw
q6AmdnN0Kurp0e+bJPDZaHVzgAcMxZUv2oobPYk5UpKNpXyRe6CbCKe8lU0yj9y+
CdlOdgs6LukDKmhOvXiBiDkmRmBvJIMmmFxx1/mkERS6M+5IbeAe1c62rigNAz3C
OIaI36Neps8LZRzQk6SziJbQ0lXD+MyhFlyYYPg84zyzvfzFGZT3rKJF/zTwE4mD
tBDBm7gwwf34zNd+isM3OpYbuNeDYoIp3vyd/qoYe+D4BhG6G6HuAxtAFLZJ+mZg
+GTRjbOPcTphv/IocSzXOX9L5B63iF0Gku9p2PMmAvNWzOKGkwerAAKDGDLh2jx8
/tJOgsFGJXsN9ciASBmnBzkx07JmlaEOEShbTyYfDoC5hX9puZFPk7x/YdtKcQSo
qCfDyFGBXP033Obf9r/zmV+OBrrI6XxlqGPKITRSwtAdKT3CBdnO/UZRrAmVF+eW
wLkh/DANo1oHxEjB5nGyeMMX5BSkkhkuT7zZwTQWKfKtz36QWKrihB1XaQNmfC4M
3kIpUQLbusDUdFb0hUR7ij8yeBNMMf41Byl5kkgG7rKL8hUlH2HQ7M81EDriSErU
fef9j3+hqoiZpYdz+z60DaOtHcuiOZ6L54exXhFhX5d6oFWJPuPm+x9u4XJaERnq
Y0zpTRgYVHh6rx7diWUtdpDpnGry5shB2CWcJQOt5UDnN9aGelQU4DOI7dWF/uoV
T+fWcyfTxivs8FFc7frSRTY3S0cDsOXiPcMveOnPhmtgG1fuXq53nm9QUaWoDD85
Cr4afgDP9JYMYKrsYhxlO6UvyyGM5m34w3x0xaW1bcfvfZC4uvWtTviERPCfXt4Q
hiaoV3vWKJkyWVbhHiSLJFhkAbuPsD879imTA62yc4JVxXg5/p2dl+RqrJAkFKkx
XroJl2ct7JcqIo5USrNxWz3WYw71TZ2aQKP/m//JXg5PIxBHLgEXG99ovqf8hn6n
Te2ohC5ETxmcgjxWE45fFADbwb/N9HRG6l9J0FH+54MDfZJ0w+JIkR0W5hvgF2Zl
4ss9MXylFimYlKiQxxb3Onsr3A+qG9noq7n3LEIcAkKqiMYzhc9bZ3vGpobFQwk2
Fn2oyvxTP/PYAMze48SYCiv681TJucTpM5VAcllXUwmJzfq5xIHnK5oHg/3cq22P
Hm3qU94kklGnRVHFtD6BDiddegDr5xwM2I8eVeRkwNcRTv8Z1gu2JorHc3l4Cq3v
0aUr+V3FmacKoZ6JgB6Izfa05sW6ObSdpal3WrP15weLMhFYp1bCSeJuhwFu8cUh
iUXIOpVAq7YccRPd2CR0fYZ5priavhAvGLyphAGqg65lfieMu9sAhuILFZLolSoK
YyBiJ34RBHel46P1C7mvvNF6Dj2jrPQm+YXBDfcB49C36Vb9XaIOHZjSlKYTZt4B
kQcAVG7f4vCgNrU9RQAFycvScsSj2vWsAcPRer26MK/+LXDwFgMQNOW1UfLKDWTJ
W/W2idbqeV21I0aIQjMF0sx2PoiJ+UDIVXNIhZUUKzvv3qBB3d2O4SfYYAHzyNJa
kQbd3xHGRNXo07w1Eiv2ky+3PjNi0C5Xso0/AlkbI8fxFa/0Jvb+kzSV3y/M8lnX
nAFEdeoDq5kW435HCEapKb66k9bfU5pqvB6uwQOYzgAvZHwlGvF8+l2IwxwPjN6t
v6phFLaZbjd6830dYFYsX0GgviBtS/OLVuuPcZbtNWJpGVHXNV2Ut3KbyPQWK820
GafMTTHBdWaN8lBj3n4kn1pPrgUjNewg+VWpMJKTLeuNS6n5LARez5t8WvnpnvFi
jQPDkw7qJjLt9WF7WKZunh1rOJFq9FGhnuX5yDCenf77cKtemhMQ4OmYg1VMEh/g
fPdpeWlohNKSXeI+BgQRK49EtfvdWD3+z9JungoF4/Pu/Ce1EmZ/DPAn71jnT7Vi
GCRXuMdd8zoOelkprs913Cx6SgwKpp1xr/fbEeyQ5bsQRqulE+/fJ/EvxRZPyP74
DBTSmZhfMs1D8rlJc1WH1dg/38dCMhVhtOElAam9G47JG7sDEe8XHg8/4EqZ37wi
R7GKAiUd27+JspG1Ec5HbSxKpKT+CyW23roNtbAenn9FqoEhoJf5Gf7DaLsoysQL
t0Uo8VM6UFNuSpMGSVlvXMow/+Z/LBP9vrWryzlT8/w9IMMe/3D1aTVVMLiPMMK3
uhRMWP4jhOmej6zrAwS8oxqP/ZAjDwV6HIT5Y+sbnQ7ATKVmjWK0eXeLGu/NvGGR
cbUogzB7Bb4RwarYm3cwTdoNJ3bgvymhwuU8jSrn5875Ee0SlQNTAa1rIG9skyKY
XAM/hQZIOqnlceFIwbGdRobfhDAZ7UqDcZCYQDsUX/uSrp81xA15cjZXAB5jKd3X
lRl82kS1WqPXk8fdHMxljNetGxeu0m00ErS3QRUJ24h/Rdw1qAS/6Og3/an0exIz
n3sPOwz5Izzl22wnRLukNYqL9J7J62qyzWRpeNbXFHAQzpxY/MMnsiJnXId38/mj
Ns2ZXCBosCTG+mqW62fz96apxB0TWLeAlqyhmtsZqsgF5WlIDjmGk1Q+ww/Qy9uu
sL7jWwrijMLGov4H8ARzYa35r2HC34A4dllJbSyK7XrKyUK8jpEkDEtZV1y/x6oA
Tnn7vgzDrwiM8RxwplbEZbQA2g87tQtxp1+GRW8yJ1yXTTiU8d31Hf9Vmb6pccjj
WvoAVAsZWigkAmf/H+n2L+r/e8FOcJAYHqOniNvt1socwXkUS8pInX7I3w+8WK10
T/oiLLmKAJCnW5WISeyHh9BoAGEXPmXqivWWfcCQEMxZlQeICN5GMXnQ1T2bS9fM
SHZHnjs0JX8Rog8kv4aNArmFrGFhkT6BGjVqwbODpDBGseIUu4fnoUwi1kTT1ZfY
CN6H5+I6ZQmA/RedApkhvp9K34t2GWBdRtXIz52dXxBKTyvxZYC15wdkuksyXUWT
rdMaKo2ntFSKcuZbF0L+W/Vjo5xGEm2YjlO51WM9Sg6GWBFJ+KBVrvXdcBs30OMf
MCEG9jgBDBGVaF7TVkp0yV4x3xImLxpwzfBu/HM5G+RllOi8eoamDe29gMzzHF+U
BOkZdUhc4TiHGx6//jhqgUMwmWhqxg/ghk3wClvyh2OJddBaGS4+VgF0P5uWSoVC
8Bmvx8Vuah1kGYJc6iG8+KrWG00XJR4HR5bTzk+BIPIwTlGrp7pdTCO3AcLA2BPp
x7GYTlg3eg78n9yZBEPXYBYNfDSvnK31W9BCbpw83bngEyBaA3pBpseT+sDAljIQ
x0fcB/CdFk0zlZdMBX1GSB1P6M0SeOgjGGi3jy6T+PwgomCGfe2KR+Qtp16xC9B1
b8Yfq4aPyhFDDQgmhNbe3IBfxDBwxbS6oFpJ7pF6v8o2L5r1H+A65/rxOJzyKARj
+/iCOJiN4rooxqrazNZrrnv1PBy9eUyxaKhuLKLSirOsO9CDW3p8X59hSy4X7qvS
eExrWbkDBvXSx1RhtNNBdw0CwW3/N9dG6sDbDugqIexCgiN+NIl/ClZcQ8RC8g/z
pnYhg+fjtqioF2A6sfxeGtfbAuqCn29v7HQ3hBV9pPAwGP9meKb7hdmaQLEFItzG
oxjBLzFW7fpY+wmkXaBdD9dBMwkwx32JlmFACUMPDweTe9ynV5vXC+fN0eOoD2mM
m6MR+y5AM1lefp0KaiZ4dOB3k1dQMFdEy3I+0YsMG6sDUqWhVcLIM19OjoCJQ5Nk
QXVCjHIEZ3Ho3FwLcHbZxX8Ji73LlJRkiA0z60K1NGH3j8vHmPOvA0j2UQ59pqAV
koF31KzHO2aPn0koUWwZW3xAoeittdH0gH9T/vrCIqkMxCDsBtEUCPGPpIWAOsNP
4vK9r1L9VhL28YJR5Io7EJLJUpuBi0PyRlrEsom7GeiCwh2jGE/ldqNHiyvJHmDg
Tlt+E6WLP2XiQAIrh9aTZW5UIRmvMDSXSOjS8pZIM3/Wlg6qHwPM9P9bPCOruRmg
BknLo+zsHBD1AXymWQC87nGJkmSTUDfMzlrNV3BpMJxH/PSsZ+2U69kRLcJDqw2C
chE4A6fijUC/gamiGgF54oHiNDbFeAIYOYxctShBxXUW1HbAMgQCBLy+Rvec9G3g
+WoAnTBwrtuLZX9AzYT0+MOpjVEhYANM9X7V2dNSn+A/VE1jWuh9CFkgo581R4w8
BMa2eG3goprRWFd+Gkm8ltogurY9b2e+Es++WwBgHKqq0ZZgN+S8x5e9P+owOL4j
Use+3VR7o4MOVRBXQ2FEDD8QL19uR5MZ2pdhhp09D2LtUx3MPWMx2vtNR+P/Bloz
UfkZXfsoUWdRrG3hGPec9FKuJYofFxoHcDyFtNnpaunbhAdUDH4wc5Vy+IVta8hG
ZiwpNfE5/nWkPpZtYRVn5iWmkcbDxklJWatnGEywNJ8poLUkHIJpkAUQlDIeOlXe
Bs95Zw8LO7xixmJFNKKv34gjBEraoCc++Zktb4efOHrzEcplXhLDrHxuHzx2iLVa
C6iVV8qBQ1jFLu4hMa14JuxonVFtHkiYsMFJHTg2X/zv4mlfQHQVVwbiNhfGZFdD
LBlJ6RjmpNbDcknyP5E0YqJQZL/oshUQu7UcaqCjEYISQKdnjNnrdHGCr20IcMG/
goD7+lZoyu7+BybcHGucMm/vUTowZ++k7rsL3QtSp5d9EL7T7CD8uwOBiMOrOSCZ
YvQ9dVYXRCD9ILM1leHX0KyVvpYJemilDnFcPp/GtNpw/OFDn++EeOBLGT+eowpN
qPgEn3bnvW2qDJO1B+PiHXjzeLEoLKgoHDtVGnaT8MicebqvxlEV5+I8/tR4P8PX
MH/Ejk3Quz5fWAg2Qs08UmCqi8CjZCoc/OrxlQZsCK7cAYb6MPPGs1cOYjhSOOiv
4cWpZz2ChcrBo2LLv7BXaWjz3k/10NyLJ1+S6WMgIWVfGLdcvul7bEKBI6v6nogK
F1UfjFUh80g2m7Xdcy+i30KAnITc2ygLPUziHH78Ntfil2N++ZwHBmrND8vRYslH
LR/tcB5YCcHf2nwCRAt3X+/seH3MqUylDwdjCLuI8aD3lDc0M0bHGU/imO+gJQpn
Urh54tQwTcQIP80/19wMCVFcyjr7Uhx0PgrjTxfWw6HjZKk73nSxPI4dtg9pthkX
cXCdmbRnsTGjfyulpjamOmNHUQPDZ8zqMFTMOuchMTSWqveYapUuqutaoKDnpTnC
6ISzl+KeOjRJugc6jgTfYnlVl2BPjocFLiIVwn9ary8xDXW8Oev5kPoyX8hRMh1j
08SHhiiRjX0txvSanxwjFimmTeXdK0i3C1gRegJVxy7aaNah2oKMDcQAvClS7pHm
dkZgQwTxOshN6xWGhCzF7dtUase8/njps/btRSxyJ3FV42f7wvVF29iBR5XdIaCX
zLtAvdoD17iLD1NsMH0foqhai7154lchcc63OU0UrxaBMHDbPnM8GwEluhHROBsc
UFy+31m8cRJ9j9oQYrsQlQxUuy177KSZ4joe8z0BYw8NiMi/Dmk5QUZ9vjXXjd9o
474aTIHBOJKKKkWIbgmV8a/q6aRndqoq9dt9w9yc8/oxUNVkkCIJq5FLBAQNzVuj
lt5oe9wK9PGMG4xxN9Q/L9y3KyZxHEX/pW9MED8a00rsBf1nUL1gLMSVg0iRfhMv
rPoIbjpIoW+z8IpMfnzjQBdMvVvMntFo8ltyoL0vDiIecEyuGk83QOrJhpWbWyKm
Mm+tIVJYJWuYWYDOBcI2ZsF8lMp+2Tgw4+00qtFBJoszYeIIj8n/YLDQT3klgSA+
77MX9dmyOonT6hKrB2ZZa2yGQ7HvnZ1EzL6gH0dvgtRlieWqHjAMH/jTmuR5FlTv
ITXOwIqf5CrIr9lxN65YlcjyzoHNItF3NXV+3rs6uhnBQFDRHIr0o/roisfGsQ4F
aUlQf8eoOJYV7GSGdZ5I/kB8W+AMJ/qTZGsjnHZiYVu0MKcjaQPs06pBi9Pgi+3w
Kw5CXhXN8sI06jRry5FZDqRwogn8lWOXfiXhfqmLQkEHcafLSSvKzRv9JPxs4dA1
8TcjrXwtpAXA5nQFAjXGbbl8grh4qDOpK6F8uSE5ePB7UtL1QMBPAx5FQOC7Y3mW
42eTaNo1FDt+BbNPW9ilWo/2p0SIgChIOpfZeEwaf44AS5KuNm/KGck4BF0BhqCO
/U77KZPrJhF+N7CHWBI5JoTiPx7DkwNT+HGETgx/YZWzJwviAAvQkwjnjOkHnhSD
o6kmAmpZhPVGOLAUmDvSTU0/HlRl/QPhxFhy9UCrGmLX0Apy2MIuwyQwo2QHZX1P
E7xwMCYOwVg/toITT1BHtMh/swG84VLJsJAGpZYoaDFda4+vCNaEP1jcqXLVEEKA
MgBXfqyAplWYGxJ14aEoqPcPoM98VG+yJZzZ0ExfHZv1LZrZtUjL6PNkkQ8A5Vb+
6gKopHfRUN3z4UQyxNjLmrp0JXfeQ/DM8pCinm1sDK4nUCKlp4ni1511siHK9xWI
O1RjWjU1AOIbVZS/HJafGwx/m1akoTtUkIvpT74Xi/I92LqMIQsksHp2vSuL+kJV
9Vfv4OKSedIFZOSbuZcZBQVvAb2gsQ7dIp/Dx9K+73Iv4g/h1Hcv+K2hCI0vtGmx
ksiHpHiuDlMtz1EaKK5s/EC3mPKcuQnSGW2NCUOLPV1eUoAfgGlfb91FTGes1tkP
HhnYNvdWBp4ZmFB6kDbHuAanxuJ0xNY3q/jp/V4S38GqhQOuphZmDeN9ERgzNfaR
fBdNBAQMpMeG8CgHet5lInxN4fgxzE8DwB+SkDKvaI9WrWoZg0gsi02Hn+dsU6GH
xMFD8a5rqDLmqicaljwJvK2Dzq4bYjv6K/fTY2g5hvmL6I0KnGSrxxl9i8XMpoNR
KMiDEF7tQg8D5u17gAAUuMy3+4pqRaqzp1ta6JTZI3RliEr2it2nR6EaFiPpIfly
oOQj74IEFKoQw1vgSqXBrzvHKuU1AnUTZPW3gBHzM5wACihJay+x7qfoWYMFhfA1
7DKbHu3ZvhxORiybrGZdDi2rw01jdTqJSU45u5rlMtDfOT5ZM9PfbSOV6clxQPuS
gPjkijLbWOKnLQna7O+Zkp0EMqgzsK83pukdj8EDhPLCTYDx75JR3Y9THscUaJxm
03KQoBxtwM4UZvIbnnabIIf88cRBj3vNuqnbiPPcoY5PTIXQ7G1Ftns0SRyLqTTk
sZIBDuM0D2yEevIH/zzU3G3K2X/6friQxEL66OfFU5LReg4blIKnnMHpluQMp/vG
Xo9TPTvLfPMvx/hir+SvWUb16Y0+jUSS6F+Wlx606j+RJ/eGZzfz3u1h2Hhr0gka
b5r/onlWsx+VVQzzzmmiWJw7fqIfi7yUM10LNZzk/vKsFoMUb29MpzP4Oza/0TvU
L7hnft4TN+ig/+X3CGRRMZEuCAAoR+zSLIxPAZWVJD3AkYND0R6j0VR21n1y705e
y2FzY/F63J6uq2zYTT0dzUugrn5Z2dJwKLzIrZQOV5N5meuh6PjAZeawrVpRLpET
HlBb4UsU7jPobCax8DuSkLkzZyhSejn1Yhwj8skAnhw4V9DozGcDSr+A0ml1UJsK
xbHOZ3v4mbdSK++jtb+fQoPw5V2Ai9skQVUWLRXQhPZ1y3OMqQxmdgsI9un9lQyn
aS0Cxkh+xWc+OQwEyeV+3FVVYH23M0LvcVB2oedMjPdaqBVYSFUuyvRiPdHdZGZT
JGaaRQPnXvknWUASkN5BrUP04WIpcrU18UA3QErcCgP09S4UR6V63BmQy0Lod7Jm
At2CpRdOosIf6LVuWWL+bCvwb++fVCKoMtiHbPX9bRnOsSDLnilAmyesGDAPG6PO
f6sETjyow7UhPqWBu83XyvN96gWh5PBYBgsMUvcYWqYYapRgBkDv/U1GADaouG2u
HaxjA148tQvdKzeOSmyA3DiX6us8Qs3GO3SZq3icHpS4OikH46unWLr7dpqpX79M
AWAvk0xF/LmQ3bkju3rsgllOjwkUDz2ae45OmBL4mjD67ETy8/NnTBOpjh/TknEo
SZI1USSNGFlqC9b+u5lwJTU7wbyU8FmqjG1zrNN2qND799G49gCPZsFoTqT4dK/s
LMUWi+hffPPRFIR139EMP6iir6HA8i+wA6eVh1ANpePBFQ+SdSob1PGU7O6JE2uX
hq0G/kpmaseeHJ2/6q0jU1ftapnPLid1c/PumDz0zXTKlFvwEckv99vxY8Dfz+VS
gUvTghDalKzKjoH+0RdQP6c+C6hZvi1kok9iffj+KIlZ+MIA7K3a+GwniT/d4vSC
f27Jmt3K/nr17V4mAKgSh7hB1liAv+PLkk+naa5fYXxalFY43xZkC92L3HCSvBDQ
J7A4ZSK6nj3xLHkM+bSiLMACH1zgz8F1Vu0ljmNL9NZgRmNL9fgb37anBSg2Zvh/
1nfoRiL1iqs0sK99Yk8MbQM+YWdBcf4ZoXQys0zChV61TJUEN1J2urBeP2f/Dg5p
WOV73NdvKkWa7Z5tgSX/EGPFx7iIFEswRDHzlsJen/KwWRytFcVoW1lsIj9FMJuE
y9mWU1gzbEqimlEpPqjoNiqjiQxWFD1unRATRaXoYGaaJfdNlm0sThE/T7iUSMHT
9P4LQNdy4O5Ebtu2JVd37gz3eIldpc4he60Q0uBdiQN+bkEJ27E7OzUS84X6Y3IR
Zz0DZotawAkXgS0cFbZVXDjwgRpP0j26OGVYIv22AkOgpY+GWAAwk7iEx3tGJ6ty
l/QnMOInDvNzWfHKvJlERz2hSpGFEjd9nikWwCpX7xeJO/EfH/GAvSIO6qbMtNvu
X650ExQwx6WbEo2kti34M//q7gomQcHsPoI0gOlPXX2qIKJMuNhulRu/5etAmYXx
4Llxqc6yhSgTtJYSARX7YEzk36hefObAnqdOqBAMNdobjIAPw9S4jEEju6Mp2BSt
dJUtYImx19ZakqbtnnxyJNdDsiuGm6X5AN7dz1FnoMVbyArddm5UFV1+TtuVTgt/
rEsN0a0VUEeEQyRq3lOiHCSb44IRcusYN2mxiSyo0S++IDUEyseCA99mR83LqB+D
TTQnTEhs91EAFTOpCITsqdQwcscIUjHKOpkWn1oBIxJUwsMB1p8ni+Xf9ddZsM08
1HKfCU9Zuhn714deaIdfklVzwpfA2zjSX8883CqrKqNX0e+3O3jGyiPeVUQwD7Gr
AbX+v+8jPWl2ujMinZV8Bbw1L/WPuKMjNOkY1btmKs79DkgeFL/CiPVEf0MvEVj+
JvLqONFWNJXd7xQFysCruZHWlT+rLxqXsmX6uID4+f/4mUKo898h/Ai/Ek6/E3iX
kCYGuIeUzpPgm7CTZJumdyq6/e7Fvs7A3Ido8XX8n6yxdJ1KeHdlrRbZ8i8OAPQ5
Ygjt+mmiNTNVNgN0ySg3wjJoZCNUVbyoWEkTiE/lQUiZTKvki50qKMFhJQUYqvfD
sIj5JzbqeLvrAhqqs7W+PNRV/HgLsAcCaiPM5vWwUQSnXtCZKiLdr2tunxgjVwyN
mIpOW7s/OmcZH46HRR7ReyQyg+DbRstbHPjbn1j7LObgPnB6bdnyfuXMMFENtDbF
wqDu6L5ZBHeFsFLzAmOD8d0p2Wrc6nXPtzsRnRLXDt34S2PdQh91tNxiqO8veEXh
h9AqQiy9HmovV1Do6UtaMLMenCXehvwkTHACGJwtw1ueUcw+NXjaa22WF7hRGHfr
C+KAN3zH0mpzeqTjiHNrh89ip1eI3JH0V2G2qmh+/iY2EU4giWbITdqgMw8Op7DB
HqHoChCeqMi8g5zZ3DdEtDwdnPUX5Ie8fnHWQaQYNX5zyLdSPI+Kap5+CnrajR3r
I6GRhPLyNyfRja0ilIs1oGNKx+vblP+s6LfQIRs4y0gdefYgeVSvZgbmclLNMysG
XvEiyawkvgGz7C6q/QOoqJqImXVKtc5qw17xISTchS/CpttFGChOcXQ/RvSlpJui
BL1zjFF73iJtJLR+LB54IDgL2nfgIKL5Qj+N5UXfIcnOwqgkhPizSmUgkCdG+zNz
Y7/mbpBEQxSjJG8eRqhTjn6/GTmg6cEK9heHp6v6E9c06xJaOsXYaNhW5pn805Az
6QulbsCMmqy8P97YcCwKHKjcree5ZPr7b7MdlydyVLxgGwrW6jNlyJ/Ic958F8U3
2NvaetgPkTBiKJHN3NIt67+1LMTGP7hhlMzlxpLgMRhPgL4nSj8HOb7A2Ybo+Ni1
WGWuH11sRj9nJKjtv4RfU+0YnqkcMCIxozvUt2Xi6DT7tiAIIXLsQIWHlxGU66uq
H1ueuagT7u1OC7kB+7wNira3acAZOL3U4Lq/NZ2up1/WAx2RmbSaJctbdNcatS8s
ubYw3zy9eCrQaYApDb5pHgTQ/CoM2MA47QDJ4NIfq4CoS0vDioqngVMC+BYseiCm
muEko6uX0s89ccLGkMoo2VKre1EjbjeVJqEFJ80gidOg6UGjh8Y2jODa0xmq9F7k
exgCT8zorH7+ZfSGoKyLOq10Rhmd52AXk8cowNNjXSRoxs55M2FDJCxWx8OuR5sI
eyWrFB37bb20E8attz6m/BlGKBE4gK38Q3VvcIy8WZzBr51yQh93yuesxunzO9JH
QFhtTZtGN4PYT+9xE7HkzSr0E9C6PYMCc351ZkftoNQXL8Kclzh6K3O2unD6ITAA
E/Gz9/jImi2BboNhH7HHwASHYKCPTrjowmf7/pTHgApECxUr/QQMKKaArG4/MgPo
uz9iFc7tIQT7Zq6gVlvAFVFTzSwezCnVokoNzbAjQuq6RDSSg6alWrdDSVz8rdRZ
lIWqfNX9iVWipYaAjOljoMMDCZASde3gF07A4M4U8ecIdQ8DCfhCp8QMu8y4kuDd
jZxDU5/+/C0fomGkqcPR1vpb8w0QTqMM78WU/UmihLCdnxLI9W9J52ybPesxglli
T/7Lj9OTbVhoU/uk2t9vSHp2A/rU6SFzt61BjxBA8qPCw9jcsAaL1SmU4F6R2zup
V6mFYVp/UhZBdwKKCRh/jzQtbTd4cVI9UCp45k/C4zOLtoSkYLfTW0O4Yn060/qX
Ew5MH4wB0DRKS9mF4zVMPLZGjQQ3RpZhxkgR4zbY7QCx+uxleG04CBpUIazjFd1v
ng73hVQ5uJ6eJycHhxpilhs9KO5HCEpZLol5EAjaGcKgWFlChraA1gVCwz8ITRR5
kpDYwnkDqqS7hN+hY3/MP0fYglL2v9WAxQrBWP/hYOiWcifkgCU6GyD2cvuJmZv8
drs1SGrDyAjQl9yGlFlGAMiwpfMRINniez1Qlej5a7OegDuoCuS1tZtKvGNUU7Vl
KNNMBVlCQ0c2DnNy7Aa/EaHHZhEL6DCnIuBNQV/x5BV15kcXtXvX24qU63AGhD52
zksFC33LDug7oca3tJzQqUzkyGEjLqKNPiMeKP62Dj/ZtV0vaCf8vEtSq5gFuW6n
RqhNYCpvzMGXK+idDHRher50vikUquu4YStc/Fdy/EtD6CGGTtDHISPApGWxAy1H
FqNCqtd4y6S1rECjlRy8erVd9RWq22hDYMTjdhUhJs9So4hXn+Jpo7LfdihY9bAG
3L7fycyaEEF8q0ekAAiHeGbb3PJt7mJ/X6O7EjOngSkE5nykIqs2ihKhblLCttWp
mkhq4hgfrSMThvj/poBalFfwwtRw0ZenkiGGOcYlzr86inIlp0iBA+1ySx47qmoT
U2JIiVzLMw7Y6/CHKKntutM6xrD7k3Jg6Cev4/FtbalqCeA57LXbs5UH88crdZYC
DMib+wUtkfAd8BK3UaxCzSpPYUwDOlwLJImKO4zreWMYeV4cuydEo6Bbmh50z/cf
/ws3NQVe6sRwAr7Lb9F3LVQwKAZets+puOPmhMRWry3HfrOAJMmFUxKDNbrFayGn
WoO7IekqPcxGw89M0ctqyV60Dp3NY77XN5xscORsLb3qqoQe6Jv9m/kk1/lJsy/P
t0kyhSwW7mjXC5UXvJ9JL0yeegWct92Yb4SXuzxtuzhFzP9z4sj5owIRsSReehU4
O90eu1+Sfaelhop5ruRcCFl3uWx35YIO+Clhvkq7AhwNYeyvsSLuMnSDW4hGOPEx
94hbUtzJdN+ASSDLhurVCiTm0TOVqTuV5zc8jJSh9kBtFN/yDHvuV2o9atwRZpnH
cs4TOrFZuL0nqBpFYMdfDDlaFn3+8sNYQhkMOpEzuzgY5U7DA1KbO4fIdixyh6Dy
AUf5Pmqcy8YNn6mXP4JC9i6OQmZdNTgybePMkzJDJndYP+hkfXkh+41Rr27k7k/q
TBTPvNgIqxKLYCZ+qIdmeL9oE519WjrXuiZ+FVUW0vV5NoyhGD0Kb0oABNmMvxl/
TEN0YEfYM7tNUnfr3zZC1RdII4nWiwnNpDQEEYs1CpG3VI4MIHya/ZZkvs/sop+w
d8IF9b5CrmLnvXccF74HLvp7iSQFIPeve/cwzFqwZ6fxQJ0sv5a4rEsUdIY5mWzw
Lrm1qKNqBqM+7FkDMto4/i3cSzKy2gJRPFO9IWHcwxLSXrbKVFkYT7Dkwzv8zzuj
5MwbyFz4VBfmdU+zPJ+Cs5BmNkYH/SYLP4u+TOxNxGhSS5FVX7uj7J9w7Zcmbfs4
H8P5y+n2RdHDxgP8zBaznCW+5E8pAbuVMbpFSu3dK+l+cvEGoWPi8KfEchXIRpyK
r0iPIYE9OXvIod/e36WMemXKZYPVid4vmvViWnB/vZ0gD3Rd7sCkbsnPGG31d2h6
HdRPEJGdf0tFQR/mymn/jtkEjF0Y9GoNqbYAgl8ikhwwbVefIHksI8RLMcTTnvT2
NRQKI9iyTSOEV/EfsyQgXku5QlLOmNSu+NObuTSyprUaSKoHZTyk5b7Y3RXt1uUF
sA2L/XfzGhtY6Kt2ZKx6U443zhGrm48MVAramI6ote3DZnvQGQTO+5CXG8B43/wn
WQJtKY0vu2VksbQmQnJYXvrIYtI5OPUrflmGciV6WiSNfAiOQoPrxoJZg2LXR2z6
VTHkGbanT3RTQW6HtEYUp9o6onbcJMgCpL9pXvOfgWeSAerZ6n+kVk1shfBXTXaG
6/tvXWp5WUTnXNNOdfUKNws6qTZQdrddMWySdHduf7STGp8+AfQHFdxK2tmt68bZ
73ftg5J8oWvXh7Tn/VmFSSK1zKBZ1DigrkB4cvJYpqNLvcQk+Hg9UtPvVMI22qr0
V0ubosaPS48oSetFE2B0rF4BptCSi4MkLHFkrWaQ3qWaNp7PWK25XgBcQinvlvaI
mY37CIT5Hutan/VhI0NRZ7xn1vy/CqgLpVWitKY4QxH0c2CIZC7AEzGEXCfOl1U8
4FklnysA4vozyaVx2u2yz1nUhUH03UErQuT833q9xnaDj+iweIC/jWY8CKHeRp+h
S8foNfVdwQemCNF9SFHJsbXinaQfvFu6+CbQDqF/37Al1+75x8q7Hl5QlBEj7edP
sS3JP7voapAYyDrbV0Nedj1Tw6pLCPTCovJ07ZeH8lnJhbWU0QmHn6pFGN5kdza2
Qp83WlZ1d/ET4OvjFmUsvDLNhNYKf2uTWPKzAmn+XU997e5tOWhuSkTWe2cBC0YN
vz4KMFB0u4tLYpkdOoR3jDapU6HB6b7gH6dGDYFtIgUKd8w/wHo4wav8rOujQ3Fk
31FBh/3STIDH2SbgzNWN1RjRJtKTk4TARz9WXn0G3Uzh+vCBh5/OUcMpaxFiTsZ3
vrkZqwpDVYosb10P7XaDrokBRqG0/v7lG4rP5neIMrXadpA6ME10N/t8+b0PiBgx
F5ltbJYZh4DyYSCXFZmFpBmXiHw0QHpAc/JLV8ojMH7f9LifBX0MgYNQEvDGBULT
AlzNkb3Wo3qKBPRagiP6CVrSB9YiJo+ZXjFVeInQQEjHMhLWGBKs79r0tiRmxgV1
GQJAl8vfPwNgXqJ1SsF1AB2U45K6nhl97VshIopM3322GR2Zds76beDMeV4wmyOM
gVKyhuvZOJIcQpKAlNNX1q+sA2+Q07lsRitMVoJ7ROPyt+JVKxcvr2NsFmDr0vNq
xIMRjAoX1lIQAAUBzivwidwm6RWEpGpcdR9HePydI1lGOL5k6hdXyCnxjyg4f2Ya
fu4qgPa+UwW2Iyj9I0AT9F4kHPT1HWIHw6tSJpmTMBtfqp8ruvW8y7FtjQeVE7OL
aT8wFBlDEMkn44gIAOAHY1iMZ1tdWCI3TwtP0JG7FdD0wVMOPVFD88excpe9a9/F
VNYcgr9tsDrx0xMJmMW44OcSAeGHW+PNsBH+VXfK8i56gCiD7TVf0VONn+Wl7UvP
H4/PxaF08Gln12xLdy2V2JjR24xZGLx2qYJLgXFGDvq57yj9sxV/xkadi3rTF/q9
c8BuRZ3STZSfdiY21C2OBi5xVY3Q/qgqITnfd3wnkzAD8kVWooP4vCn4CtKppDTw
uzmDJZ6Kg2CuU/Ee5vYWpSHPb4SdNTnOaPKkLHURpIoKN+nYNz4sIa0mY6cLKDRn
z67cXec9hfV+RkeDiSoQ4k4LknopNW5ONDwzvJEaqLsNsFYgl5mTKqMPtoLuf/W7
rcK5+vcMV6ozMfccwvSXt4bimLCo8oFuoql9aNMhYAmRRPH2AvVxUbjr8ko4QIBv
gKJ92Jl2gQuZj8H9k41FGTQ3y87gKwch/uWIqpnxpbhHKnQI5TJnD8Oh3Jlit3kX
RVv0M+VfMOWVLRjz14vxhT5SuxIDVeiKdVfNxzRAPxlmKdPO8b5gvtWMJSv+DbIj
0XUcOKhd3evJXu1T0ZLts7xCSBs0FjEtT8UnhGOTl3dXtnCcmIFlC+mBx7yUswtZ
JVCCQanWTpcKaU7J91LZZ/eaL2IzCL1QJcroqTWZOkIbrEl40atJ1MEuH3qCtU1H
UqIVkBG+WM0xvop4kFqy6HSIvibSPYZ0PVYbLMT5F2vMsbzeYrmgnL/9ImAnVXDq
uDlvsyUHDtqWj6dlp2N9BL2q3NvAAVL1lx8hnJMwYhNOjfs7+fhCA50bJhaVWu6h
kAYPeIJpML3vmHeE7joOPcQV0vHT3B8zdg/6enpVelpBXyAGfx3P5kVXNt7TT5Zi
vzMkjvNzjphgrjCPAfU9VBXl3RD0fyVR7suvdZFdYKhYSs4EoONGu7RFJOhXRdJj
goHloxBof6vN2sf2MpXfVTzuhHrUqoVqae4VcvZKrG4YPKXoy8+U8ZGkzf50c6pG
+pZdDMqhcgnYPirY/pq+JAuEz5YYIEJIIaCk7ULo7ptBwPcViz/jveseR9JH7IK9
5GUnNzvN0Y4HOTZp960DuTpwSFcv2EfHHi3+Pl9DzhiSfXJzFHrsuP4XE1v6VmTc
0d3qevhHwQ1012BXkHT3jIw2EqM5VoZOf/qHewQtXCwMP6bTUY5ZEILW6i5Cb06e
ON6ow8S+M/IgxHg9z71ctBS/iBSaBADw3eXO3ivP8l52TjkyV0DZZ8dP6aGGNKrf
XjY+Ey/PbrLBzfrcBbeiuDBfEq6Bad+OfvzK9rfEdDhMM1fE3ovBfdY05c4Ayo1k
3bkoe5UWi7ji0/K4jfjdvV46AE/pf9mnB4fa6GaTHBCYWwJX1oGG8gDuoGEFOsZC
WZ1x0KuiP0XWt6st3xxscZpazHispiZp9PxrEDFi4wf1BKrin12GdGAzvOgERBA7
ozjXC8rR1XScsceFIU7UwzcsBGjk/I+zRWlMlB4AFtox4NTB8DHTT1QAC++kgh15
CU27TQ0ql7qa4vDT/ZPuu/CU3gg0uZeWmwLR5Jb7iAWeyGmbH7tV93F2ZFYJ/N8o
yZXWQv1/dfT1nZHvnjRMufQaa/QpzQ2MIxPqnYI/8fR4P0ETBzLTl5M7IkbAAZ8e
gnauqSfBQrX+PHIfa5eY0NbdIAMUuyNoi9oORxFdzRfhY9+sc3C7EjAtL+Cts/k6
MuSAPUe6vq6IJARkH1MKdzUn3Fz30WmV1QqiC3siRdBPl5YuYTsx7jN8Ulyszl++
q5wgK2avp1xhi8l2gOD/9LUgW1OnraD/WWJqOgw/3YkqUCJCVxLIgx33HfppWvL2
4i20SjJG2V8q/WV77twsw2ufeJJLJS8CDASaB5M4LnOqGXJUtWDWGKJ1TKMZEDiL
6lQLWxG19WCD8Dbzf5OVm6u4khkOHmeY29BvNjZs2LVmtLzqxdOYw2+qOArWyB3A
fOcD/VWAAASr7v0vwLRPCZCK2H4C9L3EkkTL7ggdpMWVhcTnK6dXhujd5/BbNwOh
iy00kUes39w1iY3VZa2Lvkved8wdxmomVPK1kgckRd0BCbk7a78NcAfhreY9bOUU
pV+rivGQ9SvKsGT7zP0Xm8rjh6//AvaEmJ2AAMLyPdO2tYDcmO20SM6eSdSCyBzX
WfnztIWuZFC0dBZxQtzfZQuu1AMN3CvvIqk9fA8RkOvSvpU7eiy1YTXTTc/GbtZ3
fHvJ8OJWoGynPzl87eHUnOYHigIoMudW7vAaX3HhzsQzPQTgCkIRk1Ej/d4+1dQS
rKiDi2yUoCoO7zDGKeKlNKzJ4njAWJPMmC6ewBwabOS+EY3781sQmTDJWbE13zdi
DwSSE5Ssd3ZKyye59Y/GJwPrTevoNBNfJs+5RbpLp3ZXD+m3XyQdq4W1R04piLAq
9iS23bSZEwIPhTWc76hMeIa4rvMPdE1VxeN1+hwRns78m6da7EBgnAZnEOilHplj
4gUMtpoW0klSrPWh7S2hvi97gEpkP/TUPNi+mw+HJ1/hgoxNdCYzq5gRf/QrPj+z
jxyj0rsZvJJZDcGPIe/loS36tRrAR2L05pkkkQbx9/w8x5PQLIIidOQTyyucv+lG
6kit01sf6CMhhaV8Sh5KkySWByLdWDQqedKY8e1hqoJBQm8+gBsO5cNfnZnwqu/p
R2PtOq8pWsC9sEEtg5eMGlGMJ6/fUs9UcuaPbgJbA1905M8Mwhz6h3T6hfgOVm1E
ah/rq3VmyrNllGENZMbVqkX9Wp0RqvJYBeUQsMIHj0p9UlHfJv3potMI6lwMuGOQ
MyK+d+Ey9rKq/dtkCeuUWaCqyvRI0RauRGgt8QarqwVZRNOdmaQA8AR7w66zxztN
0J6sLizOs1ptzeKnVMDJNts/t+aC/mrimcpAhltuin7zpH55qLBMUTU4SmMWpoHE
CADMnIHal4Sh6H+EQqhxI7dlNcqCUywVlVIcxJFcB9EQGDMlqefZrvkGPcMO98kF
0u368S8gP1P4UhhWPN4CxXnHUxC93TjXveKFmx6+yiNgNDpckdPEpIOcZdl/zPq8
0LPIq9485haSKG1a2IHaZlVLMNGkXAzs/TjtRmYBA9WUlF4i9vwvcg/d0fpl5xeF
BIJ0ZlkM6yrLSUoTDoKd7Hid/HM3hKb3d1owLXwffIegIbh5rzgO9FMqxbpLw6p2
5eW3HHedfEmV7JFScdlKA8qhDlgMC9mrIuAo82irwpPY5wtFgnkRcmW0KUKm0UJ3
2vWHcB3BUARy3KeEsBKm5uzTJMnwhtzFka6LwYDZldZPtz69oIn25dKvxRszDQTY
sQ7beUhIj7cYQSVqMvxoxDVwNcnQ489F1vq1073s9a/h9aR8agiaBAY2J8GVC8sN
0UrytvpgnB7+XAv1VTSzVkeEiK2TUL+k/mle26JAQkJKFqSm+FvufW5bojTCV81D
6l4njre3++mCe1bTYIuDgdfUu7Uf5jghtTbXVSaoogjkdvkSnvpIhg1045H3nEc0
Vvshv2KJ1MMyAeUbHxz0fDaOk/b7MkPVStHHbgEsqYQrUK7bUvXUQu+PkbTnmAKh
EATB51GNwgOlutcIIM621K1guSMINqktb1Q4+W9PA1pjMjPBlqrS2DysjpbIErX9
reEyhYpYxgQy5ubieFL7/t37jeYDvXiLyZdMAwfUpz7747uCiNbeVWM/QZc/alSn
V/x+C02Qo3Hh8dY1iR0Myi0sp2Axc+qfOrDwy4UohglDM5gNC+QlWIx45bY2Q202
ARX2kRH6gWXtbPKQy7c5VpOBzlM7POce0AngX37h1P0+Rb5u6WtkmkA5iXqbSuVF
FLEc5ZYJR8LYc+dvg7CGwi4l/zgNvQbxdac1mTor6DvyJffekAdcDP7gLotlXK1t
jZAdnZvlkSauqPG6gFr/5OVVhTqr76Ap33jLzJif36EEuobvguP1f0cfqxxP+CW1
4pIiIoaITmJsNWl3wiC/SBdzZoxE6NaBflyDibf5gVO3i5I0da4elrMEDz7xWn7R
7KOk7bg8MRON5vGz9vBwt/X+O5VWAvZ041Nu49CTQ9viMsKvIBMwMIlEPhg63+em
jOQRJWSR+mzn8nIP5Ch6FjV3cj/irp2L8vtGhYfN09ye0N4H0H+JGeBGwhOGbpZD
AZIOVfZY2IYNejDNii5wxW5NMzOp2DBCVy4hTmA8vaF40u63/oIhMuMMxfzNU4lt
/8NzwXxBYFWq+y1MO1+R4RxgsxVFV3NiZU8APNln3p3nyOJ3V62qHQnGlMR4QG3W
NW8J5NVmOdP0FExCIZnsQGCmLcrCzD8hd+y/8RKGo3llukLO0J3DOLOK5Ib1nkOh
i1o+/LUeUdkjJLrnU1DNlDAXI+stbcFn++097Kao1OoGaLYZuJ8iWLLXwoyNfdVz
AFyoF8mqITaKfAZTP+R+ib61EnQY3tIaIQItrKrFaZjywIrvsCIiktZcmUvyc9n6
DpGB/IGwxdte8yDhetheGgXpGLAJuNx67Ei++ve4dAuNIRk9n23eHbf9D3+szges
GZp3RPeh3dv5RbH/yFYvbfvdWQ2MuBfZ8sZ0f15CnqmVi4uJmqQgpblZ99WJ/YIr
DBgVqw55MGMwm69vzWb8GiO9ad/Gj/pT6lHSHm0EqQ8imFlYy2CGVTguwtx1C1uj
VyLyQvLXC9ejkplIPSublUstoPUckMrUMWTezfVTswKFfLLg8Fo1tts8Q0YbCQMX
dU3MkI4juf+Xl8w9VAfPe0YRo5r6R3BdC0zBYpHjC6Z9l30lMqcMz8T5zu1hK1X6
eVRNkWMmKJ+up2j6Oe5SNtsOzzdrYKcdE3oaObTLYSihB6U70zS/YKo8igXh4Awv
64QlEx41fRE44OFwj4+Cyb2obBK5wNDSx2a6GGXVLHKRbZqeof7bImu46q1cmEiq
5jIWp5TcKHfa50JGLZe/jnFgIu6MR3Az1+1krk3x6hSl+MII+ChBTTbOQSsJOETD
GkSvGfVSoRsAqH4hvdlsTbEt7m3oadzPk00U+YXYfnt00IGQFmexnR11+wUD+isk
6iDfn1UdumGuu4AXneAfHDGVRKu61hbnfGKNWkphXaSJOQzuEcIqulG7VfiMvr8a
gTQqzvdehbJdxT0ETvYFhF/k1L5Unmq+P9K8Way89MKx1tBLnghRiTjcstMRl7nB
XXYI/6mxcoG8wj2jW6UxTrtMXNMowAwJ4gaVr1cGONXd85SQGHKS1Zh8OO/9Cmar
H6Fqnz5h5lfdGGndCpsAlp+uI0iIrtadu/OkkrCFpj2a1wJbWDFKRhFgTubVsLpD
TfMMkFoRgoKhd0RqEq5Xu+QTZiZVwq3lLRH4iq8XAUM5ZGHcCuoz+HcSmc7Fo+HJ
C4mOdcwJ5PHK6YWBg/9inSiE8Ll5UEkBH62YNco+XkF2/tPST/KVQxGE2Aj8qpm7
eJJ1WGgujCOHbZ4k5CuS+l1/FeDBc/zCtWV/BBWu4IgrZCt3kQ6WCCux8ojY6Xs/
bdCo/NQZYXAamM4s8tWlqvrWXVoZl0mFW82NrZpy+5SdkNALvVuGf2ZwybANimwN
gEOatXt2wRgqvD82NNmC6RWchvUO1ONQeVzXprj8W+pXY9AvzXw3LJeJWpABcISs
MvObLRDdqAeedFK23hC/vSsT4eY7fM2/B80tCWy4AbFcudXo4oU/sOZvnlE7D40S
5o5ObN0qArJwwUoQBwcLLubr2Ums/RiFTKsbKPeNdgSGJeiGkaMhPVlzUfmNCdeh
yH29OT5RqofX+tkWAbDV+c7ql+7sMz/GhBX4B6+0ak5UR5i4MPtdiXx6aiuK1xxk
0vp7G+0p5wta3KpaZTrhXV6sq+l4fNn9EjT1yrR9kpkttUbc5Z1KxsvdD2Xp/Z0l
MTph06JNBLVyFXeH3zfgO1xVr529FFhgvaJusPmrcegnZZg2ZPK6itPTDTgIw0R6
fC4qsUPeHrWVdqocDRuxlg7b152XrkR6ASsmYrqaWn3rFgS4GkC1bqUWpH8WNXte
JDTNPkPL6IzbtjRg6BCkYQGlbcsG4QRJhD+nyZ5fSWZMet9GED7VHkW4WaGEe60r
gda+CGCUBf3uGaNAVIaLYqBZJ4CdGAD4O2jx5mgmwrHG6GwJzUm83pUymI2d2GQG
iFduCnQ7KWsL693K158RBqrZQaQDBz/b3yaddV/D38KlQUniL+LEbhP7O9WPgndD
ELb6CqglEskRcuY7AjGK25prrMgV3KVmykUGy0PBKH0j7F0PF0D204S/nnTacIp+
0MVkDJP0qKJ7aNV+bRcXXniDW+gbwCFxxc6Uf4nXIU10alSp5Dt2uwslAfbUAX25
ky7Iin3gFo1ARx+M/H4KS3mIASEPC2J63JosGDnNPOgmW5I+uS8zDTXrIkMFZMm7
ALtzvv4cxAznLucG/HIEsz7CcJ3McESFIUuXlEaw1wlFmxIiu4Fr5eJ4dTJIKOPu
X7GCzZn0CVnyfP4+7d5WkeUs/RIB45Z/66ZSMhVrVVsc4R0aLZSSkSstDSijPtHf
gQEnGNP/Qh5ZlmVham56dBPEsPfPDB9BhvKhbz182xv2S2eUoSJQPsqeQRkydt95
Qbk9QGIfYaarqzQj8TaBewne3tID/3Snggue9mHbuRUuIILU3K8PehhPbTSEEqZB
p6E+Q1i7YKtrnMqwJXYW0UiklYFzIw6/027tN6tvaVvei0Wgpu4Vyp3dvzyMrize
yLG7gdhluDy+KH82vrBw22NjXt/px0VBgsN8OTOUVk4Wf1xRC6BWxUd288LRYq2k
2UzKr/N4VYqZ7uufhKmfYwQ84JJTGih1HJM3XzP+SvDEOLvBV+HgdYQSp/xxPhyz
m9uXcFhFFtYmQ5XnqwcaakqPQVV7PctVbtRmBeimBdn2GSSV59zgItfE0ZQqlytE
1rG3R52pD0+kBNlriQlLjlXrXk0Q+O8tK7GcCpVx8nVR0ub2UciYYiEQcqugyY1b
ZTnnEmOismr9Nn6VQURRbS8ugSI2wEOMwfV2PQVMASzzcq/ta9U+bW1LPZcjIrSM
LmP3j8ufHKF0gz2W70uLrdNdaWdIpMlxe0HO9Wa/IibLWf5wyvOqLZwFMcGqSVWd
LCAHRI7Pu0E7qBUFpKaXbtRLo5HhbTbdIz8dWU/iwiJGed3JgdPukALOgjFTIFLx
SaClOxAy7HFc65XHu7GZGljffazHgsAqcbYhjiG0fFNCg48IWjk40L9kLhRnwzWP
cdzPED7B1yL3lqgDH9E3mlXCV5RQTLJ5feM1i5/t8vlon6ua1SSgLaUXLwKoRJL5
pnH/wXyIvrgkeydyAH4PaCm+6SHAXueFTmIb9uIbrl6cNyk5Nz43cjSvfaWpPRhU
ZtUN3/kOfmZ8sKUHktVhi69Q82EF29+RZ+S93zxzy4kkCLprBsH42KQF70KFKt1i
GdOWxx+br4QgpWvssixmlFMAg+PhNo15RqKfxVnkXWXrEGeQ6quLu6ip0Mef4chV
Yuy+mlorhoZwYJHxEym6KHopzYsh5HgUi6Q0UmXr1MES6Y5f++/A3L4G1PFAjwKu
t81Y3jUM16W4iKIljF5scFziDQ6fTVzzRTvhAC80IPCT0JaHsGDYKGrJ5jv5jDUw
71izvP1AD95jLV4iWdeT+zNFbNmLaKKU9gkbmeiDKbuFBonReInQc7RzncMbx7yY
qjL9mD1a7DSH82rJMVUkRbgIoLQU7cAjuXy5TAFXd0g6DwgvwaIKE0bxpWfoxyVq
pYkBy/8R3JWQUzuPHIS6ZF91azV8Aqrca42wLuRhfHfdmMfmrIEUEv+4LCYx4NqI
9Qhfx8eStC0y8uESM2IZ675cXtjSKIzOOL9fvwqc8Z4FCgmFIEYXZBXoNTAx9ZW7
cRuha7Oh7xEBeHraTAB9LmT18hE85WjkiolK0+y6bhsiyHbsJI2Kzzq47PGfGmHc
eHSOjfcAN1je3Yym2QlL8val5umH7QquoL3sfnlXKHJ63ruWLG+aD7EfeNLhxOU/
GKA5kdjtkZtDjbZp94mAxxuL0ZlLs0wyS5DVmKcLO+wAtapd6A/5jQWEb8/jAHhk
qy8UvKOl/mMdL6nk5ETyl0E/NY3V/ftAdz8z1kpEAdAV0fRoV3FGSres6Ev6C9EC
j5zcS7TfYSvynVfXk/ZTAECsuu6XyJs9xs5MmUzQznJZaJpasvXazAliur5CT8Ub
igb8LZ/FbxgMzu5mz26K7KZ0in0ELkz41bYqbrV7KhgRDNGzZXhs99a4pyeRhns3
YNEYIgRhwlqZtLzwRvoR7FMUcs7tg6Z66qJQlAoIpFO9DX2S49Ot+4dAd7eHobTF
mHg9B8zkld8t9A8bfysoFFl1Ww+o5bKWNCcZMtLXW3f2mKkKsz8z8LOopiVLxvkR
4QRoLjrnrZpmG5yXx75+46Mzwc9roWt/5basKyRiFBPV8i/8+fBL0uyaYS0UNCr7
YDCliBMY0RnMkVuO6iDuyf6uZIe24bvoR95Ildzyf7AiCcaHeayqExDnV3KfxNl3
h9KunbYsU5aMHHJk4QnWAUm3Y6K9uOiZYPISn5qlQ82AoXxYY2PopJB8vM3ZqrUX
rVR+zh2GUfGidwcAigvDjOqEm9ysYq/oFP6lT2J8xJp+i1mAR7tKLQcge9itKBTH
hxx1eEUbS/iHb3qSH0FOeF2clJUTLaAFDcDncaQtZgUDpzKcQ+37cjltNAXd96Iw
7SUKBd2chnZUMFjEreYhoZ5TygHD7hB6NQL+JUAsjwBI6Ks3ESLkk2DSlIDH6qFF
pXjx9g3bFhi5jcmFZYEjrsLyqxllHFC53LVXQJuMoT9NSdoKM9K/uueH0CwWiPoJ
qxuciLsk3kkweOqiRqQy5MfcmsXY6IwMpHN3OxaMij/I9xJJyy0j62Z/PZyhnndS
+sqIvFTAz268ePcDHCGHHjMUV0dSuytRXeXK45iSpZBszQZLOJYkjfhtN7zdXyU/
E3mi+PNpvnxq7yyL42GAnnwdqcGBIOFt0K555eW6EJG+OkEj7w/7Z9hqr9uTf2m+
VmgLOvjdrBoeOoda5OmiU/MvoaNqEww43bWbbMhFHG0ocvktBjlyfNNYGCBF+6Wn
p8Fm10tPe6zHoHfyNw5xXrk1O1ce1netWsQ0+eh2Jvmk/20khHEVMOddROo1askI
mDpb4kKhAU/NIiVxYuKnyIMXBMdhK8TihGowGEKYmdcs49WCMOCQEp5Rpaq74VLU
gJC8Jd/HEV/CkzjETf8JGey4ya+lHtY4iO3coopx52x0EedUPe68VzAJmLOSjn3v
t0ge3QrA2aP5zh9zoe5epLbX2zaRag0ZaXN1bqOEhgPMrqSZSMlt0LUC/gCfT5X+
y880ZaV/j18LtXQDUXpznVBEjH6yD3ZvLfL1uIUgJFnUzpkM2kAtDgPnfORr9jVF
sTy9uCFkVL3tE9D0vhA4gyYgm0i7MQbYC0tpa8/pkhtJixNTeOuTT4BPCeoM351j
PrOTzbOtgri1GZwK4pD7Pe2uPvKMOncLtCZE+HHoZmZrBkQbA2vFivrGjqgD+TFx
qKk24Fe5vAGEDheXguZXFzj+iTmSKPx+MNHxf6tHM3eEjvluvUgXJNiVK6C8oMdz
BCSm3RezuBTZ4ASXT1EYQut5oU+kEL4C/sA2p5qgEH+91JQ7phbn0donFM1psoy1
0NXWyXI+lPDlkuJaqSS+I/WKs6QOmby7wwwd1Xtp0POsTgxWj+flZQDl1IAshJK8
gw3l6bT1tX7N3cKuhtiF9TP+zUzV4DYPy8mN0oJpyCpv3Kyma0g5BYTmOgeeoBZb
I48cHjdCbU5YTUKdr5Tp/ErddsF9tmq5/E9z8nF0Rn21YDOqY+SssFaBJ3HTiuwU
EcDaExG2BVvkzpiEaFOFeB5msDbK+OOBxTrnmZtYVGKp6mqogzPcMfghKSiVjzpf
wtpovoBMKJrcLltDqwKWXAPBfFPNK7E+rRGc0WiH8umX0Q9wLs1ECiRqla6G9ne+
mLEILUrk7JrOHtttqVC5J7sLpewludXBlRMLi/CWDW9Gh3jMj3CnZL028H0c9nrh
NB4sUC0pvugmKrzJkkW2XEwqPSlq7nzkbYb/34E1nwQaF9Fxz635eljHACkRJe/D
uKj8qhRkvfuO347BbvT+Pb8GxsV7hrIlt5YsZJBnQ65Cu9XfKCJ8cOZQ+GtF1AyM
Bgsu7ObigjrM/8YoP2ajZeTFzkF5C10JBbDkfvbAoBVtQuLyScl3wdm2NV5ysw9d
YZjmykmfRKYL6NNkWLQl3KhbGxm4mRYHNmhJHS/l9GcOtwBSHIi2tskmO4wxeISX
67UpTtJvxvaQEmgoIPyI7o1FswuXT2ad7tAK1rrWDF35DfUN4Wb14qRyxzLsLmAy
Skzq087VhDRcU2Gecv9A2uxZoKscbjyjtCzBAWAXriNPzBs/dJEDgGb7vMCn5HfK
LNVcJhyc87g8ZJsRHIUUAGbGfPBYccF19y7DAcZpAEGdnO+eL8DIqUpA0NcC7bLa
9twShKeOUCwbhsDBX+ogTkHTybGT9SspsVGhojnLyqpkT71slwl8pgsx0+sbIaKO
aPevhw7JYF2MMZYYpcry6EysyUgBWYzuyXEjURBMbwGiNlTY+HZgeqZEIaPG5+WT
Gb7eavDSoDYr7rFvlCjbhLBuoSuuZMURSskegOE23aM3lQDjsbAgiHWBmyhNGdfg
hEQ+V/N6QODIgzoF27wworscqDJFsEa5fsNlMulAD+a7mFPdgIKtnY/bObTxEMsJ
YHG9+IL41o2MRDe5FNjYlu16FemaPNsG/JGkuy+mvUcTlmAvRqvpOlV8QM79zlYx
MlU0q/C9I95CqU1Lufn8nl/mW43cfyFkcNZY8YSGpkF7vcvqjZIcdo6N4CpL6JPy
ml0MRjWQQO21SRJA6r75QZNugjYF0oIblgEHOklJgcKL37IYjZuMvP6vOILr0aHX
QwngwXZqzlt7awCAx/7br5hQChgbYICY3WKweJog/apzDtrJmicVlkJKf8b3Bdiz
+TbUgCdV3a7AGHDl8jSS6pZhpGUPEZKmUavCXklozggpx1UWmSsO674I6K8pNJ+g
UcwmNtmNinGzHWbuU0uCh9nUGjfBsdn1yD3tR0vcFYCud0ZCXUcqwkFpf5wCLi9P
w5W2T9Ee7I1wwQXeoG/Nlq8y1pIqBr8IOu65NfMXYZw8Ua2ZIJEVTFGlW5W+AaNM
vDAt9HpIudtSnsjgyAoHGg66O7tXeHH6TakMLCmyReZl0k4qdpExdPUGlek8SSJH
EXZnXrBHdRparCdOSjjxWiFpknC1QczI1j9HnZo8sg3fE0WiBhseFYMagbpsoNSa
6QKOhBJfeJIVa/ldzivs3XIT81s1VOjNZc1vPW+w6oAyorC5JHWm6p6pTWmzuR9d
rpyoQCV1lhbBXMqp23vSwqPmfQTa0unyyKtR6B1siDgyvLgVELZBCKVrsuRPJKU4
vLca9es0THR9xyUGOiH0jnFB+OhA2b7CPL+Orp5l8Lz+LKtyC1oVKZAYtsvOO72H
J9NHZ+qgOJiWURskyoevsuhVPFGMsQtUd9gvFL9sO4Ifm7BLHPsK6aeXy87Eo0Pj
XYcdl5hl/O5WxQHpgxkDavW1ZyCXtiBe6kjRdgACcNDOdppa4f/jk/71Ps4rZseV
RzSZBZgCT1pFdLd0nSnrNbDcJ9csGsvDr1JEpg8Pg5G/kV1MOMzAFu01uJ1kGUvY
oWW+l2KDXGCXstCo/oY+7YzHwey5Trq3Jnak0NY2m/BwGWLGpVQgzb/i+h1NiQ4d
1SEKGMnkjodBQMTFxZHYd5YeNVEgj5CqbVboC3dHDgwrC+FzefRgbc22NMAv/TEr
ZTTvVH80TPGvra6XZGM5NlZi25TYplyDkOCpaz8yY+5usiXmqRGbnuEESwdiatS+
+Nd6KRd5piMpJ2NjwQWwL0ul4cJlAZA7nMlOmtRl+VuT/hBbjZT1Mr2f//LigaYz
q9YUJ2vM2Q6o2XR1Pk1vOmA7DiGOAG+UMvV0ef6+7gckMGLxjIa+hIW9nqNZ4jjK
1VLXU4rP1OEJ8pTQtQQ4EMafV4UjSWcv8tGkh+5BAziFHN8jV3cwxQnscYNbL9P5
LZhWa25+C2HBkJhm0oTaCRCdXAlerOrrnyVpRIyQX6gMsE47ko/jmscwTU1MFWQ2
ZLNX99y0SuDaHBUlkpPaeK3hV0LG49Ttx0o/BKjdGAPAPwEgRlgEjXaPAisz5JNQ
mwaZ3Owha5X5R03XAIb4nyWUrjdQVz8Eqhc+j2yoLz3Qi4NginO1c3zm62T0YoQS
PeeR4BQj2tIdSPBpVNHvuihu9JdENOck9K8wzWzoaCISyrDPjr3YKSSOIFPdfxuq
SnQsSDBZ2CyhvnasSp26nrhB+KN2Rk1OkjeuF5exiOJQL8tVqE3H0MGETtGtod/l
5N/PT+9NK+Xz6qiM9plnEmAKORG9j9alRAO6D6XDdZknqQ8z/eN3e6mvpOYUypyv
ljmITNn/6guicjGpZ0YD8hd8XKpASr69aulI/dTz3uF73rzb4t0a8JZ+5QGtHbtO
/tMlFUH1Rx1Trwbv34bfM4NPVgV7q9Tq0T0n64tdUa0NgoXLTpxq7NgI5QrY1acl
PAb03HM6HZF4rnel0qVLA/ngER/ebSdwleQC4V8jrT6iPXM2RDayYfSl1zEEMT2M
QbrtkPFIno3ndGg8CtUGLQ9Od1aW3OdP5GVSxKnz7GvRPHpC4q0Kg8RKggqjzBwv
gRwG+2CLqIgEFtUdqXlkyNtB+6OTf5eFBMfpXOX638+oo9RjQJ3eTLR+Bis0eFRZ
HDIdSfvxkWJHqd92+rK5FlNTbLwPru9qesrYwO1akouyvCcJjWPY3SpKVdllk4ln
UrX96W5vnZf2RueKfbvfe/UiCEj9/fBqgdX0Lpbur2sdbreLCEEAKwlt7ddJaIH7
lHtjmX4J6A1cmKXo8pnehr7glXxRwEcHPnhJq7SdwqDDYf7cR0twFJG8P+f1qY1n
nUL1yT8uI+kYIgTXwxhqoMvkqf63rwVc9jsrsX/max4aOnpGv1LetSXZ61bSApvx
zrlgmKRB0JoVdme+aKXwdD/1fhDAVe9Qw18s3lDYNVM98hS5/hwcdXiUjqFl6742
ayIkuzXLlwoWGjVC5qMBkmI7vcOj4Uwc2Tpf0iJ5pNaBVM0f69LjMBGs6q5BHQ1Y
Kd0XxqwGMl9L/ubrg5eeJnRPTYPy/ZcQ1VKpMDQCGTXcaYI0YN8ROwwiTl0JjQC+
4JKUhDjD4O5PUMLPu0o7ujQnD4Zp70yKGVNJDKTk0z6M1+XPb1Vum1xRgsL2PgU0
70gREIQvmR4Sh1+N9SMDqQIQIZn1r5UlEhT10GrFy3yWW86elvN6yn+2Yc8QANGS
eT/vQGVf0eW/tlO5EcSLg/0Ox23BP0LGTkZLP/jAtIeaIN40/II3q9sHdUeZ2+vd
lU+HvUblfMr4xb0mWUwvdoJtc8J34I3TQOLHvMcdYpqGf4rMe8BYXF3llESWHHFn
355NLb9htod1fG7sYjeTtmdWfV69GP04X+BtxXlwllocWgwqmPg0KzyccIFRA+Jc
jVJ+cpV95tElOR0KmhlTPjZxK1Q78JV5x1OjTmcLuEy4u6TRzzfs0Q7EJO7Penv3
N2PvJakrkrHf4hYGh7zxBy2AeuL1vTfI8ebyE0WF6KFFf87nqHp+1gdJMGj1w5M0
sAh4EebwMPkJnfvWX88i24BpHU6n8vQW35Z2Yx3M99zS6qzhrXsZ/N2nh8+HJ7Yf
7C4wlXuFtQt4pcUWBBhm51x9iupJzE9zLt9ZmopGAYl4cTj3nUwcLG9uGNlYmD+s
c3bmd6AO4zOqsUx1/lA279MYKSlblEGQ5hTySEFEMTh/lRmo/fOKeHbZfKXiFrbC
lLwEdj6SLHMiT89sG89ioDsq+7NkCSa2UaPdfLhP+FirVLt3375t0uVyEzznbfQH
CFUautTvSNndzzzQ7mx4kw4Xrwl/Qsh9dOLVtQTIF+X2U++SgLMB4UH4DbzEltqA
V1B5ycDhs7iLWjxB4ZCEdndPYvpe6bD4aB/aHf9LbIP7NCBflwLE5a9qmPfSwsFc
3y+MFF/KxEgBUHaJNECm7JXZQIBqTHiWp7B5ApLRlcWKGTcoqIuy8ms9s31gh5wZ
RN/L1iTzMXwyNC8J6U6nNl7a4iA43cqS8zO+8e5OnyC68Zaanp0pGny+LySduR3r
b/Hm0O7/NzKP7ag3RJzeJZEuruBaJUSr9foELnv/h9uxHUPmIu2+qHZzhOgVGpN2
rB3GbBjuepO1Io25wO/tU7uAudICjhDnzklKERUF8UrARS6EL0rx0RlWEEBcXFkV
gEmN6syMKbNjfAw0YhVz3jjeDb9dID+QsBhS/fwKx0mD6rV4r5sloIkmNktwkw/X
NkeQTnTkAl37pkNaI7EhqWjZkZwF05pghM4fsVTSJz9y4MxCftTMws5mD5j0ouIb
cQNnrikqMmkTVIjUQRbwH5Oir55V/lNGKkBcu8r9gubdmqIJshdy/7jh9C1aalBu
56uJEkgi/AwMSlCE5GMerssa2AkfYlviCLb3yDPTuPM5cqvGs8V44C1pQDsfM7yX
13xNJ7mp2SHXwcFreLxHPy/1WWsBRZsckbk6Y9kMhDzQJeqohrBNIyew9Rdr4m0U
9cJUhSKv2XIQ7cOUd86sexacXe4eIL89vGOe0HmAZvz8+nyEnAUy9bS8rrmXqvyG
LJqwPAsIO23h8URacI6mddt0fdGEMvpfaDsGS356+uOqH8fQ3qmCu0ROTJ3kyr9M
DNwozVRGVGpUzjcoQd27Sv5PfuvFczKsrrhjY+iv3topEU2dg0vZZo3nSZjIytjW
6R4kxa2QA0rKQOHT/2oul+DoVHDjgt34rk+xGrx3MCMdKHhGoBBsCK/R2SAhM+Bt
E+Ed3LjrqTYnlSnwnRmjGDTy9vlzvGbccnNTIDoyYNVWQKGNHV8oiqpU+czHvNoK
SasMM44AyvxjMNGyPL2Bj+XHl0VLbwqn6swulGsyradX2kQZFL1yqgLS95CNEZ23
QmkTkdFWCY2qpuhwCExNsy8EuXJ6NPFQ8afmLATkdcFPqiL8+rFLZpdKbPal9i0a
6EWbG2uauV7JPodTN37AjP08cY6Rw3rqXdUvdT9I3wmuXoxsONtKiQHHI8Ihe0gZ
8RZ3AmaSyIGHiEpyy18PTKgihC3k4LIBM0u19xAZ0DkMj0n0aMG0Qcq59czJ2rBH
lBOE/9YbwV6lotyYj9RKJsMQWypgLZrpjo53GpVShWCYg0aa93xtdbN9O/yQvgLI
eTnGYqnH8EgVRR0tMTMDzRXKeq4Fm/0kqjpEr8yjDjv0IDZhrCFj3qG6+FEFHqxD
H8M57HKeBWIwE/s1UnQo7p2P02DwXJ20YPte6yNQDGjFxk7OfYwooD0f+SYHGUJn
5wLeRV/UbClm1quNgwJI2dVNhNapSD599kaCL2D4PeOJBuMIFBkj0RX+uakyzh/E
VqRen2urG5tMH9QKkirQAX/jUZP8wHU6zTFN+HZjERM9Ida1Zek3gn5brCEY12Ht
NkOx9KeMcyjjgY852t4hvcbdfSJwfMFSfM8HwA9YS0JPoK5fSocSjC+0IlybOVDo
QEmZ0qyLp580GJLur1QOtVUQuf3GCUeolmyycN9JoSMedJjRthy/J3o6RcLTQOpA
Yc2m2QiMnhs6/FEXC/w5ZRRPqA4hcpIkK4kjJ6irKoWwbKFFzzTBFf6oqJuYmeoE
DOi5vj7FAykLBmQ259wopCwgPPthgbnKTwYid8Xf4PlqYZLSbHmKaRGH/H19qXcX
8zZz/7owwkomG4TagioJM+6LMuDcX7G4P5pZXBXiLsRbwnwPag3uAdeqixZ12p8p
zQrsoVoKxO0N9XRNRV3m22G88dQtDIwKPQbPIBhgYtj751u9nipzWP1L/FWkn79C
bVUVgEZkuwmKgW1pgHGAcAjxwtKTWmJ/GHBs8hlQrU/SdtuRA3FBjQFCdfKj/1Oj
as/Gr6+fmN2NCjoP/H8H09f3HbT4EvnlyvfFkuKfn5U78b9zIpgWyDyIByCQOOh3
HAqa9dVUzzrPuKWjjb3oYOqH8cz5vYHtIkTxQzCacyZ9gkuoE+X89wBGNdZJbJJE
Go/VagkGpRuEBGP/f+pQ9ofVmny1kBkFHFBuSFnZzPjmolRM++SDGQHc/yeL/UcE
0gY2bMDPD0gTbwy7H1u6CXJlOh3Mzl0AfAOBZRKsX7wGCy48opthr3CkaxYynTR9
WNvcF+i0Lxr+pxanH397esFWHOPonIbEa2Tc3L8PNdqS02dyeuPaHzYSLRwTVROV
i28AKei4FxdhtUqTMJ4YpkCZf3AZzlNIJJHVULK4tWwl8d2Pdy0x1TUoMDCK8HyE
g2AYhRcuVCpui0yZQUbMQg5A0Qzau5M7vatUkwqTyZM9THi7HbI+WhnMQDX4HRbr
KIQ59+vCGmAk2YNeigHpDFXTBvwuL5jFsFVYjIqdtwJvtwHS3xvs17cHWYjVSCsA
8daaFpZB1Z9dL++gNJfyJtKYFrgL3DonAcOS37dHXZwA5Lt6evhYHzGefowObOax
H4HcYQgZzB6T5OEPxc4qL3FiAR8wnRqnZV/pUyqsr3N93d/gf9e6K3ts1aXAAOrD
ILlQgoNl9rKXX/mClPX5emuNWmF5Blr0pgaNU/Uca5MB+S+o5zTzzn0YN9j1oIhk
ZVbOO4imQef9FHBc6MJI7iMKfSIENSwgq6+QoupSpsYY12WWlOAun3ZhRyhzjGCf
WSXCur5e+LN4hV/4gRijEUZ5TTaC1m0FKjogrwpEorb2gxiB3iYgsSsvNUqHaPHX
17W5Z2LsW6TMEk05EpXg1AgwGaruqrZp8L8NnRBxEJU2LhiVkAafil97I7RjanWU
E6gHugc2iWGSoczAUY8S7GB+8WroP0vBfiRRHJrfSo2soXpOpK7+Rxsql17a+37a
MFwbCUYQgKtsvC/DvL0S/xu+aDb6nMf7uJQWcZsz8qBw47ScKPDvjXuSeXwIkTQG
WCzAOzocUF067xK8U8zKyCWmlBSVaTgSFY3sgRx0DpyNU+y4ZmJbyjGrLCRiX9NY
hAfghISLgxLW4widy6rU01/LBI0xoJ5PtR10GrNY6+JxXlrieHzK6cUI9BJWTkvs
TpXL4EFBnJ5kck0ytn+gb3wbTwNeoSeoeM+BAV+duvtMzJh6p/M73Jc+GcFPXFdA
9sECldmqVYNjzDTsfXkpV2YtDkM9xd8bC/TcyDBAyDy4O/v3MYBNW9vuP+/C3shB
hJFFxAsP9zX1z5ZQUCkkm4TLMnLj4Y1rik8LzOCUUTvb8GdN9EoPjnk+qtkWjD3+
liDMdNCWtP5JTff8uPBDmfYkGdIkjsCSCEfqZx5uBO7pOUeMKPtradVrhxkaff4L
HSLouX7cEARbL4cHBbYq9fkrhkElOMPzqdjHFMfv9r0ERcVs6YTW3BzZteysyvSR
xgSkNnj1BfdeW64J7p5+jf3/PR0KnVcI/JxPmXVRhRKOkXd8lVQepobxM4FIiCIt
dKy1LBlLOOI7Rs7NNn4KmFYQa74CsVwQ5OYDTqLbT/o1ER19dDLBdHUCTzwnS2Cb
EDI7jva8EXQICijqfXRM0qrGD3JhyPTANdjRDRd3UQ4PGuZpitexy7DGtfuNKxGK
B6oaDCWGFCb+Kj5+xzKtxNe1hpvCU9Fqifm2R8X5qIGdZziCWgt8X3iC3gll2NOS
nQHoyEtDaYUuAjJD7zIDJM6asSndK2bXRlRfs5Yjy+RVz8zntx1f3GT9+4G7E7qI
8aqbG/TyPJOKFEo8McoJE/fjFRKibccltFlwqZ4GkVmpQO0ka/KI9+FLEJ+KYjeh
+as114UN0GcbzUTNDGUtTq5k5KriD7YVB9LAjBpMP5XpG4jFaFwFpPoi0Cy55Hfo
DxGSaMpDgZkC/GoY7dbgg8szw6Ab9KY1E/HGKzBqHok9Oc6CkcmHkRrSUQNEAC86
liIwPsVxgsbejc+bIeSvBURaAB/aap4HrWaaHywEjmP8+bPgjEIlKhUn5V+6U7Fc
ZYLocwI5rjtDsy8hjKqxYZkNj6YRjnzqkY9kcJyjxpewDmMhp2Szk5NzvBfd2LNG
0TChnUq++ybmqgxqJ4meKg9HxNfn923RGS1iYZ7d1wpcgue/NEYSVplCQS2uJ0Jy
ghyvgPDPeAGbXUmwU1zKmCiH1wLjfkR4FIIPegVcsHetkHEq6pgUaqaj/Utz+g8V
dtr4u3Fk9mRcnG8Ysi+W3FRLjQI11h3VqMSvD3xuPtoK4uKTlH91MF3OoK+OrjRL
JXyh0X+4M1c+IJWzhIgHfPLDEA4JdvzA7FNljeLYgD61kYcRqh3aXTQpqikrWn5o
GvWnfhtJ9aehzdJG4fu2VuDOWdIMZeClT5wzbQefUXUPRodv6/YHzhLntM50wWcY
IGhj2XdNWWen/dGA2uDi6n3LLWt6EfBYjCf6ldCvt2pjSTlsfBE9duSRnhjmSbR3
fdouCHDOArZB6pBynGykgDfHVl+R2PXQkdWTWnOXM0bJtYird6GD/NQobuHvSkTw
xQqSEc4RWKn0+YccDz90HL4fAPIJ6Pdvf2GRM0MgKh9lqoaRlKa2c++1lp8vyg55
SCpZmq1y5F9e9QzDvu8wyFbbvgIGLfMRZn41B9JCBvXlSAUvwt3WCg5c7ZoNCwSN
jl8k59jHMqv4PG8R5bOevAYs8j5nWwD1Xs5UQcR4CSdDS2P1qea3tdB0ypKSZS0t
5yua6xxJzhlGrGe6XoU1FKevwNR7vmfuupyFRfB51otn04yHUxEN+6FuFFYyN43i
OVhGbPNDK16M204R3N1M1z377wBPnLT0UUl59K0NR4zw75OEKQvu9jGij4c/jzJc
aWUNdxm0QkR0MYfJnouLIuvN32ceFnCVfIZlsB6rZ60Qf/yAUO5lVVBvVH6cTTSq
K4QJYI2ba+HHnGtBwNBYatQA2DfoV+yYC3OyqxzkS7IPlsyWygdE86Mubg2lQj+y
qr7bE4QvhkMUpqkvYnigpklNwa8Kt3WYtCBnPpn5Z9qCWmwoY7vo9GbSkz9zbYYt
eGK6VeU2VyOjMQmRVKvlLD/YiCguQPpMG92ZQ6tNf/69BiVnKnWm31aLHKxAKYDt
usaSK/xLC02wyAPicDeoLCEXSEU7H8fTXLwHoiTWzUQ89AFAmcNEolfTOHn1dcB0
z9WNQ03uHtk+D3EOvzVT+5zkcg8EYl4TTSBIMykzX91uqny9t8K3AA063jizMCRf
9ieEw0R5mTSexhodAKIXgyjXEbGfaRzC/ZYK3y0ooITlucVWLnsTlTPJoG31kke6
tqYWe7F8n9lgjqQAPYAKnFVU5lmQLiMnPb6IAjATMPb5aATh3JABYukzNXjR5KCI
ZXhpkhgEwFpxhHl9pOwVWa8EyOqNy53HOKzgYJ+tZCXr5pwh0IspfHFcarKgkSmJ
81wkpB8rd7exm/P3IxXKA6SFG++WsuVC6356V61SwiH4ukluMgfxZJkEm+jCAMLD
yn317KE/fK38yrOAsgRgEzNildRX225uMNHOjVBmUxMXcQ2r4f7nti4WIbnwkzPx
Oz46Zn4SXmo9b+uZOZVPTEb5LJLP0B2jL23tjlW7RVXLBiDk65MLKb75gXoZKMNg
c9TuvogvrtgrJKE8aA9eDFF57IkEAI8wIcJ3MPpe5HDMqWRmNiCM5QpzbiDaBsrR
74TVi29hWjsWkyjgqB+A4sAc9o1+3dYbkESGReuKqdsIToZWUrQHJHnUFRYadHEm
gI+np34/SP1TWP5fx6sOdP6g3jvqUJYKcV/oVw/jmEzcds3N7gOfOVaR6Sn5zxky
DplhlAkJ80GJhrOjrDrhxH8a7trGt+k4cCdRm30n3G5u9TVswZ5g0sSMqyHG51b/
SzhjMNwM4e/RIbhjcQltMx/ohW1qrDuQuBmvoLvKfnbRlGWMrrbg6ORzroNZKCTa
FuALxjQhn1fxzWQtiu8abJdFWaEyNrp2/sgjVzftt8k89JmKdzgreTcWm01/Nwye
0edA4MWbh/Ub4CMT/PzUlgspQ/cCc90RIpOB0HQiEVcpbq25WV8Rn7DJQ8qRJE86
wcPpk988OrLaXMDxFz1PWdBcGw5I2set7fFK4JiFZmyE05WVTmUEzXoXmsmjQmff
W5UYJVgM4vKJRt9bqps6sFWav0QrX5/268eA2o6U/9iJ5MnV9XGXn7WdV8Kodyc6
BrWPlZzzBjgW/nBKkG9Ap/B1pgeO2ida+e37jlJIbzfzhCx8g3GmLVZqb10KKPKc
iwVwQ/uz352KnOznRvFtbUmXwS+6ejqWchFr517Er+8e4QHCkbsPkiLNpOflnnUt
VBG07pd4+A6O2ax97el0fROOko+5aLkFF2aFKMJF6OXlq0Fb578akhk0lydUYBH7
Ias8kYCl3Em8sHs7pEcx/lPS48Zhj+kJAX/sZRIS51UCsQ68l/b2TMvqOvnpW0Cn
6nvMqsBDx2yz5AmU6UGgtPJz/9eBAK2QJogBTEpal6TQNRVeqGFa9BVpAIb1A2ai
es4M3nbp+dv1wLBb2njXvU511gOf+FlIfS8fQrdtxFzPQycCXxkg2fOR6SaCqUMu
nRMLLfyiN9LNwovffK1+ANzTicyIK2EMTVm9yVtoEUHx6LC9IdxRDNMAvlionX9Y
Go5h6fw+pQmdCVkiOipFQBhp9Ej0ngVEu51T/UQuhINZM3QB8QXw4IUiWxcP7/k4
9hWGRX3s7YbhFh6DoAutE2XTvqUMJf4VKtZSLafdtLtSheHK4mEpVdANiuAxyFUo
08OiaoenG2124qHjaq/0EwyecnZzyx9kqnKsY7MJQx5weeb9ZngSxgN5h8dU7TYi
vcR4GRpalKKtEG4SaONgFn6FErONUX5McKFmDalkrkAOO+VamQxIIYChU6B3Um6j
utlWrQLEQ12+E4NAlGD/U0vqBG4jFOb2Xq9mNw7qADCaWGz1El1gu0G5/KNuptx9
F2ppTVUBuEJR8jg1WJnMuzxqJnaeIFVGcQzuoo0waeLHg3LuCKj9AmW2VWR14KAE
xyN7tf1N8iEJVCIA3lMvNPchiJOMVfPwa8yKuxL86XyhsW6cAG2b6sKLkBHPU3PP
7YtKvlcQ70AHUhUVzcmJAPqFvZdGs40G8IJVwxciMJmYgRInCt4iivbxwc/Nn/o+
PmnyESn+Xk4g4QpbBU0l7ZMrignptfo0YjcxOjuwy2N9OzvJSh94A9L9QwFwgcFM
8iJqDGRniHFSX/ybIaSZkboKR4ZiHOWx9mGfq7zIJFkEPXfKNLKCg83qTiT4L3YU
VXfJfanwcKLVeKSOkSXqPDAkegr0q36vW9ss/wC8nlzsM772Dk4wxLvgalEwpDkE
yHDUP3Ec7MSfY1RO2e03CnAfGVnFsm4A6yRX20z4r8XAYfLhE5ehe2X1TsHztL8y
3186iOGJCcJgYqpfBQ5nYuhUiYPhXfE3ttBb2qelgAWwNr7FwsAP1okH/BUhdaMH
7YW+JMvk11v9iAGhTm/tMuHHQwbHBCFA0p+wiiwlg+wSGOw5suvdc6iZ40IR90Tg
gStjoGQmL5J1UFAtwcOX5hqWrkTRprNrYGaeIzEm+gv/dtsqHdeH6/3Lh2C4TO6z
Er15hBgoQuRYypuNSP3leVMXR2ogiaKIBBS96E2MdBij/saer2yDI3TzbZGJZWAA
ItFW4bhQM5ZNVVIaD3jBFlVFxvPo7GpgDYJ7jMX/W9Q3khtNTCHY1lbS/bBM4lqB
i3jyjB6KHkHOUnxVVV8nyiQI9RoDtZDgJbynZspjUohPUdo/VeRmDzsyZQYHy0pC
cNqc+9veK4XpRy7oOYum82CGUbZQ6m1csIYek6ihjZrug7GVbp1+Bw73fsQ2CRH2
Zb9PpKebgCXh4jV1rBYYczAS0Tg8wY6t2RQul9WWLuSuPnG3HUVPCto4tizSFWd8
PhQ8lwHu+m6xxO/XFj2mbQm0HVMfaT3s8kJ797NlefkLEuRhmrgSr+am6FuSaTVn
jpNnFOllAHWunMAL8eXErsBiLdoKDoaEkano/1OHdEySsWBg46D//N5kw6cLDXxu
+tOSD/Ged4Urj7DUYMscsbLSF1FuRqwZVLYgtKuDiU1ntBxsKILx3Pg9HBp9opBo
o7cYNuAtCs2m4TqBWHjk9ljE4p4Yr0MGrKcx5yfZz9CFVjWrAH81YWx+cAaVtkZS
IfHZ6YGyiGi9+obreW0v3E6dH7hVj5ZRJE6Vdcy5negmr6156nyl4kKMWSmU0dqx
NzOxY13n9QJwNF5U04EIwnpawhjHMcl0Jc2mp3XxhYaU9TruJ6BDLr9mukuSseox
gGkZ5tj7ezbmH3uPqy9rdugE+Pdi06D14/j3vVL+oFsAIxJJZhJ3gBJP/5hAXK+c
mMXmzJDw/y8O1eY+Ok05q3KqwXoekIGwUOj8zAoHgN7N6I1DMC8eDl569SPtYPos
FpOpDjz8umRjcLnIU5S5zfjBjP6qxdisK88XmhlXsTR64aggwuDWVyoIJAn1jtpy
Cq/fgrP31evJssUo71oDU+7IrL6LGMoxIeBLK2cqZsk7quToCvHr7enffa/wRMoq
kzbgTCAfO66+1frR1TjIiNYuVEmEpuDOe9L7rlK8FT3Oo3uoceToZE/OifZ3ogB0
KyFnKuE9EaMvyCY0sEkA046VoumdmDwSlvLEYgsSeW/UeVPgaJvNbzFaedC/voAt
hJCLG3d1tyJeuw1NO6L4xu0QPOhpPcgc2d44EEMC3ZEsQGTU/o+LpUgrYCzoXDed
ZT5MzE4IJJLCQTNCc3rVhnYxQZBQF9F50YFnV6TqQGtX/PeyxLXwsFbN6ElmSwce
xaiVobedjth5wpli1QRRouBs9cgXQ6xT5nm+QSzvNFLlI9oztnzqBSb9if5oppme
qRi+KQMzBJD/WqumQWmVWyomFG8me0p1OqOdHcWtMHL9pwq5YIQipWrw4JLuzZZx
BurdPntkTDskZnljm0tMcjzOTrhJp/qybe8Lgorl16WMBDmDfKxCI/A/uTMNXZQD
Hfx972SQI9ikGvYxPtWidvuNUP99EsP2gV66qxttIZSOzuPZ6FrG4py5ok+bn0GS
RjW+2W5OlxnzI85W78syeMAgG7qXnkYWUtrd2JSPejXzcW3MTWWU8CV0ffEQIS69
u/gL4aCP6dj4/csJABbI35/ioMmeLog5X/xnUsvYxcnQZCZVUxsFD8b8MnXlNmEt
k0djEfVrVBcDQI2pWHxo0PBdxiJsL7EtIc+D5flZFPb8aB3mnrKoaP7Ze7B4tDMx
xFSUV5MvLQEf6xVrDhRXZNe73eJYMcSZGz0yYC231f8XZcL+PlXXkCB79vZuHXyA
Kmp3uKH3RuiF5qGHsLSjrNeviN3evn7ioVv7N+8YgDSQ5DrBER9r7bIl2bYjDoRm
S15aM3SBojBP4J3BEOJbjspVKvnTjRSB3VRkNEw5uclxdVz9h1vsguz6RRjin2Is
s+3cS7v3kfTOeWbaHEHzGRfCKGZI2wsEIFHPUtRM4lZGv/TVSdD9H5goCfhfPgq/
wJEMgvx132FJEzAvjMZ6yRw17ByTS/ynngA8XS1hJLPK8kOHJ7HTo89auh8ZXsVi
Vr5Hq30q+O2OmcHVBCA9n28vrPpjzA57G2WU8JOq0tRKlU9ZvCaiPoit3z2lHnDy
QiesDVhjwKtScfQtWqb17nLUaBzOIYY4B724QX5yMDPNh6Iypa2M2/3J1QkPuPTO
5L0k9ZGPTEOKTScI14vHLhfUMfKgm45zj2SPepo7JzPZxvvx+4xCPQP8LrOjnaV9
sBVSzdnKXSOr2lPMBq/OCXxpKcwkxibYEIVB3fKoRN4y1rgq++Nlfw53LuTH7pwV
7JZTs1IT0s2uLpLG7iTI+xm4GeNaUkd/j6aZ19vl+n5pYBtCAlYRyPlZ1kw3bO8g
2Al9cianAjPjLX+sHXr4sVtTuasKKLNQ67kckbLQjqLhnhY05h6LNo2KAEXaYdV6
3v8I0PvKHfdaWC3ehGBp5JOAZZLnMHeojPO+cOYRf19dcLYCSZopKJN7TwuXs586
g4vlM/pKrPNDA7oN1j1cochu8sbw1eTDGucKQunuC8HFvybYy5D8clt1ApN8rqVh
+CUEz8eE1Q5dey99LrUgNFunVThOPnxXVsZ/N568w5vQutQr/Av0Sz4z8jeGCqtW
/OIKTRS1TmVh1yHZfj7fRvnpLudI0WovPchg0zSV05IaU88jOUFUBuNprcPhVXTI
9BJZpwT/f+NaOSQiGqRSPZN9oGucvwEYqJ6+TqlXtrDXpbNC9J7WWngCfwesJT5F
DkY3Pxr0UNpT+YBz+5WyDvNxD9UfTRPHdJzl4OycfM2k8dO6Bad63NcJvrbKIcr/
C6smhxT5Y9L6pHCNfi9PYj4jQ5sm5KGWYHa8zOiKpGlhvbzYhilOn3SPVTtfb3zI
`pragma protect end_protected
