��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t�C�C]Ԃ��z�h�bǑP��v3�N)+��2�.W��܃d_�#�~�7X(�A7X�u2��J�\��m�uxL�2�j�힛Z��B�[%���	t�U��
��X}m���Y���ɛ%1�cG�G%5�*�C�fߺS�I�4���מ�q�҇���ߕ��Lm��6�z�PME�#r���o�а �W�r���n��}ru#-Z�f*%�p��A^v���K�Y@������[�گ�:�X�n�
5FGi�MgP��
��?������َ�4gZ�%}�q�rT�EK���v<�E�ln_��ɋQ�Nߓ�� g:�nɕ����̒��V��ܯr"���:��/���S�I�DF�+|M�^���vh�L�m��͗QS׉��~�zP2\*ݟ,G��}kDO��8���y4^U�~���`�F�����f����9��tԣ��܍�R���D�OjVڸK�GZ����˦N�V �M�Y:��S,S_�
�@&tZ�226�wO�o꾅/��,���i�8<
E 1��������>�B~<֍�!r�E��Cȶ��HٕUiE��>
��9�^nl��eɢy�<��
��@f��<��#�qjj^|pӚ��2���@`������ޛ<�/I+����'Ѩ�F#��U��&���D��ZFaٹ�Yvt8$ʾ�.��]I*8ڙU{��U//��|U"��A�#7������e<U@S"Cw��w1�r6�zHY�OmhM�[!¬�����>�����x6�kZ�غ��
�o��Q�T�x�� }�&ǫ�ڤl;�MB��Ӽ�qƗ��@u'r.a��\����RC�"�ٳ�5���s�ߨ\lf�{����j#c�%����V�5�ח��}.(o�Gi�c�0�'�y�>3c�e�Go��1 �j6���a�b�_N"��|5�y�@�������#�m�˒�i�L*�Ll��L�_�K�C׵�މ������͞�\��1�rT���Ô<:N�mC���]�c��GxE-�(f�EN8��63�L�ԓw��^�)Rx��Z�:5��P����� �ަOp̧L9Kck6��&�|���"jF�tI-�n���f���+�q��v�΂�,��b"V�xd[m���3���>�s�E�`��ꎐ룰n��d�V*����	�O��C$���z�G���o(�f���"Wr���W� �"d�l�'��.�}b������Y�L
�<�f�r����o}��T�>۹n����P�g�o�T�s��z�v:�Q��G�2=^��b���B��b!�{�T�Qv�B>)��y��/C�~BX+@�)9\@�B`��g�Ӵ���!��nT��"�?�]�մ������D��1V::�/�ȭ4�t<��N��t!�If���G�=�ȹ���=���,��� X�2х�c��܏�1}A��j�Z��X��+��B��6Z��6S�	�6~6�vjbJ|��3��˧�;�@��gcĘ���Zvңu�� �����=<�����B��V�vH1-�pL��s��)�q�*FYQ�8�{���XW�e&���8�`GE����}`P��	���$�HX�X��h�I�&�CX��j�{���!<���%Y�KN��Bd���5v<�"�/��sC�Z�����ep�z�-�`��I
�q�<YF�h�<�z_f�pl�F!f�`��c����M�"жnA��h�J�2&3(���HfZ����Oo�(��U�Ui��.O�kR9�L�G�*�җ�.'���~��ҝ;mY@L�I��m��;���E���:X{�S��t3z
V)r*�1>�/W���ǈ~��Ǉ`'!^1xV2�r5jk�Q�ߡ��R5��/�J1q�IY�DZz�������]`�XY��/��LƬ�m�e�w��&�f#!Z��m��S��eH��jcUrWԥ�Fe�@='�ل*a^h���Lk��Ҍ#����"���J��N�_�jх�T���
�C�m#��-n��MW	{�SI8+:�E̹���Ĩ�Ǿ����1蚄3�@�@1�]4,�۶��M�4h]��<_@"�+c
��qL�}T�l���@lJ�s����r�Č1}=���ܪ��� c�V���xO�e�RgȢv����,Y���J��S�|�K�ĝ3��}i��d�e#ڂn5��ä�%��V0S?�r�ũ!b|��9i+�|x^|4�ًK=?Q-[�B&�P�15������k��_4�]Q����r����.癘��9'��S, 'w9={k�[�H� 	�T&��͕ok���|b�a�&�A�>��m&"f��j�n I
����� j�QS����7�<� ���ژ_�~����~��oZ����S]�܂�݀]ٖC��<�
װ�r�q��-����zM&�m3�3i��@ƌf�X3�����|ՁWz��b���U��2�0r�q�*^ln\�˳�H���P$p�@^8�n<m���՗�h�Y�ۂk�e�{�~���!Vą���ɻ�W{_r%���3��Q�� �s�6tO��^���Q�@s�_jJ���ͥ�8�� �N�L�ё�h�Q�b�!=���ֹ�(�����D���PG�~Aʀ�Lԯ}�6���~P��]�r; �?K���2�S�&%�
��+8A[6vH�H���m2[|��[`�ŋ\�9�����ն�����I*�v\��Qk����c���f�t@1��äܻ 7����c�T���e�-heV����hsdlB%�=4%n1�@��2���|�k<��1�!��Џҡ�Gg��/EC�(Pv##� T��D��E����s�D�����υ�h��3@�V��Sj(��	&uh�����q.����Q��T:5�0�z��8x�&�Q Օ�v��Xʹ~�3��X%v�7:�>����%����s��7�C>MR[��"�)��IHQ�#:
(c�.����%t*�3vX��9 -:1��6�Q�H$ڲ�"�Y���C�sc1���MY{���q�6����7ݼ$�P��eJ�s&�C��u��������C�.p_%�� ��T&�#M����;�H��&$(�lѾ�@p�N�����Fe��:��_\�W ܍��u^fC
�=b�Iʕ���Gb�,���U��׽�SAx �K��qP����Ro�=��:�m���9*�>����z�x�ڞ�2�a
��ѝ�����l��֭��@]A��
���=��P��V;8���[�����&���!(O�ڊP�����@2�3<2��ʙ�aWt7���Ҩ����W��}�P���T^F�Z�l��`�x�6A����|S�9�2�.����pL����;�+��QZH��!�[�/�I��N�@���D��3X]_�(#����e�];��1���n* �L7TX��Nn��s��b��
�I�0������L+|~l>s�p��Q���V�n��=�:mEؑ��f������$����uDA~�z}׻h�������C�P��,��e{��$�p}:����S�a:i����O��g9Č5�G��H~��f.1���ײ���K�L���Z>�\���J.�b�*�v<����=^�"����-�g�b�y���#iߒ���D�5�٨�5dC����1�!�MC�
SU�`7�L_����[m����t���R8e��dS���vʗ���y�x~�_d��C}_�z7�o�J��?�����0�����_q>,�N�O��e��ڥKI�	j��*�4�o��G�[�r�1�K���rW�ึoE�Ac����u��˛w��{��A��w͍�v��!�3CW^(�NP���o�§FU�:]�R���L��ݑE2%����o���S���4'&sٵ8��YGR�Xsc���QW�����2��;A��E��;��	�h�}����8Opc2�\�EI0V8ߗ6�� lLG^D�S�C§��!|vѽ��_�,}���Uca�����w�_���\ ���	�D�p ��`���4�� �y����M��&%i@v:D��1�beD����T黆mS|	�6��$A��)|L�C��*]���Q�98i���%AL�s[��MmHy��&���z]|y{x"�G����t	��������ua�@�B鼃c�`�� O��(�R�*1��Gvo"�5��8������"M�֝?�(���\��)K�Ơ��f���s�u9����DT�l�#-G�9gZ�[cĀ=\1����؅4�nRϥ&�P��q@	�,�7K�k��W�I�_%�dĆwLڮGk,�^��җ����.m��Z��.i��\~������~A}����a������<^���(��&u$9��x��l�fb�~���X>�p��8���T��[lre�s� ��B��c��H��%�Ǜ`��,��NF�}y����*�nb�	Q�����~��d�7�wl҆�"����#�s�Oѳ#Aw}���*���w� =�T�->Ņt͎�=+�	�.��% q9���q́NO��C�u���s;*����Wn<���U���D
"�Z��O4��S_�L�(������t8�L�c���Y&��[5����0��m%�:�F���_���
gyv��R��G-���~�` ��hui%^!`]Cc�7�`�$�Q����^�aC��nV�W|c�h�\�;�.i�|�K!B�&� 0���9>	�`��7>�m�Jyk��m�CV�7LJCSa�"4�ߓ3:���7V&M1�擲��J��C�a#��%\�a�~n�Bڪ��GMrl���ڿ��l�t	�ȏ�j?~������%hP�ܛ��% ��U�)�:|�`DM�r5��N��������1�e?�7.����VO[���
�6*��%c�Ϟ�e��@�V����x��Y�/9�����]���k�ճŚ�����~�h3�K�j<��d������R���a�,;9j^G�%�ˬ�K��I�Gu;NӨb$FY�T�����HϜ�)(��zh�a����g�W%2�c�'b��s�=��֢�㲵OwM ��%�&J��G�9�D��*Z�ܖ���y�SK��-����Si�����\fl&z�;��e^El	܄���X�^a�=ෑd�t*ֆH���E����^mh���_\�&�* ���th�T��妆�du����̀�װ
��B;f�w��#AVa�Ⓑ�x�A��fЂ>Z]>�$�S�b���آ��M-$G+oЃ�!�j�xߥ�R_{U�@neǓ�-}0��_�T|�X����rp����N��Yw�i��"�5����b��2����G�8d�]m��`^����|�_T���U�Z0�b��'��f��g|Y�A\J��j�Z�a��=(b�CC��`���Y5���d3�7^�;8�T�JC`冠��^��V�����f��yt�K4�1/ϙ�Ŕ�j�R�,�6�m���:����qދ�	�
H���K�m����ϧ
��/����Ɋh�s^��N�38nw*��pvr����d��Q ���;.��ڱL؊X�U��9���.a��P�����6kL���5X�r��]��<4��ܝ6��&K(��zr�I��d1�����g&�����;�O���U��O���>���������x2�I�>�[!{�FA:��6Y�W�:�ka9{\�)��iB��U��;�ċ�#�3�_��/��|&�U{�����N�|x�2�}W6�x�*"��Z�΀ݟ����nZ���j��ZW�3��׺��2��t�>�iK�B#�;��Y��u"�G|��)g��52��_�e)�!#-5�w�[��]�"Аn �������<d��,��Q��窞�k��Cu��CP_ѝ�#���5��4YA|�bgHg�D�KF�j>Z��V������<=�߳���"_n%lvF���R�1
u%{7oG���VG���F�w2%M08 T�}��SC��o?�s�gx]Q��MF)T1����(?�[����&�x����Y���t����6����v{��oZ4�����j�U���#x4��>�6Z��g"3�֢0��/���������<m^=��ߋ}��<k�SG����=<�4){���;	�TQ�[xA��}�s'��	��ta�{��Yr�R��ͩRF�v5�G6���y�}��;��+HV(��h�u� [&Y r��=�q�?�c��j��@�K#���c�a8�Ĳ�$��8��>%nn����Ij���E��`1O��sO	#sų�J�\J���'?<A�����+�"k�\�Կp}U��13�KùhV�"D$h�������!E�E���$ GIe:�@���J�/o�]�0����@2�� �}4�ǩ3���yHY!�ێb?b槍IA�	�/��\��>�"�r{v��һHQC�e3\��U>�'	��t�9�B�0	ӹ����3�Rr>�$W��ï�d�.��|���󃺘�0�#���5�e �_^vg+��;~%vg)ݑ������PE�ϸ�7��k��T��� �]�5m���S�Wm�%���[��ݍ��À�gBO�i%;����˦I,�BW���K� '��{a�fq�� �=���x�!www������,�fɥ	��W@C��>Mx��fL4A�Sv����~��&������*~�6V� �k���;��p�&YUh='Eo��P�t��գ�x��&8�u�$Tp���œ��RU�P��Zy-t0�I4�!LBa�m�.��_���9�y�i�@�S��;�{JzTh�|�F���B0Ji�t�)	\���jtɼ�$��c�/f �U±��k���듈�C�䎀i���4%��;���<���C楌��eGT�p�Yc����:yu����ȒiC9����{xL
�K�P<g$P��$B�[����X�V�5p ���DVjHQk��zK�%X��po{_�CQ��>],��h�1Y�~�S|�^y�Z����`[�G�^BB��
��. ��J�)#)R@F���.[v�"��iL�a{�充H ,�5;v�<?F��J݁������@���JZsj�n���%������oܝ�7A�Iy6;��������Gf>P%Tw׏����Q�2�sh��7\����2� <���ATy����^L�h�-®C���`���#NN!��:b�>?��bQ^����^�`,X��~I�����X���{��!��]�Ka�a�S�7�Tuk�10�?(�:�ǬN���>0����	��j?(���
�������T�Z��P|Z�|��~��n�eے sn��h��Q해��)s╊*��F՚8�Y{��-���$"�8�4˞C��g�+��o����U#n��~�
�1Aʿ*5��c�����卬f��3������h�T��(�o�ג�g��o��^T-�Oq�<�ٚk������B���p�����+�������t%�A�ōz�O��E>��vm��k��3Lzڐk)VN�UuV��˽d��=�Nl��>r����#A�~޾0�e�����`�W�^��\a'���럾y�W�U�C2n1����˟��]$�!7�|����
+/L�]m��h%�T��ݵ	֒��'�?�m۬8=�|sXe�x?�W^،�jsl�+x�X��v��_r��OX���3xU�
ũ]Pf��d����I8� :,L�ju��̺�����H��J�o<w��M�ۯ�����#��Am7���T`���(YK���A�]�v����+�nZm���a_|�l�(-��+8��	��iǥ��"63,"��*�/���=�O0d�@���"��9�ʐ8GE:ɺp���"���__0��X �rA�ɼqj�+��t��˰d��ں�}���dPCs���B�m�^$3�����ј�)�&��3���N��Go)�!+yJց�\r�H� �t���O<N�s5^H������ҹ,헹uq9��ދ��0�XA�k����@p��i=J�	����̚������6����̬���+I���֊�H9�tuB�����k�cv��<���{���}J��$<�˅$BR�
)�� �~S�c���D� �0dX��$�����f��	E���ܧA t'FbVK�J���]�
{.�	��1���*�ۺ�Q���Nu ]gDF#�b��TN����-|�:)��$'/����,�H�����Sd��@.1e��GN��Np�#܇,O��kfls�����2�ȰS���rJ�M+����!#��=f��L�<*��%L� �u.b��$:�}���ǿF<�p��_�n1�����)=o'���<	����5`����ddI"�p��3+�6ƞ�� �jY'����'�3�0)0�+�
5YA����5,���GR�����"+g���|��>.��6�[����_�s��o�E��C��ϝ 
�s!�u=��2NF��sξ]��3��<P��
u@��IyB �-�d�aS����v���l�,���/���>�4�DO�-�`�.���{h�&ԫ1@���f�`k�"V 	��g�=�4 }�zN�vU�>��,A�e/[B�����V%�y�WP#1��qNkk/��
�ݛ��pL߶U
u��p��ŋ��r�#��֑��1�<l({鶼�9��oh��rހ9�i��u��*���*�"�ߞ33�a��<�̌s�1w��+�%����j7�,���K�"���a��HE��Jx���+SX�z���七�����T���~��0�Pj"(|��c}�Đ^�{ ϕ���@����s�9�<d	\ߺ��RG���n�!�X��J&`t�fJ'3��t�ٳ�܁����a�^����Ɉ�����3��x5N�=��U+�f�SvpY��;s��{��
�%��}��L�����6n5������"#��o����p_+��QJ ����I� >
&����c�������{��΍���<v�f&����ۂ���*[mr��φ.�ڕ;��>�X�-�Q�o��UX����l����A�
���#��\�'Ն0�`T�"������4�����W�7D��X��m?�L10_���2�9�껱H�Y9�* ���u�l8Ps0��4�kv��":��7A)����$H�-�/��pX�%$�	|�����Q9��UA�|9�Wdy�2���9\E�4�'#��6����|5=JF���D�vN !i=����4�;���M�̈́cU��*�y�m��vG �����"�WK���B�A�*rt�ͷ��5�|�T�9Pp�mpi�x.-��ibQ!�߱C[i��H��}�������,)��p�s^W����q���hA:�������~�ɜ����ld��@��>}��D�Zh�;yz��[��iu��ω)�u��� #pP0Eqb�ȹXfrj1��y�jk@�����]�(/��&,��H�a�s�*�R�������L�O�C��k���na�;�{d��7o��V՜��9�Wnef�Y�rz�i`�&rp-U����Mm�p|��{��Lq?����c�g��c5����kf�Cs8?������s���O���g�8�i�怓P*=Ρ�k��1�pӮ�΢Z���hF�6�����(�9
��Jp�����z&�'����+����͗8�W���\��ѿ��@�����|�t�9��r��'�ﾃ�Z���y���fy9Dr�,Lԛ>�̬Eg|嬭8iQFO$J2e^�_1���|"��dM�u�tTzԈ�{3�-��y[�o3�HK"S����+Y���=I�P�]n�Uv�ql��_k���hf9Lj�15Bx��W�$���;0���9o����.��ߏ�V�>�)�E��q��#���]"��~Ȼ��y�fMT�7��rL��������%��)��'�|�8P)��jB�$��w����_����A��
������2���_�u���ȩ�2�8�@մ�����lZJ��E�܉��DG\��fc+�'(�⁯5�U��y��%+ ����5Y�-b����Lߦ5�ta3b@5�����i��aڴ�F�QL� ��Rs����Z5
�cu��I���|�L�#�gme�Kk�վ��a
X+`�"E8�R�d� �-���O�I������V��,���gv �?����wz���
�O��=��X����G#��FU|� 4���tY���D�@�׏�"���9�r\�U񄱓�|��[ �t����8��h�Z�M�x�7�[O<ёm�dӪ�|�j�k_$�q����I#�� �r��ɤ�b[?Y��m"ԑdI�w��,��Y	5��iu�{�Gp_��D��\h6�&ݘ[5���hMh5��r+��b{�V��˿��^����J�9V4�,��h�hל���=�j��/D�,�'�?'1"�6�dF������mX8��o�>  h��j�`a��m4�3��kvh+�3�D�3~9��6gJے=���Gs���-hs}��í�k�D��5g�
`�H�+~I��<y�z���Km:�4�d���-{�X��2:�S0��O6���]�ٝj��_�:��3��~�F�e,B{g�}sn ��A���C����>��wt��8�k�AE0�x�^�$NQ�n��(l�ҙ2�&HV?7^��~2y?XC�I��ld�7���t�8�4~0e�y�X(�] t�9P�/�����Vz�9����;D#i��j��y�6-lq�D��U����%7��6���C�7/F�sY��6�i�����&��,���w亿-k���F3?����d�rN�)����+�qY[�ynM7���8�NG��U�1*'q�o"�Ʀض@u�^EҌ��dϢI��]F�z���}���s��9�6}>fۀ����xZ�����	����U+�F��.&8Fg��/��� �Ɍ�]�t��W���l_Ҕܸf�ć0,��;Er���oEz�Y��_3��OqU�2�郁m���!�����3FӴ���s�q4�#��^��c���FQ��	�(*����:C/���Z\��@囬5%�K���o~�\�s�"��|�1&L�|9"(���X���3%����'��!ϊ�!Ȉtߋ��������Rm�O���������R23�Yy���P���'��Oqz�$#k�9��{�g��E�Ek��ˆc`QӏȢx������h��e�I�\s����:V/@l�$�u�}�0���[L���'�/�Oc�D�5���I2������gYӪ�9'�Y�?�w�_����;��2'�6Ս��'�gS�b"�i+=ּ�޿�|̩q���r�]�Q1\2�Y�yqe�9�5���8iN�^K�g�
�Z);����c�x�t\�@'�M��c��7O����PL%���%4��Е���V��7;�'/�?),/���K���T�)ɱ�s�-�N�N��!�V�Kz�J�Y�<��ц��V*�h��ҧ�b}sԨ� 6{+WKu�Ne��`��n�����;�H�q⽭{w�����ȿ4@u�do���'Eoޭ�m!8n�@�Q�ΛQ���+��ˇ���z��5ɚHT��D ���(��DKo�g����z�n��T��|��Xrs*�Mi��f靌"	�T򨝌x���&���m����ꁴ;�{e1����bB�~xfRg��R���l��XU�������M��?�fi��4��1ОK��YWa��kt���d"c�c��-�q8��`E��Q������"���3r^��}[���T4.�(6O��b��ۋ�p�[��O�\W8j#���$9���6o�2��&��c,1Qh��.�R�����>K�(��GBO��"ݒy��R֥"d�Y��}��ϑ���(���� ��o�B81��Q�7�C�����/�|SD���Y���(o(��ݫ6�J�F�_ZQ��?9�R��m4̃嚣�Uqk�^�c�:�چ8�|��W�}�x�� �Y� LU��˕6���4t�X/mz�l����}Mε��f�(0�-���B�����%P�E�?9�wP,*M�Q�kq2~�uk�ti�­�,����\˾$�"�/&R�@
�_��(���{D)*TM38�Uq�V�R�K� 6 �rN���d�O��ƺ��z���7V@�pu��W����9�m��)8m}��X�`�p�c��B�Q���O2�k�ÒSbw%qZm���!z�Ϛ'�䫺w }��)4�1 ��g�Py�[j�vk�=3���F���g|�]sW���%uq��?F��^��n�����l.�@�����?�.� �+�!�"5���)�CfE��l��n���B@�t�0�ja�5S���M<>��7l���m-�:U�h
|�S��G!~�� S�E�Q:�Q�7Ǒ�m���9Qs6˱�FW���u�3��k.���_ͩ�q��Q.��gSc ���¿�
����ų���=����_��
���u�~���-�y�ZJqJ>�"��E��E2���}���-G�p㮘a��Oi����,��N-�yKx�5&�6jjh~P�J�R������w�,?�� ���mB+O��.�����J��gh�cW#+�
�KRu���|@gW<8�I�e��QՔ��=�_qjHk�[�8�OW�Wx�ڢv�V<�^�D~A���R�|�}D!h�-</·��p��T#�! <V�}I�`��
�����x�%��$}�@5wQ[&i�A�?�j��L���E�e��Ȼ�x��ʃ��!�����/�G��?��lc�&�>c�D����Cm@�#�Ցz�V�|7�Uf�����7�Ku�w=�o�5��d�>pg�Ƙ����Q�
0��!,(c�;LR�Y�sҫ]j�tdMG���ǐ���I�-������H=�ڤz1NN/.a��l��뜣���
Z���y0I��6�_�f�_�������g�ip��R+F3�ߘIP5��0��)��!��R�^�q����x>�|MB���R`�c0|�Y���vM�Ժe(����8Q ���-14F4�_w��CZ��/}ڟ�n\ ��
 �Ѥ�q�2Sye#b��@��U�gk��a
���n�R�{Bw���m-���i�������H�b������U��P
��R�<]�n�M�����[��=5�DN�顔�$�	i��rm��rTC��'��m�L�Z6��=�x_�+Q"��!�?8F2R��b�T`��Ts�'PEr�k�o:���)u�-��{��I����\i�[y�(� ��ǩ���&٪3��9��ﱑ ��)��6��:�$���#��3(��A'α���mik���p0Q5q;�Ee�a����l�p%�0���Ƴ��}��1���4�����&v0�[1�fH<UX�o�n�a��~`�&�Z:Mq�\/�� k���2Cd�Pt�������qzow��YR':M3�$U�pl�V�bV\������fp!����<�W���7��B1�J�5��u���8#ɻ &��T�D�$iOFa�Dݲ3n:O^r��.A$%�+��ȵ�=)20���?���_'r��Y�@PY�W�ew.�{�y5)ͷ�vyZf=%%j)6,�WV��ƒ6G����:E���Bc��}��=0�2%w�%�ɦ��A�o�n)�|�� D�Q06B^B-o B6��'*�>s�F�s�H��ۂ��y
5S�.�̿�׹>����]�ۓ�ƻ�{h��f��������=P�41�W$r��M#�4���F����5HY.$���E��t8�8�B�2�P�W���90���������������2���/��0�N�ׄt��㭢bC�fds7����er4�yr9hi�m@�����8�I�`KaS�ޢ�r�E��f����u���$̦������������CCJ�>⃸�/�)Z�W9廛���s��Ţ�3�H6z%�' ��X!�3��x�~�-e9���U�)��S��
vV��LYYg�z
�#����m���H	".�#��C��Bqh��EbO�ד�]'�J����k�J|�n4��d#`(��u��=���M�$=�����g�'W�X����s�	�Y�'X�}T2��˺C��̨�E�h1~�Co�B0�n���4R����$�v��nә!x M����a1���Jջ�o�� p��6X�2�Ʒ��^�P2tҕBձ6��dym1"������nH:D���*O�����2iEK�-��\x�4�7N��?2��,:2�B�9*�U�v�D��~��(tə��߯M�8u�S&�s@0yp�_���1?HQgF�E� d?�6�Wo�Mu�`0'�z{��&=�T� uj��ؖ��#3��`|�Tt�����X@Б�2&������K�&��Q_�vhCA("ʣi�~�%�_��[9�E]�D��ϒ�E����/��T�٩
�{���Q-���&��i��j�{AS�b5���1k?O�6�5�s-��I������^1}�R����C�-��/]ÿp�����<`���d`��ʨ�O����/@^-t%�EC�I�i�%���v�-�	5�ҥI�NP�9��TSwowKj�5ȃr�������\�h��Q�����iJ-�� �2ְt�B�����p��Ö�6��²
�20VæK���DX��-v��r���q��?�e/�POa?�,��#�ʕ�w���47�D#P�U�� �����w�te}����Z;*vd^��l҈��nz���Tm�O/ ���d�BQصW.ێ�a[7����j�`�Kʻ%mї[�SkΣL���w��b��^��O-i!^x���ڭ�����Z�5��-�P�d�������*�s�
34|v���a�N����*�H��:x�V�&=��c�{Z<V<���#�o+�F���Bl���������̣�b�0iA�'�e,�I�h8�>�ѡ��k�e�.�kŞ�"�lSKձ�]��.��,��y0�) �gP�IF��>�����gl5���}��b��,�ib!����g�s�owg� }[";1����Z���7�'J}z�ЀOd���5�8��^���7�s�θVt���+�d؊�գ4ԉ�Έ�
P��4�[I�h٩�Bl襤��95%�4u�ΪxY���B]s�a��"���!�;w��x����#�e�.�����6WR�R>�f�(�`�^^��%��Wd�Ƚ�6��GK.�S��b�y�A[Ą��h\��(% PiF��~���S@�Q�S��R��5��/w��l�F��������~)�=v�U��q�=��bR�5z���˖����Q��EX��v�n�/T��*�r˟N3�L�@{�DR`�jc�d8@����튦�G:�o��Q\��$o[�����j{Rt-W@�l9�R�ucbϼF��
�	k�R�>�P��������;p����i6�y�,;^�gp�sg��w���:h�d�(E��!�ҮBF�W��"��[3���ZS�+�ۡ�ʳ'?S����8ޖ�.�w�����m�}Q�7\mH�N��-5���{n�z嘴����I�E�&8�O��jx��?M�G�u��xͽӌ�E��K� &֬8e�:dNsLN��E�`q��|��m���ud"��Ȏ�e=�E�>p�\to�_�$�(�! ��%�ط-�O[6ݸO�1���*������GԊ�����y%��ůf�#d��֦/���=(�L#�����v	�+d�ڇ`�R��l�ö^Ƒ,N�%"oCY��>����BQuԧ�닚X���҆Kjp�k�cM�U"j7�Hղ?Y�wE�)x�@Ht�g����l׺�Ppdq��k?�x�R2~�3��<I
 �	�ޝl���Մm2<�Y�1��uj�z:1����ѥòFW|�}9�.�y�F�Uf	���-6#�z���z:�����.&飐P)"�l+B7���s�Q�8cĠ����D�8YK�����e e"�)���o���_��4����7��@)I�/��qTT�'."r⥼�yż��%��o�����R��0}Y��eWz��%^�$7D����-���!���K�15�Y�JI�iF��� �уm������9�âKb�,0АN��X��{�S
�o,c�U�L2�+�w��ߚG��Cbo�(=��M�ƝK@���;��P �2a-�vB��T�I�k�J"�iX�����ۏu��˳hވa��S��͕SR[� �J)���_�=�Љ!}��wW4�1/f�3	�Km{�΀ٳ	����ڃS�� l�����nP"�&M��S��+����9��y����$	���s�|.B�#mV�f�ǚ!�Z�L� '7�(e6Y���M����nԤ!��-9в���n�
3P �?I���3�+(�&&�j8�Ord� Pb�O���a�k朦�[���o$�Y�V��ʶ�a�;�s[Xڸ�#�=�T�������mdX6��wj5x Ry4��E�7�CҾŰ ?���G���^
&aV�S h��b�[=S��1�'�GP=��w����E6ͯv�i��B�0,��f���FMU�w�� �ƌ͹8�^e�����䧍XN�e�J��%��&���~Ft�ff�b��'�G]M�q��
�úݸ���YKO�c�	u����Е�@Ւy���	$3N�E}�"��t�ޚFY�R�� K�b�Πl3VV��ro���W��/��-�h ���U��4�'@�(��
���Z�y�f�Y�d�hޭK��B��K����b�Ԇ��5Ӊc
�����p��]��D��>IW5�q{em�P3��0w��bw�F6"�v�Tۣ��/;3�;�`�BQ��t&�ͤ�iTox�T �������"=̾����(o�P�$g�T��W���Q�ܿT<V�̄��	�g�՗�$�.Kh۲N���t�D�M$�;�e�C�e�`�nS��V�/Zk��� Y����SvC����L�o�wb���V�_�)B���3Fc�z�̛n�"�94Y(hj}GA����ͺ��1�Fy�6RCpHħ�3ʹJs¡�#����ǢRz�T�.���D��(���y�����n�1j��'T2hs$+x,w�I%�P�U���8�`���gN�*��7���g��u��MK�&�X�e��\����g6K*���1�!Ii�m�A0p��<�^���*�R&-�d��
�(��HBuG9�^� r�����&t��OԹx�?q��v��"]�$��#���mP��쌯��b���'F,�p�y��̉"oE�6i(45v&��ʗ�|U����v��'�Ά'�0M����U�!E)bb���u�;��|g�!#����}=oEWAmX#�R�w�2ەۇ�J߬<$ ��#����<Do���V��5)�H&����U�`{�dG
���y��H/;�,�ƭ$��ēpL���\h5&��'�넫o~q�<z��`�<�wOz�p�?�V�g��h[�0��<[�ë�v�����(g���?��s��/��k�#�S-�@����e���Tl	ɷD�rn&|_��2l���9�8Y��6<ޅG)'f�S��1����^Ӡ��~C��T�`#@���] �/���,W���-�k�n�,8�أ� �c�mx��g�Ѭ�����C���L��W��.�jL����F�f�x�>��^�W�.*��2�]㭅1/�c��(�O������{L�#7q.��Q�#ޙ�l�h�R��B�}TS�p�R8M���O��']GK��2�=�v �В�M�x+���ġ�3@r[�s�Գ����1&��v��f�H�f1q�hE�J�@��N�K�Z�
z��h��i^e?nD�����ÉymF˄<�,���l���#(���ZK���[Ǳ)�}�<!�Ơ�s�HP�� �n�]4\�E��ߝ=�"�}~��I1��GV��%U�hK���'����3n�z� 2!��������gr�3���M��;f���?��t����Mʾ�r�;+���G_-	����(��蓪���e������@�4`�B-�G7絠�	�E��1g��靋�����PD�2�>�K=Ic��5j�I]*�
i*���O�����<ҋrܩОBxF!���	yz��Jun�:TM�@�NL�8���p�g�g�X8x5o>���2��z|͏��oٍ�Ax���q���Ǝ�[#
���~X�˰�P9�[�^?�:WH���u�2��{���g� %6G�I�AҎBH!�\I�\n�~U��w�?��	)I�t✶G$ ���gM����Ϭ6�A�Rتc���2���zyr-0���D���e�a�DkR
A���B�t���,�n�H.:n����pɉ�2'm�gꥋ�Mƕp�鵓jk�x���z�C�ޗ���{�2-;�BokH��;x�k��g�|!��S������HqSXV��*L�G�~����s��� ���(�vlX���<n<���̸��-|(��V.̃dg�cywDhw]=0��{��>�A�$o|��pz�s�H_c��}\���T>Q|v��(u0E
�O,�Ȣ����+Z�T����[�[��!gE{�V�Ȕ@f��g���o5���8��s�tӈ��J#��?v�j;N�~4!���RA�_A�48 o���H��Y��k���c=���T<����w9�-x�=�}��YOr���e*��`L��n��i�)�s��B���*����$��H�G�Ղ����K��]Ti��KTf'�a�ί!`��U�C�X�h�Xϊ����Y�����|�@��di�FP),tf�g��)џA�$:"�Yx�a?y��E���g�Ǳ�/�A�M�v�yu'��>/[��r�ǖ��e�ʨ#m�`4����Yk�8�Q���P���C�fX����˚Yϝo1j_1��n�drϵ����S6�"6}�9������1b�0����w�>�ʿ���7���ow��4!+`v�_z�OVo&D�������B�ǠPAuR}.���or��B�^�Tt�@Y�=���^�F�sΫ��)b�6���3�KOs:xgY��g�*ȈE����v��8 ?�)�#�"@�H��}w}��he>2:�M�jDlA��{�8��s���[��2�|�>,�vr���8�"�wPh�M�c��C���$F�t��7˭�he�Ì"k��_�����dW*ase�cr���ҁ�H±WVس��ܕ��\3��!V���ҩ]	�jA�ٔ(�:��'��O��}�
�W���aկ/K헰܉�$��*�a7�VBƖ�V���j�V��͛�Y��@���|���%��7Q2����j5�˒����� ��2��{ks��2aS�(���;��V����*���rK�]��>�Lvw�&��V�̽����6���r-�\<�8��vf-j�r�8��`�nļ����i:� >�ӊӑ��ȣ�@�/M���U5R�+B5Ό��^�Wrpԛ�B�6�vTd��i���?�0;3Q�}�R���&Sg}&��8)�����ȤpF@m�q�/�nL�Y�vc���P!�|���c�7�K�ԟ�Y��C��@��y-��o�8~�&"�����ڟ1[�9��&�/톫�^��s�/�e�����Fb�HbYy��f�^	4��l��9�
yd�۳?�j��w,	���t�=��-3p�'�+@hbf~��t�pku���p;i<�F^i1[2����[�y́�iF:�����%�
�F+#M@�[�'׋2�
��qklh���I?@(��*"�V�kO��燆�W`gxhG�q�S��*,k��ș��@��T���E��a{�����.�G�"��.j�m|��C/P���E��؈��4���grR[�Q��N���YF6�o�ƅ��
�Ź�ܼ2>�C�+��j��K��h��F4�EI�����6n�m�5�	P�r�OL�Ѱ��;�M��O���j^��)"�̩�o��(�� ����z#�H?�ҽ9�ND��~�p��L2O��ԕ�g)h�;qM�q�5��	�ޔH��
��{h�7[7��Lu�w�����c��kZ��:��8�1`����#��}
�.��M�<H7o�w�H����`�q!9�_���G�V��ηpNCO��V��Y��!F@�=���d�vf�C����v<��&���4���N[��b��г�*���G�e�#i;�����F�ژ��k Ru�I�6<Pt� k�t�E؆C�,O��!�\��N�Zws������Y�F,�Z�CV�;!�����yR�8z{� q��<=�5!Ĳ�`��r�X�?1kz�_M���U[��K�5�}��/�g�� L����E�[{3����s9�G���Ԕ��a�e&N����uMlE͖*R�7����y�P,��x0��܆�Qt��U@�����	�^#�+kEߜH�g���>���:�����ks�
�|w0*cA�f�<� �"E��q�{!fL��)������ӣ���o]�.2H\
ϥWD���yFA��5�����q�)�k�4�*4�bˇ2Q�f�Q�UL���É�!���h�8��C�y�ԇ~b���3�b(�m�4��Q����D����y+�����,
�{��4l�RKY=��ĬlOy#qk���+
K�pɮ�ؚ3)5q#�$��'����W��yZ�Y���r�"��ޮe=j�K�t����Y) ��4�[in��r���!�|6b�}��)��]��l�@��,��>���޿��f�6�kia�#>�Y�ӓ�|�.�ܔ�<d���ŷC�1��Dm��U���EB��[���p���^m�|f�z���>��,ֲ�S=�%@���G\���  ?�
W\7Z2VD%�	I���>�A΋2���N��kM�խ�IU��:.�ic��BN��_�����7�-�����&~$>�#��~*a ���P�������m��E����9�u6�32��S�Z-�M�g��X�,kȋ��i��g�^0A�m�lЍ?6g$�r��a-��J(�~2��*�~`������%F����e\�z���د�fY��D"Q�����b$Q��Y��M�=K������'}���3
���d
p����m)�hx��.��RY��N-��I�����������׋�y�xL8a%�J��;���G�A��� C-��N�b�(
d�~:�*V�nδ8cR���]r�nH`�]vv���*�j5�w��q`^|A	��S0l_O�Ҋ��*���6G��\�Y��c ��$@tX�v��q9N�_$.Q'���&>���q�Ƙ7L�%���2�� $ZDzϜ�Ο���u*�nѽ��.�F��y"�0���MT�����ېs�(MϽtpİ�k���X$��ۈ,5�WvK5ż�qD�+n?z�\��<��Ƀ�~��{t؍-������,�s�(O����Xt��
�����kg݀y�i�I�`��B��G���X��ה�+#�験8���@x+��u�O����ܙ_Yɯ�-C+�*�fA7wU�uH��;P�=47��M��C������r��>G��Bi��D��k�O�B���q���1���{��ɕ	]6iIJ�c
t�,���F
�2����W��v��E%L�xtI{��r��꣥�>�s�( ��4і�����"#d�ne���W��Мa^��:EĂ]���{�A;�5��``T�:�)�w��w���j�hI�����ԡ�� h�3�Q�n!�'���e�Y� �dٟ�e ��ܲ�!�o5k�9�Y}��Ը81&����� ���G-m(D���P���d�2�ɤ�1e����b]xФ���.��߫ y&~�UYv��Y�F�,D�6��/�8�0��n��:i��xBQ�grX��y�g�yW��	�=M�YM�u݅�:}Ym��-LP=�r��C�4r̊ȟj�?4ˏ�/�� �l]� X k�n��U�eP&�Zz�OBN�j�v���k#��6���y�E�"�;�?:_4p����w6�����W��-Bj�%����p�PR;@LeU̳�h>	��;�" &y>�x�6�.�ʦ�ƅs"h�ݭj���g�ȽK��<M�Y�Ҧԕ����[�Y�PB�7�ݯ��`l��AP��Z��t1]��('H$���>���#+t���E¬���x����s��.E���.��|w��5[��jBZȇo.��1��� @���l5�3����]7����8�,��鞹*0���V���F��e�ʤ���� g�u�*���A�u�ޖ-�_�|��0nh�n�&@���=t���,^C"�kH��bBc�	y���\ؕJVl�gZ����|�c�c�^3����i���Y((Z'�ey��Q'7ɕ����!#6/�����u�UH<�5\�1��:�>���2b�.��E��o�(�4��Oa}�(��gR����I�&��7���Ŗ,��"��<�b�턬�̈�%�.H�H�?ڵ����?�Ct�Ђs.�3�U�s[�M�Jm)l�֥]vW� �Yݎ Cǎ��,���_��n#+���=kC�������e]-�EV��ɜ��7���s�^b��N�a���?�9��]����t�~M]�D�30���:K���<�&x\cT]]J��aǣq���ݸ"�z�1I�.[���1�N5<�Ǘ>S�?ΝA#�5�QD��o��%��C�HW��ho����V�^�˻M2RI�����B��t�SU�V�5
� >��ݯN JXY��ӅM���	(4��j�|qG���B	�)���m�U|-e��j36җE��L��Ԇjs� p^[ �4-p$4��]#Qw�P��Sg&!��u��Άw�+g��ڬ���T��BP����y�;_.خ��U�fi��4@Gk�66Uz��^Y���������jM�|W��y�FT�ZBos���|��󘓽��@��MJ�ڃ�0��k�p�)%����L���_)2��U� ^:����q@�[��U
�,`�H��x�(����T漯���,x,���'rH:�?��h�9s̩����b��i���Z�4�^5e�e�VG�n����?@g��*�c�ѢWE��p��m �i#_u�`0U��'�a�U�ڂv4l�h/�=�5:��DB�����2&�V8�1��PH��@u���� �Ƀk�<�~r-�>&�?��gNY��d�t��*b���k�e��j�ZR����}�b'
�IW�`I�y�U�<�9O��x���?��瓫��^M��KZj����x�7֦��i�N�"�m�f�2��|�;ݵ`r�O���V���"\E���TS�O��|§*ȨS� i����{���a��N�eǞ���q��M#�p��?4w�P̠�ڜ��Rh؜N���fұ�� ���O�L�٥A�?D���i(k���ͥ���F�3�5�4�6ol8�C��&�O����[x��2�5P�