��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t�ꎜD7���(6)oܹ�h��=$_��}�jwaM���a����J�T!\8���Ze����4�o��Q����Q���{�*� u����#L:^�q��F��Ny��V���4�K?��*UCB�M�Fb�ϲ���'*e0���"\I��F��c󜌪��OJo�T��ᭉ?U�2���V躹�$��=Nn`D�nʵ�CMέ6|����=�J.k������C��MNh�̦����M!��KBb�u���UjL��Ԍ�ʐ�o�*p��	��>��-½f���g�k_f��"j'H������o;�Xj0�ז��Wz�^`	��Ή��O)Z��:�&	d�py��L�j�̕������w��y2��(̥"+���������v�dCin��~H�4����9y�;�%*�5��I�*��, �Z�o���%�,��x�4��	u�~Q�;�(�i�,�v��:����;U^��d:��uXy���C�v�^,1B���{,�V���7 �\%���%Ͻ*�L�㇫6�ŭ*o��#×f���$��E���C2	�M��!�i����GG&�<�b���M{ �z�K�v���r�E~&w|5��~=��t����`6� }����]� �BE����b�͠���n�BD)����Sk�;���)K��\��[����a?�i_��<)������cf������f��y�����'�a1>ɭD#ab��)L%=Z`�$6	��0Ue���^E����T?�'���Y+]�5yt�ܶ	$������h"(��?P\���)X�h'\��I�vD�\��Mi�����YfA�b�U���?��'L���I����}���TM�n׆t����䋟p1���	�N�Z�}�@��L�Ƒ΋� xL[��/�����d^e4u_y1�c����\qPs��T6�h��CTv=B;TQ<���0Zq,���ƚ6Sh��xn+0�!(�Y>AYL��Ϻ�}��Z�~�� M����W�a��6ޡ=�l5��v~�jA�rD����p�;1��R Y�Q��M���|�n������5ς��q������׼���Rz*q�T�Oq,���&�HSG�f��Z��iB�q����4	ה�N�I�e�V�3S������p���a��Y��=���1��e1
���d���N0ȷ,̖�Kٿ5`�?�>	{�]
:�S��\ش᲏��ty@�w��Y��D��\J�%�0rY@�
�eŁԝY&֟s�ϫو��ۍx�J����ㅸxw��;��dk�s8�I�lk���-~���ԗ|��?}�VcJo��P�B�~��_ ey%�_^o��I&�NΨ��9l*�����m�a��x)@'K�S�A�[��D�����ٹ��dm-�J]�o��89�t<���O��`�K����^tȍ;�4ɨ�q����#@2��T����ӕA�R�\���Yۍ����s�G?��1cءK��ژ�aWX!�`�$t/h
	<˛���dT���{/�/ض%���)�:1��(db��ϒ96�D����@c�7�ue�:�������ì�B�3l�<j���	���,�~)��k�:�Rnfiq�u�g��������w�X6�ҏ�;��r�K�[�t~"�m�pֳd����-�?�b� ���z����&5�Ar��}a����O �~�时N�Lt��|f�p���� �s���}�l)�>lj	�v��`>*�0��D��v�^���\�q!�J�*�YHÉ=��������j��ȕE��my2�y���Eq�b"	g����Rd���ߏ[y&�w�%Ņ�>�xK��@>E���o�#6�`{�)�d��2�%jw���`�T�	j�n�r,t�7w,^�`8����^o�������Yԕ���G��U��ݸe�����.ָE�E^IӼ�=.א�6�5v�zl��_AܼX�!{#��Rh@�7�L5�:W��3�/~R�O%8_<�V��ư!���m>�WVkp
>���l�Պ��`h����zz��D����NA�b@�R�D.���="�-��O�|�t�.�ҹ����?��<N�5�/ʤB�k2�xB�6	�Y�N	��I�a����oI�љ�K�,Z>1��v�[?1�N�@�6�����d,���B�bע�k݆��"w�R쫼1b�V�&8>��(9U������t�(C�Q����������2 ��g)�	�/�e���bZ'A$�0�L}W��
ˇ�^�ҫ�H��Ȇǲ�tɷ�jV3���$f:�7-6�l��~��
���V���Q��!�A��r���
|m�wc�}�M��b~�=E�W�G�$�
hᏣ3i�g�ͅ'Ż�G��7����