��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t���g�l��B.��oW8Efwf�E�?w.�
3V�K��|��ǀ����~��*0�6�H�6t0|���L+�y9�rԬ����Bս&�4��F�v�3'�����\7:i�\w�*�w��'��u���q�*�/���֚�B�a^�@��{g�*g��dШ�:���q��l��2YJ\ڣ�u�ߺ�8)8���̤��+�D�̊��O��E�~2�W�c���b,[��n���+��x�z�ŜO���X�[�9K��R�w\�u��2V8�U�m*�.t��ͫ�2�RY�iT�"��[EGv���by%�i��0�
U���y�x��gx���]�G�	�
Az��xz����$u2JV幄�/A,�p�z�%�;sD�'$q���~�ա%�)}����G�^C����#�v|�S,$Mg�mHDy�	p�'..pۄ
c��;�}�⠕�z�_�%�y�,(L�/p��j�_�&�A�C��o�OsMݝ���ܾok�������{��	'����*�KuFA�C(�,�;���Rb{�����n�ثtVGyq�a����mTY[��ӲӰ�7�;(�6d�(f�-)��S0</'�G)�+�&W�g��§r�c-q��]�7�K���+P�����n����!������^!k&�Z��B��m�*?m-23Q(�*ʭB��YO4M�� V8�.�����
�8x<���61{����:���*��[zzX��q�l��I���fH�����R����7��b�2H�5XY6��#�!� �/��y@R͔%���)!J'�&t>����m�tRe"3�w�������B%���'�/�G�� *���V(�,zS:.��}�^��v0��%�EL�fHmc�}�ك�Mt_7N}�^� B�+�΍[�+���
�o��f�!����L����5���
�Ж���b<&�5{�Q\�����px֑�#*`���g�*����\���`��*�k�Cw���f	7�'� WRӮ���y�~����;�+,b������ئ�WCy�C�U_x"��i��s��au�*B��`k�§.LmŪG� ˣC��Y7��_�fj2}H6�H�1/q0��6�Gk�QR� ����m��c2 �W�9��������Ң|O��h�Ym�@dL�
=<��DOⶬ�+ݕv�/�m���|�[2;y'�.NQ�w�'���Q|��R�v�R�\�z�y�bA�Ip4B�ν0�� �e���	�J�G��/�"��/C�^�oڗ,�yMDi�H��o?��h7�D������7	ƥ�_w5n5J=S�gK4��1�I���K���Q4�$�P\P����q?���T�^RY<��kJze_��Qò�3N�T�<
#�:7�{>�!�0��4LA���a�l��������S����p|F��;���G���6�A;�>����x!8�[��*�M�T'=��'�x��m(�5��XVCC�l{���*�,�eDf�ߜ-���I�r]�Q���8#bŹQ�c(�%o�b�+�����qz c"}<Mچ?Pȉt�u���3�����}cHb�6���o�MVlX�F�=��AG�49��~��@���)OB��S����x�+&y�����d�*'=F����ܪʗ?�S<L>8�%�R|�@e{����'���3j&��o��D�����0j�XL�ޛ_��;��!�u��2+3O
����4f�y��������0\Ue��u�[�,��=4�j>�Dn����4n�#u��͘@2��(��1����~y��H�ѕ��ȁ��Nj��JY3x2���4��=�� u�T~�Z������z�ŅQ���E~�M��nx�]lR[0E4&%�3�-#���h/�Du-��HG�<Ʀ�Q-5��;�Ԏ 7{�Gf����XԒ�*�^��E
�0�3�t���.��JYvh����ä���e���S↉T��w$|�E�`���`Q���}D�D��vW��U�.���Y{&��ژ�:�[J_߿����b��\K�/��5�i%A3���B��J��e!P���J��<��ٖ���]�
�dWUy�R:��$T�s�~��s�xst�柯�x�m;cO.�6FE��˹L��nU=��T�W�����E�]���R",�����2��9�L���O���:D^������ZS�H�=�ʫ���o8 !�&Ĳ$�dNT�"��צE��ƃ��O��,�&
����}�ɻC��1�����g7
P�����u��r�Tp�G]C�} L2sӺpD��DM?�:f��Y��yB���F&x��4q H��b���R�8뎛�tӮF�_@���,�v�;	��{�E�Z���У����@:���9�D1���
zt��%�7����
0f-��2���Tr�w6��LS�A�Vy��i����i�Ÿ����i��z'�惖f�։���p�e��l�3���0��K��;�_>x��`��+��W&�	��SO.�؎'6����Rݭ��3���l�SF��mP!7��%�su`@\�k8�M���