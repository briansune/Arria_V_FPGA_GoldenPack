// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:17 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LSRtO8tsvkDA47ZPdoeLl577iZLinAdRpnmFgrngaROzBOJEM/DscMI8mBemryTk
qfHqWCEU3wesStBZhkbcBw1juxXsySOJlA6lOeVQf5YcOOH3TGPxm3mqY1SnKf37
5p1EQeqqk+ng6wGsA6sYLsXvGcm0qHKXFWFie5PoP0o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
32GFtUz6uQuSdsjQAsDnZULU1bsSQrugcvp2UqIdkvzuZGzvILlgusMgHYfkj0f6
pL6an+zVmfrvRxS9jnRQWqKfZwjEWe+nnlSv6VKOcyhJ2xeI4Dov2kqnJqTZcfox
NpJCgeT4zRpykqalSjOMvn2GtOi8KNbc2OoZ68DPFmMewafBcn7j90BtvKJ1XOTa
llD6dqHjLQwC3eS6wiW0LRfnGRw37KawBYJOcTLEQ35v923pyM0liyzcMWLpEEIi
pTx5IjN5CAV/vHHp/eRnfFP6VXXGbeifyy8lu2/knElRxstKTy6JeTnOug3tPKkD
Nlr2c5h8eIXP0iIOybOskYyp2Emmxxj+0DsXGQw4G14d/F+PGR8/aBwPoUaJENPG
dqRcZ4ki6qvDnX5/a38Zja9pEmAfT+euWQO/QOmwtMQreychZth6+dHmgOgu5axn
m4DhZ6meexotsvIaAE3g6MpwtOLrw4SgriN6OhiDqolU+8kO5IdpJUhiSp3a6cv0
bPRAgYuMspaVi16fzJSqQahKbHc1Bw820Prr3mhJAxVRnVNHbC3I17xqR1UJFxai
4O7sq7+AxwO9FrqS4IWNL8cbYXDDxPNIIuxfQoEgBuXunNP9Iys1vlszgIj0NkMe
TSwFipoMcPpYDXm/0G4SE9fiORbJtv+rRr5Ud//rju7IBO3cbo6qSfoQSfOPa+++
EMNvf71bXiThn9YgbVbF4rhBX+7QnBNfkPek+f031KLIp/YHRwEuXH2/rlbwLryD
jzsHR2BUBW8PH/07EAEaQ9EGAMGThNiTmg+l+R8jyK0YH8B+MZHx+6+P+gQUaWZ8
PHin6O97ERCBS6MyK0E98JX2TQRWLcAnOrBZN6fDD6VCCze+ZgHgsxYLKM1L3Yj8
lRcP+44i5k7e1+QAbS848wShR0qlu9Mt63EteLZa2FG9bnrePLnb8xKqhzuWm6nw
j4C3G3SCvJoLaLkaPndkPPci/Z1CYiFkPaUginR7mH+t1PxcHSF7pw9dSqlKQ479
DQ/s3PNct+m6btqpCb3n8aAFOaCy246BljnyBPEX+mMIf1fwcjWesgV+nQNPw6So
mpfKR/sVVJXZSEhRVtQoGYbnP30CEyNndpmD/3NE1Vo+kFCXF4y7A+H0lsGFyEXx
0akhsHHVk/dJ4BFjqUIoZ6F+Wx4cy3McJbvOtEJBmtMQthtiJDEcYhpiNLPVdNR5
6swd8FKOIC7l86XL0doS58HRoW94OhVE8zoX32a6wzu6m+L5nSVZbFYK+O376s3k
nbJQRoKCwKscGNeeNeazHHlOleSiXg1CqjJBMMblqQ7P/XqTf/xhFwX8Qcwf2+/V
tEsWEiXqMv1wx0484Cew1KPZax4MTGnUeES3IRWZAmiIgFojX+mOQMNGD/oXBlGH
GoSUPc0kJJjP0ozqVkQjXxzB/rSV2TbPSIhdGqai+4lR8LDAKcFWFEPR4absMR/y
+FvQX4bSsNLzbeKkBw/bue3u1KAJ72PZxzqGannajjmNTQIEupAtifQ8GkXIqG2W
g8l+L1VcPVsti5bwjLSvk2+0/HeM7pZchZj4KYmbkuY5uKC/EBMgrdowpS/RH/3P
eOKbo8MDSWCN3qOY5m3cWXV21ygBzYQsxYHCydJG27vWy1TfjYbu/IRi/xGRW44G
OPjjxecF5Lt+2yrs58Q9uMZAWA1XKitrjLYDUSm+Mf43GXa5Ps5MR8jSxTRa5aQS
q2/h03tkCQN+hifkQzx3zioWuW1ZXXYOFie5vS5ZOjpy5srUzmxLy/yElp5UeCBB
3BQeRpTlMI1lJBh+mYSAx1vmWxC5yAR5rKv/yT1X0Q9gCmiIwjPyZUBoHO4yGspH
xVYr/5lONVhWuvcR+JjUOS1SH8TalPO91SjbYKVE4AkWEVPl6iZ2IiZ3ymh30+Bw
JOKpl+v7GndrL9JfDmYRaLIBJcspgk5XOLN7c2iXV0dOj0nN+m9EdMpMANjO3x/G
02PcLg0hAqKao8McxeIG6NFzMQx6t4oVk5oTuhZF1xEOzbXfY0rey3l5Qd+0EH6z
tm+my1hD9qIErUsZwLrOABvxo0Oc8/1xATFj0Dc1j1VFedeJoURN4syCmcltqVsb
LpANcwVEIt0dlG8zjxZPoXykuP/kM2qZ3U1g4fCoG11lOWTVV0/vUGKFBa/b85G6
IrTsg/1PZ4fyKTi5U3HgYbhyVemcf5ShFlVryjDLIjHLugxgdd3CiPS3Vk9QzeFk
H6czxFXrfT6uoy7rwfKTuPHpTPoGRlmjWo6KNrpmX7udb/dzw5VFGnvmFPqNvCt8
x78WSpd5tfz4A3N/dV3egh1md6web1jkJEXja5KuUvmx4XZurcwH4KvywWdCMAIg
JFcwvjRCRePOwWPzbMz65DI6wORKXwK7V9nLEdBLDIlrruPH9siubHN/nuFOxK4T
L9ZSezIOPmmbXwsK5T6ISZasZ3Q+K/9gT5mohhgNzjrbLf8QgRKNWhpPinrM1lx5
vWiTN4Dv9SoCGmszILByhxnVqhM5kE8rYvxOZqUnjHOK5gHnblfqpGvaqzpZZYTM
dLo5569TBnbOy5ZIX7qAtIHZyUhaGLGgy8JOnStbRk8e+odM/xo66/V6ecl9YxTJ
5uojdZu7cS3fPVlKUQSakvpbG0CXXpTlcy4EslrWWD2FtizhTVCJCCKmEouTjt/T
eS9cP+nqUdwWS1EwfOfZuONxGgBmHkYPJ7luOLTRSN0KOLcfunvSBVR+/FmZ24y1
EFNjlRyhIN6jwbjHZFfvX5+VC1AwJZ3Zq40qECUuVRIJ0QykWuEyTWFMTATNaHJ8
1MBOl8y9v/oncQED/9G2DvFQthXYpC8+mXt1Vbn8WjRBO5ZSvz9M/YY9K9wAEqKl
cu3utGQ42HgQXXHmjvkzKZihaXrmwJkr6fm9O61k+btlAvuPHbQct9af71l/Phko
ZfIYyw6l8YEbgG00DEdu309wL1B21bzW5rjjcdltAztUD5e5I1z78IwwG2Wffd4l
XsMODC2KFdjF87Pe6/HGI4CadSAfjzPVfB1tO7+TCbXHSqxgR9UFEAsLpLGUc/jG
lnc4EgvyKu1L8wwpB9pmERNa5gbPAJUyQaqVk2TUdKYr/4Lr2O20NphOQaq6/hGA
sG5yEB/fdC7Mk+4I8AH5TNdLWrEwloVd4mX1w+62p5DISt9OKVMNgQMiE3VMkUdI
FogjRU5UN7vPOSQp3UVil7U5rYznpBnf8CvzpxXdovQYmPmWj+XO/xbh2h7VCBgW
/fGY5/ddajnid47n2GM0NZjTwdwE8Lp/XsTYC+2qA2J9CsXtFTMN78Ju2Zp6xBGd
7h7yFINGGHuD/kq8vEU+K0gY/Sl2SgJ3VcjYLN5TZhebjYq2yLhtBVWwcoCSrUow
ZKBVEUzE2AI6qE6uIIcz1JIpi38lH1kv54nCgr02v6irX/8iot3q3U3zoRxk9KRt
QtfhbbhDugJ6HTwCErgwUfUeKieACjBdbuOk7gKIkISHvNh8oneykxWfE5IF87Lr
/pX36ihTWzvDiuybHjFTJQT/SXX23/sw3ZcU6tCggNYgYTHtk3+B7887FE+k4AAg
ObLA/S2RUt1hK78jCAOGPYqzfGoLhZ6SE5xASGcxDEJvf5EBy9tEvkERBcaeo/JH
tmVgsSZM8+LnGXUZAHNRQnWz1yc5z/E2ktRLHSDzOLrwGckbxdrG3if3uQdmjnwA
qVrV7mPgnUbe0AsP4jPBbeGfNL+bwF/Cr6kNsaBBJvQC5jR4G24YkGWNM4jJw20V
upXhkJPT7SNuPlRNhwoUItXAbY4POcNebFGyqF9hQQrq0/rjYuGnYm1p2gyUbSm9
o04VJU+KeOtw1JGnKi7r9neJWIFGgrU6FzwKT8dzF7BW9exs1ZLd8wudQubrVEGi
/tTNPPRN66vZrnhnByosnfl+Opi4jADuHscRAUSBEPuFvi8k2ME3tlva70LXGePC
DFDKdS43UOLpW2QcoEIQp5SfOoPJkFvjLWv+v/sDJhhamnnyTb67PPwo3EKbijUx
2XQ/awfGC+dgSSyUPTzUYFG5MAbldRJHiGKqkMs+L5QP5m1LsHrYUEKq9NxZod9T
2WhXU+JrvXps9xSMUjhG+Nwi43f3a/9EYmPT1KvknAg82ZjbVct0kE57U86b76Cu
R7fWnDo7C7cORZRtSD750ii/2XfaVrDZTsGVUjDkR0OUi6YbG6NM+kMtzRc9m4OX
NfGLtUbghx+TR/RxxS5w8FJ6wSnVdBqm9D4zVLL/PZSxqMKUUNgxwNXO5agDiw+U
rfyKx2GmtETFFbbZJTs7sY5V88Sl52M3Dt2JIkhms5NEGArHInBU4Jq9MExNj/qM
wOhwv1mRDhcaoOXqRfAnsAGQS8ZIOWf9ALx2vczNQXoLvaDjVUuOWikkU6xUhmGI
3uEpajQD3yker4wcEu7SoMS3xNzr4yTa0DtdLwCJcLjVF+hlE6JR1G9pKXcNhssK
E+97+HvJ7O+fUN7NAb4CDAufzSXVbyKC85C9/ZhX1pZdL+MBajI7/QjnslG/thBY
em5IvMbMjU2XF02mucQnyGezUUBeSsabHkiQwuNIeCGp/iebsC8ih+TUpwdnmU3Q
f3++KPfGixnJ48AEYkX5NEHVEbZ9UrLIum1XJ6117k+Q8CKoXTxGUL0XO0ZRR8/1
29NAPVpZb13IOXmCBbFFNI44uiyOvzcEniVrj3gQ/7JUQ5NfytOlHXS9IzGKcjWF
rxurhhTBUFtlLnj0JOK18ipy+/ttXk0uU03GmqsZRlU1HTwmsvtYNSr1otoa87p8
/TEkGcQf0lLaltgJADk+hLdFT02hmm7+/npE8Ki3HwunoWpnF8qbXKGhaCs3Etn9
liT0ukVH2hFdpjecvi5iCdKWOPsvwlmHWvS+rwqcYRTTnhtVu/CKWeFOKLU7TSJZ
kbzA+3yjN9+ObtePiTS/D+TU1ZDEOtAlYBnGFEM4GgHLBcNIcLwL2UA2bVrtVOmd
8Ug77gfEmpF2jQTG6cdyJvpxJTJzyv38Lyh1itrB5yRNXQ86F3Mm58OP0Vxdd6HU
I2+xIiBOI0edlDwgFWMAS9qVGIedaIgCzyqXxptUoxJ/jKsgvcViEoxmy44rOCyL
8rahfwGLWIyeeAw0VdAoOys5tAOnrvceH/qJ8gshHfhsMI0Y2F1P+W7o+6+NRIRO
dQKr8gK4xWV9KL0vhNpZ+0w2hhzITUv3yAzYcKIjuW0gJPey8uClRnDr4TGAQ+me
7RwL/G0bdou6XEM1l+HOICGH0oakYvWvdNWL24C33YQ7ddyiRnEdh2GYTPTeSXdA
28KTcrWLhywyDQ+fuZr9lTWWo/SjlJ1Y3/XL8PVRtfaRgC9zNRQqFAKzAVXTdKIg
ZZYkHCMexcx7HQFTafwo8wUDzex+AMA5mdvFjcMJLNH15OTw657Ph61DxP7oRXKz
16J2+ENf/ENEaUKLmjAJDezwmYa97p3n2If2C/9jyHLBe07XreJ+ab41ML6Aa/Hb
sP5bLVrS6kVucgbfJgpX7rIxUiEU7htNSaidCzxNEtjHfOoX6luslNY79QXd8IsJ
QwuigkdjLRnO24z1QfOTERfTX8pZan9N47anQlh6wT7TEVpyooMgUcEZvTifsGul
Ft6k8HQ4rHyBmpYd69ixZPoj4qNLOlq7xyJhYxoFcJqE9zEhCIhmaY8Ck+IYQEx2
jYy5CRJZnUM7/riq/OUi+8aGrZfOKd4KI0uq/SJIyNFWcEzyoWJ/kxkRv0IL/VBN
rxNPUoVLabYfyh4Ewgc15w0uCjTk3pxhyt1boZnnFEwxp78jgjOn7Si4ILGgN4Kz
ittfnhkeQsbKcjPc3GA3ELsGiJ6NMdBHaSJTo5N1LsvWddTi/Kwh2Q1cl06J7f7u
R6OPwm87BaM0J9ztb+OOPJWAheoGo/DIvjwpBvQK4e6A4+8nbZy1diTFWcQDpSNx
aDCZSB46pH6rlY+Xq/K57dz1EtpJklTTua2WyvQQArj22Xdz2F3s4BRDtKR3Pwgh
43YDh9EbgQdAdSu12haS/wMnMV5ObLz6+IuRmZsBFmRi/HRTMFnD9SFCK6OoeZy1
dVkubzUW7byqpG048Vcyzt4DXafcPyb4iNj32/iobelV1UYQgPmHVy0JhUIo9Vuy
inWyz7LjDRTOkl+brD8JXT9D2sTrMiXIx0ex+ijkVAHuYlK9IuUqrziZWllApUDy
LemlqqcsGwmGrLTgafywpPtWnobKPaMfZkFMwhYfKeH/GEaIk0JcTQJVqX9DebHQ
mRNJkNdKhkM12Na/u7H2NQHxKXtWamjAtdTCfHNAg6wG08mUcpDDFcDol/dOcocI
Bb3F0bHSp/uHEejpntXyahAnga9+3FZoz5CWIMzQSZe1BqnPgkSO2c+dRp02ayCZ
9uGWDQ6q9HN7RppArAONy/XFaL1X4VTxSLzvQkoVSUhUYDH2wywWXiE+WVFwT+x2
dIzqJYXN4dzinN/HREaqXCgqFyAVFXIC/dlCZ7B4/lCC4ytAeMUemdNUDFB0dCPQ
XYG1k4drbzEL24Kjrdr1yWIP//yp7weuqqhSDaf/WAP8QHVB57R3ZXZZlmmXVDZG
i+VNhl30VekvhQPI5R/FoQG4CzsMlFU6hDCaUVEVkyGLeByqPwUqxLrPQkso37cu
MgODCaOCouSBSfqiusQ+Y19Sgbtc6lnk+psZ8xEd0BcUdbZ8kdDYysaFRyHVoCCz
oVlC7TIlUoYsbbyBpCfDm3esLAQQd0vdB6twqzpudDQ/Pbt6Pxn8es0UXp+q6iYM
8UH9v2x4Jj8fptylRs4d9DwVd3xyrKfJ1EcuE/34fbotfgdhlUVeJ340SP5q8f/b
iMD5tmgzHB+sEe7Byr97CkCet8UwXctwIXrKF+O/KL6HCZNM05QKELGOEfK74olT
L6YRYx8V2izrfggEvfnCJz1MXzoHONt0lmEfvvfcMZyyhO47sY5axHDMmlTb8fRu
eSD8OmtSBJ+G6K7QMSzecz/w+lbNrB8LeEvouOxxTObwNcQsxJTJ50zkbEG+6DNu
0bA33fg964uM48SjgkTuYJ8EUGgNs5pBEP8hUbVXG8niy2taIACSg9m6sl1zjZ72
VP8RJg5DcF2faidJ4SJFWU6rLC7u1B+IPWmwUoDcLQ8B0EzEK9vlpsarj7+u46GK
pNYQu6sjmUaiHKcuDAR8qwYU5TIwATxMcrlk6TT+d6khgJwp1mQl8VDuQxNqbNu+
4sdSeWhtE8SrS0sgrq3H6QacxKxDms/G0pok2ZHx/eRfdAD0fEc+HIzVuLVuVFZG
aM4oPBCnIa8n6PDe9DNMt5yiL+SR9JPF5qSe1/YQYfkd46VsDqijWyr0TzIFF39q
N4bD3safXisLkTItF5maHl/nczSJlBUgrvUdTJgjucjW2tSYidi5b8dNBRgo7JZ5
IwfS24G3rKsuVVHXDXxGr9T9rc9ePqg4nCz1rKYVCNcvb5QMdosg2U+va/0jHHBT
srRKx6a1TXHoITVXTL7eMziZmKC3s0DVDQfZWIbQNIQ1lLS8V7mg1zJbrs09tbPO
C7VvVsoa17O5TdGyYKmd+/qyGnEmWj5pt6mWa8oXP3yoB7DBFiT/JpRwkdK7Acpj
fSlkt91/KnYAa0GagSIz92ocvqvy95FgfSCjm/6V7Uj6SQjVRu9UkJ12H+ZqnGyu
17GxIcUvJJCI5ng/YANjWeRflRXmB27Xycs++ZdSzUs=
`pragma protect end_protected
