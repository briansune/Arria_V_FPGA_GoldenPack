// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:21 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C9hHMfVpR8nzRb9bEUv197MtBZy8P3FD58CMbsIsGE5IUd/JB8QodPADP8oT41H2
Pr6eWP1kSRxEQtUEBVOQzVhKpVYAVIPinK3gRANuPva42j63MxuRoEmwga4eRJuO
IiptaBMzLQWFZGBZveUG6q2yC1lS5SsGr6xzcu9SFgg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
/nkWULH0UgBMWaiVt0tMyCKimY5wlbVSpUHWSaqI8sMMfrMezNGRk7Xi9EAWeSkG
JOVYJKMs2+/tfZzCs88Jzit+U8TIwD3G6kMlBhrTqoOw2kZJtjb/xTSXFsahX4MX
yW7IaxW0VxaO1SVkJOnwDeZ4YDraAtj8odi2NdDKP6yafgYPR76BrekC5kVgEYnY
dcZiyxYqMtaWPIhOd5KQTC2dn/M80C5jMNBLXYDLZg3+bhjlLn/JTqqFgBYHe9ea
x2bjNMS3/HgV2oWxOs80crVwrmyraPOWIn6TMXnLYdEhr4mY1KQ5ztmPIPWlIuUx
CKUV6OY1AHsCMUNPBtlBd3hQKW9RioAl9YgNp6ZqjA2WQLqt5b0+80U+Piv8qNg3
EQmAyqqmNOVDfmeUioNBqh+cgR9b9fGKrEts1xnNcfRk03QdzCMivaK7eWF3dRcj
PqiRE06ozu+sTONGTQq4GvEfYqurURMKvbw1/I28x8OQpFdVyoV/WhP4E11ErpI8
cTJypKkP4IEq4ZvzC8vwUaMoLxfdml1v2TuhlJE6GQUcP4a2LyKm8aiLZX3QgMNP
aaVPHZBk1hxpOCS9N3mFMJeE3LaepPbzc23DeeQ9YhqNoZiXonnNbFbywquw3kLD
piP2PLXfg4Bhreqba3pBeexHafwDRemsSqjrL7FmFol9tdFJt7SOfk24YweM3j52
DW0C5NXLy9ovoY7pl0MYJ+U/zzZv3jm0ou/3wxMhR7PpTEog/L/YdAPa0Ftw/9gu
VWxvoofpXCo55aEav2tqdoDIKiJDCAuTAPnx0KjmpCPen5UCzdFRaF2+Zhqy4iDJ
xk8B1M9/jmCQOI8Naz3Ef0HDzu2eNT/nuoxlqInd6m33kX1XYtwKyxqRDH4LdlTb
vfHT9w2zEhW1gRM5e2wL2NiFKIroTxIHIYoBlfPwtF9On3R5CP1HO+1UejOK887m
bzeUwDnt1rWJHIwEphZOXBDIvbufFuya+R0wxIIOvCWG6sEqqv74fQtui1tvAmjN
y/nY/E6fJQKXvqviq/IqL3f4m8p+VY+BWVxVcqbxLWuQawSUbkVA7fiFavX0gNhP
EgvHmaO1fIADBp6Y/YrmTM9omDYLIco13OCN31EYy4CudJ0dOTxyE2WPQRT4bR8q
c5uiQ9/HTWE0StpJ1k+iAkZ082Rwtbn5ftCsJm5q++PY6z9F7cQ0Okt3QfJ48oal
qUPh9H4+6qygH3k5MyT3hva+lpfGnVH9Q6ePlRUod2KKuxji8LnmV8tGzUa174DX
f4mRPxJaEhU9eWf6CFae5DsQpy0s6toNMcD4XG5lF3dRY1zyp6YpcUWbFuzJa8EJ
tNOA5fKdOGP2R4zCTd2SwIrbYUXeSwfI7sCSWwn4AL6QbgrGvgP20tytjNag58bw
3nrEPI6NZ8r5VVZCZiLe1Ry+JXF0L2BqfdpHr1MbdsmPypK0IDIUz4WJEK5GUAv8
C40WV8EK8H3xydWID+Sc/7Cj2EnszaRODa37cQQsnPAiR1rVXF9Y9xm9/CoKLY/8
KPzPOiLsqy1xkPgcGWJALXxsSqrCl0I8PAzS39Om2ihuXK8NJYQiTk4hOkDjPqt/
JPtyzFwmjis8NQbVDjblAmm7Bh3ecdi9lCr1m3y8XARmf65ILFEG2Cm8HjRWaM7g
AXlGMZcBis2ij1sXIOgxYix/VHXFTMTzAQZK5rERjNTgqjzlF8/yJYkvUM0BGxU/
flvv8CGRj+DJg5HxRdqrqGq1tP3YKUzl/EUy2KP0rmBb5u1u3XmWPv+NpdvYXNQE
aWhZawTSlVo5i+I58lTw4Phl3Uil9UlsNypRxSYcxo4u5DIKnslXrQ85lV9/KkNZ
MdqmKVsuXQrTPnEuURwy6DxCzw7JESyhVDf7Qo61LH7XUolj0DDHdIxSOVRYaJBJ
FBMBnGhzoF9dCbVickPz0ApZBOlHf+aHxAcrPzSl7YCnn3UMvF260a24aCcEWIGC
AeKniAqUIpV8RPbfVkAMW5UC+S4RZTPFpewAkIvTks3yPtPNMzzPDedGR0u96t8W
oXvtP6QbM6smUvW7St7is8U+PXMBni/0xay+V8A2WEsWQ7/ZTRyXCrOpuCeJDNwC
7Qmdir/5KY66AbLKO6p3Rh8H2NslVjyTAY5kleR7HVMgXgk7Ry+2m8VXr7490V60
Jpkw4sYqJDY4UMypNqo9sbAmfEZ6tAzGUMlSDs9SQB/aqyPFWvjRE3fL1q+2+bQr
RQh+jNYV1i5WmPN6SpUN57fQ3lT6m1iH5oafGvpho3x05JSomVVjccIRbt1T/dDU
JDYpvSeTAJ83FuYhSZSq53m++0Yp9o+i8rSjFbHq1jBAsc6o+mJbcj3xprjOIbGF
v/pN3yrKOCOW+SIX6r0O0NL0YqjcJVOOB4SE05Xg6xeiPiF8h3REL/JssUIUOQqR
REuxjTsUdVEPG4nLFezBANsVV9I1eyjDx7jwp5QR0ePIa6W+e8honhjdjmqSaK+c
DaNOUSpufoe9Ih/O05xTqXmBGg2ZFIposTccppiUWsPck1mLVxpCzrdFlJ1xxP8T
WmkiZQLo7c6B3duvg/ol2GZBX1by841DePYvGiC8kneUasUcwz8lbT0HqYL5UZVa
xsPIQgMdIxF7zwTo8XfTugUAqhT/tD+UKT3Olprq/wYd1UtyWSdcg7hnQWi1mXlz
0Za4j/s64KcZ9KEUKtWuu/7XtmO2UDdPye4omye0COMDkWiE6dZTKXB3bJ/2bXRF
ccgrqgXV06QyKHnLb4+nWQMjkuC/7rcSwxebPA08L1s/tGIZV0M5ktGL6VwQqaAS
2VImSmDjGTEKWaYIv4R12+PfXg8eiA/7t/LF13yWWQNCIZUBsUT7Eh0eyhowKKjm
ZBpNGJMEiJ3u6jEXfDDytPEII7Ssqz7YYykM2QyV5ySM31nAURBfX917NUmZZVyn
3zmDSfAnRI6UgwuLH2GhZCSDsH+776DWlWLlG6bFoe4pRQWgOheJGPrZ5GbrasoW
1fFPqOZbF+NvZtUKmyplXqx3ndtc01gck16itVUvlMIFFVCKUQ2A0YQVHozOXm+6
SIOh4CXJpuqmrC5M/7QqcxwilNscGqGq0FetNDx9WpGu6C1+RGsMTyN6ltif6++w
yp40ekCvt5aVTfIn831zD+e0qRpIVLrfkOJjLJsT7qlGyl7kKmUfsZAmsiW/aDL2
6ErOo+Jo2twkQfO053ODsFewNS8gmXkfHDryFx84z7FdjPbq+4dvj5+T1+CBwCZD
gUHnhjaJQ+GPuhAFKkv/I/XTz+iLAZsIWtXBt71dU7tjC4SXhKFawVnzSBbneuBq
PXfUzY1/mFNV2ug7FJG7e+M3F1ibbmfjQ3XO2ekVLX1q+VJfCm450WVF1mbZNnWN
aA1Vnjto4+j6WPr8sqpT+CF8Xmgc8oaWT+12wf5Xmmg4JId6tOk7vHdQQ7Als7eH
Oju1S7XuSjk9wCYEItZka1VnMzchy8Qvm6taOADiNDaWhUKbnXBsDNpxY6PvdKFz
1XDP5MZ34n2SdDu3TW4G1GpMoODZk1PHiCoCe1w5KUX7m7jOW9MJw5g3iA4RZ0Uy
eoUDFUj2Ou45tKty99N42FWOkUwvmelvM3vdG17+Fv/Fm6/y9Opx0gaPz/g1C2TQ
ktPxwapxqOQq+WSwfyOZZJYACyUwUi3u9j4csjciNAlrq6PnqY7uhAMQXXsYmFRc
mcXiDUdnWb4sc7YpoNZ/TX07aYJG5dVZztuzabBL1BX3BYVuXJJRpYBM/rQgC8JJ
QVrsGhv1ATGuCzAXgNsW5UnQpAUZsLPWvj9KHZ2bvwoIoHj/Kja6givBdaMc0Jlv
hfQoPnI6TLOagKFzHT8MLwDPLlSh4rIY4bbH/7DJL/FBdEcQDE6CxvIWYrsftULM
A/5Pv67YmcMh0aGPFTAkxW4uzDhQ3/4dqMAtvX+2T3yCv9NUzUuL4t+o4uJyISH7
ivh+bcHaxPOYlDWpRRzfRC62Ze3+ihOeADKdQpyZ5hVujWoAbiLOzpTWAHov/UaQ
/vVtSuN3eSkIWdRYB8LwO+g2oqMxqjcjtKfy2MiGtWHzPyC1UhICKhsv+0wjsHz7
nhX8pZfErCylgw58493zY5ha0wXfc3v4UnT2gmUUeg2dtF0C5Jbv8WygiFq1SOI2
1FpSkfwuNaFzp1vpyJRnjsKK0fX/ILRksG+H+Asvjpumgn7+yX2tV7RQB6HRA4nY
kw4RyNd/MXY9vb0+GXD4dLPRD60LlE8j0z9++vnUtD44rH9reIKDbqT00DuzOktv
DKuOYmtpANxKmqGg54cQoALyFatSWca+UyGv2qitYSx00HdJjxQRG31N/LpgbwCA
1n+BYnPLM0qRPCjcFs/AvZHkuWHkkMq4e/h6NmWkcnie8p8dNl+4/sFrdz+jXQiM
6kGtVS/+juCLfIuLu6r2qRUUmM98P1DUsJeQYG7+RmXsnLRANTx7RZpagmepEcrg
AlbOjsTFY7V8lhWrx4w1c0CCKHDpEHSw/eif71Jnak9k//1fCWdYHcw4vHxJY77O
b4o3pQB07/6dE8SxrPE4R03NL265kglhkgEHvG8s0e/0eGAUf087uM2cBMlpn7KI
cyh2cT/yckdm1n4cszxXw8DKE5TjzqVjFWn9HHlRyxzm2+yytd/yP19v9fkh0V/w
WxB8kQAzVGNH/owS+DA8AWtSCTArgRnA5xbJzSKSmek+5cauhsGHaz/6KPiK8VjY
VGGCFZEWplptrOcYvospom+dQ+CPPOaV0Vh+10c/Kd4g6riWUMbCZwA9dc1LWBF7
NfB8NSOtgk/heCG1pvtOKewVyj/LW9g/patgRdGS+z8v4y06/Rmkd9/3PujEFhj5
+C0ODkCsmEcYNiTE9p8jbWNubWRrDTGfu083QHjpobTOPyp4zU4/aZENmbkdxqFe
0It80io+OZYOoybkfEddUfROvjAtlFe6T04o2yDn6OQGq2gBSRbatN/SUCXXOl0S
f5UzJxzfK4GXm8lR4tFBY5G3TL8v873MxhBNbQrraYmUfaNW9UhMsAxikxkRXjru
EjRaInAH0LMEACoAa4qJDIKJm6FPlKsC5E77MZ467yfQCLe4Kf70ZtGW9VZdGhU9
ECcbZRZ3PN1/wCd5pIKNbvG5jo+lG0pyy7zwkV8dxZfTsb1sHPp73tHZpkh5PLIK
UJo7TZwuHmYin0JNHOF/RR3QLW+QIgtEUE7PzGXFPpzlHDgs5tiLrY2l2PCTX+x0
os1Oj7jF8Tp7RD0giw572Ep6HdOBTNzmSYt5e0aKdRQV1yv/6W8urAsBXRcJyaku
HOcVLMc422iz27Qu/2jkkGyDoF1Go2qbfBbFZw6gHriUGgpH5x6AgxFXuzhZ/ENm
mTl2MfFhDrm2M3tHikMeN3PzZGwV4nBPrlJWW5j9MPbJYbGacN3J4iVloDQbmDAa
/kxCofM7s8yGLadbN3uqLoIVld6WF+DNHZObRootYIpCbFrVWvvLyY6/Ek0eZvBi
7GfRRmMWq49DagJVfmHmLiiDuLxVS479OWdMlPs9a4X9mv8gBYPtLp1CJ/zKgR7Y
DHIsoIS43HGQ1/LjGflgd84rXruBa4Chg5v6fpyVzIo1eUSIg3+N2MNDuTFkXxST
I85m0CqPCAWk8554IM0oPBsan7ho0e2L03dPqi/J12oidxx0K5kqt6jOi8Ny6E7f
zmHsRcyDnqD8NctvgA0/oAOxsHBpOg4L0y4OXf0VPEKu7sPt6fT9Z65K8c/MOKdL
JuNjwRyGtheTrBvfOFZp0Uk7CKuW7q3xBTHoJ07CBRmBzrvSxwlAr9Ph7L/MpzuV
ARakaq6rPzUxv9AfSzJnBJmonAN5vrMlDK7gT8m71eXXiwSQY7eiisbtaoBgh/Fh
RnsRIHGCrwpHfNECLObzuI6zkYMfiGdj1EvwX7LDtlJs2kBuGYsBDxmKtjQDqkIY
sct53gdiZbfQltxEFXMLcgx4DjV4SftCB0MYQ/8hKgEk2c2TwZelVZCrMnsMKddQ
xqSf1ZsXZ+41QqeshEeCfMqrH0cQqE9b3dsE7tXP1wgSAf0b7FNWzxuRIbbcXtM3
bNu5ByFGuf1jB7ioNRT2cpgEkdBt3ZJMU0zHC4fL/A+8xqQAvVD6clJBT/q6GPZw
a6RDrhg3QPXMwZihNUemN09SgFSBOkCzaoii+2dxWz9dozEKovbThbfUlobtEinY
duR6oGj+b6NsJiJHhzPCGZdb6iyz1mxtNMLeP2dcoPJVkakCx103Iuzuw3Ju85Bw
seI/kwH/FnCrOyw12gvYWwr3nEqfbMOXThfbKVYocx3Qiy3ATaFKoYKtYJyWKmgP
8dn8qIEMnh41R7BlJtzNCd7Pid154oFmXiz+MJAKNCEv12tv7Ao5aIf9BbZJAGC/
oBxzg/NiAZ97F9P+MeSV0Q5WByI/rLWeMm9nl4gdz2aMhWP0jsma17ZVvBBAqTqd
cfwC/CCK8efxvT+jaxSyYTqIUzKTe8iG9oWjJ3MMFsDySckUm0NZlxrEZhoUzGq9
J58xPs4xiweBwHfq2WQhb7Av8BnbDk07E+vvyfZsBBLwZeSe/+ZCD9GZ62iW0CiS
HY8xhBk6Ye++gdINq0o1qQHg3E3yeADa49TB9c+FGcRWSV2qDlout35EFu8uUhTI
hMLy2LFMOf+CQCNtMvHFmBuzZSHuCo93H3SZkPPWFBP2QrCiystPrLnkQz8wOJfs
ZAxnXLt0qV7xfX5UKIaJga1hNDd9P/95HtGT+3GxOniJoBHyDfx5DV7lGGOOssgM
rTAKkvnS5u9mRUxyZhlsAwl2AsNjmgMTPyMHMLANly0oJxiVAoDe0tSyF61l1rQy
Dzpu6y7VoWYx7lEGO1NYmpxh4gwkp0CRpjtMRGnPnaca43TYKa5zLfPpHR5WEt70
BZnvK7kfoObYVaiVhVM2e1/iMai7gmFEQMkZJmef23+lhgTZ++5fduYw5HAC7v2X
Wrs9Fb2lfK/F8NR8x15vKdXTu4iZfBXhq8QyiDklWAhRPHtmt/x37NC7ELFUVupr
gZIJUVYEFwRXm82AcosPhSKB1uqdkkdVQBffIAEmyH2hpP7nsx49ZCOwdxxBjHC8
8GNs2EjrIjJYbhB/nuOt0mbzGliWObfwxyuhI69XqcNFovHmhAtxTLEbvU7p7w2a
MI0gfqoN05VpErCdtNcNdKZBedolu+GupDWgQL9y/WomFnQcRlY/GM2yLe/NJVmt
+C0MCmxwus6ZT/86oP5u7zO9XzDlvcsdzMOLbXtsbXtYlRUrzpObk05bJuFgIzxb
cVhoanqgMKPO0ICwbBRKIb5nP91u3aH5+VwfDg6kMfl0yojvznxCauEahY5SIL/d
9HBo9TF1mphPiU082B1CHqflG4awzvipANfBKI+b9OBi8kmv5QTL2LO20mdPkk+A
bt20c2POx1H1s6WwQSAONOo8EPvXpMLRtId6yWYa6uY7DdedsqzeD3yY/as2xcyo
cbyg6INfK2dNiC8PfmPDt9EgazoXqQG1W8HDQoHkOs4sS+VRjm2pHh74g1/G35/Y
9DR44hdLhXFiRIC37DejJFxYEo+GFTWikBWoyIC2Wgq7jC2eSK1IbmS9KeHelQof
bgtALBeynwkRmk4Zh1D+/FSkt7iAHXwhK6X0cnStlNJ1X2vfPEhbyJ6yzghqPzWD
wXFo64MF8HQAfkfCoQPUrQx9MVAy10zJH2T48BbylsJPB93OTy4KMaD1kfs5gKST
J//YcW+UpsnEG1RauHLkBdsGjtmU/8VHu6bTy+FmXJPTQX7xA9beDdbTTGOEZyh3
5YIm64vjAqT2PMAOdLuAp14hnTCcgdHmaM5eUsbi5mwd9vnqteeCYQZXE3Q+Dejp
OqmHguRypFyj1x9LSSBJWYcYBS53mMa5YlQIS+gGleC8kWL7kURZL7udD7KoW1Lt
9msW9EUXnxbs37T9vlAySIxy6hQT7Fgtv9HS7d1Qc4gROlUav88WJNIh8T/sv3ca
Qv9/eqHcFSg62/TcYL8Z6VP+yt8h/DIZfjITiSomcHZX03MTMuim7rHXtmY+mOOn
MWkPl5dJX4Y7the/K6phqIqTsKkDlchrjdDNEY2n92wjeXRxdc1WQe/dpitJ0XYS
MAX9G+h0P4+dY13wX4pT9HfA+T47JHcihIigaw0IjWxztSvQ5lJL+BLe++JBG2uC
ilMoMZvE2J61oou1AErhBqCrgLHFxOrMSyr0lx6dG2EUELzXLF6nf3zIAAsCveGo
n6ZIcaMmPpOvTec6q91i69wzKwuV9+w/Wn7SWFQkTBdAokvaou3YSEwWtIj27tHb
U3xWq66LiIZZF7dajGtcUrnusNe65OOjv3/y3gnjuGJWdnGtedOj1aUkqUbaNkZ2
NZIiJY4BAywfLWZpunP60aDjfwuQw4qmIc0mB+DdwoLtxPWDiVLFVZE8fn4JNKQG
r+HmOT8YBX8pnb6TURmn+huD0RRjV6dg4gzW2yZmJEjHzQ9uGBCWx7H6ZZUk9lqL
mwCLFMDNIdUV6xXh+xxB3Nc+pzsTUhzxW+0uGskglVq56hMdn+fgzfIPoCNwNe5X
QYnC+WHw5FjRQFHoFMPxxvyt62bba3jV659cUcewSg1zDR3cB+aDweZDpca4ZMOl
ZgZ+gDCrJ7usIbQ3zKVLFe1ucKJgkkGAjXlFoGEHPsPwUpAhk8HudhD3TifVRvkk
TbYlrxSXEjQrDN1kkxAJzRxjMt/jnddWtjSK8lx3x19JxVbBcc3gJb+EMGnjpEsW
FkvBUCWM6WBY46KrIQ7O5Zljsc3cmSO71iDU7y3kftnM9Qirf3e8prWUCR47uryj
N8TA/KgFg5t9R/8sMOYrAGLBJGQ+2yUimSohsvu31y9/HRnrwZq06Ab8TN5dzMr8
1YJbTkHcV3T6Zteo3IdOF80qHFtdx7il/oomoq8m+vsoblDAnmOD+hIRBIbsHljy
npXSlmT01jmDRfOfhptLIcAMa7iSYftlYii7cN6IrvaIUUp8s18JEsnWpsHNz7lr
qSoS/JVL5CbRpVTv98nmD/Wchc2AIYCn4oZMvaC53nZLsiSyIzWaZtKIFFI0ryzE
whxIZanP2rsFth22C2Ju3vkTVJXuzuewRzx16zzg3E2hvJUMLyq6FqZ2xGCMBvzT
wZQcz38jXC7qSxQsyhd5cpm4BGWK8zj9wUI5m56jQLcaWt/PDN6DP0stbvyhd6Kg
MaFj7grYYSZbhciAurPtQza9TkOdlPH122FW+PENl7QOYybyC9a+WuLOYhhwuAwr
MvLB7TLuO53oMivA3MIRPiIE/FEcSNUDdoXgS2HUVHgbqAPLSjTHgxJ/qZ4QE8sk
eOR9CHA6lYJIIzAracDQLfqn2Fn6a675wvogC/PNhRyCYFu9GYcguNcBAg011rA2
bZd/DGrUWs8eU9TDrAmdMCWacan14SdZ0GbaK2uDwsxjY2BEvBmzpoqMv8k8Ob84
6u9pvTM4Ipkp5YQ4OVtvbzlN3YecNn7H2JW5QknYKAljPLg0QeBNj6T5K+8vUFzv
XP/X2wPjEx/Fvmo/sViZUYaosNrM5ZFN9Xpp9KrtMrN8OqaNj6S61cH9Af/iGtTF
KPfxoeOMFfZ76Og7/jo7D4qMf+SR9S4+WudU0p+/lVUn/rpWf+JEG3YBGGK8SR3h
SStA2ZLntM1tEQvBzvkK2aMt+l0CMf1SPZ8TDywuV79IYu5cncJF/NVkioNKPtY/
mYFU5kMR4XQfCnNgCAOquoG4teMt0oXw+p9/KeyVwjTVtBQwUpENEyD6X5/1INkv
LgMre2mtkRtr0lDuenlWGFV3RScY22x/BuKSzklRw/XfIxydNbKFE/K9mQ0Im9NU
6eg+nFvpyxLig8fYop4LPDqdZU1zgUT5ALrH1na3tyeTrEAlFz5NtMn6G+m8ZrP4
SnI1I7uNolCLi4pkR4I/9aHcyerD7B0DKn0rLdA3E20xK/vFUwW6rh7kU3uL+9D2
BQmfGnZriWVIQ5PU+KUJai9+CAcFqz9lOkdEsH5224/YiqMRw4EYxQ35beejKhFP
OZKHUzVPjRWKStb94vvlKkKOXXVoSeYRBiq2NJ27i5oy2V2ECSl6QchUuVwlk/W2
YzZE4B5ubipFsd4PvzlCGgYyvIDS6SKUv/XrSK/OLWiXyec8w3+8+BcD0ZouVQCc
Nrmr8PBfLiAU6BauCnpV3s7hJjyhqOM1Dj6ik1bm45l2tv9N684u+UltNgGU67VK
Z/fponQzIu1VASQqDUZzDrCEmu1V6SNd9m40044Hjhgk6C9FYAi0FWExuVq3lwso
ZeNuDNoharVBTKdwu3/qejSpg5SeECx4/SdTvFaU3fNwL21HQN4tbJla6xHGQqLH
T4+2mr4/TmnD7CPGvgBd170yLynp4s9bZvvEQX0JuRSdn25CfaIfeh4IsRO9WDK9
iu5/UT91eREqsn5XeRDQ/XQ8S3FjujLQiJU+g6O4SFt7SVJKfqgYGp12xyGuciyR
Fxb48nIX9rIwIDtUc7wxDVWy3GG9LyibkvebwjwQMBKgBs4Y9xRhiwZu8VbtcXoI
6Bt5ngLvHaO6y5FdJ2shL8YPnr24d9rMFNLwdawHYj/ndjlaXr1vH8dv23tIiYAO
aTsPQbx6k8filVv3LBpY0vfVGsGLXaEHMMkIQU5644YE9aC0ZYKOEoTKzxYD50eH
qXhCgaHeyxA6gOrq7rieRqMTr4+yCMZ/NyMSoBAD1UNOrjfe0uuM3zuzVMnu1imL
WohQI70UPVZF1gO12iobl0RtnGF3uOJKHLB2pilKXYVar8Doyv2++CtqY1HDp7v0
rMeEyHzHqUDEUPoifEFp6lPgRGLTVJzHzZfMAjsW8D9KUqFbbGeGTDVha0kS61Ap
G/1tqXxBpXe4w6rOfcpsHhT6GCZKoHCniv18TERTQWiNV6aLMktkM7FQwoBcJUFc
bb+8V4A77dnN+wbwmoTlZJ8mu4k4D1a+byOOGhdUQxsnGK4PQhrqRZXgq/OzcrLw
heNH3Hi0Arxs8JXHnoe0cw450WBCcXwDld++0jVjKTyxo84g8mjxBn7PJi8AdJpC
ZNNYlN1ke/4i6xa2LzzPdEvXx3peb2GDHc+tcwYAGbgppD0MJkB4jFki9X8Pyrod
4rbhvjlZ5cGOWymbXaJxKsJP6W5Wuoy2CoTGEW8A0CKn+81EFDDb+8lJxuxZbkPU
Jt1nNXb1e7hdcBgMYUBaXhIJXJjI6p2P5CWIs6SWgBH7vWa5jhLDHdBYG01T+Pum
e5zNlkOwKV3nukvtDduv1gFntPuovMlT8oc+FZFvAVkZB7iXifBwO8XcQDw0+2Pl
XldrSBUGIgDjAbxZQzJCttRTaO6gAQSQu2Qvx7bWH2A7BLLhiUTr+iyFEI8pNj3C
/USbR0rOCxmEbeOZfjU1nezvZxosv1n3JZuQJu/++p6tns+zBrDlEFxnsSZCOs4B
DwChkV/XP81fpLD73VLRPhqNJ6c2v5IMrDQhHRUc86HHdrVMXGYCmroMP7FUiDtm
sQFcPpVY6WWYhjxKqE2GxqcHI0a0gxaChkJYsgzWcnjNdzFUSWSWaFE+t1VngSN1
6SAVDOQualKjtOs23d9GZSxWNPtiNMfy2JHUEN8b3NlBa+7+0QRrg1bdz5067T37
0zvX2mKAsVTDCqXhz4TelYr4z8T6TaRmHNG7KK+DbJDPesAx6SZFvmq+bqAQbpTB
hQkCdpdzOz11s1q2iD17DgZtLMkl/LxAzxaTFju8EsGsr5FXpyk3s6K07I/wms/6
uDg57EgEIBvraw9PF769d7QjkIALit6UdshubwE4WG8yN4464+nfDY+dFvHWZb+b
MN9oTG0+8XluPB3sCF2h6YIg/Iz6yAadBPTRl64cTIZvS68YaEw9vmYfTIJlRoa8
WTBsde4EPzHug1z0JiTRQuuWht/D04UxC8YSTAiVsHXcZG7xwSa0UPyr+JrBETB4
hkWwJV2oMiPPl0902KcritOK+/4PlfG/EXkZQrVPU+jeX93aUZ/t+GqVoBp+Rtxl
ks5rWdiZSH1LKSLTo3fxNqfMWOyNGkGzINJZJ/L0xj7120FZt18Cis5Set96utbp
wJ628txSTBuKCEh687XmPocSU0sJW7hDLBH5Shds5stS8KKuxwG7aIEeFgrRB3Hx
zihaJm02eqNs+2BhF+TWyBqt99fICItIv7WDzrMAV+FDtEWfy4/PQjQsVi+CzJlt
U94uk3UdVtTxTd8CRz6LZDo9QaqyKzlaHCPoPQpOETUX5fwmpvsoM8Up2ak4LUlu
u3ZK0D15tXMV/7jjZwdIoob4JH7QBm0YS0oQzD179k9Sok0ygt/nlUoB3pWlT9UU
jp8uZPmXG6OEIqrJ5CuWwLRnFO5gRM4Af63yy29HT4xCTjzdSQcRDkGPcqsrDb8g
XJDl4SLK7TpyekXDd1jWlBrIyQQVY4nslrWK5tmvot2dXnLfSDH+Qnp3160hvAcC
USYvpZ8hLHei7DAUMEtIgGy9ThUEKDpIaUxDW103AhMLovNIbxUTSU+fnmkgdWrV
C1VWgGTTlAecxk5f6mVPK0776SV1Vzhqgttb4Zyd2uYpct7XAFZaY9jBeBOJ/wT9
mwBdGU/PMmmPzvwGCAbJgMK3mJri3Wzr9bRCOH9QUFE80W/ZA3SpPJqm926XJ/E2
e/CTa5FeQQ3mrNYld4DAIf3HsunzwF4urTFbZCTGyafk/Q/CE6Rqh2Ys+7Y7S9wd
ITjSklmGRRHKiGWl4HMvuxJ7brtRbE4z6zAFoh84YOS/FSfaMD3s+ecLZ9oOqtnz
R4vf/PSMTIPBxBnfpl1tEtnfcS/gHSVXh6ysw4sd3OA4WNmrNrS3AE7nwtPVIrU8
gJlCqjl5nBnGOzirwn7qWmHhOq6I3QCXxfPp2JxPvH0+cEwRqt73mMdeAQMbqyUJ
HizDtlXhkxVSynIqaNHFDrRlzTjl/IyBkvsk0+Zkk4BH0FlKt71tHKjIpnSe6B1a
Lk6yuH+KnBgQRWG29uBKv/X8C/K/NIdR+X/eXNbecNHm0DQkT1GHz58Uv/lktoDI
C6ckmbBRk8CSaFjdiIRh/gfm4t77piFALvVikEmM1CAmsx5VLED9HWUEKoOvHE+7
A/1k50iy2gPOdLygFp96hsos9AbA2CTRV08nUrKDvgEuQqWl1HpdBZUUi638vEeG
1srGgRpCuclYebr9b1kw/8iHYFruFa7WJCEdcxRrU7vK9Bi415bUyencn6aoPEod
3CvWpdS//XfFV7LymuTpKzmM4u39v6DC+INOqS7RXbpPZMyNSkw0XfhUcxrZ0e0z
U77hZUeBn/+zFEx+y18KjGZXtjOSLp4Cw7zpg30A/eHJ2cGg7XkaVKQ9Ith9QIGK
ycFOeoNGq8Il2EBNiNxCqYpP70z7Sxt4o3z0pbKsRgQT4QFBIm9PpwLd9BR+Tr+s
qgivNzbXGfCJ0PGxMosvCu5aUwWxMk7IksyBWxhD4cdIu+DFI2ksrLHPC/+HWyHH
ESm56xDa+YuKH9qT++XURcL0jEDjPZteNSSOBuPqW5b1dsBZOmErSmuqSs/GklRo
t8b+z870J3OphApepmaD/t8pUXprBju9TAtpBTfQYpA5gWRBhRZItMghUsthQ/r/
TP7a6NZkyl3n6rDB4s7evgDTTR7T44tIJSCcwcF6yRfG2XZEbA1JnXSnAnugnTlH
DQb9uOYl6BMhP9CddvmdZND3UjEwjREe94iauzuw/jailuXXoN60/aeHzJU5YIgq
9nR1FylbbY+otun5G+yOQENSHx3ltdUezeR0amYLdn67RYesBjcekjBSlFDBYeBc
1Fxp47RQaEG2TqqTd0wxPeLMXKk71PqGWjZ3mVlbAmBVvZAwq9/6UJIMunCQta+Z
I7URl+kbXczUu7U6XdJvtr3MMDtrwt5DxrQb7uX4MV3q9zEw6AdybnFXm3LbUmqu
u8DLiLQDbWg4mJtkNxImINmDEIrdkMnxa9cx6gFHWJQMOHwZ8NWGtUzqHde4zdue
VfB1aZhuSEn5dDJuxITD02NnUynW/dx8b35i3gEba4mj7d6AxDgDFil5eMy3fIyO
X/sA01ir2NPwKueGcanC10cUZABaWkToOoazKJx+7eWA1pz7ulei35wyhVjSUTq9
AGzX9keVpUcwHTKMcGhkvPSr1SU5FdiJJaEeMxmkupVGbFcO0YUhk8SS7JFzEazW
HklqTR0cEi4sGKt+pg1F/pxxLCHkiyjMPwzEWpbIm1i6ta1ZgIS7sOrW079JvPlT
DaZ9uQwgFlolC8Xst9hVH064TL0jcjAcZEGrBkiJRh43ANZVDif72WhmrEfgR715
7CThH2Q268bpvEWzHUWY1l2bc/36X6NnIRSpSdg9AwnsP5KQq6MbSA1K5wfVGYyV
vivNUGfb2ZDHkX0QmhW+ivGHhF7JA1JIAi+YCrcatn+L0+7+Dhl4CnWEpqSf4e5k
vGQhJYhyf5TcX3N6XNqlXlgLcLU0tDHHoQuvrl9ijO2FUG5RbbGdG4JE6geZi/ui
MDvdj0NkjH4FbWR6e6G23GGFyJXzmHW050xwgg0ewHhcjILSk8sPfuR4H9+H5I0O
ADoHir7chHViY3ryUugWosgJaJhmPB0LAxA6adSMGkdf0EEVn57ueUcGVGFPo7pM
AICKOtRYamLnmafl8r8D6pJOAIPsQhOBr2Z8x/5ymYc5nsvusxHGkeKp4RtFnF/Z
zW2ZdyNO9Y0fR1oz/NMmyfj+eJrVn0I7/Ik9w7J40sgtFCJ3MtMfrwiWfeDJiNKo
sGctDlXKuJwXNStGdHjz/03SD48HhMFUxsCPKTISKVhNz0EujMeFVtid/JPlmuQu
LZk4rxCbuGdmlGhx9lktrEzB0jIJ9jqNAdbSQGx7Nj2nvWa7BB6jwgKmVhyc11Cd
ofDf/0vC1AZ6QV5mb7Lsmuwxe/SPuxrOAlnMqsPoBlWIQDlWvK0WVdStMAlCaQNT
lMptn1x/6VFXPhiX5BXtA0hTFwNR0hGgRv6I2oSJ6KhT8kQ4oaQ9XxY9uA+KJNJB
Bzyh+pJgppgkjC66I7eJGLGRR2XJI6pBXqq9tUsSxDWAM00uSnTWeOFkRbTd7/Mo
tMEz8dc+DDHLTHsrBKdzb3EiOsPwwF/j91XkZnyla+aEYw5yuB+sTNG9JqQ2GqTn
VW5A0A3kGxfpav6Ix/erMnQi/B/E8mcEZgl0zfn/wgQlGLfLZ648yKq4JzZI4FQ9
YzHANb7R+ej61uiOeMgf52q3iddLR2ElRUZsTH45tJpDYBiEBt9Uq0/Kui4nLGLD
x1Hb9JvJHXwwoIPwrpaPnLXGWamXtzSTAJnB1eS8GMkHn71D0RunQWu1S0rRS0MY
tZcq1E8sjhokcZut61Bs0gIlga7l7VWA+dsCFjryik6e0oyeRMWTe0cYgTJP6KDU
4wPuphtx4XUE0BxSpr4jkWUOTT/yebotSLSo9BrGj5JIBFaeHGJG2m7Vqg/nRL0/
+ikzQCPIla7to3VArQSwBKm3cBL+r454LdVPjoIG854KxNxWyXr4BxrqvXNk/xjm
gSPTfN2emkSWLqUAUYbgAJzQ+0/2nQGP+d25OtAPzbNFkeEhQMSY8e4u0WoUxUm1
T7OcUQf9YGhZS3Mw2xIFps0XlYpXIU38GeNGWOzlty3QDzRcU9/oqMhS3TU7Q2BL
YK5MGSwn2docAzcbTMt7LvhETM/eAldboBidapXeHUlqz3t2xR072EdelfcJeqFr
zSrY8XCQELNTTOS4eTmCm4UBvpejx8yf5/WgoVubryHKN8y0sTYkovHDfjRgmf1q
l0Qi2mdjfs7rAoALc5fCJ9tf8TjgGQdkrdAwlSF/mbZ4GxGQQMt19zEmGS8KW2Q7
pMF0SKHJ5DmJ3webl3xmJ/eyPbCTrksAfymrA7av5gsP7Zf6lij/3ekHxY00Ijvv
/jC8XNXcC1Jbc6IGGZZO2FcnOPDDAQzfm+aX7Bl0bkahhXFILlwfisVcrX32MoiD
B8Kbtn39N2UhRZror+Zne3gjNk2gNmtGQ7RnE45BtvtnwzT/KeOn83m4DQXAV5ml
odvL55U8u0uuXdEbmQ5U6j1Y8CBjskrzz+K4MB4YakvXVjVNWeaxXYf5rWQ/sTqh
Pz533uJR8Nh/yykAaDIWdLCk+AsvopS3ypBgwO/j4NjbNO7/kLZTNuaeI42MLgkc
E13YwJ3xalmC09jg+FSOS8/vqzVXwpXcqWJF5jaWsd2k7mzZGwMSgEBQ3DXij/ZD
83v5aPw+ViLaBfHiEQY23NNu4U497bf1KXoOVr32YSpKSrSmvxPUPOrSqDoEGMzW
L4q5KgCQzBkQOkpNeVd/aLEjyMCpPSX/phRMi5CIozvw0fxgNzqvAEeZEo7VMO74
Z8NYGqWy+5rh9JxftPFkxErC7jqZMJS1tENKpfBq89RP7eUs17bOe0+ve47TMUds
`pragma protect end_protected
