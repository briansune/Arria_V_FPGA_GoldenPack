// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:24:07 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hpJpK4HDmpcOpWjKq9fVqhSxpR4D+TB5h0EVNTw1dCMAvWwFrYXW0rFFmtzNn1w5
0cksXqAr59QMEHuv+ZSWsGLJllzh/6kC0r9Qb8Z/m5Y6sfCi6PBf+x4wr/xcoEjI
qBfKjxlJraAq8kWcRwRnuNJ3OPt2uKEGrrxOPGppoaI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23824)
GRuGlzKfRmlCoufmAj+h+8yKMPK0sVNQFOy83fKx1pQqJQUmTec9bvLtEOW57Dr5
f0oiKzmqeuszOX2RyI6N2hZ9yGQ13NPNieKSQQUR1XXPCy8tXhHN541wpHNaWdLs
ZhAi3R6y71w9I1odBXt3uzKTWUtbmFeklthVmxou1kHWIaX/gWFiDAaLxiaiJRK4
7eG8fzTRO6Z2mf9gpYhoS7PIqELbp4MvdwL+wMPEo6uz4223c6PaCxLjDnGtKlsJ
JIItBX2nFBbFl/FPiucrF/abkHKhtfm7OtxbCHBVv12tbVnenv1yl/ZDi4QAYorg
xSXyKtLvDCzsHP/U/fwSeoMvNigJyWFHHaZREA3FpxfmWY+5ZOa2+AVkd8CupX8e
8D5mEWBdn8TohUcGRvpQrUO+0Q3Y0MXhE0XNBbfVenFz5Y1/LXL7P3Xj93aLADmJ
pmneKGXqnoZwaNoypyA30a36H1kkoyvy42GB8XWOES9TIvzL8Sh8aw9ktH0mkZ4G
or4H1kxpl8lEBbyoUMHVmaYAJQXNMB5i3JflSt8L6bx+1eF/GqNtVsnsa6pNTjW4
PTrtyxMwnlNXWgKNfc+iLcoL6E03uHsPFbpCFJbJ0x9vSf7pSF6MCtjTrb69hk7c
D2MN6bhywRqOci0K/I5tW9vUMfKctswIbvhGn2W4dZMuJvdVc5qLp/VRxyi8FxSo
ydcCbJal9FU4SqZdlIB+B2DJZMJL3MdxB7rFS9vZ0eDpKT3C8HKKLd6+GDROvAHy
/wBk8yrkdRQxOm3ZueeEbeHi5CRiIC2DUDrAgjRh/EbpO/H5+68KvXTn/y21iAsl
nsX/ICyG+i8j09JIti6rsjEL0NdgxcgBXYjlCcNr2dwoRaWF7ZYJZjDH05D/1CNT
zvKHJVWAHiX5a/08ojlOC//oTzl3ihjqNUfMCz1HqGYipK98cRPpFyF7gaD1PZR4
VRW/AIsEUPf3hdqX3ZCHDGaZmgPvNGbncAo55mx7GEoHugOqQZk/Ks3ufNuLJGd3
y9d0MNQ1G6Y/EFBZjD589PhruL/0Y4+cj8OaDGI3kZjWOTgArs1A19EEgfDzAirE
FK71fWtBBYIQ3wUASCguODAQ6rhWUNmKMs1AROd2HQg9gbQ3kcTXGzGzNiHfcUzn
BgtoQkP7sraicPE2vW1v1195SyVqu+B8R+LFPfeHTCBe+X12mzcSnjnmcEbKZXAv
R8c2Xh6VjEKvr3kf//RDmS/sd43aVKFpo0ziaMOnGh89Q4xU7/cs1EitLKGfWtkT
RSKf8kWY3neW450+Mi4OlD5zmU0iqJdG/jRmjTeARLj0owl6Zn8kFabgVwij4hjn
dFax7YAAa5JTvrOZSjLvJrvfF5FNWquevJ4efVLLRY7/Q/ULul55XYLeiFUCc9nc
nBTWPwB3Zb89jmdyc1S/sUotJyMklY3xboIouX7Zi501VZc/Dz/BQnyMqeSQ9o5J
hlg04hc1f7SAjRhmWr6bS/L32iRG2kqJBy/VKJtaghc7oqMR1pww0gXPtA4ci37i
E/hGPPMcs0ac8cSm+w9ETJ7tqoOLUKoyd+D8mXozw8JKzDYjJ9IZiaruPm+/3U36
ewOWSILYkPHo8kvtGFeXFgFNSRaRCCXqnfp5d2W0+oAa+MN6nuQ+0LLdZxuVUXvH
jzUKhb9OUwxXS7Y7AB8pEFtAlcXvmGhQkgVh1Bw4dKuN+MlEkHBMSD1RzKyAbque
JwokBxb4tBW27MeKeqNymLIEb8o9Vb4qUWwB39WN8ZY7Q40ZHFSs8+Add/ZO0ZM0
WSBu2sjajvmbzUOVJgEUzVijBEbKZQinxj8plgAlyoLk+PONQM4qSGxVjzDco5pm
XZbzGcgXmRtHz2ryIt381Ro6HyOrPFslNf4RKa5sW7miqIb8ToF9WgAFoeCrDoJD
+48DCoeUNlM0JHZ8KVvbw1X09WHelKoRpOrxNybAns6akMgez5VcLtKnahufZOVC
n0pditvA9D+tRv5RaoyL4EP5LHhuanK/Ig8O1OAchplyCcHMTRuynt6ITrfMXy43
W3Zlnq4D1Mf15Y9s6MBapGAmGn7ZcZ9s+UxrJGFnQA2SkmO5zJu8jPDaQWn0rsog
SU/kcyO2pB2cmadXktu+NDWHWWofkYKbeOgoYibSHds+oQGX+6gS0hcqgSHT0xuK
azdKc/xjEYN5E2NCBDmjLgoeARghIiyy7MPY5tMXyttR9lEgh87pQoNhPNR3EOXV
zwZGNaKtx7bF4/H+uC+c/EBzjXMH8kM0UBnED3/x11OzC0JpoOJuO0V6k3PxUwkO
hRyICGqNzqVXLdN3kayB2j+/y5/gBjBnS++Sxq0vnkc6yl13fBkGl3eBbTcQE5Nm
nwf1r1J+a3zX4Uz45gJRDYDGGrFc4FJf0dMehB3wuIG2i78y3PQ+wB5Sbt6519m+
c5LYg69sm/bk4fBFX5Sfa2X1J4dtcv0qB0MZZTm/OTxJndW96XluDXVOv5goM//Z
8LVLJ9NJowe+1doMyml+XCJhw8L+gVZUsKQAYvAFEk0pFuq25KO5yBQqc/VuWFiH
Y+lN149xqfCDvuD7BqYc+mRkyAm90MvJCekGccdesIV4Ai/8ht8tNn60XA71w1SX
9O1btqMxy/7nc5oJ1FtDzHEzhgtiapPd8jd/Kp/ot1CRiX82J+bZ2IRcx0ccRthL
sYWFwz3MXU1IZqfp8at0OifWSstVgLxYanKw5/D44SNiDBsX+iEbAEcSuovzjAmx
uDLug4l+LeS45OROreC/j97ptlFqTGS5UihbplMlhV4KjcrSUtUJqjibS9+hmsEz
oYKEDx8c8x31RQeGDo5atp57YMPm3BNqA/sFDI05POvclDj+d509PbXBPMmR93fj
p/OKxwRjyirhT8e6v33424/3veebPIJqCh2+41FEUk03l0XRwG/Y/9qMiyEm9/uB
xJKhTNKD2t//LMyMFq5g8ol9KTKj3/kZHWYegNVe+TIoRMnH5RmaKt6EDZrXjS31
armuark2w3IV2/SIlsvrU34KYwCY55C/lbaTb/5y3rNfdlncxqmJ1TKc8Cv4eq6c
RnNiVr1MwQfxiOi3sf0KQJolHusb6Ulyg9xw9HQriMk/hYV3WwG4whvyk8RjCIoT
gLKB/+n3Az04+Ilo5tlmlontPWXxhAgITT0oMA0X0PLlBPze1tQAVQOLcCZNkELv
bWoBmVrZ3S83YjATeTorquGF7Enm2nz6IF00vtU2ceJ14gOonR0rc79r7WuaZa4g
WwwA0M9FyFJMsa06FwyQegCoqhs6nDR3RypdLeoPc9lv5UjPeeDrVyjo9k5P9fH8
GW5stWYdXlR+u28ZJw2DXsBB6yJGkJjoDMs2K5OiCbgxDHVr7sK6omwz9FnFydVe
q3wOJUSpve28+8nEhCP5vAyEFbyDMfoFOmopbgqoCPAzEVKQ8PrXfad9Cd7YmEFF
MfCezcsaItRtV2GLQ+kFjUsXc5uHIRi/4S4R18xSAUIRSo3uX1x79S6yuE/JdU86
f7rWgWRacZYxGS4CWDydZxzzqTKYD+Aa8OCmmhzGclR/3GTumoTpwY0Klh96wJhR
EkXHM9YSN6eDD0vzBO2M2b6gObGWWwUoWtR8nA8WfGy2jovude5GEZcWKofpkKhr
fOhTyR2H86H5j8tQnbIHbpc7zCdzu2Zv5Lt34i8Ei5oRtkk2ncYYTDbAAQ9QNrzc
mH+pyIRDNCEL0WC5MSrQVjK7yTSQOHBj/7zrmhq+5dnIa60K2EQuh7i/jZGQ/ltg
O4VxozsZ3Allj8NVh61B42iTT6O5izjvd3cNxJOPNwnp9Kyv2aWQKZDD9+JPdqHG
fb5rquLFDpqxG3vXW9kLnGTYWCfO760KZIMULXRzfMeab3EvcmMpmiysEOrPP1Tj
fA3f8WuAIRAwkaU7eHvSnjfkJeY6WHdc/RQthutMmxOjuGtgYEIPdjONAaGcxigs
CoB28lTYc4l2EUeLeFPe52KxkuVsWpkfKZnFQsMpkMtwJIyx8IB/ZikWpoywOct5
uDE0Sc/Vpw92ttygr7WvOY6rVoOET0alZ3V2v3FXm13Yyoq43UZyPIi8Drnpe7i4
w3frNutTk3SJOa1XncLhgsypchSRR9i5ZGwJvzAbBtY/mxqOePJqzIQHA99V/3KM
QQMk9NF7nG4+yczK329R9v46W9eRiDtDeHBYL73dDIICz50IsZezvWogrunZGBNE
zG5HZzubktivl9howjErMwmHlBrTGwdxzFnnL6zqOxP6vM/PhvxSfzn6RX68k2os
Y0O7P17bUCK4QochMwkTw/kFwalqhB43THt7M5JEIzG/AvADoUf+n32rV1jwuE61
q+TaW3f7JzW0tafbezB7icDNQUpq/4587KEwUfe5RCuFDqZ6hlyukmIIX6qGOAkO
V/IhuDjRkvDRXpfJb9bPLGOZEdg1xfk4s5NdNJfU8e2CpdKg/rADOimAZ6PevWyV
gGQg3LI/LsImhg1PTIUdYauZMj5a2g7QV2pTCulG1r8ZBdHET6SGsYn2H9PZnsyG
KS/OhWRA8LARyNuzcojlT5HWeRO7y6SMlfQD8yel3Tle4jSEQsUOkD7ZQHjtWNkW
hUAZus1B29vOb6Z3lWTR1Lip+YMDHCPHOAMDLGeDH1Gx2M8MlVxsmueUFtD4nxmh
VCdUopebVXutmVgBFPzxnYgzbRpIzaor/fzXLmlX7LWegoTBIStE46goDNoBtNiI
d6/gzEViBIAlfgd8+ktKIOqmn9nqaIMBlBaLk0Q05IqyPHtc9rKiIjI+KUm2fGeM
AbxxMGYVX3QmhU44COtQ55kKP2//jHON6b4EFgGMy5I5mHzsW48rAkElevuAq10H
4ePovAlbQgrCZKp5JTPCsUJYJft3fZ5N+PBfvo2N4UxwqwVL8DYGVbKRHV8Y2v9X
6yHn85YvST/iTnzd0CHc8oPAoSbfOaB/Wq+sZdCuopF5TiulUTWoaWxWlJskd/LA
PRlVUBVTgS3v5OGyD1JBn5Sr8Uv7c7Hhs6exczz6XHOEpL6vUL8DR2n23DTycb8a
/w4TCMFV2RmCWYlxvqtrI+4Yp0YrQ0gkKziGodZQQFV11WbmpYlG89KXvvgooyLs
dqnHsLDF91lGQ0lifcIqah8lrfPm3cHVEjXT9vQgVcmqJXsn8hI9iVjOVrHmm1mU
ASm2e7+Dq51PNo9/O4YbgIx5yOomsTANxC7HLM2Lua9G+jynMGBiSaILIahWo88u
ubZg2kIIIFCvkilI74kLezP0ERjsU6ne1CuQL4k1pqgR55Lv+bew91TZ6sPDfaZm
TOL5fu8JFiCoo4XuRUjJ+ExUIoffLsv8SJwciCbd/dSW7UEKoFJ8H3yPdZ7F64pg
L8UmBojRcROwweUw8ljS/Voa2kIa1cKU9BbyujgGJTRFHoUjhrXyfqYhOGSzlQt+
da/kaD6mWPCxxZfCRsO3q3gjTWLJTeTKVpPMbFn0Kmr5RfdJ1kzjiqLlPsUTDxPp
CYA9hkGzQtPXSqO2ncxTGf5By7vFP4jbixUBp3etUE9XZtR3Ie6CwTAxQ2elNNnZ
PVmvUMC4rr9399ncoIP+W2/H6UxxuGdWliqORMTkPVBPDD1LTcnLzmKbrfcPskiK
HJc6jSWyCQc+wOU3eVw/xo4gJ8/UxGRtT7czJfYq2YcY8YGRu8Je/mK4aLqO7REG
rpVIMhE+rD3wp/ZSN9/XmoHDkmkgcgQC8zm9GLhMSPB5Cf/Yq5P3KTt5J8mVPaM9
I0crbhbg3Sj+4GO8WgXk4MLMN0gWJ1a3tuivd8sUQI5H69u8A/e6gr7xQiXQvRJZ
5JoF+qGBvtAbNUk+xr/Be/T6zhxqxH4drhl+nJAytPXywI5keuxe3TH5kGHyfyNc
ecW9iAlPgi20n4MHOn3hqd0UYQ3mf+55dC/sVX8zxGA4Cf4NJiaPPOoTHxIo2tKB
cToOA5lBUcT30Vk2DWXOR2SyplgnnQzPAb6lFeX65fGJJI87UVqSvDSaiAe4FH3I
+hHXCLG1QcF42lUx2PtabdCx3J/ZvxtHEvBG8/YnrGQijg88tIF9JYbjQYt5qWdv
+UoJASZE8pJRq3MYM2Y58p+s3RpqBrl7KpYp/Ub63GLN4r2gYqOvHsagC7L8uw/n
YX+PlMt57mduBnYe3OtRPmavuOQS0n5qr07TXUC/BRbNEo3j1/eRw3ihsDvNSoX4
Gv0wa6E6Qhr/3xMhVzQcuLEe0NIO444mTGoZ/YR9gAteA/DKwOXF6XWJklPS+zPx
801w2VmWvGrxcLvqqy0Y6eUBagWIfffQbo8FbU3JHwA3/i8q8XiOKQoL1g65Pbms
PYmOaMJeRx6e3g5RarxNUKjkZoemuhSSQd5mnrQYsSIZvabXJAabwgx4gO+HERlj
nom6sjt6thOukVWGx2ozWLH1fkjAWWVYzOIdN7Nos6J9RmX8JzpYjX+OIE+6jRs+
oZG2m9EIkQuLfZ0jw3RDjBNllkzIw+8JKRQdnQ5Ct7ND6ZPDK5FHL92wFybJ1B/S
KXUyQ0uHcnxfPa/eyLngDkvRFIiHe0OeLpZPVJ45MSl+Gg8StL3q1mlmtd2TQoWH
D4UzehtP9s8chuXl8/xRAr2pkBTObqmIelLjkb4h2GCXlp+qaY4X72eaNcmJjMer
PCpN3ucKUzKlDrOL0UmzYRfrqmE30Ewcfmkoa4vprNapgxQUCdNfDZfE0MzK4GNT
kOvtBEYiOCSSPYlAT0ZUalMHnV6GL/SvKhbUPd3LamR7SrONAhLYOHatex2wR5o3
HgBzWNhORIo3sia2cRJOy8AFTAqyPtyOvnj6baW0ODw5I0M0/JdKxtWgUcdsbLFS
11msjxPLp1RsJxquJLsB+N0wnaumkVe28fzEQ6UkS3ohk/ZJwfbLneWdEbKQSnEB
ft4UIjiW0ocyt5gWH17I7rGP7WA6OGPTQlyoSjcp2Zmogt5/WJkNS0brHKx9czeL
FXX2w6B7PbdL/yrMgGaEBNYz4SiDMeZooFkO/C++gouMJ9yQ9S79pv5afCJtmH60
Cvxg4+E5K3CAIoRF4/Uo0M4Hw9T4apZz004fH98hGpNYRk+jIg9WaroBKTTiXijo
Mvr0EZIYw6reosyXvDX/X29Uwi7siA5nKxOoP9IKFRbUfMWEF1VX8wZeboivWrus
mu+rLCUzpndtYVd+FwWULBGqPuhO59/YEsVk6psqxDT3LVHK74a1o18PkbVDNlcQ
eRMjMFItJGjwTHzMiP7VLJZsuwAwgVb5R/kAnMCiYMgPDg/dLiuZGTwE381wmcCe
HLTyubIpFQ2WtPMUZ/I2Tb5H4ntBrwQ3ZR2EEFOAntHjg7ytW9Yt75Jo0MkPKntp
dsOV5IGJRsmJHAzSaHv5likZCWj64ize4AB0BC7jQwVQ92hY+ieroN0Yd45n4S9v
AXqrcUtvS2chw6KI9xPUIkN7cw07m6oHWVGAj1quLpZWwO/A/8q45G2gnuP2teB+
T40HRSb8M7Y3M9zo7sF9vusFW7/H4FOH2y6FgvXvMhLaezS8Mr73we7ZYVAjewh1
hQ/3OampRRViDUcaBQLQr4HWoRg3LIJ0go5QZyVSdI8HdO0p83blR6DnbqvLg4tS
INwhfPdsTiUBpYKseBRpkYEsK4JtkXU0k9NtrWueGlONcOm4p2A8Bgros1qd79IC
qmsr3b1lVOShk+tCs/o6EQqoefN5nDY8mhElEdCqbkPQC6oSDocQZcMDHXkMFbAl
mAnAWIxxkLGus67GTmRjIGSMJxH5QlmO3FxWSwzZ2hBS7KqD95J2klyiM/sCHWjk
Bv+0poK1UCSe5IF0zT4naOJOlKYBFj8KIzRDlaXjr9ujByfm6XtDEEQgZ9wPBkwz
RXWVeO9iwGAKijRy5JlmpAgXWP1zsJy99C9cFyDVSk3hbfY3gRqpsa59ERDPBv6y
DwCH8T4M8qbj4L6Xmg8TnwKRQUIs6CsSaZfgSkI8s5eO3ruWj0JhHqht/YBlCLiY
bFGkGv6k3aVbPyCQGsh7sDEqb5RGByJ5lQvqFD1Zutd0mqCCaG5c9eYJ2C6BYxwA
NwicaL2Nxi3RHCIh5tQzfSR3m22gYrCiEDEBS5E1Ok+BPW/hZ6tamkUpNNhx014B
TmSQBLeVhB40PQmUnOiirgsBJIf2LMGad9zvdcoZNhT7Y9SOpmsHURz//gNBBCIP
GnBr0iIA8A3d9m0K7WdRY9nh3b8UnTtWj37e6MdYrezdjsCQGTDZN9oHzf8wzvF0
goMHVD5vJmx0mOy6V6jl2Y+HC/2jIWt/eD2j9AEBW3sPjLWMl8rgPuGJDAKt//d7
LSToXktP9k2p6ark03rkSTFE5GrN2uJmxLwDb+Fj+aJSEXSMXsjgez1ZXUHuWBpt
3i4DVbSR1dBGFu9VDmzbUo4NxRw6ePwph5Splw73EV5RAoQtx9OpjVzkNIyIMDa9
+CoMBBzm85GANB3RVlcokjjWQW8biFXvlDwpSMk3lRgblCq+qQ+40qR5SuO1QSc5
giHIeHKHPpx+GeFkWSZ3SvTzorWmcp+/R8IYO9s0gwlrQL8tq4Cri0JyZYfkJzSa
ELTotlrXZ8iBPWoJSAoSMlfjJykeH3cfV56R9571mzxyMk8+dav8hXB7Cp6IVGHi
+KWlc7pW4/FByBvHSg79feDe9jN12vTehveT2tRlwzVuQOBIBu6+rZB+xwDsBg/V
hNkOs9Dq7uxxaPd66RoV89A+k8E5OZ81EkqTa3ia9u199lBRunUoB/k0z3SOiC1n
ptS3EZVcAAQGsjjA8KFj1ZytZVmCGbWUim1iXgMUiSehoj6BPKJvxWyzThJsy2Au
ZcPy2RKN6p1WSXVNnj+clQyc70W9w/8TKJkUPUpMvkSYNW3xswm0fJdpj2kMyiit
FLXpZxF8UMYm+SMTSef5L2RKYw10AOgXrDsEfnOmT63UjQO0mgilIx7Q+vq5wHId
QQrteGyoJt2kcchxjM42ITTY1jayYKmQaIbCC3i2Y+RIo4b3I5QxB7kEe77tLKEy
nszbObD4J8rCQEJwcNqD8l81lzIGOwVNmB/Xh6r+BGo1uh6DRbyomniCKaydQ2a6
fTrEyJ2XpGEa6AOcMJn62FJGjsir7OhLVYKBaQtPXjZiD2EkyOCUY03ae6gQ02x3
Ncwb1O+a9PuWSIkl00lPHdbctG6LFZHuJ9LS+IQErikjfQwW7XBP/Uequ1v6vHNz
EHNBTA9yCc0RhQrTXz6LO1Sug9tzRpAk3iLsv6Jv2La/He2lyW6y7nXhu+JqYYAI
cYhgh4FiTgIWD+6Mf4RUkPWz5acI+rOKods8talPXmO8ZziUIwp8IcM/RwaQ84h3
cp7ztdvyF46WXOgxSrzexs/HSSRw1bNZVKkd7E0uaB76gVAobBJWtwopJiYpRQBw
zKTG/mYlBNkYXuuee9ohNK6pmNmpnHQMHdbt28ZsbjvH/db0MWg1RGG3Zoc5WODd
5CMdXC3a7T/8e3o48+OZgrJVVQLVW7OVc/7jF1ueFc1DeSPpMoNuLD4VDkQ5l1gm
rELzwK/LbkEsEk/+e1MGq+YJtNedWIrPJCKZv4ZvzspCwkSy4yKqAErMkNI2Esp3
oNiVTyFYNY7pO0HyDnd1/oaFz5VMItz8w/EPEncjEiw6s7Kuzo4rgWAHirCqRHQW
mKGdVz9RJoNRfhFnjSr76FJG39SRNtKx7PuutX+xXFKMBxIFpFMexQgLFyK7/mfX
u8lwjJmYswF4RDi4wZAltdMF2tzwdP5G4vp/sg9rCJIRCl2gbS7OelogXoNHmeMF
g73P/eUuS4BSXSgx1oM+XU3dU/Zh3IhDkViJHUXuZl6Y2Ja/XNjORLaJSFM/J4nr
NwTxNv+k+j8X1aQqWByPhWQTMOSKe0evBL7N0H9AOBO/+rpB5nyR76mCH2iGUiEx
CLbtLFOCDKNM9V+JiR710d/1f55MpCfwRcJFNstgFuQSp1Kp6/y0/QAWtYvnYIql
FUKSU9GdWnyQonKLnqyO0vooXnsKAidqlFEC3Qi2dZr2XTNw3JnIk80WQd/NHaey
TGex2jsgygWAOrarDrw4vnW6sfde8wID9LJ4nBluhm08KyaXWR/pUNcBlRZQF783
El6TViwORPdW9qhgGHNLL0gWh2p/sGJbMS0xOKTdeC9w8Qhidot+foRbtunwkaSQ
Flw+za1+2k9Ca8UObvnhBxaqlyhy4KOmxZblBDkCgF/MsKF39VKygQ2vArUxajHm
9yYHAa3tAPj0O8P+ouGB59A8QB9EpvICyYvxomhJfbfZgw+xd8xJMPan7r6MP9H3
ca/n6fS4CV/8qGUqCMBKz76Vebd9MUsN/dhiA1zwfh69vUDuVd250gGWJDSDC7f2
Dto26JTev3/xsP0HlM8fmWRhMkFMSpSaFJhK4oOsr22MsM9fNMhg/DjYasD6f3g5
Za5AV/GDrGD6nDIJft7Tlf2x22QrzAqsgiiDtzCEb7WpY/FuqjJHO7zxECwkTDpG
cVj6ZF0Ywoh9w3ehJGger50y7mbcS+a+B1+Gp/rABTnfwuoTdWn9C1YrP8bq+I5E
bxjvSP9dG3JKHLUf3/WXj2QAkRIR/RbPXzEYFMXhPgNEM0ocjT5k6kE68SPKqQA1
NLG7dkHZs//g9BWN2CyrVA+TMc4EB3D6XxUWFDVJZO9x1rcVIg3y2xgWiSnsBXld
oA9iID81FnaOt3bhppYPS8lk84ik8m4ifxIn6gvJjbYhrhP3oQXtHcNAHdv5iC12
d82OTWF5jljG33HHlJb3BKi9rioTPPeKrXPVYMHLIfTMIzH5NJSZO7F8U1iX9Jsu
PbHD096gX95wpQz8FRhL8LNkqisRPaXumgztb7nBlgyDuMeyaprO7xNkhc/4GaPA
dHR7OWhvAF3oiVCbTXht78VoHLC1yw8nzQ/BPr4zoe37SKatySBQQpymwvnmOlXe
LYj7obfSWH0o87omPVU/eyYxCKxVPHU3nrMCvdJAtpKYcAq1rnYmJjE09xXB+x/l
lPuWUzAzgFPMEfMe9ngDPh0afY2hWKc5b38/HmaojNoikkDBfWF5glVmoQCIPrnC
M69Noqhbhb1VFOZd4gvxjv5jVUYBKCR7SrQpCI3wDn0RHSz3z6lgAQ3nAwREMXCO
1oZv3whLq0goXMUkLk8eqU2Hh11SQ5Gf1EOvt214U5PG6ymXk/t9x5m1fGxQvFB4
AmeiRk7RJbLfILyzIVsuEjWWfKEBUU8FeA3Emuk2nSR2J6zNtR2OoYUv8VgT6tpl
KUA0jwvncRafGB0fTf09InyPSkQFQ7b8jEBVOKvHAZkBnN08jm0LEQnW8JY1e/zV
2u/jP15a/rJUTKV0l7o4EPGegHoursOApbrJedGN8CHU89ZNXPNJLPxq/mH772b+
fa5n+fAlHfIjP4egUQwNk5BGNbuw37Bx5ZlbMQUgf9pyyLHAOJjGZMxE35zbPRxF
b38yyDHYBQhHChisTFJsMBvaz+AizbIfpF+vFNTqrYs+cOYFBHrY99oh56jfiGqj
nDECUCUOj37EY7fBHiEPHZwaW/lmLFHihRXZrHE8/hv5OMVfOFqWfkeuCEpZl4yn
gJNib/xRZ0pXcMft119UPDxFMvxm/SLGHuRpJgQf9VCG5Su0kb7y/XOF3R5uLYNK
8uFys/OE1RQgxAsyZBFAESVB7TcfPYD664t/1Z8O6E9dmLfi+8+V2XOrK6ue+2w7
7lwnvGW8L0SXsoy0ifvRcWxfMQM+QI7Ir55uHKWk5sdfDmGaXI94Y6eXTT7qtdW1
F8SH6ONbYg42FbdUHfu9bhQniFibma5oYRUDfB1G0fINXmSPLmpwF3gLA/LAlMNK
5ZDyrzmoHcijXnE9Hk84ePJaHOUbKVCs4hLgcAHFQgXOX8Hs4q+D7IMd8ei193De
YKeXgzjYP/1tIMdcQGpdVUU7BpyLleEPdME755vbim4VN3NHqUbAHjwmMWJjFghU
V+uBJBD48tahhgI7kPqTzIaZ6cKJvp5NtzTDh4LhT9broeZtFMs2wY8G6UD06sQh
7aCS+ZUzTyVCHsse5BqT3SVTp07+ScZAKMuETd0lRdJiUfigUH/g34ovU0zgFWHB
7xnAisV7a/LIlxwSPr+/mFNlmHj3kLtXRxlVDnwNKaoN620GrKuUyhrYcmLSuWei
Rrk991fO+TqldubOfDUKqPAfzTqQ8y8wDvPRsGWD55B51+xQNSsHRZTphJ0FqZtT
8gqz7UD2SBQlLorf0GN+YoM+MO8S+m/AImCte4l7zVD6n0nCoOnYUiAtkp0Mz3NM
fTgfc0rCiVYVtL8n0OCO24NWBdUG/TcgvVs7gZjCjiEiVTGIRZKA97a9G+4mbQ7V
+EuUWraKM7kYOyzIEdtZBFm3Ez/F/1DuS9OsCanGwMBBy11prXKATttpVHciNf+Z
NINjG3Caf+otn3iS5TO0iTDpFPP/O+qhfBtXrxvMW9yjjvbiGO8jTUfeEUlZN7i/
URoygrkkaxY4AoJRTCUftGqSqAB4VR3whC1yisH6cRVn+sAtsczLwQdi7oehh3mZ
FFJfnSFkgm3VKfrQKlO7GquGUXcDqkeY1FwmeH7kK33yVJKqKwx/vUCGAEsrsd3U
UQjc8ytrKJNsSDSEUYYsvXKJ/mzp+444VjmQKSuY4B6B2ywVsyiYzLNM3dYwW8mJ
ngMurC4+6pium+YAKNe6nHHlyjVIHdksZZ5/jVwQyhYq/XmtPzlKQszBZRkenfQK
3NHozoozthlMU+ZBXmP4jCPwQwr+ThKOv79w5svMbR9jNPxPQHsccjw+uUcmyS/9
2eyk/Had11sjbbw/YwgFIyRCkRCkEs1Wa1Oo2t6aX4RCTjyD+VX8ZIKZMZCvAsMr
8PK+T0FAzbXCRlQFKeHmLcSNxTjzyT3YEBzvhyMeQFv4Q6tdGL1ahpuFSuWw9lhX
EBuIFFi82s6v2yuO3O0iqHzfT1J6rKySg99Bxuv3xZxaReT2KqLE6Ktt8P6cIOiu
bmMkyo6jkM6Lc9QfB4gTIPjvGXUpS4raXqLOEn+RQvZGSCACPZzgmx5Pcovma0p/
FuC5VfyWM78WosOi4JK2aLXXZ8kywy71qEg62tcHRNi2VhVJ/QQ5AGZDb1pHb7JN
NbqbiAmUMXyx6heh7PfaeJtqud59Alf9slzNeQWYLQla4kY2R/NeL2ahXfFayrOK
D62wGLrCIaQ4EpZ/xne71E9ABXQGI0UO10jnDmoF2sIeyPNkQ6SOXk9NXvgqJOi/
VhIH3riiDmRZUIThYbbH0nUxp0e3hHs1soCQiMP98SVaeh37WVI0vqCEnhWtSUNi
rjlv+PccEvryDye40xaWHiw2LUkbZRPWhiWioRI/RujhXpxRSUh9vL/pEM8FcWQ3
Bwkak1fTBDckc+JDV4Cz5/TTm2iysIxLQDfixnCrl8t0pvEbkKiIP20FhVyfP7TY
u1nSKGixBxKnfK+HOx295HS7cS+kH0LOU0LKS++qZ9Z5msMGNcXE4n/zLuP0qGDR
qB2Z9lWvvOcLvzX01ytLuT1AMp5BVBYwdYqd8uRAh5/FQ8fQ0fyddBk8Ykgo9MO0
skRYDg3j61uUUBxMInbUvQ2MZt/xq6ycNuk07nFeKMcs9llltxHNWjoE3jzXzhrf
BLRN6/ieZkar7KSYr9BGMYhrzh52al49wAHN7QgUtrTFbjy4ExEH5sRdSOAVCZLm
NyEn8RzIizPS2VA+9yMpPG0LOLOCxNxblk2apL1AaO6VXAvHwspkFFjjr2q2OoJa
1AUZYvfYosUJqRTRrgWsI+txMzNVP6MpsWA6orMPq6xO5NKrx++iGYOQ0n+IQFyA
guMxDFlX6h93dtR5VAyI/Sn/Rxi7G9ZP6C0ETJRovAyzPx4MLoV92mDNWFYKLG4s
6slKYDeSvXVxi+3BkNQoB7ATUpXZTBR6uA6FHS9QmL/6NPGJsiNvp7On0C0tgJZe
NMOqtZXlhXQJxTCCnwb9tKTQRBie9VAFuVmOuktsfeXIxsZM9WqUFkar+sFuRi2Q
dAE24U+kLoBAKqSgDwEezdClwRja+OnuhqiS6ep5eNqnyyvAQdi/AK1UH+ayXXO8
aE9eXHNVC2XxAWs9Ij7G1+mwvEbqE5dCIlRnW0rLMdX/ZAH+RRO9Z12ImU/VdrTj
SwKmujOWGXTaiMnStKpx/ptnboncnmTrXBC79cvC4VjOALeggwh+fYREM3xgtdh2
s4f46E6Wc/vYlf4QI0yr/feqCzZk1zvES68QfXiEv0zYBRLcjmFI0vY1uThUdh3q
aT0DD7cggYokmHI37ie8eZ6fRIWK2W7JBQC0ewNNHfwaYye4cUqstIHZeoTSQqrp
EIMPxtiaoxiZQ5eLY76Fg4NaBbfTMVV7QhOvtWM8jUzEMwRY2x1/FohOmHyqk94v
LrzBvzrgaJuvWykA80nsM7GT5LCyHBdhbe3VDlCqKoItMFGgb2+0f6fZ+Th09pr9
5bKKwDPxXLKBGJwFy3fBYUuzA3Vxen/vbKbCBTNm8ggA09oQg9ydp427yRJKCgNl
pQejmSMFd6YNH2B64ysBnTGZZKjbBUVvbHkJdfF1HSog5h0KazFkKSu1F9nnk/i7
3exNDJ4Oh82r2ChAWN/WXKejexIqllmb7H+zmVaImiFCDE723jA9yC2/fWGg0qg7
+alVjIeQB2latdEFbi7NtjrkgZwXGm3GVzT3I8hpZmldjfjt+Zq2JrYi1M8DtXLk
JHCI0BFtba55+eFgHFFJy+d/zUBnHbsQ+XK2otLR5OdhgTa7WuFhjUU7A+c6KtIT
XsJmlWfF5tA+X6LMDPpu7ee2Tm6rHuUon5k4YwjZ9KavG9elq42nEwDSBIw1ngNW
MJns0cHgWtfrk2PahP/wV8IaCwmZpcvvOpooHjmSJX0qoJnoD4ruhZWkG5y8hmiO
68yWD1ikuiV04TUhhdq4ZaWAbgTxDAhImoDEwQyjlltPUmSTKwkFx1fV+3OVXGjs
AsZ3Wl2Esc43b39QACRx6bmdOsOqBvEUIAwR04F9hHsCg5qGdXzemtTbHQGdIgBp
ccXE+cD54Ur5aaenPDifvWY3AuoTr5TuEqsi3iLPjl8HmCQEdFoPfbVqJwCcns9c
sV9e07bIN1sgpL2pCmcWrbCK0ZxFNoAU4tLcTS35E+oaxr/hf3rIDjHSm89GFHOt
32BgBArhb7PgXVMy4iNp/iJbmymQSLYFTsIGn16746nnyxAZCzPC8nQHBqIUyVpY
PVZm0lP3sjYDxmjKkXC9EOPSpRdu/Vf5DAbYksMHEffTIVleUzSbTyT5FBUz1OVN
2Fqagi3IWyIZKAVPsQ7hE15PabCswacSNLZSWfobcKcI6heRQ6ECUra2osKoJ/za
4zcDhL8tBIo4L33mIVorTKCBSgy8g3Lr6W1W+PHCh9jPyPXbIx4Uo3z7Hu8KfX1y
ksDy6F9koLhj1g1YpxHbNXgW0fVSfx465c8eb3C8+zwWBy8dK+87NdQnVMg/me6B
LHHEphehuYRvIF98MhJsc5B8i0rOAsFe/T60t7TIOcPP7OMrW25bbiNJsLzdt6xY
PxKZAf1uIU1+VqiCtQ078pG/F1luAb72COA5RXuFtmIFrC59zguFld1qARMcPQb+
ksJp0mxDZzV61vJPYuKItF6r6crviRzCI2wz7KlQb7d7cnKCZCYXZ4P7gyeEDjk3
/v8LfBLeO2+nied4WcbML+8GCPqR13RPLJkLyrqDlnz2Ls2hb4TBFI4Q3dZef1CY
pFga2PNt46KtZr93D/62A3IBMWYvxmpZ43xdYNEA8aU2Pacs1UcTLy9a4EB6EpUQ
xLL6XiTUKSZY/FmF3priubOAb8oXAz2fozwHMhE6Ws5GzqGy4rXp2A1DNcZ/uZHc
buOipAa8XJrRCsgLj1IQwPXTM232DVoDG/u2Tr39ZeOSJ2/GShPl9d2Go2foKo5D
tSpjbs0WFzMq3jWeOeAzXS/CGZaHJjY01uKAoUHWlMYf269vkTLP90AhZsl4opfg
SFCMO4J/bMYLlkf5vz1OsrhWSS/R5KIOamgXD3dCXmV/ksngaTDnXhKYy0CgFuYo
lEjjV0OQ/e3QuNRQHMAUcC1qNwIxNVGp/jMwHBQqolmh2ZvcrJuegB1Nr4xF0Qjj
nizLvVCPqq2oDJzHGlb5PnVS4eLPwlrLFIspNmowP2Sjabi9ELh+GfBHiqM98R6C
DBvyKC20iTwn927JOF0S/r6RoQcdIxdsG2rLmfD7Gnz/UfnXmEgYulQw0EdaDNT4
MVDAFQUI8V18aCrPhVNeMEQqMSmOnPoLYN1Ij5CHKKgnLaJFGJ6ODC7xkivfbR7V
F5PhfuUK8KaGD4+icO9yzMiJe880OgoMKW6PcyrU8fykveZEVxPiDV7h3Q9QyGbV
sZDn9i6/I/NrmVKyKQTt/8ykfKgUBWjS6ajap1NkUhvjoLOYlOIpSKT46+4ABbm5
zo/d++5DZJ0sKLf4D6Utuyg+eZBVXaz8amSWR+6RVG7h4G/JPnngLtakUoPzJlWi
92LCoyiTJ+EbATVZZMurnW/oxYiF1oaqoAcn/b7cI2+EZdaJzpSKuLwpdF8fUOdb
C8DB/lYXzJjmcjVNzyBmiH02stXp2Haq0qOX0W9/wVljfic8kkkaWxjJJK+SOEhx
LEYWvz0tblK6Qrz41i9n43e4J7OPlb5jLJ+mmAh+4LfVWx9y3YbXVsffwhR119eU
93U7rHnc42MfjcQl+utBVwt6TvxyDubZHqTm+GHo/8ZaUyWLQJ68SuQ8SeyL1oEQ
rHE+2tJdFUC6FMBp1kVpuawXNj5IOoBatEiML1jSVFELQsLSLo8t+gl4jcLBA1pk
OWgoQguRtMCAsHmGRzaMjHyinJkZHdCgwKD+amT+x3aMm0fWvUtEytQitF2CIO+f
XsMWU+N8J9+zK/f7jBXH9tYoP9gv4r7vEpYOQMNGZyFx1aPeXK82Obe1G0/qZYrW
zLKlWmMluK8NXnkYmJHweDJeNciwCwLmV65ZToSe+GPgulzBwNvzJM0UHQiIY60z
26kP7I5vWwrlmCb/3WFxN3XEigqA7NQ48T9KvqRNlfPOb8bjZbPEXUb+a5vF2bmq
PdqRJH5yjHDRO1PIWze4yUzEYEuweJk4JV0w3y7WvXtRwgXlFUXZZWaD8dlD7j7k
q/QH3EZgJMLo1O5gE4EYD/EznJ9hkmNNwN+9HYJQ1poZPRkR4JQgzPlrrzooR3he
RneNDc6Y3sIeRgljfpbI+iCBmnjnQDo3J5sjWtZEsDGD6UzO39q4XGZgatfp7D2N
3hCcPFRIrA8CVnHX5M7ylSwk7BzRXtwxuBxCIEINJxc7tb5z2eyiFebkFcJeaesl
kIAgK4zKYqtTlkxvhWvqmKkeqbXmaxyTZnIgMjNCZeigl/fPqoeyz1BIzclsxE/q
aV5AeCc5IxamK1qDtiORmihv3ugCboyT/+72192+vnw9RIUZBHSOov3ukwg38LJh
uS9pbyPp40zyTg9Y2XAIhXqH0zZa10TpUvtwK4379gs6EgiJXuM46NkVvR7KjbiH
9DVpmkMtEGAu1rihTUUMazIEsBjBhpfrzDr2/E7Ys453xxnNbhDBC2uUsHom69lt
nn1sKReb3nCNAyDfsnpU5s8sha5jwI6fbxFqYjuI5RSRr5+647IpzPPZMt7e55y6
PLH6KTRPk6zhvk+YLZtScz6XAhQzScstVjaOlJ4Td+UxowuUve0JBBYhLJI/t/qS
d8sqV3Icqle6GPEof516TPi7CqXZpdNgSugr7pVqMKpMfwFYeMYYa/j753dkwFSo
S2BjZWOLdsAtdPQOn24NkUsL/MrMpWxeNm7v7YdQlk3wsVctlgis9fAFZKgydhAu
kjSzV8u38vFJ5NJBU1LxTyGfFhmeTG2fDiwOPatWIzoWGxl/bID6DZMZp1QMYjS4
pj0wIAp8gXUxPgQoYOdOQAMGUNX2/kCYnjg8zfc67eHNtqMOSITSObbkrZDoauyz
5420QmgClcaRS6rQJyfqZZspzJvsXrX+bT8/eL/GMMBJJlwqg4aw70BqibFOUfgr
qmSPtsmMP9M0KdV5Zos+viRBil3xu2FTH73WTnyZbpsWMI8Dn/gXLCWPR3reYiuz
+JBh1O+EALgHAWdmBgZKrtjXw4fU1gU6htFAMFthke+iPJbdRADK54rRPAjjht/f
Z3s1QAGVPPHgW/hrqV/V0BIcKhPfL0cyNOWifckF7ce25nCx8Gv6PgjTwQ32aP+F
AmiAxKJnb79vCbuDQY7U3fZOzy5pxioM1I/rliypHvozwfvvU4mRmD8dfSC8x0vB
AhllPHV3aqeNr1Fo5jTQiVxORhYxTA0IdER/1VcVo5mLj/LwQKXjaODVNIrV7IUS
W58F3wGia2J/cOA1PW7l3lZRgTqxBIY9/Pe+FsmxVqRjRRhWBA9eBz5PUL+RbeEN
pjb/2cbUA8uarv1KPyK4pncHxM2cISLqfUMDd1T4GNeQPDS8tr5MgJvioJJUCWOH
1r+zDTOw4AvtuPIt/Vt4VOM7K+vk1iC732oTBFxXGDi3ExKV8N1pPPWxFnJkuQxu
Z+q+i2ibVQGyrxo492t+LXnxF7YwIUSyw6CIZamZKWtW1ll2ZYNHtEnp8TpCd9Py
r2ixXb3oxAyPcIAz7gBELgOyFeJfh6t/+d5RVCwcQRE/zCm8yjjl7NHenLCWJXSC
MEoqeQzf3RjUhJunWi2qXOKSuem1K77nOv9heYV4kVUS9QBcaduGE7y9ZUivKPsM
v4De+C+4TvrbqUKmo3iWbU8Rj/yjqR27hYj3Ql3WtQpAXzKPEKB0aPT6OmC2nh5x
yVK+koQhsCjZqJaWRZlBKQEIt2cObWzz64ypxQxPxaDmbPFXu7LnBa1nJeyd3f0p
L+JmdrNkX025wWLb6OmOqF28eFcm9DDYad2NF6+JoD7DDnXRWpM714wnn+vexrmf
HPHV9zAgDjh1SuPdp6Jd3gmKdEIceqsnP6jYp/xsyWWiBeAGslNurGdLtODNpRYV
GcPMmwOLhZfnZdr3DYKsWOhQ4YS7HlCSCI+m/gAhSHWC6N3AYvd3hhNLLRp1khGy
5b4RmioM+VvwrZZ+go3cvg61mfEiYw0KZkeBjHkivr6Vew+K0X04yBe8XMzSxDak
CWds7oIQENhzu0PnP2LmNlVvj+XbounG3xdCqinwUKXlHFTSnXG7FQB8znWdp6PG
UZJjE1uH4uh/yl5L5YXuIEKRtSDSPlsPvT4oLx1QA7654e8ZLGWC7Fs4w0vAcmst
bZQf2QENmBkeBqpm42F+gkK65gWUKYUVwYYZ5ZYz9ssY33JW56Nru4LvDRI824UI
gbJ4a1Q7ii8/61dan/HZIsm2WGjN0ZL8I3XJYdyr5byz7Qh80sKI0bV7E8OldK4m
hFWfFmU5LRc94E7n+h69pjU1jFzNiJk6Wpd8q+pbbw4yo7pCHZ6yN7iam5wN4G8e
7T651ReC6o7Pz/E/nJVzV9r5711zgkiAdhmoUv6nlcIJqFLfOKccFyr8zS78DaV1
oo/3Cw5iEsG2PSnf/STzSgUOJ1vtCWoWhxSpFRfsJeU2IsHOkZvgvm+Cd+8mRM0k
L7TqplqffKgt4qpXkkWgTI0JWXLgib7/jGyU1dTQntPtpiMBBpKFKxVPiy3Q1O7d
ALR2E1PwRNtqur5L3i682bupfndbSixshFmm7TtwXVfAlrU7T+IBmIa6APQ7dbHP
+55fvmUEyq7GdcoduVN5e18pb1msxEhYZMY36URBuHyS+Vdf4BM1yLy7uDAia5Ss
sa6DwLSPMKh2C7i8IwwWrs2PeaX9BefpbUfa1OBLWKub5c4NLj9EDhwuVN3aI+Y9
YOw6nUZnRktShVyNbmxR9fyxwpa3ss1de0cNK65wumJIQRpl8+T4BA5iB65srxj/
Xj/EKN76z0Hc/mnOj9jw9HKMWaYruCCW7Bj1CJm42OVMMeDO2egltGhz7ThSUmZX
A6leYSszHr/o8q7LGkHH1QXiA+AgkmMhwVvH7NTpRAfyZatwj65b00fazyxG62lA
RFTebODI65e7EjNxmkhFiH1laNLTLwyPoWzywsYQMmnmgLfT/kuFPAZwR1P/w18W
3ZwI+Mno+YBtQ1Q13ZfJjuIuVLHvJMWvSWv76ZRKiFele1A+184Kp3oudt/2Afag
3ytkDss5XqcdsE1L2rC2NBDm8i8hwB8y1bEosnbHGrTk4y6yV6gQRf8r+yiSa1vw
t2b5YVGqLvOrDhWu2L2QK293Ndir2OxMMgEWebpJHesZ0DeE+KDX6y0Z6VF5ZL3T
JuN6H3kxPrPkY3Q5RwyVal5hEd0HNW52f6eVJzHbMFvZzyjNH4kY9QFDXAIh23EU
ypMd/CvM4aoixxZHi49A4UZZd/p6X9+FBS/NplFt6EkTf7dFn0qdrfvfQiVLwtkx
zF9vLCDuiTg9z88xoabcubL1LHsiuwYNTzXWNAAfUNJszx30fXS19GaXu2KNWNRK
ezkhYPRweqIMq2w/TgKuR7RCk03Y3m/nBzv7MTU5wINLs1XUpN8iuhW7ycMT99Sb
qGiwapKW2xXHShDTiHFUVEgMYdqc+MFZQWdxX6PtPm89bPn/5+HL/mKKhLqxMfoF
59qObkxRDtzZt0hjhBUY94Arn1yRCWjbl1rHSkofgh86TJm4LE+CK5av6DJXThMW
tqZ2McDyr5mmeZKralYeI4L8LhH1KkmKTSlMSdzTtNSpM/bViswXI4gmOQ1aWG40
K8Bno6FbsIRq07zHJpgaps366dhxdjZwWm/5YBN92rIEcLNwsdSKEmSUrWkyn32m
2olbLjHia56dTXL1LDkTD9l/WeNebz5ufe+kM5zJSdJiNluvEqUA16yshRi/80A3
bs34MN8TzviSo+2S403B4OlwzkHwBHQuzIUv98MjZnt5Xb62PC8BX3cNpHEo1B1c
7Tp6ZDTeU9yR/lm68LcoAWiC3VUqSf/hD6tsv4jPCVD7XXwmIhCg5QYTWMBR/KI2
NPf6X9y9k5vs5GYT1BrW1lfKgt489CelL2+a7f3gsfnxzQUY4K4ojcg0vmPOkkWF
e3sywQR1uJ/beiDP12igQ0c8VndlmdO7zEI1B3xF6Cvf4fJcR93Y+cZwpu4oLlLa
ipiNAIe2+QKuoQbQ38r90qGhWsYKsAfWUedlUzAPhYG2bSDN5AXEK+Nb6zfuPEwa
63ZZu/tvHbB0uXOHRrwD4upIMtuRaL8ma2QdHhpQY2CL0LIKIN3jDsaI9aq0avC9
laoco/cahxmxZvUI4QmXRuYBJpJnMab8ksc8k+CYTc18ZQRptYdJOSEDAGgETX2/
G+FH8FyCDpXrri43D1mtQGLNYaeCeR4PX+tAiX+FN1WAWt9ejFgmfOy7RahBoJtU
UZB+0Es9nmCv3NbXFB/vsnGTolviaVozHQjj4ZawchNkld8K+n9UeRQwFrpP7ayz
Ee0EM8eXpj5ygaleTZeG8G/j0zPVPGEhUjBTwWyQdH9mYZ/kN3Q8OxkP9LU1n6Vl
jluv+WqFQ37L1fht9mW2EyUvFEluo+7mDGl62S5W31BWhAxpXOUV/g/r5HNc9Jgo
zqG6pSJrQwdeQmQWxeI9PSi4JUnyfBkw8FJ8eXgU3TQtDHLgFb7qHiidQqaVLhof
Hg7pRiPtahw81snVF1kH0Z7iSYLvS9duRI7OliGHfzwymXMklENz+Kh5jBE5465Z
PI3H3q4ThpBqLdnbdm3Y8u+/e6cwAZy7nj5kSIv83GyDgNfCCVyaWMgpl9pA8vJP
Abdbuy1RqZvXUEUe7a5TV3ZvNn5A+EvXVqVSByGghU2J+SzzhO2vpcS81jskHD+S
znxEN4TFwfSvvw6kO0gxxkN/+kQgvVQAqCfVa7OJHYvJxmpVU12FLY9arhn0XkY6
FsBedh8knolDPtJRM6GVkFLBhlxxcnjEEi6CMFxt//8PWjDVu9T3a3XF0nERbUcH
2qhxocT38fXJDrAU3hnNBZ0IFWFxiQcUxDsn3VH5muNXxZgT14CaAiZQEdlFlCcR
Dhm5rTJUKzWeuoihn0dTKGFTzX6xYegZTRIsV6PEnX6WmA4iw3iNLlmh3anvaXrp
t2MGXf59TiVgi0pz8UndRI6IxoqAq1VnMTjK6ySGQe3/gsKcdi+0nEA+fErtlya0
OWsOJHnAmmWKKdqsivn/G+gulnNzzrHJ/jn2QMsyK68yXuNm+fB+LhIhBrqyDjT+
hFnBJDG3Y3v8N0VbgSmjbY0+Ev3W9VlEJ6dCylsyHin6p8CwyytYXwN7do9ufkXO
AtP0/BuY/P4pOK2fdbgcwXdcQawkn0qBo+jpjGJeElbFxJuAY640200a3e0CxGMC
jw0F3OLeIjz9M/smdv/wa5JcimFi9ywjHuQkpA+A+1/1zv+4fAC0RYMbiYCFgIRx
SrCCdO5kaEJQg/V6pCP4BzSoi0eCceBO4z0RHHcm2zvmuxAuwlKRthK5OUkpyEP1
kCBHCgKokihWEHfLvjGVjDip2BxTB3y3aVhviFWZRgkN+wLica2yyGZ9+1kjTUrJ
TzsJipNgUyIgR6GSzx/D3SKobIWYtuMOCAB8e06Z3xBX0P4FwZzYoX6NOylHcfn7
Bij5qRqoC7sihzjAUfiOpEdZYs/kx9ii9WmjGmf3QXCGfzoqTHub7sOapG7vaZFl
RP9z5V/Ddswuo02hdzcJZejV1SRsoomM8gJoQ/iUfASt84G4Z0iVU7FsgxZdfTRG
iRSF0VwJOrX4F35hEUbU4QeO/n3l0d5nvibDlL/VksvZ2H22bD/1aASugzZcAVu8
ET016ZZPY5xHWrOOummoqgGN4jSllmWVGYDExa7y96sxxHw7sGfRIFLhd5zEawmD
PhlHhXPM5f6IQ9/2n2wWMhjKLf0VoKOS/71DGFZhr6RlZ9122Q8trQJf1FPDsO98
JGSZ/fwBwc2T859t7d4Lesu/KvHF+3UfrKl3ZKu2c5D8V+sBSxSOd1Ue7ID+tG4l
JB/Nh1Wtz4QTKq/1bjkuXGi4EnL+Z1jsIEXVfBwC6qXPVLhJNZUNCzL95KDOGyFv
rdpxzYYPEODFRMMP+TgQgBHPvSTumWY+XRlGPgnpTuQktJR55Zdwb7Cs1RAV7XKD
TUTJr4Kj5MAMfnWQJocN11VtQkg7+OL5/1VqdPXhs/I9Ro9qlX1T2x9Ab4LudhVC
n+6myEM4k1bW8jImXAG0hPk8Lb2M0w8QOS4T2kezfCFxJeLWfGoa1VgmJpUl4myx
B1LGMoBsWez964RGbIeNY5CN5o5xjQx/I+OmdR3gjQM/Cq296fnUXD6sjBDzRUWS
A3FERPyh9v+9ZWY/Agb8xkkIT3l78qRyII9fV4ieV3d1T+jb0sHYSL/WeAFY8wsm
pq4YQLbHDMi8iIg6TyueCyJ5HY+HRPu67hRTICnPg7lJBCNaPvcS11XGAftcreO4
u6zUShLifebeL0AM8ExcBu6+yptjyxyTPLCgUq3DdM4twp2FEPqPSJ3MyMruSlha
X9X6uDnIDPMdwb79iHHBfU+3DRY6U1gLehO8oOWZiXRFjaC+VSDYjS3PMfKeFkBZ
dp0PxGpnDgUTNs8zl0/3F6byn6LlaEEs2QOCESnDrk3MNScMlZIpqoFsbf5Mdt1G
rgRpiVmIkhA6WCDrJsoU23X1KOBsjgGWXfrlW8tTNDS6hhla6FWTrA9MnGGaBPqS
OrDaat16FXLRlp5uoB9Yw+cY2onuF/4it2TQh8/qI5ROsQ3K07aQ0Dnru2CSJ3tf
vFBZoh/3ksTcyXh+K6t95cR17Ex7yxI0BzJSzn8SzHTGs6ZevCx3DFxsvFFVtIYl
5+IwG9nRPc1Im7xrTrbvhXALV06fkEA+Etmk346GVTdtWYHYZPzfZW+1T95bHOlV
CE9ncQ2MF+diZaPKqFYTEgOI2WA04ENlAlNkn1twW/stS9NP3UijVVB/KpK+8hQn
fW56jkvZxSDjoBaUvJwA8K6ibNNNP521R2X+bFYBl7NDG3jc1GsXNWQbqXximeEE
hIO2cxOwUMJ5q+yWCOUBvQ9az6CD2ks0mQXyEMtBdepT0EpswIYetb5MKNcH3CTt
Y+otOzpdgL8DKA0BHZ9RbUC9MTfOVFPlrvHLhFm3BvQ5AlHyWJ+L9CONGyKIddQ9
bZaKBxIrUHcTwW1lrck7/JPb1uGQ/ONquC1OiIkwsAMm/gnv20nTJ53IZZFlMvLG
MYvKNEeuQ/2KYoJcaCh0BElUucVCZwLIP+IQYov0VE9wlwksXExabUHTfBeBilYi
/ZpXc/ErWZSj1UQMHdNzHDu0QTNQG6bNPOzLxMVHTcTLN47P6oMB4EUbDUY5o0Ao
/q7rCOyRhNHgPOiCeDp5Cc3QWxrVW+1BhzTw81wFmgj8Ak/MOrkA50qEULwXt+Y9
mB01MFjcTjrzcf9M0XLC6/+QGwpRowf9QHXzNNFWgF2kKxgzIN3wHMBUb7TPRr5O
5jVb0HVzHl6+dVbzuu3mP9wb+LI0Dzva3YYwzjMx4iqm8TugJStCbWPAvovOmZZH
K1NXUIBmWcOCpFcy2jjBhaPOJlDO/DTyQctPLono12Bz2utWuq3slu0qSEDa3dQb
lMqwWRRpty28SHKjpzkf8gmY4d2RZI7wkYyamMZxIz8ejssYqBRZQDWLfwWvo4cT
I4KW5MloMHpu6wdWKHx6NLkUA7yj9Q8MZ4chORpH9F3lRGwzmUThegyEWukxcpOK
BZ6pPzaeJdyqBFr7Dsr6r0z7edCqxRlo110WpEzY5mjGwla19xA7wd77RGb2qIS9
BmrRjtC0GpASbFmfwtlp7cR09tbJNObNsWX/YGyLqutBq/uVPaCC/trP/7gibAFz
hmIEuZ50f3sEkwr39oOIoPoGUvzQUFARmZ6CKJzGnCrGm5B5gC/qrsi0kFccbrpF
88N+ZiGDqQEJz42FXVld1ex6NYl5CT+F93ct1r8PMriuhV/CR55dtCTzIx8e1/i4
HIxTKLPl+FVsviEQZqUcE1RuHh2dXeWIDj7fu+6Kt6so4oi9cjZlSqNeoLHMffmB
c8Cucg403+64A9myoOoEiWKeCWS0hn8esZN7dh4XaNKyHgyg04/hdP4cKQVGRJCi
B8vEO5XmWjC1kEk5m3xFpLyhr9rrcamBqUNS/qY98U7i1NrszkMYFMQZ1eoFAdhJ
bE/leKb0CXyBhyxlMz4dh9XTBJnfJ6zI/rDELFlqJlW+C4Y2R87Fu1fehQClHCEb
UCI+cu+UnyAZu6pyzPVSEaWwsq7laDMPvPlz1Q0u4ZfSRp/V60KFqHvY74TP195j
fBvfjNAe/L1CYdYbtFuzUl5YbCI7jHJM8F4VRxlwX3s8jg+O+zPJNfn2x40tYz/S
2jNRTVBaeQ/LVMqMsnU4eCCSVHdKFMDmb+4JyUc4JSkCYBhsP+2CjksFTiHu5aqj
7z6n3+/Uy43+a28Iqc/NFPHxRg/g0nvUqPotHrHleMpIoEdosn1tJ9dxbi9oJBgt
S57sRaIKh89tomPgLDRajEChxS0F/XyzJYtXRFtHIuIOxs40UvV2pasPsCWA9zMB
xwfFKT4r9eKuCJ+R9hh7hC9PZK8g7h4Rd4MUQyJchTlBTa3h4fqk0vONaeVwkSjX
HCb3F5rzFhj3BNxWC9U81uIjdIAVC7e/FsJsis5HcZVxDNlkXCYtpXkKRzdybVzP
5imU600yB1KpogT1ciOmbb+ZXAykQ0SA3ykHDN6EVeaMTB+n1ABsmcvDvwAwsuD+
Rt1GC5Ho2Zd92Xd8ECQlEYVrg9fXJ9Q3K+mcutCpfbLeRZvb374QYOZE+ZmenlCz
UpmOKiZ1MKEZ9Fs/Gv5Qz5In3Sln6RBSyKAYpR6V1Jx3lrjF+l5/i7V6aQprSsDF
TTLJleBEf7AZTWiYNxEYoE/xF//r5TXMTErwkY8e6wpGRJkVqJQoFFlX1uBDLvvR
CdUjhsakmNbywIgSk0k41LOQLQe2m21bjrQ6ZMFvBgAZ/DOs/PZn01d39foxIZJ0
Uqq7hMyHPCgA8RHu6Q0wTbNbNZ5WWA9KlNt5gsDH9r9olY6981wDF9bMuNacoz3d
uZj3ZKBeUM88t8hfqgk3uNgu3vsqNcs9YAA9dR84aMji7c2b1xyTVtSH4z7lI3ci
ARjB+rpZpX16k7L2WZ32iiwO/ZjDkpC5IeKeZueO3/mu+XfiXlX6d4TaSyP2LbhW
Uj6cOnBpxSCvJPl2YZbYtJ4glpmK3VE3kdi7Txbki6Np1uTury9Ly3kVz4vBsI8T
OpV4+YDr4dP1b88GFoPMcb8Lt886PDtH2cLtobC1jSazObTM8ZHa+H+PqGlDsdlx
QccAgZ/Tk8OyPBefP76DoeuHCVJBaFUyuRpcSsUejZcNpi2gmK3mVz3VAUkuiKAr
Rdj1eJWuMSCQ2J4C1yJV/FqeR+pWNpKmLFCha3KVHJFIfxLj8yXl6PXqsiPMWwML
S5KW0oqUXauRhG6TztU44Y3sQG+AjRHkz6cuyHsEVd/BL5thEVrVWPVjgslNamMJ
g9yblEulwVtmnr9U3zxeHNvs6slw24c1F+lOFF/0+qSYoe3/8pJ28ZWM43JyrG7G
uDS85MxhmWX9BN2SnpfLQzt0wtMlrHVcqzDV14OnrnYyphHrL5auswhJ2iCdgiKZ
gQhkrGkuiQa38nHTJTZpn43Zw+W2iAeRTsstDQZsEBVnmWP+pdsDb3fz1tpcZWXT
Qwqy40etdUSNduKNhVZBEvjiz4jCAWyE90x0VwmAEgz1jpmdPBArnVQTxTA7J6+i
YXohasWcKxxJ0m8gDvYr91Gt9ES0yWV8szIaXObwt1l0D2Hb4hRgYOYGvDg6vCdV
zU0yhk3kvn4B3lrBAfQ+eRvgjcBLGhAuwF3d09l77V1aZavnedbLTwW68N6UELmp
eH9knjjbitabG7kZSWr+DoHT4ucyIv/MDfVlBktf3eGO4GopGr3egnNpMeLBXdhs
n2X4wT95PL1UgrG6U728ZYb1ImJ9A7HaM6E341zdX0YzZipAvvaoJX/DcKat8CWf
LxyQIPcHYaZMp/ie6IZYaX06w6w2z0V6DBI/CPBSj6/4AZ7zkcMk0gKBWVEW7o3o
5hUEVZYelWHlavtGIBBhVukmQSfZwxAuSKBtx3zKWT/mCU7QLx3euyUEml5ytROZ
kr70St3DG8LOANObzlxVVxfk1GW9Cg0Mg0XLcoX2mYfhOPFi1vuguwjuXPNOgRJc
e18owK0UsHI6OqnO36Pi/lwV3ijNKV0/PtU6QFPjPFYgX6qzBlsaeQL0pxQ4hGx7
0EsuUDresdPLnUI9pPS7w82/Rh/uWFkRQ9wbrRYOVcBW5NJtln2vgPg5fw9I+WRy
GwrNmcWzI8u6Ka8muTWHwSIMp0PWocFvCdBlha/Yj/F9b/6subBUdsCUxAjeNJrd
o5M0UCqLjhuRpOnuxDglPz01Pl9B6Ku98m2GNo4mxA2/yIxupo8fPVbY+/pcro2A
qs4i3AX50qPv1dHX1TOC2z7axUG0BRc8fkfXZELnmF0vWGQx02Q+v6IlfwVEL8qV
uhbeSiQGmnWrhgZGkSE5zwgbHrt3dRURdE/XiqPZUyvogZaNWZNsmH9jrSEMs49s
Z0Ril4AnoGrn84USyQ+bwP06Vj9yGmPhBj2OtahLBX9F56piBDmL6GA7AbleoHg0
BSXjJ35lzHv7HhJE3x8GDxfPKZgnHFTZ9JydiUUZ1J4RQWbPSfodzaAxL6zYozS3
0/c4p/rxMt3kwDS+Lml7yfvQcizsSmNpCHFKe88gC7yhjU6EBp0QfWrgnqJ76wll
yCW3nrg46A8P2UtWLJASReF/01NJemwJnrH/Q2iDCeaRf0BLzi8KorhVpeOfrMtV
wc9U6CGLAmtvdxdoWVGT/Td9ro6PzmqgidbebtFdUd5gYjMog157biYdlE4q84AN
h5+rmIZpoaHF459rX1iwXgiSAHRncoR7eDOAdCk0ISBBs6TcvT2nA/eZMftOoIs7
mA4Iw4Ppa+g2jGCNnwVx5jDrX7yUJ3pMr1tA/MbZruDAkRosv7P1fj3g2ohVnMQ+
kurCeh04BgC7KY3pJF0T9tnRG9OnB53Ahi1gkjSqGemRhV7wrAGEFzsc8CY962/a
Qv+3sFB1RHRX0jTxPPNbtxaYeT+VnNlWFl/nS3kLqJF8Nu/APw2NlIjNqZ1AAYcc
AKpUGkny19Wku3PXAj2AUwh24zSYWuywHXkGy1v5J1I05tZnDd37x4zF5hiiS7nM
noG9dQLrJt39zZkGKtNYYemIBT0NAPEa5WwXwcpXL9+L+lkTSTpgKcAaofYFSv9E
rn8iu9JmNeCyfU+ypr8ccqhIumkaRgusVFkOgF8Bjk49+wbg8ReUE3cAdD3i5ym8
9G6ceHtMFl7/X2dhoHj1Ej6OfQLenQek8poBolKh/8atu7EBLiGtSqYuvUiqGfpL
X6k/Nqs2k3f++I3K0Emktb/U4pU3FdxsbnDZZOXwWnF2IARF/REMCif1N0iFoji/
zkuzr3d8XfkRpiM7tXU51qQ/vnsfTOX3jDUuYywZmHuo8lN/ZgFF15LJ2xNq9Ec4
GNZcOvBxBgbTM1XHzVSlVt0LtpCkhY79EUA9367DjZAK2FvrxoSlapRlNi3vFYB5
vaZ885fi6M0xTARkpZhGJt1kqQhhMXGMaAV2ZAShB/C58SlTfKXFBzKYUIJjXk5m
yAhNuE1O7qghHJp4VEAdnEFUsxGtY+MEzWsPc3SStAG7R1h15ChuwfEaC9xfo21a
PQrugkRGWLVR41Wp1FJOvRveAhzARvNnGCAZmoZv7568Rn7LfKw0c3NVgBxZsHnP
DaffaZSq6lltBcBNFfDOABHvfMYqKn1Fc+SrXI+DLV2uVWmYshJ/u6gFWKnjA20p
wfxImDQRmIpnmB7nwuERZq746USE6QP/ne/kvizPqJjIbycQt+0E7mvsrRT54iQ7
z53Q2uRo2kVEinfmsKlnXf6Akkpmk2NkOakcKL0nNcDGQ2yLUtMx8zmPHrXVHoGk
FuUalPmE7Vr7tybf4BMA/nSkguoz/w2xMfvPJtJPDwBdSXPFFEnglUgrNMkVj6ef
bc3GGvjdIPEhiL+So0S4zDPp+JF66itoefqqKehFFxLom09jmizLa6PNI0AEe1a4
0/MZphtjyRqavdBjIQqUPvnV6UsZUwoNwvmSQLifN7u+BjQ0/kBQ+KCL2ec9YwO3
vU4p5o2/IiH1QE2h+8ZHSa5/l6kl8SIZvZXpMYhEriuGp+5kknYG8rnAjd4P892W
r3hdBOsHb6m3Eb1eAEIIY24TbsMDJFlmYdDvQZyqWqkc4U0L6tGEOTzrDwV+AKbJ
owW3iBPl5jl4u2hhVdGCinFQIy9IDGuuNBsl+ftFZoTFZr0TCXokolf/s0qY8Fyt
IiG617N0hOMNqYldAx807RomkIn+UjeYIFg1VhhLHkvlCgZoXfGJY9DDdp25qZVd
In/5JjULGWIoRBtYOf1RPsVR1H2Sif2UPte6QfkjX0pBhSHcOae1J69NzOotlx+n
p7T1x7HCgmwtD7Nto/OWzzdRA5RMENpk+HiSKV1jDT3C/bf5v5K0skYlrt9zmBSW
4UQAvWv9dCnnVSkl5IfMgfENOTyVr5oL5Xl5PSGrvXFRmt/u+1bWcg0wHANKIkPs
927x0BwNpBVuPudjiEl3MFLO5eDSF/s1OtlDRC9msTepRDbVF6P3qt3j0r7LaQnb
WhvJJ+cJIoFNRCtW7zLuh7ECXnurnVDpLHaEEgINTcxcZ11O8wlUEST9Vyk26Gib
ZS2TySk4CZQWRSVY2N+euEdKVulzq8JNGhXL8dp1DQQCzX4BmpEXyazg23Mqx/eJ
3V5oHfbLRlh+2+VS/bmuCrK2DiFGyQILiqtggZ1A+QjY5Km0u8OGJ+5aPj1EOirI
LG9wo8xmKUyYCoJqZS4G7JFfKmVhNlFbrfWHkIB9G6VD7POvtjf5IEyq1BIUGuB/
mIZZKo3DWLpmrHuP9VPJrpAbD/DdPhLDxf88fAQjaG9XTDeoQ1krDLSpQ0V/BpXy
ZWeTz8K60NyOvHuvoeTiFpcu7ZaEQCIvBuCs61B92UgeKJFTobNMdoQ10bHAyS94
wKSoeSzz1xv7l2ZiLpiebatg+T91TTkIW/QusjUoIdhqFezBHhqmlG5V79Ga/uKN
EyT6jcTfgQEFVtPiW+Td95NvHk8bEf12T4I5DBLPEzu6J9dDO4UONtz5dFQn2lOV
x/phvk8kTSzrjxQiOUt/2GP3+UQK7jmIlJgcOL10DfarLSjqgSKr6a9Au1lTXNPI
Hm56PLw4C5HO4v/Tb+vamV0eAgZ4FjEuL820KS50Fa4CHeH10rK9gG8Ou2ciyftY
YWobxNSuU5Vmg+yka1WYRoRPknaF9QlbXA2Al1mkHJjgk8MEhp2P+uiKkXZRwl4F
DJ6gwvTt0intUCWf9ClrzldPVq2JAtRwH1RRon1xxRYyW67tDP3a3vduiTNBz540
7Lb5B47IB9b7MwUvx11WNyA5+Rk+L6DCKT6f0xGs0OrE14OXFieZl+e+WXrG+rAo
jv8YLMCUYs0BXBak5ORb4x8JK3ZyUghs6AE2Utx7G+SUQqRGakHEYiKKyd6+WgOf
tR5GwJUHVcK952Wjm90d8C7+atWo6Q4ji709JbOyBNRoGUzllzcBBb0l4ZhVo78k
BcV1977YmjOaJFN7TyN7bIk4kHB6JS8qkec3ODGzMrvfjwxBOd7Ppl2HpvyWlT7w
9HwSiK3880VsiQVAusa3UJqePJboaKOmwm//eeqfnekoRvjlRAYhHFBvQBNmJ+w2
ZOrKFmNjSH7xeeCWysc5DMfN+UtzHAMwM4eKufKVE3BLvrxkTGMu5Wapj0vh/1Pf
S84Z0Gjs6cvLcAXKP//be+0dK5WO3RBqtG7bplFvDOllg5zuSP9oQQashDPAZ3TV
kyuzhVaFQ3dE6VS0csIro1ay+3SnZPlAPvlYmrNaxJu+Dz9sv1cqs9XBOkssqy0D
BJ2kgaHmBnSOHxR1SqqEAiVhMBLdH8MCH2RTsVx6F27nrY5xF7HaXPWHr+aB8zHl
c+TpcbvMe1IN/liFWSAu32X4mEFv+/030p73FMDhZia+F0iKOVdcR7pT9bhN7CW9
Baj+6+xXbHxkarcbAZj2/leplDSNPW4e0OQzed1rE13uIcdoNMli5eAxwNiGTA8J
dncVfdmFawnUu9/v98Acb2hNhH/1HMXx/ksZOayMEJo7gi8qaxROU2x7RSpY6rb1
sqKZObJgzxFltvT5GD9/VSt+ay20jADM/GZ/Yqq/gxleb3+h1ixvyVvWJGOD0XVM
G25bEewjlJa8nf6BKsooivxFNis393b3RyCtS0oyYkrmiTEWaeYXPOvDdSCiR5Dw
fHb0xn/Brov9baOqzzlAUFE9a6z1xgoCdLdq40njF6XCCQoqJIa2IlSKx55OMPzT
28mkNzE2Po5HjESSHOco38dFEUe+tiAwcKuC5TmlHkaYZLbFDaLxVKqXNQGHq09D
v09JF1FA7dSuCyepREqb6NOlqNMS+IJAxyHRPwmlB0PXG1cxtFUo84SPngBs+Itr
WUVoaHby52snpe4EAhuv9Y/BUSOJmXgx1c1WgXHjQcJRve61AKSXaX1uE9YFz/PV
/gh+ywS4s5u03D56h9VmlkVR4BKObSBIxCtOw7p17AP6a2B2MF+aoTotphLCD8Yc
OETUsJkecz0oBdOpojNn98lcBd8xUVEsOcLLJ5o/M5SYoMbjXB5wkzVKD4qWVWkw
8CPRREKIdiWm+DSEe5qjCg==
`pragma protect end_protected
