// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
RrGuvl9T9kqycjtz+eGK8kkesNVD55iki1nBpq9SUMF6GNg5kmH832puuHgrSa5S05a10jn+ogvM
P65WKI4vfUW1ljFJ5HnFx0zEYoTsLwQgmuQ48Ms1lf0YxZxpbLU5r4laRN5oeOFMJm3TroR3RGVJ
8x/E+uErgBFJU+u4fxoI4AEoqG3Qh4rW7MWPkedEA3Df2HMJmgu2xBnLA9pO6uWmbBGGitBtJ4iB
cgAXefJ3DAZzZJbn63ol0egWPZmlQzSHjzxgzKbvvtsW3538aJBwtu+esL8b1QHHqGIZwqtvMOcF
fIRToOp89NOkwyTo0UvTUlr50aGjmXqGHaM2Yg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8336)
IPZitPrxj057B66hD6/sRlf6SxjWIAIIrRtsGd1gUFAEAXcpqRElX9KJJoRhfYKvpEgCVNdVRvZe
4uOmkULGAVV0MPmu4S/bwN4KQkrXLePjLPPIsb4cA8PQgdhz5BN2P6y9esMRAEdATWToxfAz6dR0
7UMZ/I1GA6kGAqPuMTU5eMly8Du3oBnB90yJ2fpf87rEN1yDjrdusxp8ar2FpTHwsOqsAkGo43EI
q9KrdjEUWlAlK+SCihdw7w75qop9CarzLrzJJawmp7nwokEM/Z+qkoekDUww7Vu/yy2JC/pfufUO
KBgcl7o3w0Di6ie+Mfuq4SVpKoR+uZBo32dTwhtvjCa4H22VrV9SQLwP10S1x5HLEpvNEsqPjTHr
mHf9OheNK7L65Dp0M3MjcGz95oOtXzpjMMFeZog8wEatLKrNEubEXgBh7dBbpFC5kJ5Qaq2u3mMr
kqGi0Ws8f+QRR0k7S53wqcM2SsQEffP+ikRvejTILDWlsBOcFfvzzinUmbBdxPMGx7ovVXgdGHRW
96bhUnr9CfuBYcDLZE+CNmpWu38ABHxb5z24512Y0YVwfUoVoUw5N6WAGyrTPQVf31pSVgrKr478
2C34mn4/vwqTEbx+5USPDLHPrnMG/t9BGtxiDvDPox2VDO7uBBhKAkbX5yOdLGL1OtzicMDK+rTV
fjjYKccowoJL1RznnRehZSfxJLbVZVdik0RmtWsnfIuvwovr1waqxRicke4xzmzKkdEkLiAg9AqA
+TbUkuz9GxFZCbNVqt2aPEYYQ6WRJFZHhOH7uuvm8fJJnC6kZnWjR4NxM4kAvyevGZIZ2gBVJvwK
WCjSElqvTNMDC5yo67Pxel9Jf2j0alnyXIFImAbVHMuZ2JR0CsenBXUn7jw5L4HTwlwslO1w1Hno
+gqp33GgbPyFdrsuLk/Wj/1Djdn1jW28oMyWkeFkyW+x0Ok+sROtP1R2fTn1E/DaifM/bt9hXPwe
SIXsRYcNzRcsstLMfO47x4/nt1gpPKTQG3XQ0evqGEjHaDOUsiQjEl6X7i6Qxd31vYWN0ST362si
4t1weTMHu/G7928RBYSx4mbhZ/YmWPwH4VjCjsK6SYCOs8d0LCQHuM7XumpoxWRkYlty1e0nL1Ek
izJp3hVnscmiC+qNExqkmpoJrVr2kehpabeexOTN8FBJaiNLlnceXRz+92J9Kcfy5d4J0scWzNNx
JapBMHTMbat0ajMakTniRiU0eDmicZkatxpTDgnwTzqQfZBEUtwEeVwD4uIzFg+rzb6cqEHDXpeg
dTB5AlNl1U4yboQiu0QGpzC6yXivRH63tE+17cSlSJimlLyATcvCrUdEn9rrgrH/cMcKs4VU5pyz
ghAPWL1RrFwOPQd6AxWF48BL7ODuAKRSC97uDdtJs1ibxiBpnn32GVNTt4jqFg+AKqALFCR1oyZb
tTDsQY9ikWGIE1tKOTu7sxASRLNIDwYEi2Gsjvj+fuEXvdkDB0loy5UzpHb694gS14ryb8onD0hg
awm3hRMnHSaXz5Z8FLtP4c1dJd7H9XjanOQt8iF8fyE8TmOKeQ8+vQaUO0bUsTfz32FSyP5LrDXB
xLAPS2LrUrT0Y7a8P8LeNnUj7JQ1eI8Frq2PR+lJs9ut1IeHg6lBd3S3CHNgizpC7KPpTRwFjTQ7
ZNgK+jmFexuYkOk64pIJvpaiM5tE2aJzQRaSoRekMuYnqgTkrCrTm6fElYMS0yxobLR/yj0gd5qy
ZFC1XPwOMO+RGJyo/Em8onDXSXsEZsakL+5ithZ3FtrtWB50RfI9t9we2dHacpWkeZq7mrDUiUQG
9t4bHRGR+4htifO18nWOmEsjDOZ7nz6su4L3XbPqiL7Wu9RGWw/dlFijVPh0NDUftUImFnMOqDm/
8y7J4SMPWF4453m5MeyqF7qA4XJ0PhSFd77HrYcPFQOaJWMD4ih/yAhNyjbAERdnfDABXuSSBeIb
8vEY4Na1tTRq/OcOuejHdmiYg9vFQba9ybftKXBVikmWtBnVU+jUvslL13IOL1ZpwBm7ruIgrAk/
B+SsQ9gO6nFJd3i6W+bvkRqbXmKB3k9tzBJf/jvs4lFdVn0aTEGXuHsV76QqDSYDl82hqFegr0Z4
QzTRF+Ig6GZR6IiSYQ/bWFirUnew+dTYlO7SseQ7hfx2lmJy0xItY4rgRprj7/orC4KKIf+C5y61
+Zf36pNXSYlX5etk25MMJX1i8NT/SC9++3NyJl9i+MUk8xyn7ANZNqvmhF+Sxx1g5z54XByB5oLq
7SS/2WuPOFLxEC3PU9YCJzKf40s0zOsN8TOfoUTnqBv4CqjWDn2HUdooa74Dkz6qV3qbL6KxW///
qFENHpnThzc430LEQZxYXiPvI2ripS1BI+3HJJpU4fJ33ErSAjiXo2YUB0ZmayWfrjdmj8DQUMQE
kQcuOk8rFGvH07NbX/486q3GTnl52FxPqaZhBhdGqwKDc2iDBIrzvd09UdCeLtG9vFC5R4IPG1h3
HVKURkNosGeDow5NZkz46IYS8kMFe9FrWHFfvE/Zo7jqEd66TP17W2wCSNpPSLAyqaiX81XcvpaR
IfxDsS1CNeHW+f5ZtE8EwhgQEEw2GJrs2XECvFKZYhgt32PQlhgfMtJIs1blK/lOPLQriKbiXR6O
vMUB2RJlbLvUUtR2ACurGGoZmzgtveTV0iq9gUwd9sl6hfpT33lypD/plqq39mNCrwzei6SMWJ9J
pHAs7h9rm+qviPp+g5EevHMG7BXlajW1DgZID7w/iiNjaBlxO+ZxY99Tnl1lwHv9Lq9YovJvwZY1
OW1MQaFZuAZJyeV01HWqfrd2OL2pl+ststun47dbHA0jD96cQ6DwGtF87UJMkZZi/1rTH90r05KP
4lejJhdR9rVIGMhjWskMXAkjLemZi4eytN/GVFj30x4kTMOV5C/1iMbnbN1U5CmSpc5zbiXiX6f/
g+AWfDMUitkH+3sxPU0rr53QQvQUQ8kAPwq1Hi5er8ceFbzfndM+Tu9y6evoNRgN4RL9pafFOhnv
BkczR7bfXby8gyAD5ifAkttfgHy+KTmtjMV8KpSfkzG+/aKFFSaBP0SmSFMKaHIsXJ9GedH48tFg
98oRJJFjQ9eV5w1CNEHLl2/zkkBwxmG6RfsQpJnFq5jlAPXoAoGRxed1JrIy2f5pC/pIGp60ChtS
h1teheueFoytoNc2uhIzNsR+NDKH4d4Q/pr53DB3mm+qLuJP/IGZNCczsQR9+dbS1xnUapKOVe1B
Lfj/6mOU52z18o/y/6OduGAPPvIKCyxtxWxWs9a4vDZrBwS0SbmZUC5TW2SxYVsq6ilv/eDvexLw
rXT8YJB+l/krBoQezCclJJh1GrkalEvtMcUcPb5N5c4PTXFXrfn+MDOT5HSmDdKEzThw7zqOP4uC
NYBYSX6Da4T24ITpceiTznsSMAon7Fa7py80B1OtqdLV2uFNFqufB6mn85WQ+Y9+jPmvjJdjBN13
wMpNBTndqSb60+0vm0MwyDx2Wm6GLvp8C6tXqLquvMpgaSU3Zt7C0lnykDtkTw6sghevbiUVu9O4
iagveJRJi19eobuL0vPo/VBWGFvgbMDbZp4Guijuejos1cUG2BTzgdUx2Yd6BzfoSf/eWhtTr2Th
PxFFDySErz/vGEcYxOd4vnDKvH/hwKqL+ErJtqm/v0SYZ+RhDjwRxnNttgiUMs0qjXw3foKJHl25
e+Q3dpC8V9L3DfkToJY/D+bm/rzWldouHIT0zVKWTAn7f/3H7ZZM72P8qlwO1OFHoc5J5DsQ50P4
mjQnV53wbs2BFMSKmkE2Z+snd19a8h4fgDlaP+TEpwOjFsIEvjGPkADas9Vp4hI8jqBzoBcfq8T/
rPSgqBDuVZRkGV+q2PCh0S2vZiiFVROn8/63s9OXtQ5DNuRlaMaY+Q4R4SpXSWn1V7sD6o4xguCn
Nr9zibtH39a7iSOvbBASzrJsIEb7PIFmQ+h2rADDhr+aszXV4Wxhtsyx/gjqo/osVslVEJh+d4HE
HWGc2QTJc95d51/A1ZLogsRq1iyeFHaOB9yYlMWFYfYUtQtGN1fQL1Ge/w9qDX3SMqDyXTQ3wX46
B8A7VSGmpYyK5rNZmmISco9xdZR6AmL5LrbHBcyMTOmX8CmQETbu3lB4QcZtWlkOvYSKrr4U5TXM
aJLG1EtT14/7PzHsIv1R//qoJr3YU+1OKXAqt16b9h7YLUaiqihH9gEAoStc/iETlOyiXG2IMEze
lTdZbbehGITsyuRv1bF7nQKdEKg0lNXQe024oI0erB/3TJj/faHYU6z55etYvec6szrfKCtnEQA7
BxfFc6C3pQlwYucmC18dNFeEB9mH5gHTo9WcnHXT5bOxHCjNN9ZRxBNNpKWAxYCRa/fdnClwtwhP
FYFwMKJ3LDJYKwKk5okYNVeyv3+A5xtw91T20VWTKJ9Hl1IvhKTrkd/pAXyoQTtghKbfoLmuK3W1
CgbuHov8DhNEuzNsHV9GPLGzOYBVMV6/NNpF3wuTNP18CKw1yZDX5F/yZ7d6VUgatK5E/xKSyrIX
Kj77uz3XD8G+a8CIJHgSxmXIbmVSJ56ONlLGgONtMzUdF4Pdkn4oMPPUqSLNG5f2wkywX7iB0QW1
fNtnFKyJommsXvRmLqeGhXAx3iEgS30OoxaSZDVRjsCvKutfNXButGPAXPOELvTudh9uz4qcR4Dz
ywffUT/ngpWEt/iYJF4KYpcG1EKpGOopnng84v5pMlxJQnPUOyrtzqhTA9m7OovryIu86Pa7FYrY
mrByGp+GzSHrXObT49AkAoeOm5GOdnDXub2vLnval4VddNsblG/cLyEgdt2P+NaMHy852IyJpoVZ
3B9KIT3yRw0HXU7VgFcCWb1bonIkd6RrhjWyRQVyedJ42r0gf/kcTx6EQCvyY9RfLiaZHYbaR0wS
T4Scsb2+qnlwL2yRxKpbHKBqnnEZE/3Nj9TS2aqnTkPP/B4bZ8Bn2ekUAHWdz9PlLo+/SJYqAZdU
W9smaSECcM5ww8+19lhlrmkljlWpBBh/1cPAcuMkqIfhadxNFaO4vptJSRKtgOjjJ39CPzFiJ9dL
dRmQiu/IsX/5RJ94XS2yDhiulPQxpXc6RG5NwiD9PmhHgopO3v0h9b1uFUlhg/jJEEzVz7EjaxDm
utfgc/RYcuhGKiAu2VFJ/L13CrH3tDa0nmaLTyeH5/K0Mo3UjGIv6mJJQXNc7kX66UHpOGoEYVrf
Czr+uZ4FeFHB1YQCJ0ERgobsvJQFnpTCD/0DaSYM1cCVXRF3HGawsDv1pDcsfQWPVSon0ArD0rFt
ux1+qIPP8iaew/wLcROaAJm573T7rYOWid/aJGJTUVkGNBGKrY2FsOBLiu51wW9zjQGnhx2Pht1K
KevwaoWbV1ewu/0YsWMf6NzyGO5LRIkhexB56+ohni78YOoQxJbujE9dg3P3EMvC7w1X9SBhAKB0
0GcVzioDTbOI90A3f1Bqz2yfFj8wBLgRVECWnmw9la0SQVgeDd0RqXxwu2EtbGUjL7AG9XViij6X
8/fURfIhU4DvZTeUS7MdoEjWYuUkbPhcPmqfVRorjtiU+B1LNFIPqlLOcV+aTe+N1Uncf63fRy1y
V8yYYdNvmHCV9tG2YgAE/cDOM0OdkLAAA5BONJXCpfeoe9FwGQHGB4C1OS0w4m6tBETSJrqpFlcg
KKin5cjaJT0pCVdjHR1SM0CJt3vBDJj52VqjTIsi/xm0ZNpoSwZX8eWVLAax/3nGXxH3D1ohbo9k
267+iwDoIKjhCrcXOru++hAgy9PeMwtVqpir2vgdfnoH+8XfpJnDS5KcfNCRH0ccYSKDCXXUrrGQ
MgUYRsRDsiNJ972Ebc99Y3fVxaGLXUDPVBaxytEOuwX3ROgv/AZMycOuYkpQkuKYU8fDjPjwcVcq
6uzMv/+01jQPENubkWBjMY5DNowpDYqeguh7HUlsUWq7aCwXFFQiou9oeeboJM4z3/cxyIYkhsAj
bkzDdG4ZIhGi9B/iTFcT0U2duEd8Hhiv5mleqoUs6HSxTfWAwHD8yhkI5StOYZ7SFLp4rycDkWh1
lwuAcdhHTaD3nAJk2Y5HDs1Tr2uZDZLzDQ9iXG5V98Stoh3p9jUrTPRAaw3M+4SocPn9R4j44JRC
M/VjD1t9c0u2MKmrFlHFdYPbazsAp0paBtYWLlXGYJ9AaXY05fCtta2fQk2gKzYTU+TDr1MJw1uH
XRZA/p4Z38sEOrFNoOZ9zartp45GF68ka3V8snMj/fLbuUZeJlG6QWnU0ML3tPKHq4QEuM0d2QhE
i6IBMYZbTV1gojON/mF4r5TqS58LUKye2qmsWL4nVP3+K3aLEYEUVv03vuBmXKDWG/fUPi0zriBT
EHdOc1wIBMP9Fs0nbBNeVdJEDV3eACIPa4Jhhord+DtMgRABDhlDk5wwBkklwIjHGhZl9arOXdxD
ZtbtWByF1fKwCEfxD0vyzFwtywqE3rWTzfF24Cjy2vSn+yXf01HN0NeNdAhAXPuUh0ppCyts7W/M
dIKrYRkgLKDEGCj045mVuJ2mIINNTWE23hF8FTWpETLfiIlnnsbQX2mY4vIjr6APHKT3CsUq6hvx
aFXBUczcsJdaRvxgL+vXg+cW5ojJvI65D3mxHWCS3AxrljlAFj7eSFr8+wGdMALGis195usjpChs
WY7w44NCUupgdY65QvCcPEsGk6CyeZ5//MGyKpaSS+B3BTyonJ2SYsKLC7YE48rfjnk1t6QxgcoR
t3eA4PjH9xl/ltYdr+LT/zGP1BFY5neuV5lfduxsojXI4vdAooUbkUEWhp+7WCdH+KP0qzmtgOW+
tw7WOPsPdU+RVhHm8EjYJRRqGZf7f7sPpNMCvEBUTgLeHfXo7uxTEQkw3fdJNCsvOZUSEAcyqgqi
z54Nwth2tHTdO4ZlLI0MERTzt6O0C/l6TFZEEJelsiT+1BNjiWVdarFm8Ee3jv/nL9tp6dETLPdI
JJqv8sfO10LzHmSQlHPvF9njqmvABJlHhMmdDImijtrF0QYQMPpe/+8n1GKgbpXDRhnwqA8tH9Yf
XvClA7T000dW9JpQUI7DtFjCtGE0y4M9kDkzQsRerTldCo+MFGnEcMFvpiJD0FvvBJlb0vJRdmFP
Rh+JHhOVrKtO3Zx2knjaUU4t+6bt9ELZwihE/t4wSTKklGPJDli1nbU+Vclyykgk6m1vmUo8299/
vQy1FQ+hrjMpIYydhjCxeQjYLw3UfVV2wBkJ3zHbG9nV3BivbHHvINYpEltuwBuhC0005vD5YpjV
FEjk+TPe/ScLfPxU4Q/szjD2HrLoxIiHmDYOFGnGFZd3uQfBTnw041uAsMC21TvdEbzAFc+a/C2i
goAAuc5TuX/dS3j4prRB7SiwUnwETXfJlNfexg8zj1UlZ8uVPXR6udsY4mqAvMG7LPVzg4/EKrBN
iPn3nvRdKclTs7PzXIWXh4hpA3pCvR3w+FzRSOhperXaddVTsmEEjSviEOHDDbaLxAgyzmKZlJAf
/6DHGEQkX0Pckyt2i1Fun+Yzl8cq/9IkBrFQLW3wegyaTa0wmbqKoNGXEjmwRvvIYqKoeQFQ0635
Uv5L6aA5TKPXOnEIbvtq6owXsBTqoboO4wij2tKFS086YJmrFdmUOlkgNJw+M6fyb3o5NMKX8BSV
Zsk605q3IBLGX6P8Xt0bUNdYxy0JWCuRvkgOjKPjwM2xCN7+jnHWWBMlRDH3z4Ta9Krl22Z4RKqr
m0Q2ZA37bdnrU3GnvX0Y2gY9puRXY79tIl0CtsV3Bm731oC2ThH6Sqq1pEJObQ/Hgfzih7e3JfmU
ffWafu9loyXV1WCqFECKH+ZQ3izT5olbt1rdAocQcJ3J6LNqAbRFe12q1G/29I7k6rtEivRWnh1t
1vH08AU4Jibvhba5fGM8+ImHGIFRlS3xWYOWXS+W96F1VwoOuMftaX4jsgmrnXFn6s3ma93Ahnh5
+1/WV55pwHXqLplvQzPv1GyKL/2qMMm2rUJ1bv/2YOYSxQh0ZF3jxpuIiP+AVh//Z941+rASju2d
AnMMTaOZAYli9VAucTzLQYm9P9Z2dcIns0SvSLdAWJBGWg5AZkmegW65VELerlr5///9hEV0L5cJ
4+vy/gb8QCEyuVx4cGEIzjyJT/be7NUAcjifZ429ikxUHroj58GneyWZf/EmwPrCCmCjUzi+ik+j
baWRu28L6xv/IDzEp/KaU3wpr5ZAV2vwcwWCWVl/vltizDTJXtJgnEtqQdTKkvYLjykEaATOwDGn
xd0DNjk1fyUQHhyEr77YMcajmcLRPJhbSHhCrjdHcsaSnyi+ilTPdJU53JU+PYWnxznOQ+APmAYc
MImai8tLKi/jaoUh1QR7Jn5jRxRCUCT6BG5uGnSLuBEkSHlZOmANZMz8lv5EFUn1vZge4SMLjb3F
E0lnRgxgRPkCa8AxlNVLHljiMdlzypbmnzBWE7LUVP+q8vAp6cQOgNNba2AFswGR9IvYrpjDJh6H
Q9uZQUo4DY2D7KT5NwkkF6VNabhSao+zcl+E4lKqiZ52iV7lDiyYXqhHD4bhDzsuuixU8z71xT7S
U9N4m5dg0fOaOr1+UNo8B40BN26ksuwOmMf5uoKMuOtexzJ6pyL8tg/+y2rhkjzlJqaz8HPbnOYI
ag+0iLvopPG4rqTxDmSiWKJ44rv4VQqiMb1s4VWvXnimVm0aTreywhuLhEmSn+7CKtaEvILmUbfX
KN7lHqiKGOy7tV9n6LqrwL4JcN9kqcB25rJ6qNbQgQsc0eNE44vl5KrAAQKAYKm7Y7p5Er2WmS98
PxCfrWvqKFRXs8SVlfvAVARvg86y6mheHZG6f+1I8HtuK0uhvEaPHGZiSxsL6SJhCLjA1UZDcOXU
LUJn9qAgBVyj3EAfVlaJrZ6xmTMp/eTKyWBiJkr3T8Rt63iCoYNfHaGnOlx39uphBuqTurkmaH9F
iuKw6gV6r15351D9rDAm5V7zvGdJ2TLyc7sjX+EgHufR6Ux7n4xgAGEMG2eAq023Ee8as7npacfW
wJev3FIgspvEre1+BCHSnj1U1iu8lObzy0yi+cwvO3uYtp+zE1+2jpC8jQHCe0ih87Fqio8ANiOz
N6ErO/d4RL9DaRIU4iu0D9KwrqwY072YDvK4VAB0li+G91TSZDAPhFY0iine7QD8cWqZ/5bTy7nB
YeRYEgotpN5+ZEcodJ1A2yn17ZVsQu1SXc2uG+WOHxzcvDEoP0S1UoYczQxXKZb6zc2r7vZs+ZtX
gyo2sbvFO2p/VWSvb6EmhgVMtzCexW7iiblnIhLlllRmKcYA13SnpMVMhN6bios1FGWjCFKUiNeu
eH7iFg9UkRalskfnppI+zlFxg/TL3chZanQkCDohGWBoImKYuBd2/5EDz9/fXDB+xIXgj0bwQ01B
jUk2DCvpskKYj5WtFWUglMqu5830Ya7hxuihrJpBL7VUX9fm+9HbFSQtjzR9hbWe2LVo9YuOq6fa
Ylzwoy+k3hUMg13d8Aqs84pdukpTQ8ANbS2BELf7xO+2fJbKOUX37o8u77nhtQnxGLOEmPIGy5eI
0joBKQBd21/QUiQCa4w84xHgp9R8vj6mMVl8xnP7lC1Uoz6oaR/D5yAHAQcqDlq4aKFrZV6j7eus
mANyMqPBqqjiETQhddmha1tDciNta18HppIk4BQkJfl/MZTpI0xpnvwrc6/GtZ9+to3z5jUDbicP
0cM0CdJngxDBVSY4PiMY7xvoDTzNabln/Dd004gfaawECNACdUTfP/lbAwjybZ8IDrayUeRxyz3U
hSvnMN14EgwNAqplDU18tk3RmayN1g5J1ii0jSQgQYOizUS124Jujh9dcYcShqkzk5u7/Z0c6QmV
/3HCLB+WELfkACPOa2CutVJNVtXql9Tz3LiyMztXlGUGFxHcle+IbrGVfvZVZaUxR7GE85mG+V7L
uCGFMSWcAjz8TsYXXWanr4ga85LdbGJxZ7qz2KcohfPsGCX/DJQeETMyQGeW3PWh7jMO71xQwvDt
NCHGib3eu8EDYUVs/5tIuNnkNSl+UAfPBpH3cg/GwbYIeCpViKiiPGK6HkW847C7GytjbYE7q2Ez
a6aCWaJB5Bg4lDhr4MPAX9yvLzmtzlYxLBkPOvHBgEYCzaunzU9NOhcEiFahrrNI48X4zirvqp2A
c2o7BB6dPYurNVQnsavjRzLuWwkUM7HhF1TXhZzboREeEPUQ60beXGDCC18JJ02katg8V6LpLgOl
i/Ia9K/gylDKiGKbMqNH/9b9Fk/KMC70IdpG9MZTpFAQCHnC6DH3MH1SJEQbsU/d6bgeuBb2tMKe
vNqAiTXzXDiRbddPyQVgrlGLnqNhyp3IJKM5BW42sz044yMC0SEHubEhiI/iAKqyLvVCtH8guFGv
mailw+9c9Y2ITX5YJN1kOm5JDK65h77iCQ82JSvccxLTtKb6Kn8wm7FAMVUbsf3NyPqOyM7WQ/J2
Fu4BnwCheQ0T8QSk94Ka4NK6bMnsqRZ2FsA9raEdLWpNal0D/5SGwOI9eCszWfpZOlCIKXeyNFR8
gJ7SnRXtQDdzXeo16VsUC4u7Xt856cCm+hAWGKFSYiFRB7wqLUydBlKjIteyBbseJnzloxzGy1yC
M/Wecsknt7nSmeNaW9TTOS1S0PoImJjsr97sKKCV60VWh7PrC+jS2cUCwmsQ9dAfKqu+1Abtr8YH
ylJ0+HZw760AoRMzBrz8PjYBDYqDKLrKBWT0Tnc8N+GmDFh3NMarwuAVwO+SD+MjMKwJzy3+zpMo
VQu2CeqaUvVg2M+ss42c9lf6j0UCs21FKyE9CSKJ6dcXSfj2D41JpyjNE3dSON7WC3quBK+oMiV/
ibI26ur7gVBwdACWO6dgGFr1tWWFxRalbG3eeEUEradQZuFb87WKWRLPRQd6GQacP79PEKueexlM
ZnDtlYgfyVysvbQoOmMuj0vwE9sfIM1ktls4XhbBx0exuodspmEz/CzSJdu7FGuMjh8/3YjKgUGb
h/1AlVtPHMESSjF46wYrDeUswl5sKTGi8JBRzlyyDTMBQmDkhriDUbCymvcmN4h+VDNUC497jXXa
ibKe1C/nHm33XWGdBMc=
`pragma protect end_protected
