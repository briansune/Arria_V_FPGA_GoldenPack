// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:28:05 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bEPf/ATPdlIgmlIoZEyled229/UCToj6A290ezsPIyeu72Fm0Df7XrMmX/Gewn6O
N/nw5S5005Uc0lobATivi/9eyoh7I50HLR9UVaf0IT34I8sAz4SZAxUO+afiwHMf
vTMz5uPMbrBFU6WwSa6VLFnUWGxg9J6qcP0uwff6LAw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9664)
bfWs7a87g8DJ1EQnqcidM5T0Nz423YNwI2sbYDGKejMJctfmW8nNOy+ICPySUe7F
pHRS9UjnTc0/4JF3xmi8gU1fYCh9qDYR6a8+fMRx2LjTtOts3E/cNknQUL+nyjJu
JOSJ7XJ5OA05BldXVWT8P/AZuJe9czSCiQUyPYJftqbS7tPFaF5LJ22sW84n9mMu
eI7qVQPWb3jFbd2fvMRcO3SL9dDJnUa8ZY8t1dXYzv87QOuIYkqc3wS7m08UFFay
zfsXk7ML16sXIvmCIdPHScNyiBPayM85ab7wHpFHXvcfGEfBqTE3Qkof/NmYG6vM
Q61RVf3CSoNz0WxOaycXLmorYHpPgH0vDslBWZ0focWBSN8Zl3KrXNM0CgO8azka
hPf8B9p98QM6UcenD3oNQsBn7sj+rfFuY8LcZBAsx5KK0Cp/0hyjYb0fIHx5MrAV
AYiXFuZCL/Vv0hWqehBI+iCEt019VCFv+iupudavXW0Yod9st6JB/NPINgG3kdl2
zo1t8DN23/PJ51bcCPuVY3zI/5K1um4YWQa/ek8pni/lUf06xJz1BoRA+tJxs4kN
jcjGfw0ltN2mIOLA+jI3xqsWN9Is77vjGL0WXuMkdp6DUJRttdmz26v0GPWIkpT8
c4x5Y+F5Q1WR7RTNjRLF3h9zFazcuo2l+OU50JmTkKFqBo7G4hA3tDFsqZT63GmO
lb9Ui7w7syrekuMjXRkZ35+ABsHEu14lyKpwCWhi1Ry9m3OWq+vi115Bxk+TFw+Y
jIm7tVehRUUkUwxroDzSpAF0/oHsXsMpyMX3Ae/aqlp766Bl+HSrb0Dw+o0My8M2
vwkPsIEvzwxl55WkDCIQFZMWXqZLbV/+Sse34dOfAXHZbv/hLPM1uXdPlZPPh+K7
C8uL7Pm26G2xy5WUqMvOuNuPLYFU/H5Hgo0+R1aTzCZh3DNEBRnTE7R8USdANWen
ABl/gY5geAUZyViz5n5bXU41owucajXOkhcviGcHdO8ZR4EBGN7dKMaJOLDe0m++
VajZVRkqhkRdMf7Y2Q8WA3HCtaKXUMWsoMenp4xLdL3OEgXVwADZkSA2otYCrwKb
c7a2o4c9VhebAFbSsrkiZXp7BwDz8J0xvV6FSnc3DrxVVow04f/SyaMjUNxr7XpT
8lTtrj3ItFcWXD/kppqL3VEQcKuCB7Z6/BOz52BcwLqUVkM9zI3sDDtm+jPTOa7E
uMUps+RKYQ5bgMQYYSm/iB6TxEXOdpbw71hKeOYthd0eABIotT7fuxVKVNErNEJH
A3NZOdHsTNk08xnOZMQH4pquqMv26O+dQVUQIwBJ6ZLFuwz1bFdod/uVRYyO/Qdr
XT6eCq1a9BWilyHvAdHqlMrlmgpkmARhY9g/FApV5DSy06xSOE6W5baD86sm5WjB
1xLXbEnq/bT/ZjL2Jv0JQA1ksaA+iYVGvEKI9mc43nH779ZtAfFfZSTsIgPz+Z8b
bwUQSY93W8i1YWQ2vLWCOi1t/QtHHr7l89f5oGbo9oyJ5Lww+Sv6u2zGs+XUKgBd
8jdLOH+7oa190Hb/4RJTUPhJpVR3qQWENO5SuGZE3AiTQh5odx8nTiyQEnb0LgAn
/zjocli2lBvjeMMY7WWqT7lhIsAk8MAu1BP/IjZ7BbrYnCXL7z19lGpysAQS+ejF
5JvIOHC0F0YnwzUxDpWp54bnI7SFifr2SZ0QzGUdajWCJP2FKb0q9XDYl4w5EXEb
38qDNnNPirsHwwteq7N1hL3P+I9ZDi6J1+HusqbgWB6AZOEZ3jqfFzoMUF6PmjDf
YEH32c7yxx1X4+GQ8kel23t0F3qT7Q+3sZWGn6tpBVCDC1vnKFhEUtIrrK56KCBW
8mNchUHQbJODBMFC4u/sty7VV0NSqhtx3K0cjje3kDzDHDA/bDbycbrVTqLM8grK
sxOzT/Z8gdXGAeHB+FKKj8R0Ff2c6CA6VCSQYwrR3gpzqEQAzS/8y0vvQm6Pjb+R
5eSqmA9c35PD8sTbHiC+rcxi4fCvjyBnqT4c9n1NcAQYrihwAhlU/2DRJanlL7C8
VYJVWFgjAq0wJeM7uI2A0y7EBUW5yaH8w/ev6XYtWwL7K9xk20ZHDl+a6tTb4tcw
x7WXwlArDq3C0Y7Z7qC9AqVqllB+peWn2G4aBIfDKyTYpMHx2TvbW1HPOImsxisv
j2ba8/VwrC4SRsa0aNckCUOSGPJjyjV2qfu8vZPKTo8iEfMC+5kZOdII3I8TeHf7
gCT40PNg7VImm8xsPQ7dEBYntOW8Besna0YfxjDmHkW0ljpj5Hx0p3Q5Wyek8/pG
0tdxUNcv5O5vVRcbe44qlhab/F1L4X2jDXhKx6k2VvInQGXxGup8bPhyTk/SCVKp
1NHsvyPHg0WKh45EXH+WLXY+L5u3YPTKejfPtLBISiIIlDjvTQGdME2SntTDsQ2l
su+IVN7PfGX2m1hfD2p2eCPa2fzwqT/KjQbbDSGmE28zO7mvEnwE02JErw9FlRzo
CFPGzd9qPJWIl5pbUZ0PvwlYgtyBlt5uTNII4POgm6AXSYHqxK/IsdlPXZ02amgc
gw/LPrJmNF3k7FvuA7BLTzz6YfeEQWkmDLCzuww1DQEoFIZnMXxT7dfBiVvFYyKA
/IEct0ovHuq9i8REIDJo/jixLlAAGk4kvnkjxkh24cP/iBsmmJPggDOMV4YbtuYD
bHfVOzkbE8wvdAhysl6j/VGIE5H9eIRF7Ml/Z8/vjx3JCkpzao/o+OjnWISWspcu
E2+JGhPtw/WlAYxG+QizUSUTnywvpV/crWdmrhj6VULUFbpSTurODnbiUVe70UiM
YcZKVZJOebNX/XwHfLGK613g9Qy/p7RDVuiGChvxq8Nin6fvbhEpSwKhPZ/joElL
Smv2Tr2YxbY/10i982DZppGboqsDSpo6BEq7nKmLj4ienF+u2N3i+k66Rlt+Rnzs
eUyJ5B13ziQ5BUghgLdZep1v/b7zDKy/sLuinEu79kGeJHFT6nj/dOHi33HtBsQF
xj3T8khR98SxAx+FAdw5PUYyreM20cAIDSbvYte3ePrn0vygouB2hja8Ggq6LmRa
BhHEmgOjbkU673gUaHulaUpA+A4acACFygVlmefbaI/8rhykYCvld4zXwKgy/cJH
SjI/cZZyIG0KWi8j3GvaagVic+b8pfFQi2EyjEYzNGqplenjlejMT1FbitMF4Ncx
376Rve/KRo1ofBYvwN7doH3S56xOkd+BO+EFLJu9OvhOdqfKamwQMtlUATNXABjR
R2xV1UIdjaYhgFto9BJSKDqfnlc0AIjrKXh7Np84luhmOIIX/cs6iwMZFHieyuhv
3YTKGK0bS9Gu5KswkbE3Gh5qMElW9cBF+shliCnnwAWncL3cJ8oBp0Qf9s7RcOol
98MGCwU+sX9JG43mt9w1CSRmKKX2ByUG1bMppKKP0iRXFKaSCoBnekV2dZBEODWd
d25bq0NMc4E0+SaKAaLObxZX+FQhZrkx4Bfy/t9FLMru3bgdVM44oLug+I3oPN+k
QjlEXz0/vqO4yzYccLA+iREqUzVqBXR/ndJB1K33FZYG3jYwFu+2xBjvfdzEx85s
CTMfBONJunW8Pswycmwgam7DtiIpT2YXnZnMJPczEG7stdcoe8H7sSXFeGlp/QlW
Fle9DNejeA226wLaGzy49MmmIYdvupJLnt8OyRQ5wlfvxkrrpq5pKvYpzSvLUz9C
QHbailDaVUokn2/WXVsmToUgmImcSe3iJ/N7GG7lOVjByP28T0BiRC3edzV+GiHo
dZcLLPNSvZBa6La7FbOu74sMGWNUFuwwz6fcLoMwgE1+5dHB5B3DcCDrdksG9tWa
YjAiB/OHGtGGROhvjCsB0LIW5xpGyeF/y0B1VS+qW3ZvGD9QAjTmrNyh89bTMTLB
51YF21+zf3AUtnM0LhwLdFCOXFplD7SaKuuHXZAEUJ2Db9ftaLc1xzd07kK9Q5wM
r+ulx/91cVnblRfVz+LIrvK5uSdEWyNa5jp4b9CiBz2hF7lLfZ2FqlUWV4KmXsLQ
rRS1t7jY3i9YkK7tTbLRN/v022E2UkwjZqEM/rhWonOPdqsLyfABNtUrlWLsd/zh
pbyVP7cVs621HfspAi3rCd0YfRI6Tfzh6l3vjlC7Lg9QlKwD+KIBVMqMwgSVLZOg
bDtuIee+iFTDIqDdkVAUVKTgxC8gCkDj4YTjOgHcEZcK4O2/nVq9laDI44tS58KQ
SSiJtniniPt/aT7Fy/gCEFZW+gD7JWEKPHT4nQMk7jte5rJswYvfhXl9+8AtvuYf
4F77sD75o19dhg75cRLFKyzI9zYX2lgNF+0YfHveinLhTXQxqwLElFnulbqxATBt
oiiQRn13bMzc2/JmrXDpwvg0un6lGc4ZeinYQnt58DdfGUQxEZBaSSUPfZ5pgksk
HWc0HI/SxTKprBpX7E+XzU0s+2mKRZ1A6VKQkVWWmtnaSbE9sWjuw46agluQTnbb
BEdaKMw2Mq5k1fW4+le4OAebGXSLNhIyQDWNPSCNiBdG2nncvKLiheDPF02dfZL+
hzaWJyEq149zL6ZjuMnxCV3AGKe/phNo9F8ce/GEhj8Bw1oCguNFLsxXOUIxAhhT
z/Xn1hfhvdPjIocXtAYgJ2QmGFg79kaUNasDwSdBCQ25821CzUzzcs68VpUHoJqV
tB/sbOwozo7IQJ1kddIkqVRwtoQ0OPLMztm6+SLYDWlQrYdjDz0iJ+IiJp4y2sM6
hkC6okcEBFVtLcwwOT5/ZAkqKdpCsQqxEEBCHZ/Lbs67XDKggMzluHxh6NMrcMwW
rSqLaiRoZLYdTtYemYQpjVc185Yuo2itngDZ7ZIJk1SS7KOks4BavXkMKz6YdEv+
TqOM5dlivJO+5anlv2OPnrPA0SZyF3bqcF2zvDft0FakUxvX6TA0xQhbnXV35YkB
rN2rT3h3I+6enpC3NaaFvN6juTPkrYmPDnN+qXGdaXc0sN6ryaDUIOcgAQspfD7B
z61H6H63YtF/0hKkYSrLxyilgfr0r5X4mB1lXyXZEvdeOi7vV1hG9SFjudrHDkHI
X/xNQnFjfNuYnW82WDVDKb2O6klzJ4IlLj4OyRkyKJSVGCCkbh7/TDwMb1DFzg1Y
H2Oga4lAnwHgB1/Xa0yD+ctirV1I3JJRrdVjilV6kTDHxcmzg4qtUFgiDESspZ1N
a9blFnGidZQnzLeYB3X04eii14B7lymTeP0KeXPEMtoqo+wShj4V7558g0YDJ5Ut
ji1t4/B6N0nLVvSHcGfo7Yp+6PLZmmjxDQC665C7cEPJjo+gsZEXTJOqmhPqJM//
jObVUE0gb2x1dvkBIKeVAdw31BpmlJL+K0R6+2fJTvQe1XOMeidfit55o7KLpqLS
x8jgZ3KbmON4NByZas0Y8FZvz3rdRKlJioDuN7S94GlJWN4KBaAJS34BtezjyUvQ
o015YaClnS2tKPQuEMA5Bc2tW1CzL1rw4MEoZp4Hdj5C//qQzVXenfjFHXox88gG
qnjPE/JCQLNScasIOF6hXnbqvEtwj6HYKkhCJ3ij489UXmZoERTULcp8wXyL9rNE
+4peqdwibEE2qkFbhBI/7W9rk4jDALF6kWt/geS+oo3wh8as6CUj739E62yPTGGa
I6DeOQwx0MT55F/Op69NDey7R7IQlf36x3yBTfaE5p2DoSh/mIRX3RFKObxS9KYI
g34vPnqqYlruvrQCUtEOd2kA1U31UtTxXxwPrzY5Xyp5mSjLSqbY6YJycp+hayU/
zAtgV5+hQwEQ5tBOy7LRarvfgHLwhdsG+AG5umTN2JCefsC6qoa+2WxVcvRtahQ7
7UCU0S+zN7GVJUiZrgdn7dr7RgYLrkLopesIHBHimONSClt+wdnnTh4znr5KNFNB
01XLmsYGk9zBf2MpW7YducGzCb3ZTmAQDeFtkmjNX/VcDPHeW77dvXKXeGQvJ/tI
yF1a7jJfrBkP25VaPnNh/cFPaFz5faGms/f9xN/ROpAdEi5cfbVD7PBmzsIflW/h
Ry9cgQ9nK8eT7ZQlJ6Qm3cxKnJAtnGGtSeOVYzei97L+yB3Vb9Vwnjq8mNPAuwS4
0nU2Fh/HAyu/TuSSQDKfsD87ONrUODvOwsyNytg/gujAQ8xg1yD/5Guv5/I1/dJI
dJY8iNHOYWszoV8wKK7cVc2rWVDm2Qr1ZPCbSg0TXSbEujMdaH9RzQkkQFGHd0mk
KjfJqkppARsN53gubaoTIf55i+M20DALcvpz3aqwrKxaC6UVvv0MDc/0cRhB+j/Q
IA5Ui4D7IKR97IRbZP1pENgkMfuhEm8QKf3F7cOS7xAIWgukpUW9cOxBDvnbrdOL
KyoPP0rHdLrbxJ7W15eq5Ar9M9LZeTsczT+GLIGnEXaCDR9J+ZzPXloB++NeDmjG
DDMFdaJosZksSBUfk2m0w8ZpMxwMT+cdKn5fMTOhZbMCdaiLGUHCPFRA2IdsP/3I
jydIVYUDB6StofkboM3b+T9lzZIJz1sb6gYPGlQlFX94o7VWvXwGb7JJXyf/Ehik
6jdTuP8KTRbmk+HNUbPT+MQMpz25Cb7h6Dre5GfPGYSyHraYOogRm4ElteCw9ogp
NUA0FIr4R39gvgp669HxkeupWx2kuyg80/xqYgCAGfoqWzwunMguHt4ECkXLmThL
KSviCihtbfLPmtc/lGT1GEs3gPgyaCm1xQ1cKYKYvbYFhX7jfJez8uDn6VSjDFst
mdbR29W0w5DhAxICxW3Wjh8GrjjE8yyH7pOUlsvQeyMZYry7ZATgfuJGhRcr8cSo
AV/SJw4mlEfRym7ODZOCbjqmnpipnSj300Qbh2/gB4LxT6DSL1aNJKbF3BYuIGWE
C0+hvmLO8D9is9eCwBFUE1XL7Byq94/YegaN2tBY2jfr1zg++Lecs2oJFKP4VAXP
Vh/pXyQRcBSJB1VYfdQz03JffkWHrQSOE+1gXJSeTv7Bma57E76dS0IbcB98RR1W
xKaSpWUFwqfIe/H1YtablL/0WRmhTTlj5zOSNpoeJltGq7mthp8nOfhWvFNkJKOr
B80+yWK840u1a4hyf5DqeMrVB3WWj+1YF+fKMNbTeOXbHQRWoflwvLvb0fyDuaLo
GBRIHZsrO7uGTiNTJEPcNO+Zrr+PR/KjItfEuAMmE1tuRMkIagXh79Sk+ILp2COR
giV/LpvSHT2TubwtGD8I6euIBSJoS8jzwWgTr2SF8UPTqPwSQTgdUKhADM+jLtzn
UQAQKUZzMMt1xb65wZkCQjwYaRYj8SCXfkKCkSzbouFI/r6jo0lL218WStMA1sj7
2FoVJ96XgcfblhWVrxLHQOl+0o8wytEChLEK+AhmJxR8OY5Ct9Cc5fmqWveRWFDm
Fc8Tsz1E9HdQlFAI5z5ZacE/OkkUSuvheFeajeBBQ+y9pSAaiOZsLWVDwzP5pXRa
ExxpOwb8HWETAQNgxqyq02XZcdYCLtcEcXekba1RyPxN28pKwQgeNzsaG3Ew7+Ib
rZQQN2oA93PGCfpzPs184uh3BattjolslhO0jeKKpInAb+jUGJUjA8EYSesFjW3e
B5hBF3kW3qurG08KCv7t/GLXRBIzMvZvm4RhA2EfPp2Tbgd+XPv9MDN/buM2Z2Nv
3hOvURTxIfRGNjYmzreA4qhl+wd3B0OiJsOZFH7KIuy6tJQQHPVea1xqZu0+X8Fp
RJMVBGyl79DfgRwWExW2V4b36HYgwjxaRaYVDM7SVS0zKZOFjRzh1kowaFjn+XbN
Fqtx3V2zPyxk1Ans9FmSxQ3XcyUt0IXb2QiFTufiYDfYvNcg6aa7kMK5ZUf8oGkP
ck+8tWI0vrR3JQP7ILe4qJ38gygSy1+tIiZyYuC9PL6Ch5FNW9suc5LiLXC4/us9
9loA10K2bR8Wl4RpDJeQz7ChQgWLHRMYaf5CpVXJd11NMdNVoL/MJ4OXEpFP3QW9
N54uUfB0b7OkNjZ2GTAaFMOSRaQVEMVsSM3kQd8cXx1lqxrGVrUF5eSYAZu2uRGY
0iEDERiFC3K+8zpf8o/NLYXvX0AqoVZq901W9rHwq8gaqpCWynT52IYMfdce/Wnj
hpCTa7tQ9VaA/K4TdevcZECeymxwA0oCDO/JS4AoTtHhalSNIEkZ3rca+aXY7Hxz
kt8LJphKZpJ6ydnBO1wHGh7pRiJDiqnYNpvcZEr3oGaYHRtWOoQn5GW8BAAMsZo6
lNqmtMCxDpBLHGhAgYQI6710K55AqnjaWD3WDMwM5sf2rmfotM5EkFTT0/FFbI1J
fjSlc+cw5Ii7K7Zq4PqAYnVUQkbZEGT5Fu3KwcLqTgZWI5n3KYD7Y2um+VLUziBA
+XZDNMLlbzYxHgMijK1tVEHqDpsE08hWc95n4DeSWOABbM8WJg6WogLAqTqjzscl
SK3fum2S2zVPSnrXXQ6/i2sNiPPDjb7bXy4UnG2lrxU16h34G1W91wK2dttPTbcV
j46kBn4GU2IWiLKB/X6KpcIWh98Zqzlb/e5KDtPU/fnYgQc9DvEGOwVoNgvfJdYy
kZFKw9Zt64OLTS+ktuzI/JAk5bUIT/Pj42n48/JlVMtgfyGJvM+Dd+G+P0DbOP7t
jT2nkhOZRF6mGnZvTagA6mszWVkgI92kiei5brbBS1hC7hyZ3Zblu6GDucWuilVQ
QXD5TyhBQ3LO5bVRjPE0v1PCso3ejgr2r8jn9BSFiOoRsYKxwkXs+nsQa+3I6xEh
Y/iAzM4XCo62Sw8hM3bTD0gy+oBCh7DcF5fpTWb3z3WGtcDrTlQE9jkNvG0+7oKH
5S9ve4zhJMPfHYG+e5A5Q/nVgv2jMhw+FQz9aUeoY2tKIhJDFTohERv05JKJ/KwH
UPgqcqR+uFZQqQrugFvUh8NwLu5T9vqW983qL73cj0HEDvsxn/sA8lj9VyIrHHyv
sPaNsHgSPr08LTHuRhpP1jidnLxJSPnS1C0BeFnqpXXnhAcNY/jB9FY/xta3avFb
Gnr+Oiy1N3NbCm4+xb5aVcc8ApaJUiAy6um8qjzANsJTeNqn1oz9nzySGuaZrXO+
XVxfJm1Pn/QI3GELVXGbiaJir4Vhuri2qdzlwT9DTI0k4TRztnTxJrSt505yfmIB
M5BhIgJB4513Y6yhMlGrELo1EckNynXIoSrcSkarIYs3iAK+0cBHAvAqXLBz59NB
h3uW0mRz3OEuo75Q5vk4n0lqCMBi2D4RSD1VZSE9eokAOcs54sDfiNhkbJrBNOl0
EaEDEouKKyfI1hiPVw6ztdJmeuGcwXOuh4GWEu7YaqXzFmVIU5baO8Rtotsdtaj5
YlCAM7Bf7c5RA/zhFN6orG37flWV7WLdoHYH6kVlTTBnN/l865Iw4f8T/G4gsa/E
2ZyuUcp4HZABgEU/aSt9NhL9pJqrORu2C2n2PGTSvVgZdEeYVE3QGJWgJeUMDQwX
hPFDfz0F1KAfyGshgY8XocPmilVFzvKrG5J7gAFX2nzNEPDnLygUzlmNI2kKjKDC
8o5M5KKKwNViR/Pb39pUTewfmjA6ElNYVqAfJXdcZJ9QvM1QvR3ebVaH+XyXfQsY
qO0cb1YiNDdpi3soVQheZYqn602rhNlxYeBdaOZZkc52TuZCSLZiIF1zx2MnhFr+
zuvAlX5r0noXAqMb2qR2UJzVuBsWKX3IygpdW9TDXWFLwBQ3QDaeYB45yO23Am7s
cbAGzlIMMsFfLlo9clg98B7VfzIuTd1/H0PMXZTSgYlRmC8KTHEaLcsrynQcEM2f
OGzHQxiZvCJPpUniqXHvZonPz9KQ8ZAO0Fd8dFX7IAl+MZethL7GNPECWaa2+po7
kd72fzasIjOQdQS/nkFV366oFBlpI3xyeKizioiaA6QTHbAD91nvswdSOYHTk+HR
C1b5dqkS0UWNv/LehZwLed3TM6LfGDqtMR2yHioKuUz+Xgao3vmS4Tg2xTBNUkEQ
QZH5PJhf5FoxqE61QNwBRA0iEEozWXHjUiBi20yClqgczaJbdlTEO4cHi8OnBHcH
aZAO27gD91W1D3RD7OJ5LUHlL8opkOUHGHrFasQxQ01xdDFjecYG8R3DX1BxlT3k
rZzd2mkM/Br3j4KE2+aI0dQQtKzI+2BZhTzsNa2cs3mfO0Jxy4qtPl27oDHqFFuw
ILFVSQPoEIJAukTfjZxoG+3RQRY4Vs4VNmA6zWJpBEd3Vgr228S70usQsXZraNEW
xcvYEwIGhi/AHKSSW9uzjViDv+Lldk6SQm7QYQP+TnYFEGV7TT22QKgmGW6xrZI9
cWCRMO7Gv1g0WZRw02oqFqoSlRJnqE1uTGLQrf3FzuZoCJtfbmQgNgl+7LXce6mq
S9dxw7WzWQsLUESIQGH2ZM3/2KSTOoorkcpGEConnQESny2P0plhLAg+Pl6dAEfu
qzyMCK38tOpmNMgw83ybSU3pvbdxAdo0h3xV+qz6EK5T0urbbByvLagVd9C7aF7B
Xwvb805HfLWIi0dAU3irXVSZPLHkRpVw75O7fjV7jVQJy6gEXP4oBN0SzihTA8Hb
dTzHunnVjB0rHZaoPWjXhLy3+dSeJkjXTZgh32eyfHIufkSkIzNHIK2f9STlLl7k
sAaI+jyKk0E81a2lz70J+oObroFQTZmVD6VJq/3jR85BwG/Iwaju6fKd6daXejGY
adRL19JNWMeAX5s/0AhGlVXEVS+8MO7khEN//vupccEWOxkHREDyE5WPiyQOi+Jm
wfi3hTw+zOy08vZggwhaNucz5/vX7ngFcQsNiQ1PEqDvEd8k8iSlrEV+0p075jBV
nsWYlYvy3bjX9SQwwnI4dgR6wsMhxZdTpz3vrfKjWYsdC8+7Nbk4JbcOzMQIK4y9
zs1ItA7UFYQPA0HSjNYPt2AbNwNvCHbGF0UhaXWc5yQit5BiKcelu2Qh4XMwINc4
NBQ4eRb5iMgJwEXFfxG/CWlqTZpYlbLN8J6cdfS2wYv+o7zhA9oazv6VVlXZEJrc
xbK6py98sgr0OsykSM+l61Q5H1g2dIiDxdVn0tGtoP+h8HklxtgO26k4kEo0+5rN
NOJSkoC/mLDiHxmUeAc/bxfn+b4Fu7XO9yJjP77UD80Mpuf7RII7/GurnqiETcAp
CMz+w2lkSweZPYWLj5uxplAIHAp6HLX86NDQ3S2cNN8ZD4fcsiZqnBiKTlhcCJBp
HVklAfTa3kKgbAtlfk7naESZtbjWl/GBVlZndal1DxudMZYsH43M2+ecjgLQmcpu
6+l5o5vulk4KmBkMTFPqjz3IbE15Ghi0jO4AXfu4m6rZqgx7/VKPvW7vyjRtjC0z
RarCBkKc0Qs3D515/nUS472P80HxrXAcdXF4cPTX1blxN6JFzyXKTj5nhYd5shxb
IWyNYl8N3q9ZQ1G/Ti96w/PLyzh6rHi5luqeUR06C60uhGo2CuWIJfs1yVH6TFeT
FGTKvKB3EbsQObk9Ck6MTYAPIilF08a3MbTSar0AW1RPPTYVaNarAYFB+qFmUuRh
X1kIkfifIbfPbm2uGlG2y32vSYhvYfZ8uBqUIzmEUC2y0bBN54oQZ99pB1qByNON
Z+3YiwJsAae8ciSBmPwAU09k8Nd4Aw3kZWBIVgFjZRQK6kPZi4f0T5xJ8ZIxEakk
BSZroLVWZL9CZjDfivvrLfmHOYldNADcQr3kFNXIJeQZGfe+tYmrMO8T7GjcMxx/
k9JPmhZio/6uGg4iZL91LbCtikG7bBsqhggmhnaA5pFf/yMNZv9OC/p/tp63n/Or
6EAIWw1D4UwUx/+9PidvI7j8lB83M9PK/cEX1xcp6zug0QtcBNayOL0PsdME9Ofr
L3cTFo1QuU8xo+g37CHKgtNArVkv1QJAK+/a5v+hPDeodCATFb/NqwFyj86dLP8m
f0gITlMUzNbL/ZlxbrvfjQzmIL1jEHP4baTyDRCnn7iXTrx27y6bMxabcWxw6TI+
F9zCj0D/6Vs4p5gMA07LWhcNGOde4tslAgFxNpaB+8Gmf9QNUOtCX1yAGLgIxFhe
KEFbg0JWcsqtiA4E8rYdWdTIr1wo3JzUeF6fwMGaxTtHtBOQIfQCRNfw0va1GQEy
OPl+uSkVGrP9wxdjgDwLBNHYJc9NVjVCiQ7prDE849zLJdslKh0lL30e8fneRV/4
MDIofHspUxIgi1gPRDY7F6MBlnfK5uUcumTrf+J9DqfL4LC4WL52XEHur6oNvCHj
RNasUMAVjQwED/mHwDIz5cay0Cca0d2ht4zk5d5kOfjb+ILTyps/TDgXXoaSEOPB
7S0qYPted5aL/CjeR28bcBfQQ6D4h5mxiLcNlgmzogMygIm0EPzFI1uOreZzKbOh
q5XcV2ly5b/2bAw9cynEiKEVfS6ERLlgtz2NWnltwRHyx8Riw+2tVv/RMX+LqDjo
jPapu/7NgGQANZGqx+CnNUrKegIy/fU2i4smYC6X7L9/6gRj0LpSKxyreOA5dCSr
mUYIoCgmZ5ujHip7WSD/SROnHg8iW55q0CnfAd/hGwhlGXvNAvSmPhfoyCqFnl6G
UFmNhVtBhh2/HcseQyHxbkjTTKcEc4OixQqDjkke+JQAQRf3bFf36HzH8jFkM3VK
Y4viOiy0IF2KiZ3XzwJI+hXAhVpjimIEzexU/o05Z9qk1gHMIosXvUvA4hSw9YAY
dClXQDlKdbKgBnzBDumXqETUe4Galvz8K3MnbyS2BiebQNDquPtyKUMo17pOBTWx
prxXCtDhZSYeJeaEyfS/jTOU/Pd3msIRIO/8YVbpSp+dVGS5BDfAs/0Gp+2hWZZa
Ecye5tDr+LWoDjDygAJIDoY355t3TjhWzKkyLFeHIzJ3Cu1qJZr+L0I01g6EtejO
Dl7fAg8M2idGJhymEuSolgtCLtx0QCs27BsIAe20y45kUY53H9Hy3YhN6mGkW5DC
RVO6CGuGLEA2q2iM65Zxnw==
`pragma protect end_protected
