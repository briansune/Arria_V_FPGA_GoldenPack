// top.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module top (
		input  wire        clk_clk,                       //            clk.clk
		input  wire [31:0] dut_hip_ctrl_test_in,          //   dut_hip_ctrl.test_in
		input  wire        dut_hip_ctrl_simu_mode_pipe,   //               .simu_mode_pipe
		input  wire        dut_hip_pipe_sim_pipe_pclk_in, //   dut_hip_pipe.sim_pipe_pclk_in
		output wire [1:0]  dut_hip_pipe_sim_pipe_rate,    //               .sim_pipe_rate
		output wire [4:0]  dut_hip_pipe_sim_ltssmstate,   //               .sim_ltssmstate
		output wire [2:0]  dut_hip_pipe_eidleinfersel0,   //               .eidleinfersel0
		output wire [2:0]  dut_hip_pipe_eidleinfersel1,   //               .eidleinfersel1
		output wire [2:0]  dut_hip_pipe_eidleinfersel2,   //               .eidleinfersel2
		output wire [2:0]  dut_hip_pipe_eidleinfersel3,   //               .eidleinfersel3
		output wire [1:0]  dut_hip_pipe_powerdown0,       //               .powerdown0
		output wire [1:0]  dut_hip_pipe_powerdown1,       //               .powerdown1
		output wire [1:0]  dut_hip_pipe_powerdown2,       //               .powerdown2
		output wire [1:0]  dut_hip_pipe_powerdown3,       //               .powerdown3
		output wire        dut_hip_pipe_rxpolarity0,      //               .rxpolarity0
		output wire        dut_hip_pipe_rxpolarity1,      //               .rxpolarity1
		output wire        dut_hip_pipe_rxpolarity2,      //               .rxpolarity2
		output wire        dut_hip_pipe_rxpolarity3,      //               .rxpolarity3
		output wire        dut_hip_pipe_txcompl0,         //               .txcompl0
		output wire        dut_hip_pipe_txcompl1,         //               .txcompl1
		output wire        dut_hip_pipe_txcompl2,         //               .txcompl2
		output wire        dut_hip_pipe_txcompl3,         //               .txcompl3
		output wire [7:0]  dut_hip_pipe_txdata0,          //               .txdata0
		output wire [7:0]  dut_hip_pipe_txdata1,          //               .txdata1
		output wire [7:0]  dut_hip_pipe_txdata2,          //               .txdata2
		output wire [7:0]  dut_hip_pipe_txdata3,          //               .txdata3
		output wire        dut_hip_pipe_txdatak0,         //               .txdatak0
		output wire        dut_hip_pipe_txdatak1,         //               .txdatak1
		output wire        dut_hip_pipe_txdatak2,         //               .txdatak2
		output wire        dut_hip_pipe_txdatak3,         //               .txdatak3
		output wire        dut_hip_pipe_txdetectrx0,      //               .txdetectrx0
		output wire        dut_hip_pipe_txdetectrx1,      //               .txdetectrx1
		output wire        dut_hip_pipe_txdetectrx2,      //               .txdetectrx2
		output wire        dut_hip_pipe_txdetectrx3,      //               .txdetectrx3
		output wire        dut_hip_pipe_txelecidle0,      //               .txelecidle0
		output wire        dut_hip_pipe_txelecidle1,      //               .txelecidle1
		output wire        dut_hip_pipe_txelecidle2,      //               .txelecidle2
		output wire        dut_hip_pipe_txelecidle3,      //               .txelecidle3
		output wire        dut_hip_pipe_txswing0,         //               .txswing0
		output wire        dut_hip_pipe_txswing1,         //               .txswing1
		output wire        dut_hip_pipe_txswing2,         //               .txswing2
		output wire        dut_hip_pipe_txswing3,         //               .txswing3
		output wire [2:0]  dut_hip_pipe_txmargin0,        //               .txmargin0
		output wire [2:0]  dut_hip_pipe_txmargin1,        //               .txmargin1
		output wire [2:0]  dut_hip_pipe_txmargin2,        //               .txmargin2
		output wire [2:0]  dut_hip_pipe_txmargin3,        //               .txmargin3
		output wire        dut_hip_pipe_txdeemph0,        //               .txdeemph0
		output wire        dut_hip_pipe_txdeemph1,        //               .txdeemph1
		output wire        dut_hip_pipe_txdeemph2,        //               .txdeemph2
		output wire        dut_hip_pipe_txdeemph3,        //               .txdeemph3
		input  wire        dut_hip_pipe_phystatus0,       //               .phystatus0
		input  wire        dut_hip_pipe_phystatus1,       //               .phystatus1
		input  wire        dut_hip_pipe_phystatus2,       //               .phystatus2
		input  wire        dut_hip_pipe_phystatus3,       //               .phystatus3
		input  wire [7:0]  dut_hip_pipe_rxdata0,          //               .rxdata0
		input  wire [7:0]  dut_hip_pipe_rxdata1,          //               .rxdata1
		input  wire [7:0]  dut_hip_pipe_rxdata2,          //               .rxdata2
		input  wire [7:0]  dut_hip_pipe_rxdata3,          //               .rxdata3
		input  wire        dut_hip_pipe_rxdatak0,         //               .rxdatak0
		input  wire        dut_hip_pipe_rxdatak1,         //               .rxdatak1
		input  wire        dut_hip_pipe_rxdatak2,         //               .rxdatak2
		input  wire        dut_hip_pipe_rxdatak3,         //               .rxdatak3
		input  wire        dut_hip_pipe_rxelecidle0,      //               .rxelecidle0
		input  wire        dut_hip_pipe_rxelecidle1,      //               .rxelecidle1
		input  wire        dut_hip_pipe_rxelecidle2,      //               .rxelecidle2
		input  wire        dut_hip_pipe_rxelecidle3,      //               .rxelecidle3
		input  wire [2:0]  dut_hip_pipe_rxstatus0,        //               .rxstatus0
		input  wire [2:0]  dut_hip_pipe_rxstatus1,        //               .rxstatus1
		input  wire [2:0]  dut_hip_pipe_rxstatus2,        //               .rxstatus2
		input  wire [2:0]  dut_hip_pipe_rxstatus3,        //               .rxstatus3
		input  wire        dut_hip_pipe_rxvalid0,         //               .rxvalid0
		input  wire        dut_hip_pipe_rxvalid1,         //               .rxvalid1
		input  wire        dut_hip_pipe_rxvalid2,         //               .rxvalid2
		input  wire        dut_hip_pipe_rxvalid3,         //               .rxvalid3
		input  wire        dut_hip_serial_rx_in0,         // dut_hip_serial.rx_in0
		input  wire        dut_hip_serial_rx_in1,         //               .rx_in1
		input  wire        dut_hip_serial_rx_in2,         //               .rx_in2
		input  wire        dut_hip_serial_rx_in3,         //               .rx_in3
		output wire        dut_hip_serial_tx_out0,        //               .tx_out0
		output wire        dut_hip_serial_tx_out1,        //               .tx_out1
		output wire        dut_hip_serial_tx_out2,        //               .tx_out2
		output wire        dut_hip_serial_tx_out3,        //               .tx_out3
		input  wire        dut_npor_npor,                 //       dut_npor.npor
		input  wire        dut_npor_pin_perst,            //               .pin_perst
		input  wire        dut_refclk_clk,                //     dut_refclk.clk
		output wire        pld_clk_clk,                   //        pld_clk.clk
		input  wire        reset_reset_n,                 //          reset.reset_n
		output wire        status_hip_derr_cor_ext_rcv,   //     status_hip.derr_cor_ext_rcv
		output wire        status_hip_derr_cor_ext_rpl,   //               .derr_cor_ext_rpl
		output wire        status_hip_derr_rpl,           //               .derr_rpl
		output wire        status_hip_dlup_exit,          //               .dlup_exit
		output wire        status_hip_ev128ns,            //               .ev128ns
		output wire        status_hip_ev1us,              //               .ev1us
		output wire        status_hip_hotrst_exit,        //               .hotrst_exit
		output wire [3:0]  status_hip_int_status,         //               .int_status
		output wire        status_hip_l2_exit,            //               .l2_exit
		output wire [3:0]  status_hip_lane_act,           //               .lane_act
		output wire [4:0]  status_hip_ltssmstate,         //               .ltssmstate
		output wire [7:0]  status_hip_ko_cpl_spc_header,  //               .ko_cpl_spc_header
		output wire [11:0] status_hip_ko_cpl_spc_data,    //               .ko_cpl_spc_data
		output wire [3:0]  tl_cfg_tl_cfg_add,             //         tl_cfg.tl_cfg_add
		output wire [31:0] tl_cfg_tl_cfg_ctl,             //               .tl_cfg_ctl
		output wire [52:0] tl_cfg_tl_cfg_sts              //               .tl_cfg_sts
	);

	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_readdata;                 // alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> pcie_reconfig_driver_0:reconfig_mgmt_readdata
	wire          pcie_reconfig_driver_0_reconfig_mgmt_waitrequest;              // alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> pcie_reconfig_driver_0:reconfig_mgmt_waitrequest
	wire    [6:0] pcie_reconfig_driver_0_reconfig_mgmt_address;                  // pcie_reconfig_driver_0:reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	wire          pcie_reconfig_driver_0_reconfig_mgmt_read;                     // pcie_reconfig_driver_0:reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	wire          pcie_reconfig_driver_0_reconfig_mgmt_write;                    // pcie_reconfig_driver_0:reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_writedata;                // pcie_reconfig_driver_0:reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	wire          dut_rx_st_valid;                                               // DUT:rx_st_valid -> APPS:rx_st_valid
	wire  [127:0] dut_rx_st_data;                                                // DUT:rx_st_data -> APPS:rx_st_data
	wire          dut_rx_st_ready;                                               // APPS:rx_st_ready -> DUT:rx_st_ready
	wire          dut_rx_st_startofpacket;                                       // DUT:rx_st_sop -> APPS:rx_st_sop
	wire          dut_rx_st_endofpacket;                                         // DUT:rx_st_eop -> APPS:rx_st_eop
	wire          dut_rx_st_error;                                               // DUT:rx_st_err -> APPS:rx_st_err
	wire          dut_rx_st_empty;                                               // DUT:rx_st_empty -> APPS:rx_st_empty
	wire    [0:0] apps_tx_st_valid;                                              // APPS:tx_st_valid -> DUT:tx_st_valid
	wire  [127:0] apps_tx_st_data;                                               // APPS:tx_st_data -> DUT:tx_st_data
	wire          apps_tx_st_ready;                                              // DUT:tx_st_ready -> APPS:tx_st_ready
	wire    [0:0] apps_tx_st_startofpacket;                                      // APPS:tx_st_sop -> DUT:tx_st_sop
	wire    [0:0] apps_tx_st_endofpacket;                                        // APPS:tx_st_eop -> DUT:tx_st_eop
	wire    [0:0] apps_tx_st_error;                                              // APPS:tx_st_err -> DUT:tx_st_err
	wire    [0:0] apps_tx_st_empty;                                              // APPS:tx_st_empty -> DUT:tx_st_empty
	wire          dut_coreclkout_hip_clk;                                        // DUT:coreclkout -> APPS:coreclkout_hip
	wire          apps_pld_clk_hip_clk;                                          // APPS:pld_clk_hip -> [DUT:pld_clk, pcie_av_hip_de_hip_status_0:pld_clk, pcie_reconfig_driver_0:pld_clk]
	wire          pcie_reconfig_driver_0_cal_busy_in_cal_busy_in;                // pcie_reconfig_driver_0:cal_busy_in -> alt_xcvr_reconfig_0:cal_busy_in
	wire          pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_sts_wr;      // pcie_av_hip_de_hip_status_0:to_apps_tl_cfg_sts_wr -> APPS:tl_cfg_sts_wr
	wire    [6:0] apps_config_tl_cpl_err;                                        // APPS:cpl_err -> pcie_av_hip_de_hip_status_0:to_apps_cpl_err
	wire   [52:0] pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_sts;         // pcie_av_hip_de_hip_status_0:to_apps_tl_cfg_sts -> APPS:tl_cfg_sts
	wire          apps_config_tl_cpl_pending;                                    // APPS:cpl_pending -> pcie_av_hip_de_hip_status_0:to_apps_cpl_pending
	wire          pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_ctl_wr;      // pcie_av_hip_de_hip_status_0:to_apps_tl_cfg_ctl_wr -> APPS:tl_cfg_ctl_wr
	wire    [3:0] pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_add;         // pcie_av_hip_de_hip_status_0:to_apps_tl_cfg_add -> APPS:tl_cfg_add
	wire   [31:0] pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_ctl;         // pcie_av_hip_de_hip_status_0:to_apps_tl_cfg_ctl -> APPS:tl_cfg_ctl
	wire    [4:0] apps_config_tl_hpg_ctrler;                                     // APPS:hpg_ctrler -> pcie_av_hip_de_hip_status_0:to_apps_hpg_ctrler
	wire          dut_config_tl_tl_cfg_sts_wr;                                   // DUT:tl_cfg_sts_wr -> pcie_av_hip_de_hip_status_0:to_hip_tl_cfg_sts_wr
	wire    [6:0] pcie_av_hip_de_hip_status_0_config_tl_hip_cpl_err;             // pcie_av_hip_de_hip_status_0:to_hip_cpl_err -> DUT:cpl_err
	wire   [52:0] dut_config_tl_tl_cfg_sts;                                      // DUT:tl_cfg_sts -> pcie_av_hip_de_hip_status_0:to_hip_tl_cfg_sts
	wire          pcie_av_hip_de_hip_status_0_config_tl_hip_cpl_pending;         // pcie_av_hip_de_hip_status_0:to_hip_cpl_pending -> DUT:cpl_pending
	wire          dut_config_tl_tl_cfg_ctl_wr;                                   // DUT:tl_cfg_ctl_wr -> pcie_av_hip_de_hip_status_0:to_hip_tl_cfg_ctl_wr
	wire    [3:0] dut_config_tl_tl_cfg_add;                                      // DUT:tl_cfg_add -> pcie_av_hip_de_hip_status_0:to_hip_tl_cfg_add
	wire   [31:0] dut_config_tl_tl_cfg_ctl;                                      // DUT:tl_cfg_ctl -> pcie_av_hip_de_hip_status_0:to_hip_tl_cfg_ctl
	wire    [4:0] pcie_av_hip_de_hip_status_0_config_tl_hip_hpg_ctrler;          // pcie_av_hip_de_hip_status_0:to_hip_hpg_ctrler -> DUT:tl_hpg_ctrl_er
	wire    [1:0] dut_hip_currentspeed_currentspeed;                             // DUT:dl_current_speed -> pcie_reconfig_driver_0:currentspeed
	wire          dut_hip_rst_serdes_pll_locked;                                 // DUT:serdes_pll_locked -> APPS:serdes_pll_locked
	wire          dut_hip_rst_testin_zero;                                       // DUT:testin_zero -> APPS:testin_zero
	wire          apps_hip_rst_pld_core_ready;                                   // APPS:pld_core_ready -> DUT:pld_core_ready
	wire          dut_hip_rst_reset_status;                                      // DUT:reset_status -> APPS:reset_status
	wire          dut_hip_rst_pld_clk_inuse;                                     // DUT:pld_clk_inuse -> APPS:pld_clk_inuse
	wire          pcie_av_hip_de_hip_status_0_hip_status_apps_derr_cor_ext_rcv;  // pcie_av_hip_de_hip_status_0:to_apps_derr_cor_ext_rcv -> APPS:derr_cor_ext_rcv
	wire          pcie_av_hip_de_hip_status_0_hip_status_apps_hotrst_exit;       // pcie_av_hip_de_hip_status_0:to_apps_hotrst_exit -> APPS:hotrst_exit
	wire   [11:0] pcie_av_hip_de_hip_status_0_hip_status_apps_ko_cpl_spc_data;   // pcie_av_hip_de_hip_status_0:to_apps_ko_cpl_spc_data -> APPS:ko_cpl_spc_data
	wire          pcie_av_hip_de_hip_status_0_hip_status_apps_dlup_exit;         // pcie_av_hip_de_hip_status_0:to_apps_dlup_exit -> APPS:dlup_exit
	wire          pcie_av_hip_de_hip_status_0_hip_status_apps_derr_cor_ext_rpl;  // pcie_av_hip_de_hip_status_0:to_apps_derr_cor_ext_rpl -> APPS:derr_cor_ext_rpl
	wire          pcie_av_hip_de_hip_status_0_hip_status_apps_l2_exit;           // pcie_av_hip_de_hip_status_0:to_apps_l2_exit -> APPS:l2_exit
	wire    [3:0] pcie_av_hip_de_hip_status_0_hip_status_apps_int_status;        // pcie_av_hip_de_hip_status_0:to_apps_int_status -> APPS:int_status
	wire          pcie_av_hip_de_hip_status_0_hip_status_apps_ev128ns;           // pcie_av_hip_de_hip_status_0:to_apps_ev128ns -> APPS:ev128ns
	wire    [4:0] pcie_av_hip_de_hip_status_0_hip_status_apps_ltssmstate;        // pcie_av_hip_de_hip_status_0:to_apps_ltssmstate -> APPS:ltssmstate
	wire    [3:0] pcie_av_hip_de_hip_status_0_hip_status_apps_lane_act;          // pcie_av_hip_de_hip_status_0:to_apps_lane_act -> APPS:lane_act
	wire          pcie_av_hip_de_hip_status_0_hip_status_apps_derr_rpl;          // pcie_av_hip_de_hip_status_0:to_apps_derr_rpl -> APPS:derr_rpl
	wire          pcie_av_hip_de_hip_status_0_hip_status_apps_ev1us;             // pcie_av_hip_de_hip_status_0:to_apps_ev1us -> APPS:ev1us
	wire    [7:0] pcie_av_hip_de_hip_status_0_hip_status_apps_ko_cpl_spc_header; // pcie_av_hip_de_hip_status_0:to_apps_ko_cpl_spc_header -> APPS:ko_cpl_spc_header
	wire          apps_hip_status_drv_derr_cor_ext_rcv;                          // APPS:derr_cor_ext_rcv_drv -> pcie_reconfig_driver_0:derr_cor_ext_rcv_drv
	wire          apps_hip_status_drv_hotrst_exit;                               // APPS:hotrst_exit_drv -> pcie_reconfig_driver_0:hotrst_exit_drv
	wire   [11:0] apps_hip_status_drv_ko_cpl_spc_data;                           // APPS:ko_cpl_spc_data_drv -> pcie_reconfig_driver_0:ko_cpl_spc_data_drv
	wire          apps_hip_status_drv_dlup_exit;                                 // APPS:dlup_exit_drv -> pcie_reconfig_driver_0:dlup_exit_drv
	wire          apps_hip_status_drv_derr_cor_ext_rpl;                          // APPS:derr_cor_ext_rpl_drv -> pcie_reconfig_driver_0:derr_cor_ext_rpl_drv
	wire          apps_hip_status_drv_l2_exit;                                   // APPS:l2_exit_drv -> pcie_reconfig_driver_0:l2_exit_drv
	wire    [3:0] apps_hip_status_drv_int_status;                                // APPS:int_status_drv -> pcie_reconfig_driver_0:int_status_drv
	wire          apps_hip_status_drv_ev128ns;                                   // APPS:ev128ns_drv -> pcie_reconfig_driver_0:ev128ns_drv
	wire    [4:0] apps_hip_status_drv_ltssmstate;                                // APPS:ltssmstate_drv -> pcie_reconfig_driver_0:ltssmstate_drv
	wire    [3:0] apps_hip_status_drv_lane_act;                                  // APPS:lane_act_drv -> pcie_reconfig_driver_0:lane_act_drv
	wire          apps_hip_status_drv_derr_rpl;                                  // APPS:derr_rpl_drv -> pcie_reconfig_driver_0:derr_rpl_drv
	wire          apps_hip_status_drv_ev1us;                                     // APPS:ev1us_drv -> pcie_reconfig_driver_0:ev1us_drv
	wire    [7:0] apps_hip_status_drv_ko_cpl_spc_header;                         // APPS:ko_cpl_spc_header_drv -> pcie_reconfig_driver_0:ko_cpl_spc_header_drv
	wire          dut_hip_status_derr_cor_ext_rcv;                               // DUT:derr_cor_ext_rcv0 -> pcie_av_hip_de_hip_status_0:to_hip_derr_cor_ext_rcv
	wire          dut_hip_status_hotrst_exit;                                    // DUT:hotrst_exit -> pcie_av_hip_de_hip_status_0:to_hip_hotrst_exit
	wire   [11:0] dut_hip_status_ko_cpl_spc_data;                                // DUT:ko_cpl_spc_data -> pcie_av_hip_de_hip_status_0:to_hip_ko_cpl_spc_data
	wire          dut_hip_status_dlup_exit;                                      // DUT:dlup_exit -> pcie_av_hip_de_hip_status_0:to_hip_dlup_exit
	wire          dut_hip_status_derr_cor_ext_rpl;                               // DUT:derr_cor_ext_rpl -> pcie_av_hip_de_hip_status_0:to_hip_derr_cor_ext_rpl
	wire          dut_hip_status_l2_exit;                                        // DUT:l2_exit -> pcie_av_hip_de_hip_status_0:to_hip_l2_exit
	wire    [3:0] dut_hip_status_int_status;                                     // DUT:int_status -> pcie_av_hip_de_hip_status_0:to_hip_int_status
	wire          dut_hip_status_ev128ns;                                        // DUT:ev128ns -> pcie_av_hip_de_hip_status_0:to_hip_ev128ns
	wire    [4:0] dut_hip_status_ltssmstate;                                     // DUT:dl_ltssm -> pcie_av_hip_de_hip_status_0:to_hip_ltssmstate
	wire    [3:0] dut_hip_status_lane_act;                                       // DUT:lane_act -> pcie_av_hip_de_hip_status_0:to_hip_lane_act
	wire          dut_hip_status_derr_rpl;                                       // DUT:derr_rpl -> pcie_av_hip_de_hip_status_0:to_hip_derr_rpl
	wire          dut_hip_status_ev1us;                                          // DUT:ev1us -> pcie_av_hip_de_hip_status_0:to_hip_ev1us
	wire    [7:0] dut_hip_status_ko_cpl_spc_header;                              // DUT:ko_cpl_spc_header -> pcie_av_hip_de_hip_status_0:to_hip_ko_cpl_spc_header
	wire          apps_int_msi_app_msi_req;                                      // APPS:app_msi_req -> DUT:app_msi_req
	wire    [2:0] apps_int_msi_app_msi_tc;                                       // APPS:app_msi_tc -> DUT:app_msi_tc
	wire    [0:0] apps_int_msi_app_int_sts;                                      // APPS:app_int_sts -> DUT:app_int_sts_vec
	wire          dut_int_msi_app_msi_ack;                                       // DUT:app_msi_ack -> APPS:app_msi_ack
	wire    [4:0] apps_int_msi_app_msi_num;                                      // APPS:app_msi_num -> DUT:app_msi_num
	wire          apps_lmi_lmi_rden;                                             // APPS:lmi_rden -> DUT:lmi_rden
	wire   [11:0] apps_lmi_lmi_addr;                                             // APPS:lmi_addr -> DUT:lmi_addr
	wire   [31:0] apps_lmi_lmi_din;                                              // APPS:lmi_din -> DUT:lmi_din
	wire          dut_lmi_lmi_ack;                                               // DUT:lmi_ack -> APPS:lmi_ack
	wire   [31:0] dut_lmi_lmi_dout;                                              // DUT:lmi_dout -> APPS:lmi_dout
	wire          apps_lmi_lmi_wren;                                             // APPS:lmi_wren -> DUT:lmi_wren
	wire          apps_power_mngt_pme_to_cr;                                     // APPS:pme_to_cr -> DUT:pme_to_cr
	wire          dut_power_mngt_pme_to_sr;                                      // DUT:pme_to_sr -> APPS:pme_to_sr
	wire          apps_power_mngt_pm_event;                                      // APPS:pm_event -> DUT:pm_event
	wire          apps_power_mngt_pm_auxpwr;                                     // APPS:pm_auxpwr -> DUT:pm_auxpwr
	wire    [9:0] apps_power_mngt_pm_data;                                       // APPS:pm_data -> DUT:pm_data
	wire          alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy;               // alt_xcvr_reconfig_0:reconfig_busy -> pcie_reconfig_driver_0:reconfig_busy
	wire  [229:0] dut_reconfig_from_xcvr_reconfig_from_xcvr;                     // DUT:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire  [349:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr;         // alt_xcvr_reconfig_0:reconfig_to_xcvr -> DUT:reconfig_to_xcvr
	wire   [15:0] dut_rx_bar_be_rx_st_be;                                        // DUT:rx_st_be -> APPS:rx_st_be
	wire          apps_rx_bar_be_rx_st_mask;                                     // APPS:rx_st_mask -> DUT:rx_st_mask
	wire    [7:0] dut_rx_bar_be_rx_st_bar;                                       // DUT:rx_st_bar -> APPS:rx_st_bar
	wire    [7:0] dut_tx_cred_tx_cred_hdrfcp;                                    // DUT:tx_cred_hdrfcp -> APPS:tx_cred_hdrfcp
	wire   [11:0] dut_tx_cred_tx_cred_datafcp;                                   // DUT:tx_cred_datafcp -> APPS:tx_cred_datafcp
	wire   [11:0] dut_tx_cred_tx_cred_datafccp;                                  // DUT:tx_cred_datafccp -> APPS:tx_cred_datafccp
	wire    [5:0] dut_tx_cred_tx_cred_fchipcons;                                 // DUT:tx_cred_fchipcons -> APPS:tx_cred_fchipcons
	wire    [7:0] dut_tx_cred_tx_cred_hdrfcnp;                                   // DUT:tx_cred_hdrfcnp -> APPS:tx_cred_hdrfcnp
	wire   [11:0] dut_tx_cred_tx_cred_datafcnp;                                  // DUT:tx_cred_datafcnp -> APPS:tx_cred_datafcnp
	wire    [5:0] dut_tx_cred_tx_cred_fcinfinite;                                // DUT:tx_cred_fcinfinite -> APPS:tx_cred_fcinfinite
	wire    [7:0] dut_tx_cred_tx_cred_hdrfccp;                                   // DUT:tx_cred_hdrfccp -> APPS:tx_cred_hdrfccp
	wire          dut_tx_fifo_fifo_empty;                                        // DUT:tx_fifo_empty -> APPS:tx_fifo_empty
	wire          rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, pcie_reconfig_driver_0:reconfig_xcvr_rst]

	altpcied_sv_hwtcl #(
		.device_family_hwtcl              ("Arria V"),
		.lane_mask_hwtcl                  ("x4"),
		.gen123_lane_rate_mode_hwtcl      ("Gen2 (5.0 Gbps)"),
		.pld_clockrate_hwtcl              (125000000),
		.port_type_hwtcl                  ("Native endpoint"),
		.ast_width_hwtcl                  ("Avalon-ST 128-bit"),
		.extend_tag_field_hwtcl           (32),
		.max_payload_size_hwtcl           (256),
		.num_of_func_hwtcl                (1),
		.multiple_packets_per_cycle_hwtcl (0),
		.port_width_be_hwtcl              (16),
		.port_width_data_hwtcl            (128),
		.avalon_waddr_hwltcl              (12),
		.check_bus_master_ena_hwtcl       (1),
		.check_rx_buffer_cpl_hwtcl        (1),
		.use_crc_forwarding_hwtcl         (0)
	) apps (
		.coreclkout_hip        (dut_coreclkout_hip_clk),                                        // coreclkout_hip.clk
		.pld_clk_hip           (apps_pld_clk_hip_clk),                                          //    pld_clk_hip.clk
		.rx_st_sop             (dut_rx_st_startofpacket),                                       //          rx_st.startofpacket
		.rx_st_eop             (dut_rx_st_endofpacket),                                         //               .endofpacket
		.rx_st_err             (dut_rx_st_error),                                               //               .error
		.rx_st_valid           (dut_rx_st_valid),                                               //               .valid
		.rx_st_empty           (dut_rx_st_empty),                                               //               .empty
		.rx_st_ready           (dut_rx_st_ready),                                               //               .ready
		.rx_st_data            (dut_rx_st_data),                                                //               .data
		.rx_st_bar             (dut_rx_bar_be_rx_st_bar),                                       //      rx_bar_be.rx_st_bar
		.rx_st_be              (dut_rx_bar_be_rx_st_be),                                        //               .rx_st_be
		.rx_st_mask            (apps_rx_bar_be_rx_st_mask),                                     //               .rx_st_mask
		.tx_st_sop             (apps_tx_st_startofpacket),                                      //          tx_st.startofpacket
		.tx_st_eop             (apps_tx_st_endofpacket),                                        //               .endofpacket
		.tx_st_err             (apps_tx_st_error),                                              //               .error
		.tx_st_valid           (apps_tx_st_valid),                                              //               .valid
		.tx_st_empty           (apps_tx_st_empty),                                              //               .empty
		.tx_st_ready           (apps_tx_st_ready),                                              //               .ready
		.tx_st_data            (apps_tx_st_data),                                               //               .data
		.tx_fifo_empty         (dut_tx_fifo_fifo_empty),                                        //        tx_fifo.fifo_empty
		.tx_cred_datafccp      (dut_tx_cred_tx_cred_datafccp),                                  //        tx_cred.tx_cred_datafccp
		.tx_cred_datafcnp      (dut_tx_cred_tx_cred_datafcnp),                                  //               .tx_cred_datafcnp
		.tx_cred_datafcp       (dut_tx_cred_tx_cred_datafcp),                                   //               .tx_cred_datafcp
		.tx_cred_fchipcons     (dut_tx_cred_tx_cred_fchipcons),                                 //               .tx_cred_fchipcons
		.tx_cred_fcinfinite    (dut_tx_cred_tx_cred_fcinfinite),                                //               .tx_cred_fcinfinite
		.tx_cred_hdrfccp       (dut_tx_cred_tx_cred_hdrfccp),                                   //               .tx_cred_hdrfccp
		.tx_cred_hdrfcnp       (dut_tx_cred_tx_cred_hdrfcnp),                                   //               .tx_cred_hdrfcnp
		.tx_cred_hdrfcp        (dut_tx_cred_tx_cred_hdrfcp),                                    //               .tx_cred_hdrfcp
		.reset_status          (dut_hip_rst_reset_status),                                      //        hip_rst.reset_status
		.serdes_pll_locked     (dut_hip_rst_serdes_pll_locked),                                 //               .serdes_pll_locked
		.pld_clk_inuse         (dut_hip_rst_pld_clk_inuse),                                     //               .pld_clk_inuse
		.pld_core_ready        (apps_hip_rst_pld_core_ready),                                   //               .pld_core_ready
		.testin_zero           (dut_hip_rst_testin_zero),                                       //               .testin_zero
		.app_int_sts           (apps_int_msi_app_int_sts),                                      //        int_msi.app_int_sts
		.app_msi_req           (apps_int_msi_app_msi_req),                                      //               .app_msi_req
		.app_msi_tc            (apps_int_msi_app_msi_tc),                                       //               .app_msi_tc
		.app_msi_ack           (dut_int_msi_app_msi_ack),                                       //               .app_msi_ack
		.app_msi_num           (apps_int_msi_app_msi_num),                                      //               .app_msi_num
		.derr_cor_ext_rcv      (pcie_av_hip_de_hip_status_0_hip_status_apps_derr_cor_ext_rcv),  //     hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl      (pcie_av_hip_de_hip_status_0_hip_status_apps_derr_cor_ext_rpl),  //               .derr_cor_ext_rpl
		.derr_rpl              (pcie_av_hip_de_hip_status_0_hip_status_apps_derr_rpl),          //               .derr_rpl
		.dlup_exit             (pcie_av_hip_de_hip_status_0_hip_status_apps_dlup_exit),         //               .dlup_exit
		.ev128ns               (pcie_av_hip_de_hip_status_0_hip_status_apps_ev128ns),           //               .ev128ns
		.ev1us                 (pcie_av_hip_de_hip_status_0_hip_status_apps_ev1us),             //               .ev1us
		.hotrst_exit           (pcie_av_hip_de_hip_status_0_hip_status_apps_hotrst_exit),       //               .hotrst_exit
		.int_status            (pcie_av_hip_de_hip_status_0_hip_status_apps_int_status),        //               .int_status
		.l2_exit               (pcie_av_hip_de_hip_status_0_hip_status_apps_l2_exit),           //               .l2_exit
		.lane_act              (pcie_av_hip_de_hip_status_0_hip_status_apps_lane_act),          //               .lane_act
		.ltssmstate            (pcie_av_hip_de_hip_status_0_hip_status_apps_ltssmstate),        //               .ltssmstate
		.ko_cpl_spc_header     (pcie_av_hip_de_hip_status_0_hip_status_apps_ko_cpl_spc_header), //               .ko_cpl_spc_header
		.ko_cpl_spc_data       (pcie_av_hip_de_hip_status_0_hip_status_apps_ko_cpl_spc_data),   //               .ko_cpl_spc_data
		.derr_cor_ext_rcv_drv  (apps_hip_status_drv_derr_cor_ext_rcv),                          // hip_status_drv.derr_cor_ext_rcv
		.derr_cor_ext_rpl_drv  (apps_hip_status_drv_derr_cor_ext_rpl),                          //               .derr_cor_ext_rpl
		.derr_rpl_drv          (apps_hip_status_drv_derr_rpl),                                  //               .derr_rpl
		.dlup_exit_drv         (apps_hip_status_drv_dlup_exit),                                 //               .dlup_exit
		.ev128ns_drv           (apps_hip_status_drv_ev128ns),                                   //               .ev128ns
		.ev1us_drv             (apps_hip_status_drv_ev1us),                                     //               .ev1us
		.hotrst_exit_drv       (apps_hip_status_drv_hotrst_exit),                               //               .hotrst_exit
		.int_status_drv        (apps_hip_status_drv_int_status),                                //               .int_status
		.l2_exit_drv           (apps_hip_status_drv_l2_exit),                                   //               .l2_exit
		.lane_act_drv          (apps_hip_status_drv_lane_act),                                  //               .lane_act
		.ltssmstate_drv        (apps_hip_status_drv_ltssmstate),                                //               .ltssmstate
		.ko_cpl_spc_header_drv (apps_hip_status_drv_ko_cpl_spc_header),                         //               .ko_cpl_spc_header
		.ko_cpl_spc_data_drv   (apps_hip_status_drv_ko_cpl_spc_data),                           //               .ko_cpl_spc_data
		.hpg_ctrler            (apps_config_tl_hpg_ctrler),                                     //      config_tl.hpg_ctrler
		.tl_cfg_ctl            (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_ctl),         //               .tl_cfg_ctl
		.cpl_err               (apps_config_tl_cpl_err),                                        //               .cpl_err
		.tl_cfg_ctl_wr         (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_ctl_wr),      //               .tl_cfg_ctl_wr
		.tl_cfg_sts_wr         (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_sts_wr),      //               .tl_cfg_sts_wr
		.tl_cfg_add            (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_add),         //               .tl_cfg_add
		.tl_cfg_sts            (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_sts),         //               .tl_cfg_sts
		.cpl_pending           (apps_config_tl_cpl_pending),                                    //               .cpl_pending
		.lmi_addr              (apps_lmi_lmi_addr),                                             //            lmi.lmi_addr
		.lmi_din               (apps_lmi_lmi_din),                                              //               .lmi_din
		.lmi_rden              (apps_lmi_lmi_rden),                                             //               .lmi_rden
		.lmi_wren              (apps_lmi_lmi_wren),                                             //               .lmi_wren
		.lmi_ack               (dut_lmi_lmi_ack),                                               //               .lmi_ack
		.lmi_dout              (dut_lmi_lmi_dout),                                              //               .lmi_dout
		.pm_auxpwr             (apps_power_mngt_pm_auxpwr),                                     //     power_mngt.pm_auxpwr
		.pm_data               (apps_power_mngt_pm_data),                                       //               .pm_data
		.pme_to_cr             (apps_power_mngt_pme_to_cr),                                     //               .pme_to_cr
		.pm_event              (apps_power_mngt_pm_event),                                      //               .pm_event
		.pme_to_sr             (dut_power_mngt_pme_to_sr),                                      //               .pme_to_sr
		.rx_st_parity          (16'b0000000000000000),                                          //    (terminated)
		.rx_bar_dec_func_num   (3'b000),                                                        //    (terminated)
		.tx_st_parity          (),                                                              //    (terminated)
		.sim_pipe_pclk_out     (1'b0),                                                          //    (terminated)
		.app_int_ack           (1'b0),                                                          //    (terminated)
		.app_msi_func          (),                                                              //    (terminated)
		.serr_out              (1'b0),                                                          //    (terminated)
		.dlup                  (1'b0),                                                          //    (terminated)
		.rx_par_err            (1'b0),                                                          //    (terminated)
		.tx_par_err            (2'b00),                                                         //    (terminated)
		.cfg_par_err           (1'b0),                                                          //    (terminated)
		.rxfc_cplbuf_ovf       (1'b0),                                                          //    (terminated)
		.cpl_err_func          (),                                                              //    (terminated)
		.pm_event_func         ()                                                               //    (terminated)
	);

	altpcie_av_hip_ast_hwtcl #(
		.ACDS_VERSION_HWTCL                        ("14.0"),
		.lane_mask_hwtcl                           ("x4"),
		.gen12_lane_rate_mode_hwtcl                ("Gen2 (5.0 Gbps)"),
		.pcie_spec_version_hwtcl                   ("2.1"),
		.ast_width_hwtcl                           ("Avalon-ST 128-bit"),
		.pll_refclk_freq_hwtcl                     ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl               (0),
		.in_cvp_mode_hwtcl                         (0),
		.hip_reconfig_hwtcl                        (0),
		.num_of_func_hwtcl                         (1),
		.use_crc_forwarding_hwtcl                  (0),
		.port_link_number_hwtcl                    (1),
		.slotclkcfg_hwtcl                          (1),
		.enable_slot_register_hwtcl                (0),
		.vsec_id_hwtcl                             (4466),
		.vsec_rev_hwtcl                            (0),
		.user_id_hwtcl                             (0),
		.porttype_func0_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_0_hwtcl                    (20),
		.bar0_io_space_0_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_0_hwtcl              ("Disabled"),
		.bar0_prefetchable_0_hwtcl                 ("Disabled"),
		.bar1_size_mask_0_hwtcl                    (0),
		.bar1_io_space_0_hwtcl                     ("Disabled"),
		.bar1_prefetchable_0_hwtcl                 ("Disabled"),
		.bar2_size_mask_0_hwtcl                    (10),
		.bar2_io_space_0_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_0_hwtcl              ("Disabled"),
		.bar2_prefetchable_0_hwtcl                 ("Disabled"),
		.bar3_size_mask_0_hwtcl                    (0),
		.bar3_io_space_0_hwtcl                     ("Disabled"),
		.bar3_prefetchable_0_hwtcl                 ("Disabled"),
		.bar4_size_mask_0_hwtcl                    (0),
		.bar4_io_space_0_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_0_hwtcl              ("Disabled"),
		.bar4_prefetchable_0_hwtcl                 ("Disabled"),
		.bar5_size_mask_0_hwtcl                    (0),
		.bar5_io_space_0_hwtcl                     ("Disabled"),
		.bar5_prefetchable_0_hwtcl                 ("Disabled"),
		.expansion_base_address_register_0_hwtcl   (0),
		.io_window_addr_width_hwtcl                (0),
		.prefetchable_mem_window_addr_width_hwtcl  (0),
		.vendor_id_0_hwtcl                         (4466),
		.device_id_0_hwtcl                         (57345),
		.revision_id_0_hwtcl                       (1),
		.class_code_0_hwtcl                        (0),
		.subsystem_vendor_id_0_hwtcl               (198),
		.subsystem_device_id_0_hwtcl               (8560),
		.max_payload_size_0_hwtcl                  (256),
		.extend_tag_field_0_hwtcl                  ("32"),
		.completion_timeout_0_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_0_hwtcl (1),
		.flr_capability_0_hwtcl                    (0),
		.use_aer_0_hwtcl                           (0),
		.ecrc_check_capable_0_hwtcl                (0),
		.ecrc_gen_capable_0_hwtcl                  (0),
		.dll_active_report_support_0_hwtcl         (0),
		.surprise_down_error_support_0_hwtcl       (0),
		.msi_multi_message_capable_0_hwtcl         ("4"),
		.msi_64bit_addressing_capable_0_hwtcl      ("true"),
		.msi_masking_capable_0_hwtcl               ("false"),
		.msi_support_0_hwtcl                       ("true"),
		.enable_function_msix_support_0_hwtcl      (0),
		.msix_table_size_0_hwtcl                   (0),
		.msix_table_offset_0_hwtcl                 ("0"),
		.msix_table_bir_0_hwtcl                    (0),
		.msix_pba_offset_0_hwtcl                   ("0"),
		.msix_pba_bir_0_hwtcl                      (0),
		.interrupt_pin_0_hwtcl                     ("inta"),
		.slot_power_scale_0_hwtcl                  (0),
		.slot_power_limit_0_hwtcl                  (0),
		.slot_number_0_hwtcl                       (0),
		.rx_ei_l0s_0_hwtcl                         (0),
		.endpoint_l0_latency_0_hwtcl               (0),
		.endpoint_l1_latency_0_hwtcl               (0),
		.reconfig_to_xcvr_width                    (350),
		.hip_hard_reset_hwtcl                      (1),
		.reconfig_from_xcvr_width                  (230),
		.single_rx_detect_hwtcl                    (4),
		.enable_l0s_aspm_hwtcl                     ("false"),
		.aspm_optionality_hwtcl                    ("true"),
		.enable_adapter_half_rate_mode_hwtcl       ("true"),
		.millisecond_cycle_count_hwtcl             (124250),
		.credit_buffer_allocation_aux_hwtcl        ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl      (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl        (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl   (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl     (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl       (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl         (0),
		.cpl_spc_header_hwtcl                      (67),
		.cpl_spc_data_hwtcl                        (269),
		.port_width_data_hwtcl                     (128),
		.bypass_clk_switch_hwtcl                   ("disable"),
		.cvp_rate_sel_hwtcl                        ("full_rate"),
		.cvp_data_compressed_hwtcl                 ("false"),
		.cvp_data_encrypted_hwtcl                  ("false"),
		.cvp_mode_reset_hwtcl                      ("false"),
		.cvp_clk_reset_hwtcl                       ("false"),
		.core_clk_sel_hwtcl                        ("pld_clk"),
		.enable_rx_buffer_checking_hwtcl           ("false"),
		.disable_link_x2_support_hwtcl             ("false"),
		.device_number_hwtcl                       (0),
		.pipex1_debug_sel_hwtcl                    ("disable"),
		.pclk_out_sel_hwtcl                        ("pclk"),
		.no_soft_reset_hwtcl                       ("false"),
		.d1_support_hwtcl                          ("false"),
		.d2_support_hwtcl                          ("false"),
		.d0_pme_hwtcl                              ("false"),
		.d1_pme_hwtcl                              ("false"),
		.d2_pme_hwtcl                              ("false"),
		.d3_hot_pme_hwtcl                          ("false"),
		.d3_cold_pme_hwtcl                         ("false"),
		.low_priority_vc_hwtcl                     ("single_vc"),
		.enable_l1_aspm_hwtcl                      ("false"),
		.l1_exit_latency_sameclock_hwtcl           (0),
		.l1_exit_latency_diffclock_hwtcl           (0),
		.hot_plug_support_hwtcl                    (0),
		.no_command_completed_hwtcl                ("false"),
		.eie_before_nfts_count_hwtcl               (4),
		.gen2_diffclock_nfts_count_hwtcl           (255),
		.gen2_sameclock_nfts_count_hwtcl           (255),
		.deemphasis_enable_hwtcl                   ("false"),
		.l0_exit_latency_sameclock_hwtcl           (6),
		.l0_exit_latency_diffclock_hwtcl           (6),
		.vc0_clk_enable_hwtcl                      ("true"),
		.register_pipe_signals_hwtcl               ("true"),
		.tx_cdc_almost_empty_hwtcl                 (5),
		.rx_l0s_count_idl_hwtcl                    (0),
		.cdc_dummy_insert_limit_hwtcl              (11),
		.ei_delay_powerdown_count_hwtcl            (10),
		.skp_os_schedule_count_hwtcl               (0),
		.fc_init_timer_hwtcl                       (1024),
		.l01_entry_latency_hwtcl                   (31),
		.flow_control_update_count_hwtcl           (30),
		.flow_control_timeout_count_hwtcl          (200),
		.retry_buffer_last_active_address_hwtcl    (255),
		.reserved_debug_hwtcl                      (0),
		.use_tl_cfg_sync_hwtcl                     (1),
		.diffclock_nfts_count_hwtcl                (255),
		.sameclock_nfts_count_hwtcl                (255),
		.l2_async_logic_hwtcl                      ("disable"),
		.rx_cdc_almost_full_hwtcl                  (12),
		.tx_cdc_almost_full_hwtcl                  (11),
		.indicator_hwtcl                           (0),
		.maximum_current_0_hwtcl                   (0),
		.disable_snoop_packet_0_hwtcl              ("false"),
		.bridge_port_vga_enable_0_hwtcl            ("false"),
		.bridge_port_ssid_support_0_hwtcl          ("false"),
		.ssvid_0_hwtcl                             (0),
		.ssid_0_hwtcl                              (0),
		.porttype_func1_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_1_hwtcl                    (28),
		.bar0_io_space_1_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_1_hwtcl              ("Enabled"),
		.bar0_prefetchable_1_hwtcl                 ("Enabled"),
		.bar1_size_mask_1_hwtcl                    (0),
		.bar1_io_space_1_hwtcl                     ("Disabled"),
		.bar1_prefetchable_1_hwtcl                 ("Disabled"),
		.bar2_size_mask_1_hwtcl                    (10),
		.bar2_io_space_1_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_1_hwtcl              ("Disabled"),
		.bar2_prefetchable_1_hwtcl                 ("Disabled"),
		.bar3_size_mask_1_hwtcl                    (0),
		.bar3_io_space_1_hwtcl                     ("Disabled"),
		.bar3_prefetchable_1_hwtcl                 ("Disabled"),
		.bar4_size_mask_1_hwtcl                    (0),
		.bar4_io_space_1_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_1_hwtcl              ("Disabled"),
		.bar4_prefetchable_1_hwtcl                 ("Disabled"),
		.bar5_size_mask_1_hwtcl                    (0),
		.bar5_io_space_1_hwtcl                     ("Disabled"),
		.bar5_prefetchable_1_hwtcl                 ("Disabled"),
		.expansion_base_address_register_1_hwtcl   (0),
		.vendor_id_1_hwtcl                         (0),
		.device_id_1_hwtcl                         (1),
		.revision_id_1_hwtcl                       (1),
		.class_code_1_hwtcl                        (0),
		.subsystem_vendor_id_1_hwtcl               (0),
		.subsystem_device_id_1_hwtcl               (0),
		.max_payload_size_1_hwtcl                  (256),
		.extend_tag_field_1_hwtcl                  ("32"),
		.completion_timeout_1_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_1_hwtcl (1),
		.flr_capability_1_hwtcl                    (0),
		.use_aer_1_hwtcl                           (0),
		.ecrc_check_capable_1_hwtcl                (0),
		.ecrc_gen_capable_1_hwtcl                  (0),
		.dll_active_report_support_1_hwtcl         (0),
		.surprise_down_error_support_1_hwtcl       (0),
		.msi_multi_message_capable_1_hwtcl         ("4"),
		.msi_64bit_addressing_capable_1_hwtcl      ("true"),
		.msi_masking_capable_1_hwtcl               ("false"),
		.msi_support_1_hwtcl                       ("true"),
		.enable_function_msix_support_1_hwtcl      (0),
		.msix_table_size_1_hwtcl                   (0),
		.msix_table_offset_1_hwtcl                 ("0"),
		.msix_table_bir_1_hwtcl                    (0),
		.msix_pba_offset_1_hwtcl                   ("0"),
		.msix_pba_bir_1_hwtcl                      (0),
		.interrupt_pin_1_hwtcl                     ("inta"),
		.slot_power_scale_1_hwtcl                  (0),
		.slot_power_limit_1_hwtcl                  (0),
		.slot_number_1_hwtcl                       (0),
		.rx_ei_l0s_1_hwtcl                         (0),
		.endpoint_l0_latency_1_hwtcl               (0),
		.endpoint_l1_latency_1_hwtcl               (0),
		.maximum_current_1_hwtcl                   (0),
		.disable_snoop_packet_1_hwtcl              ("false"),
		.bridge_port_vga_enable_1_hwtcl            ("false"),
		.bridge_port_ssid_support_1_hwtcl          ("false"),
		.ssvid_1_hwtcl                             (0),
		.ssid_1_hwtcl                              (0),
		.porttype_func2_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_2_hwtcl                    (28),
		.bar0_io_space_2_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_2_hwtcl              ("Enabled"),
		.bar0_prefetchable_2_hwtcl                 ("Enabled"),
		.bar1_size_mask_2_hwtcl                    (0),
		.bar1_io_space_2_hwtcl                     ("Disabled"),
		.bar1_prefetchable_2_hwtcl                 ("Disabled"),
		.bar2_size_mask_2_hwtcl                    (10),
		.bar2_io_space_2_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_2_hwtcl              ("Disabled"),
		.bar2_prefetchable_2_hwtcl                 ("Disabled"),
		.bar3_size_mask_2_hwtcl                    (0),
		.bar3_io_space_2_hwtcl                     ("Disabled"),
		.bar3_prefetchable_2_hwtcl                 ("Disabled"),
		.bar4_size_mask_2_hwtcl                    (0),
		.bar4_io_space_2_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_2_hwtcl              ("Disabled"),
		.bar4_prefetchable_2_hwtcl                 ("Disabled"),
		.bar5_size_mask_2_hwtcl                    (0),
		.bar5_io_space_2_hwtcl                     ("Disabled"),
		.bar5_prefetchable_2_hwtcl                 ("Disabled"),
		.expansion_base_address_register_2_hwtcl   (0),
		.vendor_id_2_hwtcl                         (0),
		.device_id_2_hwtcl                         (1),
		.revision_id_2_hwtcl                       (1),
		.class_code_2_hwtcl                        (0),
		.subsystem_vendor_id_2_hwtcl               (0),
		.subsystem_device_id_2_hwtcl               (0),
		.max_payload_size_2_hwtcl                  (256),
		.extend_tag_field_2_hwtcl                  ("32"),
		.completion_timeout_2_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_2_hwtcl (1),
		.flr_capability_2_hwtcl                    (0),
		.use_aer_2_hwtcl                           (0),
		.ecrc_check_capable_2_hwtcl                (0),
		.ecrc_gen_capable_2_hwtcl                  (0),
		.dll_active_report_support_2_hwtcl         (0),
		.surprise_down_error_support_2_hwtcl       (0),
		.msi_multi_message_capable_2_hwtcl         ("4"),
		.msi_64bit_addressing_capable_2_hwtcl      ("true"),
		.msi_masking_capable_2_hwtcl               ("false"),
		.msi_support_2_hwtcl                       ("true"),
		.enable_function_msix_support_2_hwtcl      (0),
		.msix_table_size_2_hwtcl                   (0),
		.msix_table_offset_2_hwtcl                 ("0"),
		.msix_table_bir_2_hwtcl                    (0),
		.msix_pba_offset_2_hwtcl                   ("0"),
		.msix_pba_bir_2_hwtcl                      (0),
		.interrupt_pin_2_hwtcl                     ("inta"),
		.slot_power_scale_2_hwtcl                  (0),
		.slot_power_limit_2_hwtcl                  (0),
		.slot_number_2_hwtcl                       (0),
		.rx_ei_l0s_2_hwtcl                         (0),
		.endpoint_l0_latency_2_hwtcl               (0),
		.endpoint_l1_latency_2_hwtcl               (0),
		.maximum_current_2_hwtcl                   (0),
		.disable_snoop_packet_2_hwtcl              ("false"),
		.bridge_port_vga_enable_2_hwtcl            ("false"),
		.bridge_port_ssid_support_2_hwtcl          ("false"),
		.ssvid_2_hwtcl                             (0),
		.ssid_2_hwtcl                              (0),
		.porttype_func3_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_3_hwtcl                    (28),
		.bar0_io_space_3_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_3_hwtcl              ("Enabled"),
		.bar0_prefetchable_3_hwtcl                 ("Enabled"),
		.bar1_size_mask_3_hwtcl                    (0),
		.bar1_io_space_3_hwtcl                     ("Disabled"),
		.bar1_prefetchable_3_hwtcl                 ("Disabled"),
		.bar2_size_mask_3_hwtcl                    (10),
		.bar2_io_space_3_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_3_hwtcl              ("Disabled"),
		.bar2_prefetchable_3_hwtcl                 ("Disabled"),
		.bar3_size_mask_3_hwtcl                    (0),
		.bar3_io_space_3_hwtcl                     ("Disabled"),
		.bar3_prefetchable_3_hwtcl                 ("Disabled"),
		.bar4_size_mask_3_hwtcl                    (0),
		.bar4_io_space_3_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_3_hwtcl              ("Disabled"),
		.bar4_prefetchable_3_hwtcl                 ("Disabled"),
		.bar5_size_mask_3_hwtcl                    (0),
		.bar5_io_space_3_hwtcl                     ("Disabled"),
		.bar5_prefetchable_3_hwtcl                 ("Disabled"),
		.expansion_base_address_register_3_hwtcl   (0),
		.vendor_id_3_hwtcl                         (0),
		.device_id_3_hwtcl                         (1),
		.revision_id_3_hwtcl                       (1),
		.class_code_3_hwtcl                        (0),
		.subsystem_vendor_id_3_hwtcl               (0),
		.subsystem_device_id_3_hwtcl               (0),
		.max_payload_size_3_hwtcl                  (256),
		.extend_tag_field_3_hwtcl                  ("32"),
		.completion_timeout_3_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_3_hwtcl (1),
		.flr_capability_3_hwtcl                    (0),
		.use_aer_3_hwtcl                           (0),
		.ecrc_check_capable_3_hwtcl                (0),
		.ecrc_gen_capable_3_hwtcl                  (0),
		.dll_active_report_support_3_hwtcl         (0),
		.surprise_down_error_support_3_hwtcl       (0),
		.msi_multi_message_capable_3_hwtcl         ("4"),
		.msi_64bit_addressing_capable_3_hwtcl      ("true"),
		.msi_masking_capable_3_hwtcl               ("false"),
		.msi_support_3_hwtcl                       ("true"),
		.enable_function_msix_support_3_hwtcl      (0),
		.msix_table_size_3_hwtcl                   (0),
		.msix_table_offset_3_hwtcl                 ("0"),
		.msix_table_bir_3_hwtcl                    (0),
		.msix_pba_offset_3_hwtcl                   ("0"),
		.msix_pba_bir_3_hwtcl                      (0),
		.interrupt_pin_3_hwtcl                     ("inta"),
		.slot_power_scale_3_hwtcl                  (0),
		.slot_power_limit_3_hwtcl                  (0),
		.slot_number_3_hwtcl                       (0),
		.rx_ei_l0s_3_hwtcl                         (0),
		.endpoint_l0_latency_3_hwtcl               (0),
		.endpoint_l1_latency_3_hwtcl               (0),
		.maximum_current_3_hwtcl                   (0),
		.disable_snoop_packet_3_hwtcl              ("false"),
		.bridge_port_vga_enable_3_hwtcl            ("false"),
		.bridge_port_ssid_support_3_hwtcl          ("false"),
		.ssvid_3_hwtcl                             (0),
		.ssid_3_hwtcl                              (0),
		.porttype_func4_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_4_hwtcl                    (28),
		.bar0_io_space_4_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_4_hwtcl              ("Enabled"),
		.bar0_prefetchable_4_hwtcl                 ("Enabled"),
		.bar1_size_mask_4_hwtcl                    (0),
		.bar1_io_space_4_hwtcl                     ("Disabled"),
		.bar1_prefetchable_4_hwtcl                 ("Disabled"),
		.bar2_size_mask_4_hwtcl                    (10),
		.bar2_io_space_4_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_4_hwtcl              ("Disabled"),
		.bar2_prefetchable_4_hwtcl                 ("Disabled"),
		.bar3_size_mask_4_hwtcl                    (0),
		.bar3_io_space_4_hwtcl                     ("Disabled"),
		.bar3_prefetchable_4_hwtcl                 ("Disabled"),
		.bar4_size_mask_4_hwtcl                    (0),
		.bar4_io_space_4_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_4_hwtcl              ("Disabled"),
		.bar4_prefetchable_4_hwtcl                 ("Disabled"),
		.bar5_size_mask_4_hwtcl                    (0),
		.bar5_io_space_4_hwtcl                     ("Disabled"),
		.bar5_prefetchable_4_hwtcl                 ("Disabled"),
		.expansion_base_address_register_4_hwtcl   (0),
		.vendor_id_4_hwtcl                         (0),
		.device_id_4_hwtcl                         (1),
		.revision_id_4_hwtcl                       (1),
		.class_code_4_hwtcl                        (0),
		.subsystem_vendor_id_4_hwtcl               (0),
		.subsystem_device_id_4_hwtcl               (0),
		.max_payload_size_4_hwtcl                  (256),
		.extend_tag_field_4_hwtcl                  ("32"),
		.completion_timeout_4_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_4_hwtcl (1),
		.flr_capability_4_hwtcl                    (0),
		.use_aer_4_hwtcl                           (0),
		.ecrc_check_capable_4_hwtcl                (0),
		.ecrc_gen_capable_4_hwtcl                  (0),
		.dll_active_report_support_4_hwtcl         (0),
		.surprise_down_error_support_4_hwtcl       (0),
		.msi_multi_message_capable_4_hwtcl         ("4"),
		.msi_64bit_addressing_capable_4_hwtcl      ("true"),
		.msi_masking_capable_4_hwtcl               ("false"),
		.msi_support_4_hwtcl                       ("true"),
		.enable_function_msix_support_4_hwtcl      (0),
		.msix_table_size_4_hwtcl                   (0),
		.msix_table_offset_4_hwtcl                 ("0"),
		.msix_table_bir_4_hwtcl                    (0),
		.msix_pba_offset_4_hwtcl                   ("0"),
		.msix_pba_bir_4_hwtcl                      (0),
		.interrupt_pin_4_hwtcl                     ("inta"),
		.slot_power_scale_4_hwtcl                  (0),
		.slot_power_limit_4_hwtcl                  (0),
		.slot_number_4_hwtcl                       (0),
		.rx_ei_l0s_4_hwtcl                         (0),
		.endpoint_l0_latency_4_hwtcl               (0),
		.endpoint_l1_latency_4_hwtcl               (0),
		.maximum_current_4_hwtcl                   (0),
		.disable_snoop_packet_4_hwtcl              ("false"),
		.bridge_port_vga_enable_4_hwtcl            ("false"),
		.bridge_port_ssid_support_4_hwtcl          ("false"),
		.ssvid_4_hwtcl                             (0),
		.ssid_4_hwtcl                              (0),
		.porttype_func5_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_5_hwtcl                    (28),
		.bar0_io_space_5_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_5_hwtcl              ("Enabled"),
		.bar0_prefetchable_5_hwtcl                 ("Enabled"),
		.bar1_size_mask_5_hwtcl                    (0),
		.bar1_io_space_5_hwtcl                     ("Disabled"),
		.bar1_prefetchable_5_hwtcl                 ("Disabled"),
		.bar2_size_mask_5_hwtcl                    (10),
		.bar2_io_space_5_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_5_hwtcl              ("Disabled"),
		.bar2_prefetchable_5_hwtcl                 ("Disabled"),
		.bar3_size_mask_5_hwtcl                    (0),
		.bar3_io_space_5_hwtcl                     ("Disabled"),
		.bar3_prefetchable_5_hwtcl                 ("Disabled"),
		.bar4_size_mask_5_hwtcl                    (0),
		.bar4_io_space_5_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_5_hwtcl              ("Disabled"),
		.bar4_prefetchable_5_hwtcl                 ("Disabled"),
		.bar5_size_mask_5_hwtcl                    (0),
		.bar5_io_space_5_hwtcl                     ("Disabled"),
		.bar5_prefetchable_5_hwtcl                 ("Disabled"),
		.expansion_base_address_register_5_hwtcl   (0),
		.vendor_id_5_hwtcl                         (0),
		.device_id_5_hwtcl                         (1),
		.revision_id_5_hwtcl                       (1),
		.class_code_5_hwtcl                        (0),
		.subsystem_vendor_id_5_hwtcl               (0),
		.subsystem_device_id_5_hwtcl               (0),
		.max_payload_size_5_hwtcl                  (256),
		.extend_tag_field_5_hwtcl                  ("32"),
		.completion_timeout_5_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_5_hwtcl (1),
		.flr_capability_5_hwtcl                    (0),
		.use_aer_5_hwtcl                           (0),
		.ecrc_check_capable_5_hwtcl                (0),
		.ecrc_gen_capable_5_hwtcl                  (0),
		.dll_active_report_support_5_hwtcl         (0),
		.surprise_down_error_support_5_hwtcl       (0),
		.msi_multi_message_capable_5_hwtcl         ("4"),
		.msi_64bit_addressing_capable_5_hwtcl      ("true"),
		.msi_masking_capable_5_hwtcl               ("false"),
		.msi_support_5_hwtcl                       ("true"),
		.enable_function_msix_support_5_hwtcl      (0),
		.msix_table_size_5_hwtcl                   (0),
		.msix_table_offset_5_hwtcl                 ("0"),
		.msix_table_bir_5_hwtcl                    (0),
		.msix_pba_offset_5_hwtcl                   ("0"),
		.msix_pba_bir_5_hwtcl                      (0),
		.interrupt_pin_5_hwtcl                     ("inta"),
		.slot_power_scale_5_hwtcl                  (0),
		.slot_power_limit_5_hwtcl                  (0),
		.slot_number_5_hwtcl                       (0),
		.rx_ei_l0s_5_hwtcl                         (0),
		.endpoint_l0_latency_5_hwtcl               (0),
		.endpoint_l1_latency_5_hwtcl               (0),
		.maximum_current_5_hwtcl                   (0),
		.disable_snoop_packet_5_hwtcl              ("false"),
		.bridge_port_vga_enable_5_hwtcl            ("false"),
		.bridge_port_ssid_support_5_hwtcl          ("false"),
		.ssvid_5_hwtcl                             (0),
		.ssid_5_hwtcl                              (0),
		.porttype_func6_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_6_hwtcl                    (28),
		.bar0_io_space_6_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_6_hwtcl              ("Enabled"),
		.bar0_prefetchable_6_hwtcl                 ("Enabled"),
		.bar1_size_mask_6_hwtcl                    (0),
		.bar1_io_space_6_hwtcl                     ("Disabled"),
		.bar1_prefetchable_6_hwtcl                 ("Disabled"),
		.bar2_size_mask_6_hwtcl                    (10),
		.bar2_io_space_6_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_6_hwtcl              ("Disabled"),
		.bar2_prefetchable_6_hwtcl                 ("Disabled"),
		.bar3_size_mask_6_hwtcl                    (0),
		.bar3_io_space_6_hwtcl                     ("Disabled"),
		.bar3_prefetchable_6_hwtcl                 ("Disabled"),
		.bar4_size_mask_6_hwtcl                    (0),
		.bar4_io_space_6_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_6_hwtcl              ("Disabled"),
		.bar4_prefetchable_6_hwtcl                 ("Disabled"),
		.bar5_size_mask_6_hwtcl                    (0),
		.bar5_io_space_6_hwtcl                     ("Disabled"),
		.bar5_prefetchable_6_hwtcl                 ("Disabled"),
		.expansion_base_address_register_6_hwtcl   (0),
		.vendor_id_6_hwtcl                         (0),
		.device_id_6_hwtcl                         (1),
		.revision_id_6_hwtcl                       (1),
		.class_code_6_hwtcl                        (0),
		.subsystem_vendor_id_6_hwtcl               (0),
		.subsystem_device_id_6_hwtcl               (0),
		.max_payload_size_6_hwtcl                  (256),
		.extend_tag_field_6_hwtcl                  ("32"),
		.completion_timeout_6_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_6_hwtcl (1),
		.flr_capability_6_hwtcl                    (0),
		.use_aer_6_hwtcl                           (0),
		.ecrc_check_capable_6_hwtcl                (0),
		.ecrc_gen_capable_6_hwtcl                  (0),
		.dll_active_report_support_6_hwtcl         (0),
		.surprise_down_error_support_6_hwtcl       (0),
		.msi_multi_message_capable_6_hwtcl         ("4"),
		.msi_64bit_addressing_capable_6_hwtcl      ("true"),
		.msi_masking_capable_6_hwtcl               ("false"),
		.msi_support_6_hwtcl                       ("true"),
		.enable_function_msix_support_6_hwtcl      (0),
		.msix_table_size_6_hwtcl                   (0),
		.msix_table_offset_6_hwtcl                 ("0"),
		.msix_table_bir_6_hwtcl                    (0),
		.msix_pba_offset_6_hwtcl                   ("0"),
		.msix_pba_bir_6_hwtcl                      (0),
		.interrupt_pin_6_hwtcl                     ("inta"),
		.slot_power_scale_6_hwtcl                  (0),
		.slot_power_limit_6_hwtcl                  (0),
		.slot_number_6_hwtcl                       (0),
		.rx_ei_l0s_6_hwtcl                         (0),
		.endpoint_l0_latency_6_hwtcl               (0),
		.endpoint_l1_latency_6_hwtcl               (0),
		.maximum_current_6_hwtcl                   (0),
		.disable_snoop_packet_6_hwtcl              ("false"),
		.bridge_port_vga_enable_6_hwtcl            ("false"),
		.bridge_port_ssid_support_6_hwtcl          ("false"),
		.ssvid_6_hwtcl                             (0),
		.ssid_6_hwtcl                              (0),
		.porttype_func7_hwtcl                      ("Native endpoint"),
		.bar0_size_mask_7_hwtcl                    (28),
		.bar0_io_space_7_hwtcl                     ("Disabled"),
		.bar0_64bit_mem_space_7_hwtcl              ("Enabled"),
		.bar0_prefetchable_7_hwtcl                 ("Enabled"),
		.bar1_size_mask_7_hwtcl                    (0),
		.bar1_io_space_7_hwtcl                     ("Disabled"),
		.bar1_prefetchable_7_hwtcl                 ("Disabled"),
		.bar2_size_mask_7_hwtcl                    (10),
		.bar2_io_space_7_hwtcl                     ("Disabled"),
		.bar2_64bit_mem_space_7_hwtcl              ("Disabled"),
		.bar2_prefetchable_7_hwtcl                 ("Disabled"),
		.bar3_size_mask_7_hwtcl                    (0),
		.bar3_io_space_7_hwtcl                     ("Disabled"),
		.bar3_prefetchable_7_hwtcl                 ("Disabled"),
		.bar4_size_mask_7_hwtcl                    (0),
		.bar4_io_space_7_hwtcl                     ("Disabled"),
		.bar4_64bit_mem_space_7_hwtcl              ("Disabled"),
		.bar4_prefetchable_7_hwtcl                 ("Disabled"),
		.bar5_size_mask_7_hwtcl                    (0),
		.bar5_io_space_7_hwtcl                     ("Disabled"),
		.bar5_prefetchable_7_hwtcl                 ("Disabled"),
		.expansion_base_address_register_7_hwtcl   (0),
		.vendor_id_7_hwtcl                         (0),
		.device_id_7_hwtcl                         (1),
		.revision_id_7_hwtcl                       (1),
		.class_code_7_hwtcl                        (0),
		.subsystem_vendor_id_7_hwtcl               (0),
		.subsystem_device_id_7_hwtcl               (0),
		.max_payload_size_7_hwtcl                  (256),
		.extend_tag_field_7_hwtcl                  ("32"),
		.completion_timeout_7_hwtcl                ("ABCD"),
		.enable_completion_timeout_disable_7_hwtcl (1),
		.flr_capability_7_hwtcl                    (0),
		.use_aer_7_hwtcl                           (0),
		.ecrc_check_capable_7_hwtcl                (0),
		.ecrc_gen_capable_7_hwtcl                  (0),
		.dll_active_report_support_7_hwtcl         (0),
		.surprise_down_error_support_7_hwtcl       (0),
		.msi_multi_message_capable_7_hwtcl         ("4"),
		.msi_64bit_addressing_capable_7_hwtcl      ("true"),
		.msi_masking_capable_7_hwtcl               ("false"),
		.msi_support_7_hwtcl                       ("true"),
		.enable_function_msix_support_7_hwtcl      (0),
		.msix_table_size_7_hwtcl                   (0),
		.msix_table_offset_7_hwtcl                 ("0"),
		.msix_table_bir_7_hwtcl                    (0),
		.msix_pba_offset_7_hwtcl                   ("0"),
		.msix_pba_bir_7_hwtcl                      (0),
		.interrupt_pin_7_hwtcl                     ("inta"),
		.slot_power_scale_7_hwtcl                  (0),
		.slot_power_limit_7_hwtcl                  (0),
		.slot_number_7_hwtcl                       (0),
		.rx_ei_l0s_7_hwtcl                         (0),
		.endpoint_l0_latency_7_hwtcl               (0),
		.endpoint_l1_latency_7_hwtcl               (0),
		.maximum_current_7_hwtcl                   (0),
		.disable_snoop_packet_7_hwtcl              ("false"),
		.bridge_port_vga_enable_7_hwtcl            ("false"),
		.bridge_port_ssid_support_7_hwtcl          ("false"),
		.ssvid_7_hwtcl                             (0),
		.ssid_7_hwtcl                              (0),
		.rpre_emph_a_val_hwtcl                     (12),
		.rpre_emph_b_val_hwtcl                     (0),
		.rpre_emph_c_val_hwtcl                     (19),
		.rpre_emph_d_val_hwtcl                     (13),
		.rpre_emph_e_val_hwtcl                     (21),
		.rvod_sel_a_val_hwtcl                      (42),
		.rvod_sel_b_val_hwtcl                      (30),
		.rvod_sel_c_val_hwtcl                      (43),
		.rvod_sel_d_val_hwtcl                      (43),
		.rvod_sel_e_val_hwtcl                      (9)
	) dut (
		.npor                   (dut_npor_npor),                                         //               npor.npor
		.pin_perst              (dut_npor_pin_perst),                                    //                   .pin_perst
		.test_in                (dut_hip_ctrl_test_in),                                  //           hip_ctrl.test_in
		.simu_mode_pipe         (dut_hip_ctrl_simu_mode_pipe),                           //                   .simu_mode_pipe
		.pld_clk                (apps_pld_clk_hip_clk),                                  //            pld_clk.clk
		.coreclkout             (dut_coreclkout_hip_clk),                                //     coreclkout_hip.clk
		.refclk                 (dut_refclk_clk),                                        //             refclk.clk
		.rx_in0                 (dut_hip_serial_rx_in0),                                 //         hip_serial.rx_in0
		.rx_in1                 (dut_hip_serial_rx_in1),                                 //                   .rx_in1
		.rx_in2                 (dut_hip_serial_rx_in2),                                 //                   .rx_in2
		.rx_in3                 (dut_hip_serial_rx_in3),                                 //                   .rx_in3
		.tx_out0                (dut_hip_serial_tx_out0),                                //                   .tx_out0
		.tx_out1                (dut_hip_serial_tx_out1),                                //                   .tx_out1
		.tx_out2                (dut_hip_serial_tx_out2),                                //                   .tx_out2
		.tx_out3                (dut_hip_serial_tx_out3),                                //                   .tx_out3
		.rx_st_valid            (dut_rx_st_valid),                                       //              rx_st.valid
		.rx_st_sop              (dut_rx_st_startofpacket),                               //                   .startofpacket
		.rx_st_eop              (dut_rx_st_endofpacket),                                 //                   .endofpacket
		.rx_st_empty            (dut_rx_st_empty),                                       //                   .empty
		.rx_st_ready            (dut_rx_st_ready),                                       //                   .ready
		.rx_st_err              (dut_rx_st_error),                                       //                   .error
		.rx_st_data             (dut_rx_st_data),                                        //                   .data
		.rx_st_bar              (dut_rx_bar_be_rx_st_bar),                               //          rx_bar_be.rx_st_bar
		.rx_st_be               (dut_rx_bar_be_rx_st_be),                                //                   .rx_st_be
		.rx_st_mask             (apps_rx_bar_be_rx_st_mask),                             //                   .rx_st_mask
		.tx_st_valid            (apps_tx_st_valid),                                      //              tx_st.valid
		.tx_st_sop              (apps_tx_st_startofpacket),                              //                   .startofpacket
		.tx_st_eop              (apps_tx_st_endofpacket),                                //                   .endofpacket
		.tx_st_empty            (apps_tx_st_empty),                                      //                   .empty
		.tx_st_ready            (apps_tx_st_ready),                                      //                   .ready
		.tx_st_err              (apps_tx_st_error),                                      //                   .error
		.tx_st_data             (apps_tx_st_data),                                       //                   .data
		.tx_fifo_empty          (dut_tx_fifo_fifo_empty),                                //            tx_fifo.fifo_empty
		.tx_cred_datafccp       (dut_tx_cred_tx_cred_datafccp),                          //            tx_cred.tx_cred_datafccp
		.tx_cred_datafcnp       (dut_tx_cred_tx_cred_datafcnp),                          //                   .tx_cred_datafcnp
		.tx_cred_datafcp        (dut_tx_cred_tx_cred_datafcp),                           //                   .tx_cred_datafcp
		.tx_cred_fchipcons      (dut_tx_cred_tx_cred_fchipcons),                         //                   .tx_cred_fchipcons
		.tx_cred_fcinfinite     (dut_tx_cred_tx_cred_fcinfinite),                        //                   .tx_cred_fcinfinite
		.tx_cred_hdrfccp        (dut_tx_cred_tx_cred_hdrfccp),                           //                   .tx_cred_hdrfccp
		.tx_cred_hdrfcnp        (dut_tx_cred_tx_cred_hdrfcnp),                           //                   .tx_cred_hdrfcnp
		.tx_cred_hdrfcp         (dut_tx_cred_tx_cred_hdrfcp),                            //                   .tx_cred_hdrfcp
		.sim_pipe_pclk_in       (dut_hip_pipe_sim_pipe_pclk_in),                         //           hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate          (dut_hip_pipe_sim_pipe_rate),                            //                   .sim_pipe_rate
		.sim_ltssmstate         (dut_hip_pipe_sim_ltssmstate),                           //                   .sim_ltssmstate
		.eidleinfersel0         (dut_hip_pipe_eidleinfersel0),                           //                   .eidleinfersel0
		.eidleinfersel1         (dut_hip_pipe_eidleinfersel1),                           //                   .eidleinfersel1
		.eidleinfersel2         (dut_hip_pipe_eidleinfersel2),                           //                   .eidleinfersel2
		.eidleinfersel3         (dut_hip_pipe_eidleinfersel3),                           //                   .eidleinfersel3
		.powerdown0             (dut_hip_pipe_powerdown0),                               //                   .powerdown0
		.powerdown1             (dut_hip_pipe_powerdown1),                               //                   .powerdown1
		.powerdown2             (dut_hip_pipe_powerdown2),                               //                   .powerdown2
		.powerdown3             (dut_hip_pipe_powerdown3),                               //                   .powerdown3
		.rxpolarity0            (dut_hip_pipe_rxpolarity0),                              //                   .rxpolarity0
		.rxpolarity1            (dut_hip_pipe_rxpolarity1),                              //                   .rxpolarity1
		.rxpolarity2            (dut_hip_pipe_rxpolarity2),                              //                   .rxpolarity2
		.rxpolarity3            (dut_hip_pipe_rxpolarity3),                              //                   .rxpolarity3
		.txcompl0               (dut_hip_pipe_txcompl0),                                 //                   .txcompl0
		.txcompl1               (dut_hip_pipe_txcompl1),                                 //                   .txcompl1
		.txcompl2               (dut_hip_pipe_txcompl2),                                 //                   .txcompl2
		.txcompl3               (dut_hip_pipe_txcompl3),                                 //                   .txcompl3
		.txdata0                (dut_hip_pipe_txdata0),                                  //                   .txdata0
		.txdata1                (dut_hip_pipe_txdata1),                                  //                   .txdata1
		.txdata2                (dut_hip_pipe_txdata2),                                  //                   .txdata2
		.txdata3                (dut_hip_pipe_txdata3),                                  //                   .txdata3
		.txdatak0               (dut_hip_pipe_txdatak0),                                 //                   .txdatak0
		.txdatak1               (dut_hip_pipe_txdatak1),                                 //                   .txdatak1
		.txdatak2               (dut_hip_pipe_txdatak2),                                 //                   .txdatak2
		.txdatak3               (dut_hip_pipe_txdatak3),                                 //                   .txdatak3
		.txdetectrx0            (dut_hip_pipe_txdetectrx0),                              //                   .txdetectrx0
		.txdetectrx1            (dut_hip_pipe_txdetectrx1),                              //                   .txdetectrx1
		.txdetectrx2            (dut_hip_pipe_txdetectrx2),                              //                   .txdetectrx2
		.txdetectrx3            (dut_hip_pipe_txdetectrx3),                              //                   .txdetectrx3
		.txelecidle0            (dut_hip_pipe_txelecidle0),                              //                   .txelecidle0
		.txelecidle1            (dut_hip_pipe_txelecidle1),                              //                   .txelecidle1
		.txelecidle2            (dut_hip_pipe_txelecidle2),                              //                   .txelecidle2
		.txelecidle3            (dut_hip_pipe_txelecidle3),                              //                   .txelecidle3
		.txswing0               (dut_hip_pipe_txswing0),                                 //                   .txswing0
		.txswing1               (dut_hip_pipe_txswing1),                                 //                   .txswing1
		.txswing2               (dut_hip_pipe_txswing2),                                 //                   .txswing2
		.txswing3               (dut_hip_pipe_txswing3),                                 //                   .txswing3
		.txmargin0              (dut_hip_pipe_txmargin0),                                //                   .txmargin0
		.txmargin1              (dut_hip_pipe_txmargin1),                                //                   .txmargin1
		.txmargin2              (dut_hip_pipe_txmargin2),                                //                   .txmargin2
		.txmargin3              (dut_hip_pipe_txmargin3),                                //                   .txmargin3
		.txdeemph0              (dut_hip_pipe_txdeemph0),                                //                   .txdeemph0
		.txdeemph1              (dut_hip_pipe_txdeemph1),                                //                   .txdeemph1
		.txdeemph2              (dut_hip_pipe_txdeemph2),                                //                   .txdeemph2
		.txdeemph3              (dut_hip_pipe_txdeemph3),                                //                   .txdeemph3
		.phystatus0             (dut_hip_pipe_phystatus0),                               //                   .phystatus0
		.phystatus1             (dut_hip_pipe_phystatus1),                               //                   .phystatus1
		.phystatus2             (dut_hip_pipe_phystatus2),                               //                   .phystatus2
		.phystatus3             (dut_hip_pipe_phystatus3),                               //                   .phystatus3
		.rxdata0                (dut_hip_pipe_rxdata0),                                  //                   .rxdata0
		.rxdata1                (dut_hip_pipe_rxdata1),                                  //                   .rxdata1
		.rxdata2                (dut_hip_pipe_rxdata2),                                  //                   .rxdata2
		.rxdata3                (dut_hip_pipe_rxdata3),                                  //                   .rxdata3
		.rxdatak0               (dut_hip_pipe_rxdatak0),                                 //                   .rxdatak0
		.rxdatak1               (dut_hip_pipe_rxdatak1),                                 //                   .rxdatak1
		.rxdatak2               (dut_hip_pipe_rxdatak2),                                 //                   .rxdatak2
		.rxdatak3               (dut_hip_pipe_rxdatak3),                                 //                   .rxdatak3
		.rxelecidle0            (dut_hip_pipe_rxelecidle0),                              //                   .rxelecidle0
		.rxelecidle1            (dut_hip_pipe_rxelecidle1),                              //                   .rxelecidle1
		.rxelecidle2            (dut_hip_pipe_rxelecidle2),                              //                   .rxelecidle2
		.rxelecidle3            (dut_hip_pipe_rxelecidle3),                              //                   .rxelecidle3
		.rxstatus0              (dut_hip_pipe_rxstatus0),                                //                   .rxstatus0
		.rxstatus1              (dut_hip_pipe_rxstatus1),                                //                   .rxstatus1
		.rxstatus2              (dut_hip_pipe_rxstatus2),                                //                   .rxstatus2
		.rxstatus3              (dut_hip_pipe_rxstatus3),                                //                   .rxstatus3
		.rxvalid0               (dut_hip_pipe_rxvalid0),                                 //                   .rxvalid0
		.rxvalid1               (dut_hip_pipe_rxvalid1),                                 //                   .rxvalid1
		.rxvalid2               (dut_hip_pipe_rxvalid2),                                 //                   .rxvalid2
		.rxvalid3               (dut_hip_pipe_rxvalid3),                                 //                   .rxvalid3
		.reset_status           (dut_hip_rst_reset_status),                              //            hip_rst.reset_status
		.serdes_pll_locked      (dut_hip_rst_serdes_pll_locked),                         //                   .serdes_pll_locked
		.pld_clk_inuse          (dut_hip_rst_pld_clk_inuse),                             //                   .pld_clk_inuse
		.pld_core_ready         (apps_hip_rst_pld_core_ready),                           //                   .pld_core_ready
		.testin_zero            (dut_hip_rst_testin_zero),                               //                   .testin_zero
		.lmi_addr               (apps_lmi_lmi_addr),                                     //                lmi.lmi_addr
		.lmi_din                (apps_lmi_lmi_din),                                      //                   .lmi_din
		.lmi_rden               (apps_lmi_lmi_rden),                                     //                   .lmi_rden
		.lmi_wren               (apps_lmi_lmi_wren),                                     //                   .lmi_wren
		.lmi_ack                (dut_lmi_lmi_ack),                                       //                   .lmi_ack
		.lmi_dout               (dut_lmi_lmi_dout),                                      //                   .lmi_dout
		.pm_auxpwr              (apps_power_mngt_pm_auxpwr),                             //         power_mngt.pm_auxpwr
		.pm_data                (apps_power_mngt_pm_data),                               //                   .pm_data
		.pme_to_cr              (apps_power_mngt_pme_to_cr),                             //                   .pme_to_cr
		.pm_event               (apps_power_mngt_pm_event),                              //                   .pm_event
		.pme_to_sr              (dut_power_mngt_pme_to_sr),                              //                   .pme_to_sr
		.reconfig_to_xcvr       (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr), //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr     (dut_reconfig_from_xcvr_reconfig_from_xcvr),             // reconfig_from_xcvr.reconfig_from_xcvr
		.app_msi_num            (apps_int_msi_app_msi_num),                              //            int_msi.app_msi_num
		.app_msi_req            (apps_int_msi_app_msi_req),                              //                   .app_msi_req
		.app_msi_tc             (apps_int_msi_app_msi_tc),                               //                   .app_msi_tc
		.app_msi_ack            (dut_int_msi_app_msi_ack),                               //                   .app_msi_ack
		.app_int_sts_vec        (apps_int_msi_app_int_sts),                              //                   .app_int_sts
		.tl_hpg_ctrl_er         (pcie_av_hip_de_hip_status_0_config_tl_hip_hpg_ctrler),  //          config_tl.hpg_ctrler
		.tl_cfg_ctl             (dut_config_tl_tl_cfg_ctl),                              //                   .tl_cfg_ctl
		.cpl_err                (pcie_av_hip_de_hip_status_0_config_tl_hip_cpl_err),     //                   .cpl_err
		.tl_cfg_add             (dut_config_tl_tl_cfg_add),                              //                   .tl_cfg_add
		.tl_cfg_ctl_wr          (dut_config_tl_tl_cfg_ctl_wr),                           //                   .tl_cfg_ctl_wr
		.tl_cfg_sts_wr          (dut_config_tl_tl_cfg_sts_wr),                           //                   .tl_cfg_sts_wr
		.tl_cfg_sts             (dut_config_tl_tl_cfg_sts),                              //                   .tl_cfg_sts
		.cpl_pending            (pcie_av_hip_de_hip_status_0_config_tl_hip_cpl_pending), //                   .cpl_pending
		.derr_cor_ext_rcv0      (dut_hip_status_derr_cor_ext_rcv),                       //         hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl       (dut_hip_status_derr_cor_ext_rpl),                       //                   .derr_cor_ext_rpl
		.derr_rpl               (dut_hip_status_derr_rpl),                               //                   .derr_rpl
		.dlup_exit              (dut_hip_status_dlup_exit),                              //                   .dlup_exit
		.dl_ltssm               (dut_hip_status_ltssmstate),                             //                   .ltssmstate
		.ev128ns                (dut_hip_status_ev128ns),                                //                   .ev128ns
		.ev1us                  (dut_hip_status_ev1us),                                  //                   .ev1us
		.hotrst_exit            (dut_hip_status_hotrst_exit),                            //                   .hotrst_exit
		.int_status             (dut_hip_status_int_status),                             //                   .int_status
		.l2_exit                (dut_hip_status_l2_exit),                                //                   .l2_exit
		.lane_act               (dut_hip_status_lane_act),                               //                   .lane_act
		.ko_cpl_spc_header      (dut_hip_status_ko_cpl_spc_header),                      //                   .ko_cpl_spc_header
		.ko_cpl_spc_data        (dut_hip_status_ko_cpl_spc_data),                        //                   .ko_cpl_spc_data
		.dl_current_speed       (dut_hip_currentspeed_currentspeed),                     //   hip_currentspeed.currentspeed
		.rx_in4                 (1'b0),                                                  //        (terminated)
		.rx_in5                 (1'b0),                                                  //        (terminated)
		.rx_in6                 (1'b0),                                                  //        (terminated)
		.rx_in7                 (1'b0),                                                  //        (terminated)
		.tx_out4                (),                                                      //        (terminated)
		.tx_out5                (),                                                      //        (terminated)
		.tx_out6                (),                                                      //        (terminated)
		.tx_out7                (),                                                      //        (terminated)
		.rx_fifo_empty          (),                                                      //        (terminated)
		.rx_fifo_full           (),                                                      //        (terminated)
		.rx_bar_dec_func_num    (),                                                      //        (terminated)
		.tx_fifo_full           (),                                                      //        (terminated)
		.tx_fifo_rdp            (),                                                      //        (terminated)
		.tx_fifo_wrp            (),                                                      //        (terminated)
		.eidleinfersel4         (),                                                      //        (terminated)
		.eidleinfersel5         (),                                                      //        (terminated)
		.eidleinfersel6         (),                                                      //        (terminated)
		.eidleinfersel7         (),                                                      //        (terminated)
		.powerdown4             (),                                                      //        (terminated)
		.powerdown5             (),                                                      //        (terminated)
		.powerdown6             (),                                                      //        (terminated)
		.powerdown7             (),                                                      //        (terminated)
		.rxpolarity4            (),                                                      //        (terminated)
		.rxpolarity5            (),                                                      //        (terminated)
		.rxpolarity6            (),                                                      //        (terminated)
		.rxpolarity7            (),                                                      //        (terminated)
		.txcompl4               (),                                                      //        (terminated)
		.txcompl5               (),                                                      //        (terminated)
		.txcompl6               (),                                                      //        (terminated)
		.txcompl7               (),                                                      //        (terminated)
		.txdata4                (),                                                      //        (terminated)
		.txdata5                (),                                                      //        (terminated)
		.txdata6                (),                                                      //        (terminated)
		.txdata7                (),                                                      //        (terminated)
		.txdatak4               (),                                                      //        (terminated)
		.txdatak5               (),                                                      //        (terminated)
		.txdatak6               (),                                                      //        (terminated)
		.txdatak7               (),                                                      //        (terminated)
		.txdetectrx4            (),                                                      //        (terminated)
		.txdetectrx5            (),                                                      //        (terminated)
		.txdetectrx6            (),                                                      //        (terminated)
		.txdetectrx7            (),                                                      //        (terminated)
		.txelecidle4            (),                                                      //        (terminated)
		.txelecidle5            (),                                                      //        (terminated)
		.txelecidle6            (),                                                      //        (terminated)
		.txelecidle7            (),                                                      //        (terminated)
		.txswing4               (),                                                      //        (terminated)
		.txswing5               (),                                                      //        (terminated)
		.txswing6               (),                                                      //        (terminated)
		.txswing7               (),                                                      //        (terminated)
		.txmargin4              (),                                                      //        (terminated)
		.txmargin5              (),                                                      //        (terminated)
		.txmargin6              (),                                                      //        (terminated)
		.txmargin7              (),                                                      //        (terminated)
		.txdeemph4              (),                                                      //        (terminated)
		.txdeemph5              (),                                                      //        (terminated)
		.txdeemph6              (),                                                      //        (terminated)
		.txdeemph7              (),                                                      //        (terminated)
		.phystatus4             (1'b0),                                                  //        (terminated)
		.phystatus5             (1'b0),                                                  //        (terminated)
		.phystatus6             (1'b0),                                                  //        (terminated)
		.phystatus7             (1'b0),                                                  //        (terminated)
		.rxdata4                (8'b00000000),                                           //        (terminated)
		.rxdata5                (8'b00000000),                                           //        (terminated)
		.rxdata6                (8'b00000000),                                           //        (terminated)
		.rxdata7                (8'b00000000),                                           //        (terminated)
		.rxdatak4               (1'b0),                                                  //        (terminated)
		.rxdatak5               (1'b0),                                                  //        (terminated)
		.rxdatak6               (1'b0),                                                  //        (terminated)
		.rxdatak7               (1'b0),                                                  //        (terminated)
		.rxelecidle4            (1'b0),                                                  //        (terminated)
		.rxelecidle5            (1'b0),                                                  //        (terminated)
		.rxelecidle6            (1'b0),                                                  //        (terminated)
		.rxelecidle7            (1'b0),                                                  //        (terminated)
		.rxstatus4              (3'b000),                                                //        (terminated)
		.rxstatus5              (3'b000),                                                //        (terminated)
		.rxstatus6              (3'b000),                                                //        (terminated)
		.rxstatus7              (3'b000),                                                //        (terminated)
		.rxvalid4               (1'b0),                                                  //        (terminated)
		.rxvalid5               (1'b0),                                                  //        (terminated)
		.rxvalid6               (1'b0),                                                  //        (terminated)
		.rxvalid7               (1'b0),                                                  //        (terminated)
		.sim_pipe_pclk_out      (),                                                      //        (terminated)
		.pm_event_func          (3'b000),                                                //        (terminated)
		.hip_reconfig_clk       (1'b0),                                                  //        (terminated)
		.hip_reconfig_rst_n     (1'b0),                                                  //        (terminated)
		.hip_reconfig_address   (10'b0000000000),                                        //        (terminated)
		.hip_reconfig_byte_en   (2'b00),                                                 //        (terminated)
		.hip_reconfig_read      (1'b0),                                                  //        (terminated)
		.hip_reconfig_readdata  (),                                                      //        (terminated)
		.hip_reconfig_write     (1'b0),                                                  //        (terminated)
		.hip_reconfig_writedata (16'b0000000000000000),                                  //        (terminated)
		.ser_shift_load         (1'b0),                                                  //        (terminated)
		.interface_sel          (1'b0),                                                  //        (terminated)
		.app_msi_func           (3'b000),                                                //        (terminated)
		.serr_out               (),                                                      //        (terminated)
		.aer_msi_num            (5'b00000),                                              //        (terminated)
		.pex_msi_num            (5'b00000),                                              //        (terminated)
		.cpl_err_func           (3'b000)                                                 //        (terminated)
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Arria V"),
		.number_of_reconfig_interfaces (5),
		.enable_offset                 (1),
		.enable_lc                     (0),
		.enable_dcd                    (1),
		.enable_dcd_power_up           (0),
		.enable_analog                 (0),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),       //      reconfig_busy.reconfig_busy
		.cal_busy_in               (pcie_reconfig_driver_0_cal_busy_in_cal_busy_in),        //        cal_busy_in.cal_busy_in
		.mgmt_clk_clk              (clk_clk),                                               //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                        //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),          //      reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),             //                   .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),         //                   .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest),      //                   .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),            //                   .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),        //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr), //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (dut_reconfig_from_xcvr_reconfig_from_xcvr),             // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                      //        (terminated)
		.rx_cal_busy               (),                                                      //        (terminated)
		.reconfig_mif_address      (),                                                      //        (terminated)
		.reconfig_mif_read         (),                                                      //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                  //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                   //        (terminated)
	);

	altpcie_av_hip_ast_hip_status_bridge pcie_av_hip_de_hip_status_0 (
		.pld_clk                   (apps_pld_clk_hip_clk),                                          //           pld_clk.clk
		.export_pld_clk            (pld_clk_clk),                                                   //    export_pld_clk.clk
		.to_hip_derr_cor_ext_rcv   (dut_hip_status_derr_cor_ext_rcv),                               //    hip_status_hip.derr_cor_ext_rcv
		.to_hip_derr_cor_ext_rpl   (dut_hip_status_derr_cor_ext_rpl),                               //                  .derr_cor_ext_rpl
		.to_hip_derr_rpl           (dut_hip_status_derr_rpl),                                       //                  .derr_rpl
		.to_hip_dlup_exit          (dut_hip_status_dlup_exit),                                      //                  .dlup_exit
		.to_hip_ev128ns            (dut_hip_status_ev128ns),                                        //                  .ev128ns
		.to_hip_ev1us              (dut_hip_status_ev1us),                                          //                  .ev1us
		.to_hip_hotrst_exit        (dut_hip_status_hotrst_exit),                                    //                  .hotrst_exit
		.to_hip_int_status         (dut_hip_status_int_status),                                     //                  .int_status
		.to_hip_l2_exit            (dut_hip_status_l2_exit),                                        //                  .l2_exit
		.to_hip_lane_act           (dut_hip_status_lane_act),                                       //                  .lane_act
		.to_hip_ltssmstate         (dut_hip_status_ltssmstate),                                     //                  .ltssmstate
		.to_hip_ko_cpl_spc_header  (dut_hip_status_ko_cpl_spc_header),                              //                  .ko_cpl_spc_header
		.to_hip_ko_cpl_spc_data    (dut_hip_status_ko_cpl_spc_data),                                //                  .ko_cpl_spc_data
		.to_apps_derr_cor_ext_rcv  (pcie_av_hip_de_hip_status_0_hip_status_apps_derr_cor_ext_rcv),  //   hip_status_apps.derr_cor_ext_rcv
		.to_apps_derr_cor_ext_rpl  (pcie_av_hip_de_hip_status_0_hip_status_apps_derr_cor_ext_rpl),  //                  .derr_cor_ext_rpl
		.to_apps_derr_rpl          (pcie_av_hip_de_hip_status_0_hip_status_apps_derr_rpl),          //                  .derr_rpl
		.to_apps_dlup_exit         (pcie_av_hip_de_hip_status_0_hip_status_apps_dlup_exit),         //                  .dlup_exit
		.to_apps_ev128ns           (pcie_av_hip_de_hip_status_0_hip_status_apps_ev128ns),           //                  .ev128ns
		.to_apps_ev1us             (pcie_av_hip_de_hip_status_0_hip_status_apps_ev1us),             //                  .ev1us
		.to_apps_hotrst_exit       (pcie_av_hip_de_hip_status_0_hip_status_apps_hotrst_exit),       //                  .hotrst_exit
		.to_apps_int_status        (pcie_av_hip_de_hip_status_0_hip_status_apps_int_status),        //                  .int_status
		.to_apps_l2_exit           (pcie_av_hip_de_hip_status_0_hip_status_apps_l2_exit),           //                  .l2_exit
		.to_apps_lane_act          (pcie_av_hip_de_hip_status_0_hip_status_apps_lane_act),          //                  .lane_act
		.to_apps_ltssmstate        (pcie_av_hip_de_hip_status_0_hip_status_apps_ltssmstate),        //                  .ltssmstate
		.to_apps_ko_cpl_spc_header (pcie_av_hip_de_hip_status_0_hip_status_apps_ko_cpl_spc_header), //                  .ko_cpl_spc_header
		.to_apps_ko_cpl_spc_data   (pcie_av_hip_de_hip_status_0_hip_status_apps_ko_cpl_spc_data),   //                  .ko_cpl_spc_data
		.export_derr_cor_ext_rcv   (status_hip_derr_cor_ext_rcv),                                   // hip_status_export.derr_cor_ext_rcv
		.export_derr_cor_ext_rpl   (status_hip_derr_cor_ext_rpl),                                   //                  .derr_cor_ext_rpl
		.export_derr_rpl           (status_hip_derr_rpl),                                           //                  .derr_rpl
		.export_dlup_exit          (status_hip_dlup_exit),                                          //                  .dlup_exit
		.export_ev128ns            (status_hip_ev128ns),                                            //                  .ev128ns
		.export_ev1us              (status_hip_ev1us),                                              //                  .ev1us
		.export_hotrst_exit        (status_hip_hotrst_exit),                                        //                  .hotrst_exit
		.export_int_status         (status_hip_int_status),                                         //                  .int_status
		.export_l2_exit            (status_hip_l2_exit),                                            //                  .l2_exit
		.export_lane_act           (status_hip_lane_act),                                           //                  .lane_act
		.export_ltssmstate         (status_hip_ltssmstate),                                         //                  .ltssmstate
		.export_ko_cpl_spc_header  (status_hip_ko_cpl_spc_header),                                  //                  .ko_cpl_spc_header
		.export_ko_cpl_spc_data    (status_hip_ko_cpl_spc_data),                                    //                  .ko_cpl_spc_data
		.to_hip_hpg_ctrler         (pcie_av_hip_de_hip_status_0_config_tl_hip_hpg_ctrler),          //     config_tl_hip.hpg_ctrler
		.to_hip_tl_cfg_add         (dut_config_tl_tl_cfg_add),                                      //                  .tl_cfg_add
		.to_hip_tl_cfg_ctl         (dut_config_tl_tl_cfg_ctl),                                      //                  .tl_cfg_ctl
		.to_hip_tl_cfg_sts         (dut_config_tl_tl_cfg_sts),                                      //                  .tl_cfg_sts
		.to_hip_tl_cfg_ctl_wr      (dut_config_tl_tl_cfg_ctl_wr),                                   //                  .tl_cfg_ctl_wr
		.to_hip_tl_cfg_sts_wr      (dut_config_tl_tl_cfg_sts_wr),                                   //                  .tl_cfg_sts_wr
		.to_hip_cpl_err            (pcie_av_hip_de_hip_status_0_config_tl_hip_cpl_err),             //                  .cpl_err
		.to_hip_cpl_pending        (pcie_av_hip_de_hip_status_0_config_tl_hip_cpl_pending),         //                  .cpl_pending
		.to_apps_hpg_ctrler        (apps_config_tl_hpg_ctrler),                                     //    config_tl_apps.hpg_ctrler
		.to_apps_tl_cfg_add        (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_add),         //                  .tl_cfg_add
		.to_apps_tl_cfg_ctl        (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_ctl),         //                  .tl_cfg_ctl
		.to_apps_tl_cfg_sts        (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_sts),         //                  .tl_cfg_sts
		.to_apps_tl_cfg_ctl_wr     (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_ctl_wr),      //                  .tl_cfg_ctl_wr
		.to_apps_tl_cfg_sts_wr     (pcie_av_hip_de_hip_status_0_config_tl_apps_tl_cfg_sts_wr),      //                  .tl_cfg_sts_wr
		.to_apps_cpl_err           (apps_config_tl_cpl_err),                                        //                  .cpl_err
		.to_apps_cpl_pending       (apps_config_tl_cpl_pending),                                    //                  .cpl_pending
		.export_tl_cfg_add         (tl_cfg_tl_cfg_add),                                             //  config_tl_export.tl_cfg_add
		.export_tl_cfg_ctl         (tl_cfg_tl_cfg_ctl),                                             //                  .tl_cfg_ctl
		.export_tl_cfg_sts         (tl_cfg_tl_cfg_sts)                                              //                  .tl_cfg_sts
	);

	altpcie_reconfig_driver #(
		.INTENDED_DEVICE_FAMILY        ("Arria V"),
		.gen123_lane_rate_mode_hwtcl   ("Gen2 (5.0 Gbps)"),
		.number_of_reconfig_interfaces (5)
	) pcie_reconfig_driver_0 (
		.reconfig_xcvr_clk         (clk_clk),                                          // reconfig_xcvr_clk.clk
		.reconfig_xcvr_rst         (rst_controller_reset_out_reset),                   // reconfig_xcvr_rst.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),     //     reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),        //                  .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),    //                  .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest), //                  .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),       //                  .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),   //                  .writedata
		.currentspeed              (dut_hip_currentspeed_currentspeed),                //  hip_currentspeed.currentspeed
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),  //     reconfig_busy.reconfig_busy
		.pld_clk                   (apps_pld_clk_hip_clk),                             //           pld_clk.clk
		.cal_busy_in               (pcie_reconfig_driver_0_cal_busy_in_cal_busy_in),   //       cal_busy_in.cal_busy_in
		.derr_cor_ext_rcv_drv      (apps_hip_status_drv_derr_cor_ext_rcv),             //    hip_status_drv.derr_cor_ext_rcv
		.derr_cor_ext_rpl_drv      (apps_hip_status_drv_derr_cor_ext_rpl),             //                  .derr_cor_ext_rpl
		.derr_rpl_drv              (apps_hip_status_drv_derr_rpl),                     //                  .derr_rpl
		.dlup_exit_drv             (apps_hip_status_drv_dlup_exit),                    //                  .dlup_exit
		.ev128ns_drv               (apps_hip_status_drv_ev128ns),                      //                  .ev128ns
		.ev1us_drv                 (apps_hip_status_drv_ev1us),                        //                  .ev1us
		.hotrst_exit_drv           (apps_hip_status_drv_hotrst_exit),                  //                  .hotrst_exit
		.int_status_drv            (apps_hip_status_drv_int_status),                   //                  .int_status
		.l2_exit_drv               (apps_hip_status_drv_l2_exit),                      //                  .l2_exit
		.lane_act_drv              (apps_hip_status_drv_lane_act),                     //                  .lane_act
		.ltssmstate_drv            (apps_hip_status_drv_ltssmstate),                   //                  .ltssmstate
		.ko_cpl_spc_header_drv     (apps_hip_status_drv_ko_cpl_spc_header),            //                  .ko_cpl_spc_header
		.ko_cpl_spc_data_drv       (apps_hip_status_drv_ko_cpl_spc_data),              //                  .ko_cpl_spc_data
		.dlup_drv                  (1'b0),                                             //       (terminated)
		.rx_par_err_drv            (1'b0),                                             //       (terminated)
		.tx_par_err_drv            (2'b00),                                            //       (terminated)
		.cfg_par_err_drv           (1'b0)                                              //       (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
