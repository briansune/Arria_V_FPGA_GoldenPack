// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:28 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XO4dLKE+ItKSZrsBN1AO6HMPS8+uncxH1CpdboqT6lVHjNZNtXCeBjpVBDqSpbYk
tl7jO4v/WpV6BohvT4qs+X7VCC11fDMLIPXyyfGXMh60K22tbHd66TIJFAREtpMZ
Obtp0SpBFJDKgDN1EzyoYZrfdxWiGsgnSZih2T5O+/c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18352)
pRuvsvntvxuSoM/o2qbs1Y8iQKBc9qju+fW4Twb8nVhOPVXmfd+vMg6sTk86hNvL
Chlpb9lynZ9rNR70dPP5BpisDjDmf0mu4xHXEO/em01/qs8RuV447WYC4JcF7min
yj09OCk1eOtaUt81r8HsOO/wxoFqu8rnkzH8Xn5CB7aSY0gmc6IuG1IdKod8/Hgn
NQSwWK2QKhdHZsTfw2fEgBmYL5zH0BZ3dcFpJnaIohdWqiXO+9YcPOhQ6pygACUM
AicwwBVjhB40KdWwlNYFdbwDjGJPW+6AulS2gmhyOU1k/E99B1P2tb9FPsKSRzFw
SfbLgt2EkA+WXcCyDS2Fv/kaehvupIO4I+ouN7igvSlrVA90gZwky2YhRFY0vsZQ
qqQyWr+20YV770YlXQvpEQe5O4cgkhqUbrql+Q6ax7D9P7B8GaTNkehmLgx221BT
Qhhj+GtvZKAAwR2Unrn78hJIYF2w4olKK6yqJPiZWzFj+GFv8EPHCCLY94coqYN2
ooBVzadhWZL9/0PksqOkZijhPsu+c7QngwbWqutt4/eG9eTnxJ7oKzIG7MTPO4Ot
S45BpstUnZy+kRsxxeeKaqKytGyFQbe7JmM4dwXOj6FN998rEn5q36SK/oNQLJJu
+UHRtNrBLZ9qN/0YrFSeBwHDf51nJ+LXY4WUVTZ7yn5DEs/gvxlozNh/UCMwTU1l
L0hl/VVOuM9itzu708k+LGuU9auRtuw4du6rwLlp1iHKI2tI8xuseNf+BL+wSSlO
029V3PY5sT0tmH4X5swEYOVnhwgMCeHVxomLaBCAO4VL/T0BuR3X9Rc3WBsqWW0B
W3JSkyib4Xssi1tZJoZXINgSaQkr4LYAu2SV1r5W81YreJ4quGeaglPpK3y/cOIH
yS0SxRWQ+a/q1nZZzXkyC4IWAJY/p3MEHKmSn9NPsv9ZC0YfLWiqUtm1yvbWCfB1
11nDs09OROEyvoU56ajjWP7NpZWDj8FntvxymL/I0fdVRgNoP2//m7MttNYcp4kI
+VUOjUyyvTCgaQKNhf7AAi8QdAzwzrKczPo6A0efQCcEI3Txp6fnl07qkPqJ8lHD
w+HesGcLneQuYlKl7bR9YgQ9aqGK83bxb8tNA8RMVqiU3bnKB3lnOO/3PTbBoe/o
Y6MVKj+UbacsrT85OSemFgtgCgeOL1w0KriEIRy37ngp0aAVl1uGO4wBYbRB/ueh
hHOIvuoMEFdZ5XqNpUh22QzaNaYrZ7nf3XvfoHN9B1QjMGLBrs1c9o/tGdxXr5DH
b9S2EnlNNbq81l4gJoSyaoKddiEAGyCBnfJkcyElh/JoSO9f0oTZyD9Sdb/ACqja
xekVxNoQPvQX0Q9Qbzpdcoku5rKUq/rbxBtLjR2yTJ3IAe+DJPPLGwfjeRm+BCQp
oe6yN5eywEXu0SR9isZmnj+gq4Dl9zZsDjE1eTVz6rAHWKcY3Sj3LL9apZZ+yk0Q
Em2uuBq3NGeek7JrJOZfXHNAeYqLGefTCyF8o+8TvjQq0/PDk4sXFifeiUAPDQl5
r58W2HUz8TDpC84Y9k+wO1GSpjfF6FqtlYV+vub9p9l3Iuu2QzriRgOZH0l9EPao
xz11abtrfEC0/R4z9aUeau5li0Nl0dPj6d9SKAvU+Gk24cVNiCZikUpqz2SnOSX+
syly3fybvQtKFdxLUILL1uUdQ2tmk+ehFGfplH7A/7pvNMPTUADlaOW8VcmxPhCM
JJHVJfSEERZaVd0a/eAjVRmQg6LwDlxnWfzoqc4aVe3ILuo/NRM79B46zk9CA9xc
UF8nHI0M9pRqZSOvgBNCn00+vJ2EGVjQIC75IaoRYAKK5FxVClhLn9TBPDw9k5kL
GY2G9Ndx4Eap3T4dZJmmbzshef0+uUn2H8tilBFUlSOTWbducMX89gVyDEInabBK
ubWdre0KMiolcp9qFSelwqHkZj1lt+ks0za7DMHXEWz9X2jkTJkxeaULqwt2ky70
yA02KuYq5C/VBgwteakaa+mOXlx+qoHPAGPbznA9hue+FhGwy7w1v31v4LGpZg+C
cVpAXYwW0OPnSvULokUTWNg7p3L5uMvS+D56+3hVLt+if2UIlMJuP0v9ouO2vPE1
mNy/T9HDf68xUiEjQIKXlAEjMidJS1r6LNosBx8JJIfvXw/8izYbdZSrWMYv+Tqo
SWgxusaK/FGHfOnEF5xQsKmG2rOeDGqwf4NbJx4t3JHLqj7Fxz6WV294aG71j3sm
8t9KS3RaKAe6ezdSmrFeNV8mndF6vF/8mFwuSRt71vjTc3DSXyfoO8PfuGkfaPmV
SqKxGvUtlSF81/wQKuCx1rtYTEX4wOcWaVQZU7Hp0ajoRZcMpUgTea8z1qWN8bRh
/MqXGlK9a5XImEziRyJ3ab5o3PPvFDVXy+q0bGk4SN8IPIuDdI0VMgGkyGBlCP7W
8dKpVoOZR8UsMOGp2Qxzv/TbFNoPZiUAVAqvXg9YYya9fyRuawgGd6XEevXHIYCF
elZgJ27jwC1/C0RMu7K4jVqZt8apWFuV5eI6dkzOXT+iSVNU3QDUnJcDfpA0f9dF
l7161eaVJhF6vepwgw4cGRNT3vPFOj2NTSgQGav+qQndDW42QypTIS65DJFl8D8x
Qleof1ikVANXytsFt0CljicYwKHk0vmNl3QSriR8kTqdS6fK2PehjSo8F6zKGDth
4KErrFyCPYwSySXFreEzsiIxC0Ii1e5gyCCrVUHoQ48PKgNdoettjy0SJ87t/T6f
neEuIPeoayf+20N9u7GUj2g7w2zzsnjAIFRhACwDRmNvswTewCoYyiREOWsWzbfF
QNNYVCSVdqRRensGqNl/A9YkLcIZSL4OMHTzCMMqZrFHjUsaGQ7mme+t13SPPWFJ
qQtvM4aIGOn4NyQy60r5x3Mv9VEBm/serv2i3BXza/bHX8McVvXF3HuqJhWuEqv/
7YwrAkK1iSZEPGMVznwh2xR2bI/Mzthu90cfufRKsZLBah8CMLl2f5xMCjxPXmiU
GHXdDowfwyhvK+qppGkjnUdUkctSoKeehuT27e1Sp+SWpaZ5HXE0ytSoEaF/ca8i
gQ8vxs9OwDZGjhPh2Y9pKXYLVR24WWV9ClabtwEhw3bqZRBWe1gpD1Pg5UjrRygo
aExD1K/bpT5ank8GZXPKxnx+YMWSr5O82aB0pdzlEKoLMyWKP4EPPvT0cBcGgw0Z
VT4gjeojGhlmNZlDGODynYLrdtS7A5HDA5AMh8rYorT/aQggvTsTcWZZeIcIeU6k
DkpHCa4qcgINTKOO9u8i5BoKtK8WTX0GN4Ed8m5po+qRKZ9zaCC/ru9UfrnvwwyW
cVO/hL65+YLAwstKhQTJKPDyTv8Qo2YvVyA/ylo0zjjiQb0iW7FRDnd14uMtP6V3
ZlKeJpDcMDnFHPY8dTTJ3/MgJ7uTbN/KyCq/y/GBHdrYNVclTDJlgX8N132LDY3y
8av0tD2sfQs/ptl4FkDsW1HD8e0wdoQsoxaaETerm1Y8CKb+bruEWRtqaBdsV3cn
NpWMp+hjanup1JvseN9hCpkFqVvvIOCIpPek+J/yAua4n4rNN3s/0ckORXRrmMZv
xNsxQjFQgtYnQ1al5hh5alVdWwkYF4gJelRNe4z+k5O0NyV5FdIv+3tN3imMnNDX
JCvK3txuIFZe5vAYNjmojc1wXy9yNwNY+aBOgId2DVEfRBseOhfeLTUBF6pWjEjy
rIcQr5eo9A/va9GFztZuzdP0WmyQP9MetI+VkmOTLnvHSnnTNRsjjIiIdMlE8Ybi
pKZn4XuAay9x0UC3xA9x+x9m44gSSY+AEL1k65lzMAHz6fVUNtWpTE22gqFY3qMK
WAOGix9AoivK5c9uhgJR94Hf7OTY55eEhqNe816T72RS8s/J6ntJboESlR/6wqbp
iAxvRbzwMsBoBxpEloGJnjU/9jRqQy3qLJB0wM2lYKMNtSkmoXK59mP5lkpPkZnF
/Oh4yuua8ktdT4NwSXn1A5qdNkX9f02oGp2EIiwVA525BlOBa1gXTlo3jCIoyBhY
2j3kcOFJ1iz+p/2Ew5rOGs7eAxtfgG6XowecAugaEAV6nh3bXitKc95GVGTmo3BV
wuRCqiloY/eAFuPnjJeBv3rmXn93x6iYef+kkJFYR6FWMri9Lle7DP4bXe99tYR1
XFgukAHODeoBar2hZY7p4MwSeb4C4LZTPW8E4GmSFIi0WqLF3JfpD9Vdk8zLo0y1
tj8HJpkKAYS7g9JJHzW9YeIaweFYNonOZwny9ow1fBkw3iKRrPmo0OCwmi/LDOsg
C1kzXb/JBEW7gTLokO5QyqBUZKyWNfxijsaKUEfyrzhiwjqI6ZadshyMCP+MvKmG
/A4ZhcSBNvQ2j82YVuJZz5DO9dM3tyi4nb2uOQ9xZ/UIHLW0+qIp0V76ruaw5CSj
L4FGUJuowgB3COca1sAKoj0PyJdD/z07tAIyq3QQFxKg7pcLmvF05i7yNA61Qiky
1B5xMtLg/bkvxdt3VZhGigo/uLXjkcEqRQPY+8O/KzwW5zotj9Z0ykUBSGrih5OK
f4IRoZLVrNR7dnkX8W1tu2nXMzW3xsqVuAN2oJj8+p48+l3wyJhlqvAeEhKe6Y2g
TN00QRuuY7jJRiaE+kKR6q5TnqVxP070SmnfV0cpwmTILaARdP82In/leveL4MuA
sr7G+LKZIhPYXfjpu2JDfvF0i1baA6VUQFRL54DxJiA6bST+FQ35Ypp3G2vl+dt1
BIlJh7a3FjCvA3el1HoaQy5jURqrPi5MgECxGwslwSv9aYhSZUOWZ1OxQrva72ZE
2a09ZgI1Cj7iKX6hn2SmD3YZw2Qzp7npVeb4iHSjWD1Hz2MZM9K6296Lp3yr+IPB
o6g6GB3jrxxSs4FqiDXnjH4I6wUwwB/N0JYZwP0JbhoeZ+5SW4yd6pr2s0+27ypx
gpMGI0dKF7ixDfyGoFFy7X+C6CUxZ3GGY4DHvaN9BKBjBffBe2WSHdCZJpofFfqc
/4pkKBUY/rbw0W7CBZzPM+WQYZKFlMXVA67G4EjY7OGGqdWIncvy2vP8NLTv+hrH
S3u8DUBOsEYStll/E+nsBJVHY1qbkykKIiUZhdPNNrQ1pjhGqFplsjONhwn+yH8p
GUbzHRMLhRW2TK7vHboB9qS5qFjOjqPRA6BywwcWfcHQsIMM5YF8rVvA48dZ4ony
v44f4ecCEqDf9ugmhffop/0v+RRh8Xkqe2IVR+2YsQQBxJMA0zZyKGX2bJnUMPHM
I6nbmY7YG91Jeryytm2uycFQCd7Qt9XKaCfTFGV6mA6hVmQF7ArT2CxNlNrKD5kO
PoD1khLV2Z+DAwfu87l2sRxP52DKSYkGvOhha/K0LiI9QjnWa+tVEUrRBFJN0sIf
QnVsmMTu4UQhNHQvBXGhHwli0grNoTDpaWS6APYJbXI0F1Vpgux3okeeQw+FxWRY
Q30JgInh70jnVdTVRslfATzqFjuQ/uaAMADid21EWtgCixQ7E8XAaX5IXMAozfsq
TAGdBrgLv+jSivybWETxEuA6AMyTr9Z1xtMAejpzpzPTi/D/RtlE32IAiTiuJohV
fn+kdhgd2FnGnELd5sTr4ovghtXtMxh4hSQPiX8Dgi0lMqssNaMa2vsL4Ud9EeaB
CHjb+6QY4wbeBfoBqYoBJ2uf6Tqha09jpv2HyAp9JiC3tvp7Ok0dC2igWh60BsP9
bCYMQVjaIxtvi8T7nzQd9Cfjr2xGUmf5h3X2Oh4s8kJmX/bvSehkf7UAf8zIJail
GZEGIBl4TBqAh0vNyM5Xg+BkPsp/XYkKaMXYW2NuUV8nTKZ+QBn5eBwqQWvB5pFi
vetYuhcKO19a3tTAOfrRJRMP8PfHRfmlxhEIdf0DvlFdLOusMD1vdr6znUuSaeoR
0O3k4OTzGoDLDwWHh1zF0quycBSqW5764xy0z3Wc0N7up0O2Ir3uwIJhiwc9FD8I
U7OAcrg9sVaRdGVVjnls9SuZ1mOSO/9oi5s55oBSVbiRSXEzM98pjrcoQ+luo6qJ
PjVHDEFGI9cnz+nqSft3NzwXho6IaFNXa9k4q2Ez9BgpBGX6eiohW6EG3eAORDX0
GUyaWR0yaZmOap8/y3gHacjS3Q6RUXowuPbrhSQCZC4pb2V/U4ceVAGCaz/ZAy/d
3Y/CPJzW/wVuJV1DWVmmugLuJRGjUYKfkwHBMeE09aqa5Pcqd/2qEi/STarnNF0Q
n1gz57AveYYRUOSsiTS3pLwx6qdDlU7MBer4XLnCXN9k65iHX5sJ4rVgkQerJVHS
GAzV+TAyYLOx1I876DkH9HZau++L402Y7QHA3ICtGIVw99sPH9yYdwMEuwuv4Lp8
DDsZuD8zwgzDF80yRuZw6LQla8711AToFTjadTyiSkVbOeUgvlNaxR4AVLIckk8/
y60VdNLnM5X9ltrvcFZNiUMFDmmRwBbgGECXsTxWY+NoM1Ud8aNWotbnDXmevLfK
alfG4lkzNDbZVTFrLv2lsLTyq4Z+9W2ppI0vjpvNggoQNSv+838f6zTBY5NGdzL/
qEkqNQ3k/6GZ59KGJtlu54CgbH1QPis5QW/Iyi8SSjalLdLx55QFgn0AQee5SjdS
FdkAS1ql/HROTkH5VoKY4oFgz2PPplAsMQMyDwonTv7pBZmGDLr/n2MlyB+XxryV
cI1f4ekO/gdk2a/S8NkWXt4katsJ6neVdP5aAX9n6KZk5dlzgaqbgKC8hBkKur/x
OOkFeepTxq5Hladmd/1NqLWK8oLdx4F63veEYNw3n9u4gxZUHqR9wRHulMl8ps9g
6tcj131RQMobDKmQxblnhlelDNAr6++p2UgwGJwq9wEeh++ShR5P6xsWtejxFUnR
yhd4Gn3yk7LfHANHPCXKGxOlt1Mx7Amjz9ENFQigDbAZMnbZ4IqK/FzCPTaK77YY
dPDY0EZvsRqjMhZDgv0GKcKxiYiJVDmNYqRb8F7guvomfBGEJmuMrcznfhWAL5bM
y+qsBnuGYoDn3TsPYM0sRSTEVZ87oM8gXl4bG5LrYsrwesF68Hqy60uzXaw+phE4
aUZ7aJPi8dwKHWj8d4Rk5v0mRhF8FyCIGCrySuWUZyZg68VvGaG5ULuaByI/Snff
SdMNkvotRGGljryATRqxHfht4dqPYbqNLRCa7MGKzNpkaok5C5IP1wzfIL9SQyuh
nMeRaALD8eo7SWmfmkPVvRuT/UfpakFbPVnszwu9RxnGH9T8HfTTQT7gqjG314q9
wEaBX2CgYJc4F0IXIx6coPd88jVGd2GtLx/TAtTMX00HkRx/MrKNVIpE7hp3Y4ie
u9Yy310YpLJxCvy+jxCycrY/QWu48E9R8+Gf29PygOXTozlaNItUYl5+5114CVgD
RNZO9eRUSjrfxJehXuTgObn6MLPp0dadIR2EBflHbU9UcNTkN6FehnvAGb8cybA4
OKLs6IcwFHyt0+ZKuFfcaxc5Lyq6GZzp9GsSM5EoYes2xA42BqsY5H0E7LIf701S
iLwiDyT9LLf4GjeJOBOqtbDFoQ6plATrhYRRe5Ddpz7jZ6JOC/T7T8N1j/EVh1xC
WIkBWjPy3sIGOO4f7f3jSaKxakyuD+ieMTqYS+GPq3R0qzCsO0T26UC/PVLf4GSq
kt82KgN1CWsJ8qndt0DRBUsMiUHCwm4vGDLzy+tMLuv87XLhPZAQCMSCDYSlMvj+
g4H58qZxZmmDpb68R+efTPp2AKXS8ymMmTCboog1NQ/UmWf7qfCM6BQn+Nt84/23
Yihc7R1oEKYRE+4KiLpj9dmPiPuet2t/BCyhdrtkyAFCzYWNpEpozb+AvvEgiSti
2yBApJv1aHZZyv7KSZ2kJWDMflFHEaPCKTzp1mVRt4tkaxHAWGZTJhJ0ppMDmdv9
pAO0UGuauB0GBn3GAtacHO+qp1smx47pa4LQyjgu2zWIQ+4uBWCOCwmhIhHwsdhK
m9Ra1xXWIf7DNWsbRV4SAroHnwQiTr/o88jz7Gak0bM30vrtjxSgZXMjNboXeIif
oSsbWtTEHmNbPLUeC8WKybyAaEzqJswdUCV+AtrUfakPqV93cwr7iTU9FaXlNi0R
gcW+UBKIKLEO0JiY0PtFfWMLI1x2SljjKCwlswsT0swGc1RucLJcNZQNstXBeZMj
Lk7brA3HjXEN1M2bkv9EQmAHvBDA/s1GgF4sc5l90p+yx/CAwRUAQvAkrbr8z/2u
JLv3+19VMrTLxbTZ4PaeeHPt82v1IZqOAl/9aOjn5fAVZvylg51FI4WV7hZvuWOF
s1WqDWLzLMAXHdngZf09aaLHVa70O9kHb/RDxiLIX40p2zZTo1xSVt31ypjXcuEi
nSFXFKrJ6Zegt2jXptfEI2yHocA83fqHdZuGyShXNg8V2Ihk4T/s/vsM5LMMgmlW
YboV4Vy6iUs2MLBz0apWaQF33oS31MAnFebHED/9CZ+ngm7UzTbimJBE7ywtPU8Z
BnUDa/wliENEv5acja1m+W5R5vCqvPPJ0dH/wsoDjY/U7jd2I4xhEHLQiDnTf9dD
dVgUv6w3yg0GuI1EyQQ/4BrE3j0gnsylJ37NNvFK/ftI1nIOkaM/aKgFd/LIBfP0
ZFfA8/Fmjlgi//4B7tpawDXicuAh77KRFxbMA6X10iQhHUpv5WwbIfYsyQ3Lc6FW
Zxw+bILxYuNo7ELceTsRvMeGh+M0kXW+ePO1Q1JV2TeftzA8rfnmIR4ku8Pet+D4
gCJ4z+rWQkm++4h/dgEN1mYeOiB1z7hGq5wj1Ze0+D9cIWIznDotS7wCYRYq4nHY
iX+Nffx0l9lawPDo3YVf4PTTJsmP6HbOZ7+R4ZjO23fq0AuiHVUeB7rsB51Ol//+
LQzltPhMQ8Qz0PCcUkh9h0GHIMCvphQjqbydhaG/fm0S9g+4iQVgEAV9giSYXxIm
u/CeHUgeluDNuk4cgN8v3RaBFlhESHMBqXt6mRBf4cWrorLVJTHDFlAv7pVZTEz5
qPQSyPl7lGZMzXNkoIqN7jk+hcp6MJc10rTA3WsdApi1CsJTJnQQKPw5mRFc6Df/
4H4oXGB/dzT5Eb75zNoC7F8ed6jPmRmVWqVeXrvfG9XLmmvGBArKSCjH19Y+fe6L
k27IuFKIY2xisAeNr2653urKRuAUOBm1C+Ad4ceiD0Z8sGJuI61CrRpAVZxrDTd1
uimrPMCTBV0E/x0m12V/ZAWC34KFIgzlWi46iMcgN9yV8qeSpFd6AiEG+/AvBrGY
lqsSd1InfG96r3Fo0VWDriGHQKv9HztGJ1aZcRFlxpHmKU+3b3tw6SdIfU9s7PjG
yZ/nVVd+r2jkICWuloe7X8dMaC2eR08QkE3goZHXVihCPfU4urn83SM7rMyzKujw
OBBOBi/mAGac94YLeYUHIiqqIDVMPeL6QumK4fWT9D7S8Im0bobjUuVSSwmMcjTJ
lAma+qZsLP/DlN3X8yH+mW5hGaclIATFcZ6g4/DVk1cxfpP3+vy/EdjM75+qDlI8
6N0k56j28weHEWaK2k3/aSAkj8oiJVT/loZCsK+rOj8mlsQQuO5IEL569xDQIAqt
1gJHNT3eUMk6gjn06PnSg84RhQVEt6Q3FeiMF63xwOk+LvVIAZvKrMEGGlz2JVjD
cu8Y1m8+bAlGAl/E68/PYQbD62FqhMePwwUDt3bZx1uSy56sfEXr8dAVRvBTkUJE
RuWZYRTnrfznelnPStIwYYOMNNScvNNgvkT2FkAvBD7MQVGWvwYeyrbWERvtcY5i
WC1xJMLb2l+PQzE8fniOiBL2nTD1AdAk3K0o0Zs28xGDrh/bpqo4rIcS2gbYnTD4
P4biUCNZQXHt6Tls+yp+0444p2JSAiFoxyk0JusjacYpIPJOLlna7gva3K0gG39m
RsiKu/ixebAeij5SoBtx6jpja+/V4ARMizrdyz6zMXht2BSrfMt4XpIoETHsaDhU
0SH/0jQ1CGa6fWoDrBFfcxPydERt5FWBf9HI0jg3Wug+kGgLajD3/bCacS4anxq4
dZ+UIdttS1QGJ5NsTTinceuQ2BdL0s41lOnmznF5k6QtI81scQbD+SIoqg23vLRv
QNUYqEVZLYgGAp/tkPxRYBBOL2+yxwlYvWXQH/XwjwX3UmRTcXTy6Xrvu73m4lAX
mdk3YXfxw6Y/xTQqKpLb3RzdPUibe9RypbL2wSadwyXQ2F1pcSQLH91RzagpNYVg
5kupnKejwmhGnvB4j/wOhKpQmIM4ZVJkPNnZ3byDIM07LPWLCUptM3kzDNp8yerK
vlB2y73Bw2/74j61fnHlSf+kEFqhJRNmG7A5TnrXaRck9UeltPU8HPDaHTIKKUGW
3olYY6XvYOoNIfBWWaeU84W/BHrYi/VsvJ2kZo+NbLBLM5DDrVB9pqxMcD+Qdvwi
JJFVI2ewo3UejdEz29B+gedYJhlIUp016xu4K0C62zQTZHqn5Mi1TDENpyYBXNoF
wujpmtQn/v8A8ZAjSQFQ+wQdVBMXiomFPpyn2+eOQ1vE1IOst+94EhoDX23yy19U
777Gyzgig7b3tMYPAxx26KtJIZXOshu5SLyEzM/0iRlthCKkWAoz8LMGjAd5vL5/
9jiVXlE+XPnhWsZwIyWo6BaH6GdwDrAQAj7bKfWGLsLFUZrhHPNRu7i+pJw7aFE3
uCdO9HiHb/UcOLERRmspgqF5GNc66GI5jaW+ssyF6qMVYQgRnQHuaozTbSQrc/UB
9tm6q3xbl6GRS7smbrjpn6tAEz37aIUAiHSAQHUS0q1VVL6RKZqjBFFz3+MsV4dn
gfW45UPKB49giqXBuVTObbaImQgORRJWeYcDRnFKvFYbperkvP78tEH3QDSzQjz6
B2FMn6bWjVvfxsY0cmMcEpFY/JhonH11Dkh1YWyUYCYJzZJqHLku+uwfBwMyB0f1
SE5Wn9d/VOF01Y9KvdA2ln/aP42oxt1Vi2WqZgk0Jb03tFhSgn5xRa9YM+nA8FbE
JODMOtVG5dGjeZGuIhs7EAfnNi5j90uBkwpKJOWFLeRqtkVNoDv/JcAuNNxbfEtl
ojJiYU0/H3MJp5GRrsswIqxMjdH94a1ifmgp4uRsR12j6xkPQLHQh253PBZGGXgw
euO+gSb8GPb7F3nmu7I8CETKEUj4YU3zbky3x2+dY17butrL2Z4xgvFRk0GWPU4d
zLySTGXaUt7GoEP513AL2jnzBUiag2BkP50atjC+mR4SBsOI6ir1RtDKb8GUOXFn
WYBeDP7HkJ9Hhnk8K72NXr+ellPv2+n3F6nIJbngft9yxbz7qMKWTzdehHrPtzmt
Y71QrnG8haK5BVSJ7zMxCwfx3S2YN5Q3KfwcuXExHDTsJg+eerZkHmXrs9jVelkj
AkqhSjPcGNkhYzH14QwJjyD0iJRC7hFvFCXfVeRaQZajeitj9U3CfRP6a/5nGh7t
gRTQIAN/33ntM/Jjw5C+5do9gN9/lql+CcTpOQDf8GC68ZCScRtVBXS5n1U6HOfQ
gpKD4X5EfeQUv5ipE6NlmSyBCy1oVan32XtNwYHMxVcnRaOtx28uxXV079GAESCy
+VgQ7I4JGDOPKjvC2x2WADJZoEKvTyBRR96Eo9w3JgLT9ivCxln6ZCkZgIS/W/AJ
tbz8NBcwDiwtK+vqiqgltEkgw3ByF3CIrJez3YaaztOySa7Bz+SdIDMtkcSlEkGQ
harh/Stkwz+DsE+PNUaEwmI6fC1LS+ZG9gnRZQHD8gMYaD6xYqJ02pq1EMhyZgTh
ArGnZ9mYdRyHCpmW2fYNcy1gQAjBh26eiXdDxFkDIbv5wA3QVrreYFtu3Zu3TaGv
MJf7g/MHNvDllg3x6TyNdrb6LgR70066uWMni8jDbNWAio6YFtrdgP2XvtOZMAM/
LGMXIjpEIWi7DocYQurq7b75Pnq0U+us4IoPZ7d8TJkvJDV1Rc+L4SYVTItyh6qe
e9cVwK2GsEl2On/0hzYIb3OTdptpHOvVLv61XQ/ZWdno7xRW0lFWCK11/5YZHpBz
FD81KBsopKvY51On5Ns1vUlngyFb8rAixztH0AQEFO3f1xzD/z1fRxC+x7xrXuUQ
DSKpLVUVFpnt/RxcL213GNnGIVrVP/f/HRXbOtXhv91l5+bwYgjSXsSXHEpP+1bT
HOeoY1jM7bJz9Kgz2JTfCuonwqWGkfcKMNxeo6ccHYUqjTB0HkqZSL+1AxOAYOoe
grbOLdu70SnvmWgXK7x77EdzjPgol7im9WornUJBcH3dr/zP7B8PqM/dVLA2pQ/e
Q8RDZ9vBG5YU8HHMtWXzeLqYojf97YftUqRZPfclMMxwmQbDGMTXJgq6IxIUsSpF
AgI/1dnrMgwzDjSw0SPSwoD7V98LGfqrB4p6aEirlBeIW7wIR3TalHg6qZglrY1B
2uHBDNikI8utNdMmyFP4h6e/oI5BNlrgEBHIHcK/Lh7oBO1kED1M6m7KxHQDUTFv
o2tkqYw1FiXBOJgM1ftXH8yzdm1pQnclUPh+Rovt4XRECVJK6tjddWURmcup6tYM
q39tk8aLRepZjgl7+tCohxxHXmIvwH8eZ+tUgWglXdQYE+3FHOMGOon9M9cJbKL/
PPtSmc+XbLafqrUG5Eg4k4IjZvStSPeaM1r7MdnJnqQNTp/z+nJv5LH+51P96P8/
aGZ9iBBIksoSSU8cg9J3wh30tJSYlHo007lnvgGVrTFM8TX4addYm4aZkjwsHt5t
MJGQVozCRE0P/hRsX5EJ2j5gxBJbvIa1/SKN1GeemmMH8EXhhUqqLDrFHkayfGwi
e3/4fotxzW0Q94uQzAAB/7Gl8bHHlyq/hBoFvnObDwrMMdzaOdT88FeoFL5pSSoP
ROnhjmlYrtyQTXRiSirzIIz2VYt7ZMwW2OeORLtj/QsQik4a3UPUpQ/MwBKnnZXr
ii09zHzOQLrd7fLw7mDw0X6+b5+KVTCavJDVOqHSXOil64rD/Ukb8kZYl5qmOCgx
OKNOvHmoDhX5aclMeNqIwsK/+WvXyIMOm0kxlxbgUK2IlHceL2BURk5CY3FTFY2y
9J0Wvezd+T0BHh6l6j4UUaVnMO9aHJb7yT0Exh/QlQaxt184nBd6VxLtgerx2IsQ
pF6BHQ9sQyIrSaLvLHJoHveXzemjdRr392CLURTkR9LzAEo2GUTwihP045wfZQfH
1NvPCmFuoIlHZS/7jpPxCKUs3ZPnKjT9iE1XjXvAOUJqZS9tVOY0IhXFEIB0Qor8
Y+Jb7bO6LoKwgvqhNdLrJ7Pcbev1I67LNQtgWpiHzLzO/BScrXVJV49+sNqQi+Xn
9l0x1Z5QFhu0HKnBB4JTrsVW19WscVs2TRIQgmYF0+IFbIYa2M39F+mo7wvbOxxm
5bYPL6kwZqodxb3XBulJVI/UYPYHL6CSWJqodrcCKym+uTb4k9Mry3cncTjI+Olw
j+bS9FiK76gvdsM2ePFox7j9K3D4l6ckg26maXd38dBh0t2XQipcTC8mcqr9HsEX
4GpeZRkdixzJwH9adCN2tC41wHLkPLR+y6J1iYAVII68Wthho+W2NcQsFUicmRcF
MC5bcsEJc1lCTG+9GDUwXZf+t2EN7U8eJeC/1xi9s28lwLSkXW4oAV1yvhp8Q9Bi
7PCPBSQNjHNvoKKFbf4ozjx2bFh4QvOrflsxi3bOQwA2hs8qvHtfD1+DU67CQ1Y2
U2gXm4al/Ynh/fcjkPHtR+ljMe7DOcyUtX2syFOOSXNrDafmapIZPGmTpQj1BJOb
WPH4LB2CpVQqzeLEtC21eaQWaHqtpw6fV3R2mfYs0OYurTnLdg1xr+gdiX7fGrUY
hbwA4I5V7k/UfbZY8KTEzkchOnxsPGfCe9vXBYzKay13bfnJB5/ucebTciCpSOwi
z4pJkDQ09LM6BBLUMd6ng/B9F5v0lduNVBR+wa4hv2lT7y7qJEZpzMjFu+XovCJ8
YRMvZTVCoNbZJHhgu3sEcNaLyaS5EScBiT4kKYdHm/c6XDXEv3CbdAuPrL70HArh
ZQsMzOPoQBRd3BAJ+uEfjDmhA/bGyyrz4njmxPfF1vrxFY0OgNP/Yl+hPAmY05q9
iU/ZNissnL9Zz8eTKOzE6N249Jcbq3Fl3ckqB1S6FvuGusjw/v94PvQahmrA+CLM
ww+W+iDYtIz5W4atbHBZ/WhfInJYr7u5xyXL80SFdzSqUzbTW270VhgI5IFiNE/k
zklQwyUwPH2o49j4p34MvmJDIGEokB62xSezO9x6/RMQGjbFhZJgd5U5hqtJX9A/
/degBaQD6fIhzHeLt+89zFI0lWlR+WhQjnB5dcrADullbFd9o++ypVzm0tMJNVbp
XPoWkdvmmmUIxlUEVjjIldzhsiDYKZVVyh3Amn4rlRGgKilAwxhYs/1+jnJegVxC
xe2bnBWzPBaA+U8c8iJjInhEUe7ryOWZaBcUdqUw2nzRRGkhctnjpfWr1SKq9240
6MtKg+rJIwbmsKJL814MgvGjhTce1GnGeFr5bQtvChyZ3f7Ie5cCbfatJk8FT5ww
byYS5bM7CdMbZi0e42vBOfvLh0rxhYUXNWheHUPim3gkZdyJa0g7e+l4lgY86WWF
2FigTaI/fi1QhW+YQ2vI76y8QfR0HTQefQAmifjjrefEmnqP6Bp5ZzxcuG7SvKwb
kSSzAGf4bd6EHOckqvIQkyfBvFbH+JWydgjA12mJW6ou6n04HZ2O0KMxlIO9Kbtk
HdlsBU7ByiZmn2CbMEIgOZgCjAGfZOuCaWEe6C0q7O70pFFNM2PiShXqyqYXQR/k
21tcgGLVKvE9lJjWtbAp0rTU/PIKtWDIPzd18iZzi8ZXBQLnJEDr0Sp7QXf5Cq1X
3MF7q6KAp+xmnUWqSwLznv4uSC3JYEej2gRHHnci7tL26timGiyrVtaDe1Ot4WxO
pEW5weDNaOsgJE7fQlA6AnvCeLS1EuHFjuPm4JggXgbND16h+em2MYDm2QxJ6gRM
0+HNHn2P7zRKCEf6TVAslB/ab0Ty/ZBL2qgZDoj0YN6vTg7USggBMYkA15X3aI43
jDoYvnA3AgRl8oOX/ayIUtuZBqp4Hmvu9Aik/mW49wAIFFJa5GBaUPipP1VGN2NP
DkCr2cDRJ1OSyZql/L06Tv6xaT54XtgLT4xoet0cTXOj5aXg0ORhVVDkmZ93T1yb
PqWvKwK75oTXAsGFzhZifkO5gdtAKvbUm3ISG0KrGRGB/UxFFItrRe1G4AV2pflf
B9E6ipj36TEN4lUxXbQtOHDcKL+H+tP2skHgxahqDfGUJ3ZDNwxEKlTG0t6+Z2vj
WQrtsE/YyNnuq4ZBlk32UCISr/wyjGeccYnYZVE6wV45GQ8k60H3D5GfsnI0qE4E
w0TulkhGpRjjWM/fwCQymsmmaaL5d/4vwG2uZ8ASuwcfNFtFujg2vTGFVkhPkY+w
WxqI/fjI8XV3mee2hEQURf/Cbs4COqhUxumZABYZ9w3tRTDm4Sdg5JSrtZ4k/Lab
D7/cBfHyoPzSokxPq8D7uJzbmYwug+AtTklcrTJ7vCSmgZe7INbo+xoRAJYs42ZX
xi7Gx0wLTGf2x3zSPUo4t0086msnhxiO5JtD/cguG78+Q7PsylsUYqE15Y3QCDHK
uruZPJWhtWmOWQKyWzLb1onZvPDRWMnKIux0cXNajYEiRpMfT613d5xy/G7B+Izn
uuk9HgG4uViVDk/QI9Xvbdl4Rp4f6J28tCt8FtQDpabBN+uE0Dhv5rNdIVgFlAwh
fpsWSN6aR2qxwWTpAb1JJmlVZC27EjKqfWm0WZd18VDdwbLcHAj3xR38e5MlnBbR
95wSP3L9Ihs5KgsBN5RM0p5+2XhTQ3ef8fl9X6xwSARWWdjsZi2vRDLo2Oz0vWVM
/Mix2BTlEBI9nnZxqArAoeDs8GjUy/imdDiFKz9vhfnOQ2VH6hvthXyu7EZ1cQnL
13CcGrIV6QEdwh8rKPcdXempAzxpbfFz6UqCrAq2SBF+CP4rEHoSPk2DvulFV3YC
aTN6bfrw0wNoKbWdzEhrOFCfwY0L5H5t+A7L1zO9x/S7KbizCF0VpoXJxJy+N8cO
eqvXjhvk8iRZLDXBTLq7jlXPeVUpx1rOKWU515YDTOzL4KzjYssRj/7X+zDiJBiz
1BG8a98yaQusvIix2d/mYFL+BOLCCrhb9z7spLJ0btoV+yxOkgTELu+BaLU2yrbN
eGhR3DzKK+qDpeUalp8X1Jp9argOdPVghjYSnS3SWKs5wmL+Y6jZDPCoep1rdata
VxsvltfZ67LFlY1w9oT5KKJ7Vjsoc9rCf8K2wBIO6nFge+2KGtrSZCpRXxwwuQB2
3R/zLLA+x2bpLnJ6J8Uq3BhMg1Vn3xXZX8gr7pMGZF/+aoc1E50Ex7iS3jJccLxy
ZB/XuxKoaefyadCydTmE8olGXbtHygHGWRn8IoyBePjuqtg/MPU/qZ1luzkQqucF
75s5e6dO3QTk3j3WDDtBA4eD8LRm9+z4c5uFANuG2u0USfAn0gtYUnbPs8Ov5qmy
JwUtupl4zMW7uaapslujo9UgXpWnDgN3E2t/wtnjr9Nqe9T2SPRMHhAQ09at30+z
fBdEJwA75L0Fe1wWVcInAyWTJykmzaP1cl5sHfaE4Xb7Y+uhT4l/rIaGI58MWykl
epJtVW1MOCJh760v+UjqoUaCrEcvBbvslLdEyZlrh/AKWnQf3acDG6FVDXrSC9X3
TJgO5zzr6ZEirB3/5BTXscGgnnNNXQBJLJKA3XgMpjzNutC4gnOjRhLgy39h9quO
sghtFJOKLWxjtNEDR1g46M3ysIYQ274FjKNyb322edTOpsjyoFaiboNe6TBQ8gqA
SUJxmizPwz8rpGHrRxcIaGdvgB1yIDlEKMxCJ/vgF3WwIVI7zryRfU1ZZyrbk/ee
AH8bjsk4WobTO7CXaHEQzRYGyCd3Ct9W8kCEe3U5DZjoQehmvnNbOb8DdJkpfUBe
vDQRdp2MyoVRQpOJ+Jy0KOokyfIm7C0vL56mw645Pl9bznoL6ld2g7EHfp7D5LnI
9rIDkg0qyNs9aAztCl8uqI5SLj6sFOdywcMzxki5+yVqUcHgFxV89HTBBkg2PuLx
iB6MNjqI0QA7zJ+CDFGnJxMg+2IpQ3vPvpdygyFOt/8jKsduVh53MoaEtmLdhvoO
O1HiO19WwZIBuZqDtv2MU/QwGwgUIAfKNTAzQszW9oQnYjCtzroSzeVoWrtep5RH
voR8YYFOEkIRYnxqCWY4QALJMQk7urGpJLEGtJUvNfi2ZBwpNS44A8qfIFHhbWIx
ebWQgxIcC2JWf/ybKfVLwbYGl1Cblp8u/rLEA8RFBRv+lGNTcmIm3PqCM8Z8nbXk
o9uD6Kqfg5J3ACMOtYLd2R9p04BBY6fETt7mb3xBqq2YM3UsGxCdpwiZ8d5KgCW2
ALZyH5BOFlcf8B1SsqcQfeyzPJJFHXNszj/AAqKrac9eSZykUlUoEF+Q56yIM06j
WvCQFHRo+Ys3XCoCahgseyZocY27Br4dPXaEPlLJlq3ruAaQzEqCC64MsPhBmUgQ
IptvEAUhzz8U8lcKo0pV8r/EEgKUzpAdVc/14I0iPTiexR/d47YHgsD+wuN5fuq8
RAWjswiagwHJAWQ2wxlWiYpjtUO6ZBf2X8A/79sgLFEAtSBpwEm4rPqIHFYvRUEn
NT/zZXzGPqn3s142/PFIDYtUp1YJ2J7Hn7Tx21C2OsJ5q+kpR7mgyHSGJQUGWtjO
qZpqD/QCMMAtb5A2ZJ5AG1llMI1vmDttMk1mEsv6soUXiMtPt+6SDL97fICXU9q+
2+Tl9bo5bMy/7h27/EJEv52Xh0qRIBdHTN0m0gV/7U3/A6jFGM1kmSGMDNTLQ+gT
dbqK1h7KnV8V3ZAGvzNhIjCHI+SbiLHi5Z5AFTpY0w3DxpoqoGzJok8pocnR7cOn
M6FwsvUaZBJP9CaMgPaea2cTO7iJkpFQSqEwBQG2ZwjOle/vyr0IvnZjiiC8b+RQ
kIFYsegR390o1CdOqvoJL5AhmF981ZGY7TWYvvqGxERWqx94FFCD7EAGq3g0dsOS
j3nFbdI4ev8Cpcc2YATvPtc5lwJ/EES/Ku9x+9vHbKd9wGjsvIsj8XDzGfJtyfvK
vyUgKAwZi/vtq7kSySvuClw8Vpidee7AOW1IdSLaus5S4YNQ0ft8xX5rJ/gIYUmf
b+IpSuC5tHSPjQMbCUs7qPwAwHmQNpzrCTPQ667HVrSYmtceeIMvZjuMzNA2ao0p
MBC+vfIM22HwRLZXLmL0E0yWApeKlhIopggSMLaK4G+FTzMaa4mygitXVw/Vn1Xq
GtJGRYjTBFsWu6QUZd84doqrVqZ7lBbDPdG8aeott8SwwyFTBTqdSeBgFFdaDdVN
AOZ5cciXwXeDBMpvYKqBYFCl99J3BAwwD6R/ADqD22qTupPhIe5LT9oUxblhf4D9
MVBETKY9gc+RvQXzvxPB5JoDLOHsv4PQ9Mu+3mRA/9k3XhWgqhbvmWPXN1eAxasR
FHXk3fV25+vQb6HfvHSAeZ2/0h3Gh3KX6tMA5UlQwpkjHk0kDZyCEGbQv4F/vk+6
HblDYevWEi6ZRom5oSrd363uZ2Gr9IIRUviI/6SKzXOZb14sJac5HpHBn1mbrDSQ
RETNDKDv3MJ7x/NyRwFkRo/aMJmgwJB0J8CC8bwzUOmtfIGd6m8oa4PtdjvvWqiX
x0MWlOvG3jZneYQ7vjlLkyhjxpHEsm4YXM2plS0RufTp6qI/M0U2rkAIpovJSScf
uUSG9rO/tYzDAyfrTsEsDVae3lFQawH7tDdantsmuOeuWeAFV/BQkSsGzl1SVCYm
VlF+eG6lPol4Z+FasLdQhSQE3mOanpIc8IaqSzwLliKKPqx86kM7FZikmTnf3vRm
E9dmuXUNTzhyGs9KkR8GoUK5K826vmkgzmsH8N90LQhBEtHpe61LEDGRYxyEL8IX
epq8TU/jGrF2BEu4WDpruw24DRCLC+foHv/hTdhCHh7Du1uWZ65fBaJE7SN4Pw5v
bqMoQeLtu90KLQrkTs+uSQb/d4UtBdqLYWFup6z4a3yHW4CwjpzXYH0/mFB6vNqi
taSxCKzvOXQUj16pKvhQNpsoWlE024M3azAJBsuS6GdZmp5wChpZ1Kt3SCdNnvqn
bIZ16AJw5yrUTM+96B+nQVq5tJ6hraG5XIvthdtq3X/WNT6y/L1DxPvAM5cL8N38
KuTPy04oZ/Z2kV55aNnKJLKJ/GZCe7K1cZ8b+bUYo1ES680cbZBI4/yOhfpOeibF
llaeAz3ZgRQ+a1/f1ZpD7FQQvRYMYntP/OzFlnOyXsbCCljIdL4CtBYA6bL4mIgv
oSBYwG76+D3UyKNB23fDlnl6r4aRUgDCx9YnILqbMjYCC5/IqorZmGmCvJpET0uk
9OW5tAaz9tQ9hh04Cj8G2cGYEYwoMHllf2KMN7F3ET9jQylOYEqIHyXmQzQcBjB2
aOyaKm2Lf2Il6nTfCRzvKauK7muVY1O1qIkoWVf8KqVExUZn9bAqrBkF+Ha87ydS
CJPwojgNW1C1/K6uQmOFp9NNL+aIvA4rfVEa6q/3pgqBlT8cdfzcplf/lxm08ugL
M5+Qu41ko4lSVj39w7BAyRBjS46FHf+pM3pHtoWeHmHMjt8ZO9neRexd7VFHSS+O
XbZlwN2OqZCgbQUCaQmDn2N5wH973O2JTaIgTzwmo8f10xCa6saoKk8Es2j38FTS
kAT7p5M0/tVyoTBDb53GykbmXM5sueAigffbZWl2V6t7rQm0NXNmE8ZurYyOTK5c
tKwDoUHyeSjeEdTHmMs56+s3+Z1jC93Ke23m/PYFQHh4z21vjQoo7aLlB01F0cCm
CDhqvdGW+SAQ+X71/qlnmcI3/ieNjiwMfK47blZatF0TNWrBVuC49iCS6T9JcFkr
rGRa+g9ahbXO2diuf2D9iFz345AQW31ixy/WuNLi+bE/G/d9iC7LiE/xgh6j9UNY
mI+2OS+7O9e4RqQjIfd00WawfCOboX43/iRnOIJJYraxA5vKPv3FUGeE3P+HPKft
mBohnaeQRYRUEn7Huobtufb3bVLsHPZbrZQ6P9r0mvtWIOMUx1RwBDxcm5dMAg3q
js6mRCUKI0FU8DxNiTwqvKHscrKezttpaoO1qjzxR+hyD0znR7CIxlwSeYfWLSFF
ItOww7TmMfwSP4dtozCLhy0GCDbDqJeJ++gIvKPaLwHxAUojTrqLjolWs3xvk8Tb
+0gHh/lsVSc6Ges4sjh499lrLFA722NgTZ4fmH0v5nxswzQHlOr6kKxyNs7i+W1f
XHy5MK4b/1S6VXWlImmTiANt2swp1Q5f1ZgXU+srSz+I8osV9gyGshzVKA8XJION
CpQ74s2V6OTL/K1EanBEbuWvD4RegGWgyK5JY84mBoVy9jW+/NfNuh4B3lX7NNmA
bm9MewGV8/2rGwBUKFt//Lin3fWWMR31jNHxlj4LxF/Cly/eBE7DWKWjh+UyNXCk
RTBY+ibu71DFwjWewRPqEzTrgbajwD5gEXSyBFprAAFyxTCDcQHj0Ebl0QY+jKRr
4TKU1hdAiXSGpBwhTGh9FNRdIMKwGxN35i0J42D02WaVCAZgQE0um4TB1wnBrdvQ
/XQuaphqiw7SuMVCcjAd6FTGjMyPBvV0bKu1LfSvCy/4rh+Xjk2wnisez7JXOj0K
YrmLIk9y5vZxh9LC08gE8OYr/CfjZSTLIXLNHHkR39JkiKjv8i11XQN0lR99086z
wvM9UGSErtXJcta+BkK1udH0U7vg4EazBGl8z2xu11ibYhyZLvvqIFa1VJTjPi1O
mVU0HPlsoOS9Mc1aMj0p8dJ3NAOfmfvFoyKKd8pHBApLfw3nU7nAlcGWH52uDul8
a0mJSHScrk8bNYEUN4iC2JfZ77pm8lIPUeLrE/YB1My8BEP4ikzOlOd0/q0dEKrA
VsyzFU4Frn2eEjc/6WQDcQB85W/v46vk9nd9uDRIQDHom/f2BIsjJFDuDCbk8y62
ytpjHtXeKb1sg9clfYbXexD/h9xR/oTDiRITE+Kelm0r1Hh6qXOsIYP9ea5mT9OD
1mnvfITRH7wH04KW1bFCzPwRVuNfO+D0DipdCmYl5Su31KTXc214D9eLy7oDWwK0
V2MLA0Z80AiWF17cG/hdla2ZLNzGVr5bK6ZY5XhMNVl55aIo5E1g9gIcOL51Frvf
yW90FTt/QuWMSLquSnwF4TAghlgHM5IuXAAz3GReJI/CVJqO9yusatsYUuNh8fy7
koajXQ7eJbwd0KNtNb9LvZKkjZ6w2kmZm94dBN5+0DOHZCExUiDU2/OGokF5cHri
/K0IkdJNQUHWThN8JPtMQSWEqTjmzW4fd3QL/yhaYMOmoOnuOtIqLIMWkYYs+5Uh
tfYrJGD/wlCQlx99at5KEqdqK7f/otmTvnTzOWLsohtfu8Oj6cMH20DCZfM7AQEA
tN3GWmfXVomBuV0wxhX65/KwTyOqZ6BYF6Cn+xAf+7H9uVwg2U3Eczu/8dXS9rGN
jgXiqXzWIqtOhbFF73SyIy9pU1/pw8FNzTNYvulHYGS4xJfuTFPIOELQ/Cbc80te
0XIeXvOkwdKg91BQYKXIGS+6NEHaS9dUJQaRTRTbyQ98OoLILzS+ZHlnEbw/iltC
McPMaJ5No9hYmqMfyfNc5pVQwi9nCPlP2A5e1EYzo8BE+MrN0UgML6G/AJCvyVuE
L+Obfw1LSLImyWTGo4lg3p+Cldy1HrvVLC84Ss7PaX9tKagtD8DaXZLnzre7w1S5
5mwm8OZjyJDIFcLYWJXsmmdeKEsKyNKRIUbvSQqC27XRym6/KoDScg0fFufQ+eaH
S/wQWK5fMYAfp5JjkmDAl58D/dbt88FV508UVhK0NkXXG4/bPtH8vrj05WvrkPAU
IFBgli2MyD0Lu4/RtmI6713mvemJx08/2V7QC/didnc5z//AsmqUBHhJRauDxOjy
cwsfhDKmIIYLGm394aF+ehKS2o7LG32qv9Kv0tAsWvMonGyXk30VjzS9PxqR5Gcv
YEEn1aA1f415xlhFciHJJLP7YDo43MkgtKY5EhQqHskjVVLBJf38BG60ZoQ3u3x3
u/u9vy+TRJ0FvYV5SVPVL5MjFQ1ARx+MrebCJAsibqLMJzmMBlT+UFXCaW+oIppj
sOtgd2rLTfUNb/EG9j2Ri1rNBxp26WpZNvVhGcnCEc++Zq8/fLfKDOofLv5suCvV
hhNmTo/0Z5xovXJBxdeLd+rLTluoaWp82C7UT7+uOAF1E1g832TPsBXLjRAcgoXU
G+3ekO3rlzx2ygfhTszY1B93JDogRJvQGAQxNuqifx2nYRwJ6EfGjbEMQjREZOAH
jdGAKJaW1ZD6xM7SSg7LMPDOb31hdzgIEk/BArlZTXcUlyu08k1p/XQdnVQ65/6c
JBifrdjr1RU4KCjNbpfq56iTgBmQbUI0gwUMIaPrwVuvELKFjPVnUDilL/nLbnW0
441JVIFNdF+cfr9ALxIAfM4+3rslnjDI2w7UHqPRslJpGoUU8Ku0u5es+o67EKJi
u0DxmfeXp2YOfBCrGAT3u+XGuoAD7EUgZQyeMQspUvJbV5RJW/JlOK0j0Ez5cOH3
m7CjXhOZS3PbOsyRmmRyjniwcNXq0k8crq8iO2iliS1tvfN3wD383YhRiF1p3YTe
wC+Nb/e/jT2BoK1jk/l5NON7XFopwdywUnnZIwzyB4SqkS6y8gqzUFZnICfrZT3K
gB3lz7XKitm6AacrWrbb63tCO3/1Exn69IiLoUQw/ikdkSMPv+Pm7kqG/ooJD+EG
Ub+cmnPaSamRDcjVrAYRYeHAndbHMpvrTWChPHPT/AceaWA+NgZB/APfmnreFtWF
bXKCWPNc5+mGcB/wLTk2gqzDfkmeMuQ6VdVzOeH6lYLNQ8ASb1TdYjv2bkpyU9At
vnNjHET6LM7xntEooRVd/6pKVZTuwCpb0byloFVMGIdtekWOMTHKNX7lyGRazkPS
QY8/2nUnvkCOjMMbZYo92WD284Q2Q6NE7JbcQuJZa6LhaugdxagW2+7lhxM+Ajrq
AJwZgsqDYvHGShHu88gDLwGn2K77+lWlmJzoSsrDuRUlOuR+Gtvegc7nAArV6Cwy
HLXgO/xaojGdAkPhJFsHv7u+IHFdkbYQFfDF/oZ3TX4BQ1tf3ZV1o4FSBSFrARly
S4gQvxGx1KfUPllxg5hNW1BS2GphUCS5BSu6ss4epOLvUuNW+Adp2iXk7YALv+61
VL42OEb5w6i6UD+rP2rkvPsiShzhXoqRv6C9epm+cjAE2HkZCuSMaEoqoZXdNhIr
ty5RwTKxZ16M3NylwWRB0XMWQgz1bWr3vl8kBF0K1BY23Ya150NpZ2s30qwL9TRh
HdY9mPT2M3hBjj0ARqmaXYJfpRLKNgJWWyLD8lTdaGs17rKfUIL18vX4t5+RsP4l
s+jK5sHIIQRvLS2dFNizu5LLVCzcSGZ7X6eS/+f9a6L1a94r3Vpt2nPBGYm0LFya
5R/32TGjbzbjk4Ay+sMQvoFNqbKvXhbg0af5fzvl0dxZqPgy/Pvdl1rKJIPcO7jg
gxHi8VL1ny8IqAg8nbDDujYyllPlRPHfcCkdCqEyxIolEfLrh9TXiZMLKTeK6mRp
DIt1eLNBKdm9KuwrgkLb3iYh4QscPVDES/sdEgbUZ2LK2Lq1gBN/J0ADGhYsdNV2
nOBJkegBkQXtPEFxmlqDw5bcBeGWcnDGHNdPNgZ2ifLmFhvzvARLggIQTlEjJjOd
0pjMnMEdSiRqFfMH/eFjdS+rV5Z4ojla7k3jW/pz2LQQ2nN9OyqZq/5OaQ5iF+5I
YlJPmNP4+SPFSo/iY+qwKNw1Jg6X8FKBA31y9p41ieogTb7VK3loeck5wf0Q63vJ
iXP+KZIiREqC+dyhjuQmY2pEcat1WDBEoQwzP7McH0E0C8v3HANU6ajmpOBZSMs4
xekFOPokp6PQSoLzVTnB847eD9zQKOXfGy5t5vcmalOLNYgX2fTh5cBFP9IDn6A4
fEXWUtc7i29M/pYBz0NyQJFnvssvbPvTLah0WOOTolGRsZIqptfTZE3z0nRXoOJB
za9CYicrSV7hrW5tN64u6QE535tZTCQPH3Mdm9G2+OXRUs//V408gxiCBxZ9uJhn
LTQCjeS5KnK7PukThrUtq3Y2shVKvu8H+6gxMrtkjzT3fyeX2qlVPNCGzIz/1Bi/
iAlAcDXGAE0H982BpoKUvLTZ51khtCt/OkB8P0jUdcoMB/ueHGDj5pQoc2Fn8dJ7
fis7keMyruvTgSQ5AG4Q4jrt6rqanTlvmDoIsxY6yZrsC0DGyRxvpxPcp68AX2to
yBnJCtaz0Gl0DxYQ/bbFWK+sqw2lxN5RuVzFV66tVkyQKN8UElK7nwQ2wHb+/WJP
FvpNe3A/k8sR5/N1+vzWkiDs/OakgfzVU6pFe+Gm7c7NN6i7eHXxgYCuwYx2wwvA
WHsnsTmv3hDC5VWMf7rNlJMBFM4o8FRqlF/qbWm/CatePws7NFh4vZDK291yJqKe
XwHJqZbCRVBF7xahReQv6w==
`pragma protect end_protected
