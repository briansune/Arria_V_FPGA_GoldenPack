// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:33 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
a5fMIqJvf2UqLq4Rzz4JzJNS+nlRoonoUrXctqSyuiRBp1xKsWCmAkojX8HRq8hg
GbegvRk0W0je/nvgd1zSfAwMap1n8HEFK9dbj8EK2Pqf3umIUO0V1kzyYskxqiam
lKY9/46oqHwkg5gTeIoW77BMHNivbGaZeWUQ1AuYq20=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
tw/zSgkJgQ0h1ozdD52UNA7cW/Y0P15SC3fKGuqh7wZs3FFmlHRmEpLZx+vYQCUB
4v8XnmyzGbGcCO8ki/uOWBC1Pme94JUaaJPaZHb8fRiWXhvWwheH56Xq6OvX1zxO
UkP2ro9UCfX/sXtwuNJZy+GZVEcxzqF1u3I4z0a9LfahbDImPda8y5QvgAjKhQ66
WtD4TM7qSHv93uJIRBHPV5O6NqeLYtvr4t/0CbxgVyDkOKUUXjAEg8VGStDBk3tx
mWP9IW/bzpTnbm+MZ5EdFZfzAmHz1ylhB6xhKYroq297Z5ymyxTxo4ZbuXuq7O7q
EbmilTJZrw0VIjB3E+ae2dEGnne2NupzKw+GMKikswhbFCVWVyaTTbPcYd3qqcet
MtEjJagVITi4f+UR6YdRmQ2EON29lXFTBPtlA3XXxvoLt4z39SD5PXXFVYTTH1a1
j8KN3yGDwxeRFvjc85Sl8Z85vhTJm+YXr5nGEYMQFj7gg+K+tMLZXBElUpB8eHTH
JsL4ULjmdzXt4fY/cVOalofmIaRIIfhA9upS+HiDS+CxUDt36jEHkVMCVbBtuM1x
wPgwk8O+A2xj3jcepenBuzT1sif+XhfjzF4Q4f9dxwF5ZrZOEJXvQ5ZezJB7Z8ym
N7h7boVYXOAXhViz0GFGOfnTFfuIN87zhk0WiYVoh0v7ylhV18XEDfFUaHI0utv0
rX4fFpSIX1Y9qrYXAVFHMCrceSiC/w6D6YKMj6p75oFLlGMkh2ZTh6mGhikraoeS
hg4aM7rv1yXTiFukWNpmuZ+UujD6Dg/Q/Zxjw6LFgbmSRSot9F+epHb5ihsjMITj
nms5JJpVGkXOHOlMaoDO0lZMh7ISyp1ZycOq4G3s1neL2XA9MWoM9196qcnLKAtv
4NDhtPtgfZ1JbHEQZthHqEuWiubWuRx6S8Jxj1k2VCisTYKKqrq968dRDvXs0CQu
APr+epq5nGi5M1jEhi9cIny9YQpA6Iwf4pPM3CLS7oi0I5osi0FLBYoWkll2OuDp
U+d40YHGolV64u1q87fer76tWBAhoIZhUYMil9LbagjJAlgpgyNARJVPymDx34q5
He/f+BTAqqQuwGK6yV6itMyyqXluJy0ytmleStyDeJVqJCOQDvv4nHl46+KaNqQb
4J4y3BMteyRe0kGGeYBYM/hHt7jA++BCGTyhDLBFRiFIqhYBLhqIPlCGEGfqDVSP
2JOzubSXgkg+NuBY5lw5zdw2Rpg5LS1leAiLemS3MxfbmiH5REKsm/jQVm1jql0m
eGeLwd3HxpOAeeoBI4R3yPnwX+eJQp0nwSukn1BU0326QqTfhmbxtuKoyCnxnfzh
h9ARjWtW2GJ6dt3Ujh9ZHmZoQmKS8GHan2PcmgtG5IFqL7itLlTgHA7r/JxsGHVT
cEEUjxcLncfehnUOS+0FH5j5k8kDu49tS1W6GESgkON3+FUb4lANfp/GRh1lzk9p
KsG8hmiPWS4czelf9raZKuwF7I0VCz89wn16BtD8rjcugKdVyToRthfRwg5AU/c7
E722rC4xF1q8nV8uSOWWr9JlmPS9CiiIor6VgRjLAcdFic0hPTn7DHWO11VyXnUW
tE/1ndntwyNzcKSalmufArsMyG1uxfnreWgGQr6JH1+iImr24MVMShyGsgpnGO5z
ic93s7J+2fx6qhw/m84JY1i3mAiF1qhNA+jRuh3IE/bdpfMEMOv41kfOEdbOIzdw
XAlxvvsJ0f6wjm7hCuZjajWfh5aVfQDuL2MGF61JN3YZW1FAb/WXTVNbTbovIm4p
FFUTVl3iE/dVOSpLp2YTdB5iKl27mFUiRYihziKN2IXDyi64sp+NIaNkKVu0BuFH
hiypVXbeiZa+a7DyuY+wHv6SlFrVrjn6PBYdQqKTEwSpWEP+D4lkq3xfEcaC+cdR
uKlnCMcxSXHCivnZExC1PPpQJOZVOlrdgyuTHEGWP8bcM9lbqh3LPNYCQOQd82GI
wUmmoSb2DBgFvfKp2B135j6BzQtvs4BQIN9BUTvs4XwvEBLxdUwRORfpDjTJFMKr
o43iRsQcwu5MGFqifv20AmelJWA8mGIK8/LDO+y0g6XpZm+1vfUWEwAZj1aw7YE1
iCkaSKHgjCBfdyYjWSef0K9KqGDQ9yAgIyqHeoxusPqk+xHGF8bEJKMNGtvW4WBu
jFmbiNNgDhRCQmMgdxgZkDuedFWjlqyfwl7CCC5WRtk1F/uSOfJBHS61cPFPcZLy
UKIgLqJuoXQTF1z/gNzk8D0FolSoV7JQNRRdiVOz+fGHBk3Eg2nFkTTUNl+m+U28
dm4k+xySGZC/xHTqNESHQVhShKExyQBXNyWXDVYjvmIAD1bWjzSGwfKCHDoXUufe
+O30H3xyd2ec210YB2yb3N9QLnomL7ufpSpON3bYLoTeKhoWrNdzHBNptovGmiKz
JkghsEOeaYVcuXqiHyHr1g5XBrXOBVJSbf6UFiEy/g7Q1IGMH4uvvj+QqyoucPdf
UJE7COtRxcQ0l3v7IX/NWNzssDZ+DvgDK0T/6vUfob8Psmd/+7I+xHB7b8TYmHa9
6t0osQ6a8GXJ2l/ZRfYh4lYcHGNKd4EHIiBuwKRy7/XCV27JM9KwVqt7sahpoOgb
qK6MtnXoqf48oZOHm6hO0/GbyCv/21hHNVU3+e6uugSYnOjZRSeKuZ9Lb3ualhpY
2c5xULsynHzWRacsSdODpzWFI203Ebotld6dOi6nt11pgFF35kOmGbbMgFqwEq+P
qWvHK5DQ0qzKgbXqWEaof4osEffF+GOdsjusJZLs13BPOG2ukh6lELF5YDebCs2s
DYRQeYft83yhe69i75+tIM9lDf9n8DDZl7Qe886OOgNCG/DUhzbUn4r+ZNsMe3DC
QxcDOoEMePfIf1wt599kbzu32QvMsU2v1Hho5siEHTZfDYzWTVVqzZghzITNAJ4N
t6TjFVeSuBXE85BJspy3INFzlO9R7ymVUsDOPNBecz4LuTLH/Z3QKORXmxaeR+4K
rzIBQhmqZeA68boNoQnSx0jF+7XYTEzU6rdfX5EzvLe6vsLARloLIuyGaMVOrI0x
7CjO5RuPHVKlaFTTDGE34KcORgkK/0JUhv+ic8kqCSDbVKVl32VDLKTwMr/OtOWC
09kEKYsRv68Ok/oO+jXLOCfOhHG1Wg1sUrES//y32doXyFxPIUR0YHy0xj/VpP/7
Q2dDl5kSUW9V80HkUhRmSwWyiJnl+gVCwxCa8a5JES0EOxY5qW6rSP39xEHBbAne
0H4VjQXiU8uc3UG+JIbjcsyTn2hQ+yMMa29srqyH1I0xS8L7cIIT4wz+gEVi4+38
ZaSgKc7khMS8mqXnX1QC7XfdiZ5F25KufRWoytHCf64yu1J8YIzg//HuZ1uzUv57
BG6xd4FhfdqHpiBhzSN7xUkKtsmnJLqx9lgUdK/mMsr4KH0OxWz5kha/vNerUnYC
hwY4TS1HMfZYrYbsryNUA+Df5E5rM43gp57by0gqmSxpSSzp5DoQl/aVJIL+sX/j
7PcAV1GRnpSremOee5H/EMigxXx3dJJEOWB8k+YLXHX8TzbQXzij8eRE6Uvp6mEJ
jaMGzWF5hKG7gF4ovS+t2z6VYQ4DdjMtSns7vIvRaXt/Qop8l3Bna8MAhO4WEkfk
OTOtH0DMENYEfplGyQSCPEzK1OuQ1PD2w+KvSticsmih0IgE83v3W2wpzr6cWeJq
kvhQpO701Y4snfEQ3bJ0SukgTU5tbxi3zHZm+fiwKylUkIvPyr47BNVc/bv65XXS
YTF054zMULdOF3Fz9Kpr0mYGooLTlLuyKYFPvTubhBexFwJp8/wp5FoVl7fKUfpY
6lcKOQ1lGac/VatmE6o0QjfCsHbhQ/SBNsxnhkPUof9cJlaulQLViqybeBA+baFz
X/myAOG1NPvNd89GF11961L7TrQVvp5jJB6SKR4UJ9bFRFOWG82wL/kFvfY6ww5a
b/dYkm0866A5fBuB0HrBBsx1stfNoo1r+a24t2dG2mrZo7RgBF8sRVuyMW1WccJg
ArMnNHmn3s8hd2vS+1UjFWQWwdI0TYCzdl45n11B87CnTb6Ekogg8C0/poaCM+a4
fhMl/uGrare3Zhcl1slfvt6Rs7bzIWPl8lIvH1lxDNdqnhgZn28nLYHtjKJnGqIO
4WRQzDdWKRnBAxlfOujFkKmjbOay0XPMtLgViEUf929EQyZZxr3t27J1NHQPLWoY
+LRABdcnjDkooFfxe2u4VMMYVxVaC15PY/BweFlnbgurXeBfGQ+XAVV8IrhQExmH
Z7MiD5knhBxtfwcJLqMoWjtJAYBu/KNErposA2T4QaU/JdyeW9inHo6AOJEkkozi
auad6zAD023v79hO5ex+7iM/IDC/TXbvQmsSqa51pfEgLbtaBGCqWa7H6sm7aL7H
cSn4cC8U16A9VRkKpi4a4oIMm+8YKkqkEmODi8eWUClrobwDblNZU/YwAMhZ7Iyo
HxImAZeXva/a7hFbXgV56ql9/ZCFqmTk06ivBl0ZyOOEp2w2G279uEvfaerKdlE7
tkhpzt9Ph2OuvYa7/HpgRNhNZ/fGhACcHVFIVQj4cFkc+2J7egez+MAxk4xgmaIE
O3aWqRkbPPFmxQVqN3MYFeSzNd7X6G25KRLqCPmBAVll7SH30aHETxhI0NshimMK
Mfi3joI22vAR16UptdXZgd9Uhi95p+Uw5jFVtIDDMXd55xc5B9n8PxblHxAYMScn
BfJw2eBTGvWv0uemLUEqNZ2n0/8cYIFCfu/0ibPHGIkuJPBmjubML9nw/vVB798F
wuWaAV4H7hmSsQTDlf/+wTqaLKBuRhoRb18Lw0J9sjgd4Zv1LdGK4Zr4wR0AjnvP
bmj188DODbNWjIzZIGgfYYIPNhfviq3+ktbHwYaBoE4fyxZHjHUU0+krlu85ti8b
ykx+FDSre8EeGkKUeaLLVvZGbWIRYAXQ3eYlqTMv2pRqvVeNnWXmMZl0LjPzXSoM
xDmbOfH4/XnV4Gy/X3yxTTZjJuEcFr2mzVs0MaQ5db3yqG+4ytBCZPlyHBBVK/Yx
FAa1sL33HVOUcqNx0X/bhe8AwJs80x9Qfs3tve7qTy8FxOgRbHbmcRrg5JcQsMWf
9iZTuShmvNUos6jNqHP6eXKMAzeHcHqHWSKu5XMqPa/8YIw0qB+76bkbikA4uenB
V0q+1oWqBhBwdfki9N2yd+vlrg7K0AY82PloZ1yIBsJ0I0gnaAIYn0A00AnwmCEd
cQwg0Lga2q0NQ1Llj8CwRccPsPoh6Detrzuc/6EbojWutlK138IOSTFJKvoORwpa
yzkw56oFTXqzzX0N3oh3doxa/UJKD+xzMoSiX+bOmWzXvqgAakUIO6LMOuU+tIrj
LD691ZPFTsO3K1kTAFYaag+H2t2op2HuALlSxfberodXOdEZ8rcwLuYUegObFiU9
d6TTPXBtNWaWnH8gLTx7mgX1nrjR7Zjqkul6Ih5Fy+TjghoYKui+rEocNBCMHkQS
b9DG4Y/Wgi8dZGc2IBplIa1/olSuJwCj2NxXHj5CYo3xJiIavFPlxHAL+XQ6r7Pv
DKtFuj0uCbP6gTjaZmsvw72EwnS83dgEFV+aw224VduKyjZummpT/4p6Cg4UFLZi
7hUxjVcQrUjLETrZCb4UUfHrowJAGdiV4h54CbdGVJhLpF+1ekXMvGmZzw5thci6
7SFfVHtGzIIatRoAYfNAz0QjFIY1y0y/uSIwaTkR62yd8mKhHVcdaPj4FG5JeCir
o4XuDGrWiPO3b4gUGnHLomU3WpeuoqWTZCeUMXMibzHNAZZRpU5qS6LU2QjL8s6+
W1kXitdRIPvEMUFOVqRRCt9FTipCY2NTFbNxSBDWO8jKyx4Nuv5jN1iiMe5S6r8u
75w+T7NoGqNX8q2VcHKyv3NfLRqk5JqV5l8mM59dfynFSTcCAtyHgKZovVbNOhRb
Ik1Lk9zC90R9vkCzJ8dnbmrRpRnO3L0l9Qqw0NPkzVzhTTpPAlFGB8SJd7FDWag4
P0VepwuBrWgT+2C15oOFRPzULj4LlW5pij8N/arh+HCNN0UUfSIvnkmU+PKxLwII
qry7XNCDi5WsEfVei/BUy7ydI2aNJBLusyMfc8NoBpJ9rLFlDCrsSVmoC4muard7
KosxBTh8HSXjWg533zvbOJ8EmvR/VIKab1OUnpUmL1wzAiZwx0k7wyTrfN2ihU0M
JVdjaTQAYnIpYydi3QhdTqmvN8bm9TwElPbTBHK6GH/SnjyMoJze5RvtgRJ11+2z
jogVZAUE3mFW8of3SSAJUm5M1zheen/Wfz7FSYhquk6HGbDofASxt6G/Hbvsz0lI
5mlVKVyoUgUNihFh7k9SYKIOWz9bGUYLhVmshOvbjBnvE3zgtB/DDG3TRaB8MIea
9K+/JFoTkPZG4YlfVfspyRY4t0Uel+oPAKY5OU9KDDKXNnnkRy2u0fSx2KMDrvd/
hS35G3nng8e5yHxsCf+NsOXuyCtwQVoRq5nhZlS2erruFNYJ67f6OwdOWd7gu0+i
DI+C1PFCuFSNKfNm+jZ65hulmjWFyNpkpml17G3xYisE7NPCIg/GpOtfpwWtamjz
a9b1CN0a42zRG9HDs4MHMWO+7pfMINLGf+PQNGnzjzZs4As16iftmP2CHl6ePgSP
3kyLIjoabGkMz86aiNM9LmUUh41HHxuM4nwCOFHM7THWv1v4Iln/SXKIn2R5C7fz
SJHOCtBJDldEC8AErFTqruEAxpxRZpCEYCnFu/a8uo9gWSOyHJrNGvT4puf6as9+
vFcf/3ua/qZNjg+K76v1O8IQ9H2rxvrOpRBQimNTYMhXI6t6+6Z7P3K56PE0R9gA
ABiD9+YAU2TGNSuFdkKDrt7A7Ky7rRvrYaa9mufP8i1N+iCZPCl2Quy0QqQP78nw
AxsKK9P7tjKnrRncqqlOGDopXMwO1kc3NIkiB+IbXkTxC38Y0jRSHCpneRdpCrM0
c5GSjswLa4uROfS0tNrIRKA02QbQIL+Khu8BSIEiTNxjXGlWnwNGkMQ6IIph1LQ+
vag2+gruuLaPywb38gn6wbJTEVHyQn+rCJdOCY36zKoEOf/EDXKYPUOW/3byygSR
snMhW5cOnmydUaEdiL3V8sQE5vkTHYBpw8nPofh1GFrqmdD92ibqkprHas3tToUf
pZ3pRdcf4vEq5vNrBInkHv4ZjFIsRu+AUgvko1Koj5eQAlN0MVxW2fF1OnHs7Y6t
reOXYvQVAjnrov0JRBjPgFwp3pW2R0CPbyruMEItS/i08GrYk50cIK7aOAwfBfwR
e907b4SWl0JNYZabLKCmRfsG6BL6n6QCCKUTBMB6nDwdE70FjaCfJObrOTktn7Vv
cmmDIJhh6gmGduLvkb6W/vq++DumH+VcGVzZs5wQTkJ1EhfuiRRU++y1PINgic7y
XM+ybOmMLJ+84faNP/Gkc94MR7tWsYz2vMChDcgwWrY=
`pragma protect end_protected
