// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:36 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RX50I6chyO0qC0XpcVKj8ul7iLcnZwXaqv8P9GDEgzUNpW2FPTYJOmYDSlqDUrPf
3zQr5pCfz1o2dLQsiUc9aA3Wt2Mg5Jpz9Q3NzT4vBrEvD2OhESGNOy/S5HvhXc0b
qmLU1+paQE55irxSaG5LHurQTE4fhns46ZGTxQKjn4s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16304)
moBJHM6Vas9FgbnCib5qMUFsw0Oi4pw7MtxE0YWr1XMFyM2RdKhHZ8Wh8+J5tNzb
uf9N1eQc48yhiIf8zO64s9JAT6BAOOfNNDiFhMhYwpUQgFtXKXTH0S9lYfkGtTU4
ZxYEZdMRbToAKNxOPMxyFH+J9d+lFdWEgSjeK3CZdI1sCxt98zQOMYPUogHCou1c
EyvgegczD4KJ1tRZOhfZQay+U/+4zN84ZbaUEWxbT+XeqH+sjDe/ILHLQilCKJG1
dEGOOoJ3p2toMpBZURw8ovelEIbfjJpRPpoG2RQOp6eeOYZIM8xs7q7ezbiAJQhL
3kgKGbSHKjQyJcZPUVedLfZt4Q+FflOG5jdVkkM0uu3SWwwaP//yFsohMQStRlAc
FSaLEPnbnQjPXDEJH1tHkHiCKpn/XmIWz7B544YtoTLZGxKjqfwmGslAM5Cv+T7c
nbGMVp9PKhfIxoNmeC7q/EP9J7lS/VIRcbc+mrJwc1cvjKYWLD2+Cfmu1SCOMka8
zTyZqXQLdAIEdEntwUqaxuEeV9dm/OM9Uy5nSej6LFB+yjyUnmzjfwq8ndcDH0F9
9MiRclA7vCycOnmMmgmKyYGv5BkVI4e/7s6hIh2lqC5Yhw9YbkBperL818HVNYrl
bGTxeQwtURI0zXPRgvdHnQqsN9AS9wgbl1edGU8lcMRzY64LlN7HL9l66Dg7ue1K
/D4F7DsN1JUYQMv0t/5SmD3uwylhFbZeA9kO8uUdGuINCHqyP8eFaTTF6WOW7b7a
n4+mwo6gWd/SV0k6JXSf6GDw8Lczcucxt35Rt67zF2wsLewS5C6qvOVRU+DFM6Nw
npGvUdOTq00gaEX5uj1QuIongZZIii1M5ohHTLYiU7Zfw+BR04fYAzDagDfjwnW3
DQH5RmQBOWIqL2Q9r8wyVRwy37WaAaWCz56IHHpJnOyDXd/b/Cb8QeUKKsINACWU
bT3aiVZIRgi0b9VKzVgCmHy6mh32jD3J27fgY2JB3lRQvs38JpxoObspVb3gCHxH
fTorpJZznAGWGjryqsgViy9pV+0iUMbXE/mUk/7D/9FO7bU8rt+ndqOkSqo2sMck
sJv6h1wEYSo7gROGrBfnapMhgTEkCMOESZJ1o6cGPRvZKiQOF4HZ+6xJkn8myHrS
1hZdFg48vEGHDuRW4Lmn1mZq38eK3zvBJDthJplFOV1GgaZZqoUmUkaVjkn9kPJR
l8A6SyV6D+YFRUGT0C6gnR/MIzk7Bf6Beo0PdRYcJZZdW2StEnYjemgL8qlKHEUP
YWe2h2le5II9ZN9Zxf+eq+/KbeCM2AJ+42DWiLCN/HiqekH/arubkq6kIF3KDyZD
n41gLnFm/U+1moSVajw7ZBvc06ubw69a0SfttorDH7dxnbV+iZg8imJv6QBgGmn1
Q1nJxYbcYNaHtgfau5m5qKKiJX0eYdgHt8dAoKwQ6YiIpso+N2ZqVXRbMoysfpLS
bzqmsnPghuE8BkPrH9GiekvypX9jdfsQi5LuGuoGTIu7Qxt3V2yxX/AaQtGF1LOr
eX8E3fl+oNk4pJUEeTp3WHAHQw7RR+FxwiVYy0J1+gDBWIEJ3P6PihqU24X9LQiS
BUG2r4Dt3LboUCVFBc/hI+rk0rav875QVn38ZA6ZDX3t/D8OQCzDiK63/sPpnrVy
RSptgkPNFR4Z61fLiz58yIVf8zpuONeLXMonU+doHBQZHy6Cdo67hzRKxJeEDqkQ
zbaR327nzFh7DTsL8kl+Fca6CFQ82RmXV3X2O7sa5liwT+K373QogmEER6hTD2Qp
2OAdmj0VAjtEICrD0XoCuGSCBcLVC//sXSo2h1EiSXlar4enI16J2aHMDVdunJc9
tJ/dL2sKgcS68/ZPIC3pxp94by4WmoPFgg1NMzDPtl03UX2byRGio0q3wJIcJ382
pDSOGey0AP2gki9FE01OvwbF/FzPWDVNEFxqGxYKTsvsd5g5tMqaQiPxJnvVtuQT
8LV5Pba4BrD+g8ZWNBDFE9JCDeT3ykgMaueZv3/ZNL2Q5eNkgA90+mi7CDJHk8ex
5s2CNEFjfS2ugoXAh7d01wPORdB5qGOYIVRqKW4q/MiNg47Io3tiCZ5LoRbIrBE7
cqwFso0mguV9sNx7zeTF/Q3RndcOAP/ypiJ129QBr/DJkjzho0B8KJShx4nFZQH4
aYwnvxqVpCeBgBpB09RfAOiv8hjcaElTm4SHm5mPwS5mkezuaIrsMD2FQSpg7NeF
Qz6Nbj7DiYqosC+63MBnZ+therkvBU82H7MI70oHgTZlER74Fr75A4IsyUqHNrHx
Q68XhqM4IbYU7d7XLSitMz4bNr7SchkH+18GEZhDwDaWDJ2YyjSWxZuAEITi/heh
Cl6QTGoAF6KQ7Qh2b6o3bJh1UYG4jeBKnxISnyNVNQXecSb/+NEtfVgtBbKkjCFZ
tvvfaua7SSKfFMVTg3fQ7EjBN/HLBjJ5INyKJr78M+O6/F/jZL4Vj/tM62vh+vZP
XX7K6BpErlmaa87JrQ8kDIJ+75ysgD+AvjnS/L+3f5+lpm/Ye4cQfdiJL/c6cGQ1
XMnN1ZqomQvD0InPE4umHj/LzH9gjbV86t0cb3eLvn8jZAVPKful3mceZAadhYvV
F+aVWZryELv1M5UlZ1ccGllgvFUCHzA6O/vZ3FRF3/OLMPWABSjhpnwbwAPzLeI6
lQvLgfE8zW5Gi9iGoUQZkPGmEj05IyaZWszH9bS1FYEDaV9jGQiNNsstjihRKBMx
zYDKE0z+H3jSvdLuf8IzSOaSI+re1WKY0urv61Dqf7itIxTL2Q9v3gphdzh1ryqH
fqOinD6Bqu8+xahfHwnNgYZoTFkwJL55R3NmyfoeceCK0rMa4PyXOf+Zoa/goI5U
+0cqkjV7E/rbfvogSmv72GIZubQO+2Ze5OQdPMCoATQ2zEgUN4UOsAQcTfovcpIa
G+q5H/1EPUxB8ctUwoD5aLsuY6XCIefqllUzgxJDyQy460Vh7d85ZUPIiES5iRVf
nNEACIpDSBNhphDXtNP3Yjo8hDSOtXgbNW/HKoK7Gh48CdY3KkR1Ir4uWr8Rw2wH
vPhigtWXD66xW11m0eiXTyhVaAScm1guL49eXqFSJ9iG8orYCIiQBbwbbtunWwef
EDRzDFTp8L5X/oAl+aNx/sNigTckz4k7PJSkDGonrFT4yB+GMq3cixG4jQJiChnG
4OAWGd9ZewM1LWzpZpJ8WCQQsHcppvPhZhKgkzTJMCO9PkVF5bD5fS0gP0dLY+IU
QBdiYVErLLFOlpauB25Bum+4CoQh2QQSK9Rd4qcPqRcidazpGxzEOsC8bwINvU5+
3kDsVly309AjxIxIFBilNvd3mnfSvnxZivfpC8NZ5rwJjgmUPfuGx8IFFkzev6Cc
G6Yt9b14GEugxO6MUQ2UsXnwcDEhyB7V108nKyXpnIBQir0XbUw3aRpg2l5Nj8UZ
U3hxzOJ0nRt/nmzomYxP5GCT3bWzjMZF4PxeriG5AgLYScdmC+YV5E484XM0yN6w
5e0/aVVg+LAFx7BCV2k01RB9y8zmUhjjdsyM5DRQQDSUOPWWqNb7dDue+Fgg8G0I
DdYwIwE38gNUH45cYTBJ1PQpaX6h90h8Wsu0kRBnNyRCJeh9D/JQgr1xsBQ9Inqz
ezGQgKBL8vfbf5DexZ9NgCUSZeCuJHkB7b8XryTkxGY/khUb5JhJwzcmhk2YA82W
BxNWtid6KxZgZPilYJ7s2kSO5OKI//wQ4a93eKd//XIg8MIAvN3jSOnCvw4Lt9rJ
2RffovPFOIS/00Ppf0SvbXq82I7WCCQU19r+5KNjv2vYlHB2hSKG1cda6ebIupD/
xmItJm8Ner5g8axsN+l2ZgJye/G+IYPkzKH4+bRL0uSPgFmUQvq45gOqMhbTfDk1
RwYaI36T4Yjn1vALNLecN5fgfaidf8Jq5/BnWDTOcrjZ7agJNpKzxZySHyOodvEa
26tV+IAQ5BwEtGHBZAwuzl0pdinb4cvT3iwWjvgYBOEOaLwZgvPuYGfOXkhzhQSd
stvMW36bs7iJfJPX70X45sl0+82KSHqzWGR27sKgpZJGMTIM8oNK1xqCyfqHTHlW
SqACu2oiGdjAd1hKvGRXI1McGdbo5JFWtEJYRwScZ6j8FlXzCc3V9VlqMBhRW0dy
c7PTMZ1ePyWLtNTnRkUZo5KpXj9sLv+MQLMBiV2FTrYmdEtmrN3QNZzIyNhGAhlv
9G4LyZhu/s+P7tQGB0O1G2jsewCU+WUB2zOMQctQptqbQwkd9y3I41so5e9aRSYT
146/02R6i+o1eFVgMeEHVxzv4/rACqfzL4V0HuTz2nB5slVFwjqPo5sY6ZfezeWE
jGIlsZDm5ToqHqnugv3zXnabwcb+dBHaSfS5dHzAL4cwWP+XekrFZ/W08lS08/ku
zZODb+/9CxEV9oT1A+1HgIX8wArEuCyKLLkdmC764ZqyYX4BoDpP1YsgcDt92lax
9vrLKC3FfncNkmstwT8R9pUKf5LVb3/ysPBwbsnAyQ/lfJZk9wk6ag9/yhQ0oQS3
9JvMAN/HtLdrS1QDPCfjJyS/2KsPCVFet6Qypt18BZgx1SkALLa0auLhbvqnmeMH
LqAsUohinry/eqgc3OFNNpsHbkKqy+qJVnQQObaGMtgKPnmajrAlsUjuQW5gecT9
6B32EBMeU3T+gPfGT1c5NvUGIhBlcCxfbwCpmz7PVdaDXT3hip3RyNxQWBwZV5dU
ERFCFzcPGRZCYrsORnOztYgtztVzjROKYhE49BoeOvaNPfN3dGp00LoUbjYrbXxk
yguKqRMRizNZcfdbQ/7ICDDiltm5feCEUA9j4tuZAer7OWjdPCSZHOKvhyePDGn7
KhqSBnXnAr4esmfU/zJaKF+JCgGSO/jJc8eGGjD/RrKNIONhwGp/Yf0NrWRvLezR
F0Y3tAFGMC35i5Ao1cKlKO8OM129l3mSdYTsEd0E9SqqNWavPFV0/jxOGoWGOHig
kCpKONmwOkW8nMLETD4TfVUqBCX+dKUNAAJg1huHpRECJnATl2qlx5vszJB7EqJA
hAwELU6MnLBh+zn0T6RoX0xx7M+7KCvEjDgpyzY1r4XXr8HSYrGZldZNqafPoe7i
EBGmRRivrx/ED8QDGTvfH7oW8MOF8KRUeu2afDdfBg8sH8KllvZiP524EV3igAka
MiG/sqNWQNZTkG4y0cqQGYzyQm9kSsTzUxoJTQqEbZxHXzeAyChqBSrFF69BIjAY
NA5li/Jc1kCVC2xbeAsFSvL9MutY5JB1WYXz2KW6m50Pj5x1tmxA6/QOXZlTt0Q/
d+TLV7ilamQx3gB3V+un1UN3r6xODlxEfxWmbmVAglR81qtetqEq+m2o/URyWxce
dNl9zIQkEDG8DH/WmK93ksjIsL3Yl90/DEQ8w7qCibIx1NSgYvKgYke1n5J1Gv7g
RD5HVLHX5xf9CGOz21wR0O2WupuD+I0mYJiXbHSTwgph/0VJopcFFmoj9nZ5GH3s
DAe9J6VSGT9BvJ4EEOH1Q3Iex1vMMVYTLfpbksOizRHfzZjuHUaiygaaclbCY3yk
WZfoJe9t6dpFrTmdNdsx5h3pk86OCXQmv0Mwchk0m2FiDMlblXuhJFRwSbH23DhU
R2q7Lww6ge8NLSOATt3EdlyzRB6CKyZkpsk7ICsZX+AEn4svOs8EKW3lU2Td1bcy
vOXGqLFGiskt1eZLF9EGP5eVDHzQEXWeA1nLy0IMKvECkaIhSoqzOD8k//M1MsyN
co6YBDqC5rgbd1Nc8PADogJ1Ce3Z550FzcxeztQJTZFtagmm8vGsLmhDUi9AfRMd
YVjcL8iJE6LfHjiqi1GIZcEcwtUlEUmE/up4X5L2Zgaok/uzLSIUx90ZLBC8YF6g
dpXcG66zc66aHysob5k4Bvvdv24OT8BYj9x6TZIDFKYvRIcR5yOgph+h6QvCSgnC
ulyw5M8w5aLUuuC1wk8TznvmqTNjPz6w6w0QkV5AYhCYC0iL1fc0STN6BGggb79m
FY7WvmB1l+FZxpyiByoKOTafP5xJBC4/votf+b/yUXFDbdzuZ5htb92Iej3ehFcP
PdeinFk+lry77JPmRl5x0vEFc0E/azEJWzJ0bpOxsvRApIF16Y2QSASeoO9UprbK
3Ndm+rDTo378kXvsKeXGGjpB5r2kWQA6KNeLU9PIwfqmTDbOsoFHinOqN8Ctz1cP
I09NxA33tD6pZJX6VLNsJ7qJc+H9XZQFbRQTNHCuJtIojbRX18yF4I7KMtg7kaTp
yHvblKLAwIvyxV/6L8AmKr7ZQK5g4ISugIbAvDa82gpNgvx4G77M9gKGrqrUAkoo
L2Y1H2mCCvbDHt4yWwQE3ISdJWwC2gXUxLl55sDQY/FQnZBqgRpokvu5os988jmS
kZv8Cwvv6KL5O9V/XZZ2wdCRPY3k+kDW3RadTK/ZHz3FGKHpbN9rbA0b44YFsgky
w6WV+7GL0mLajNxCbqKP84y24c5GSrgXE7yUgUgPVl3PB5cetu95oAbwKnJ3vnpe
wRRasNRhFRIPcSbPdHqxOVBQt8ouifWy2KVDb2oGcdyyF44tzvxv4pDU5x4oin13
GZMDTdPDe0tmbDlLZULO5OY/DDhX9vdCJKtVV5CUt2Q5jc7ASOk8Kle2EojnnaKk
ecrqQqmMjciU0XYV+/ekKXuZB7RXQCH39IQAgZFvPegBkaovUzcJj9wToA6zbSOm
SJmsAM1tMjoVKoGYM6wCH15+gibJy0AG/f1ayIzW7zuoaXqkq6buv9vugYt+HQJs
CiXIIKvymJB5rHYC7q+sWsTEzy4/JXgANlP6XEF1DoXdr6p3KVH1Mgqnc+SSEVi4
hk3qHthb+V0VSlUgZzKyHIdEojpGgRJnduAPZPh2wMVOStURIdgBouQ5l+OjVzEr
sZxpI2SziqfdAy5B5wUbygohq+8S/d+cins0t3dpdeA3LrmKY1CZF3+iLekONsYg
JbJDxO8G/r454liwVLYTO+rM83Rsx6jiKo059eXVJ4xrSWfCo/Hk4whtSU9+ee0f
IZhkj9ndQjwGu+N3b1jILYlIUKLM6Lxw605NLG5MsEqtOsmhE4xkWJ9+R5lsH5DU
iJbf9ddIeO76AAQRZQVMsWKl58Kqqeqp0xIukHlXvvFilLyqOY7G7n/qNN5l2IV9
hAE/Pwx3ujWCimFbohwY2Zpw2U+FGx9rJRewN6zObJ8nh1Z1IiaCVbBa58TlfzjD
Ixf1f1GWQ1FM6WkyY2VzHg9pMT/Mmw6beaGv1VAfUB28Ldy2Mtdn2Q46uH0lQiR5
T/XxXccyZPnVkZ+4I/20ZjqWKAlrcTP513nq6UHgw/o1MD+NTp1mvSHpj5TRloX2
jPGHJxFzLBB4MC2QdIQQycI1oi9slU3/+ekVh8t9iblO3WfGO9AU4TDey7N7UTvW
x56BVaCxyOnE+yOgxkw9BZE2ADDJoDJbz5fHnVyfYjfStAY4YSDjI33MqVCfTi/p
352IR1Ru93o4qIAgaiaQOjhdP2Xhnk5E+/nOyprpDj8gcglYWdlRg7a5MjRvjaLQ
TkYGg77S9VOTJYU5J9Nl8t80sE3j/o84gA/y3Ptew7ejuLvvkWzt0WYMTT3xdJf2
kp9TLmlMU1z/1AebuJkD2O92i8YhlwYRe22vsxP3m41Mm3v9D6tql9zhRzhiLzOf
hc/7pqTgkOFFneMPecD+lnYYq6Ev49Ij5/Lr5Kokp6vuop9L/aa/5xu3292I6/gH
LFyDeDc4sQqRmKWJXvq7N6ecfNn6KDzJGjdDfHCncQECwJS0FYcrUVVfP3MthGkL
e0SGuCAPIjQXElyLfsvGCmm+HyiW2AeB2q2prqFFHnThjpBH+8jQw+UNZ01IWXDU
gHk5S7XUnLEFiVtoHqs4XYQtcW0Yc5kopv4GkAg7uQM1FodbZHpg/J8k91Ip2YUP
nHXSHX5nxLtW4jsPT47F97hdXqXt7oMZB3O5/X6cXad0Fd4JD0+JEJ1ZjGKe5sTK
2LOZoCsAsH2B7FIcFf+4CS0WdwBCrbGyKT5aORyKAlLP9vuc79X5IFcfxP0JKs65
csXZ9QZoGcCfQMjb1U4UA15cst7h54F4a3PEAPe1Lr1HltIOFJEmevgZzNylIjwR
VGt2CHBGoeggkrG/GnsgDYhzdrtbY6t/wfM2LvG959qBc7Xe0qslaJygtH5m4l1i
dTcoQ3DUVcgbvUlsDL43fdSXrzJPV52w58xklWXGyeutEoMzIg8t/8sTOVTRaFX1
NprprMXKuOftUviqzccAzVS4RMHlz5OT8Spj2knPsOVcCgNjVxIVh62yahL43n6o
CxnVG6hsTivxWI9ZXhSI8K1K/D2cnq8aIVJ5jCRAqbC99pUuujtXRw0GaqGEjW3k
5SOAKW0Q4BK7q4fGHCoTlzkQ+lO6su0rhXMeXKGHKcaxu/5RITew/5rhR9S5qizV
nMaWYY7QPAgGuIUslk0U7UqwLlNYtLBo9hHBsmQPNXDMucT+nnfgsFod69Fjy0ve
Til4+bOFaJOjZSSf9xtAxJEpMrrh9gzhJ6vWyjUIa7E8GzZ/JZ6jli0gBqiI2tR9
CNKQNdv/8wLFruhgZLZ6xVMTFcJupEbmRjRl3EF4Q2uAGb1gLEh7A30wW5UFdXQX
Hk4n15mScMDtUfDCgKJ8U/X3S67J12LERkEnah3hYrjaSr1G0AhIiin1PsXeG3Fc
1cAdIcb1sDeN4lmnyamaNOLRVgDLymK1WSdCOQ4eEiRtL7gFwpIPK1j1fwAvk8xJ
N3FPW0TFloJyc5Qsa/QtFbNQqYCDIaYdKesAoCVG/RFgp/5rj3bvdRFXjvuykc0o
9aZ3SkvOR8yQkkJbvNp1uIGbNN/lh/d0dmyN7UxG0hoWnwuP0Hyv0SOZdXsIMUJh
ZRMrK+wvuio09TODiujcRqOjaWbshNLqPvBP8ckwXLc0TfItY0kEhXNPh6m803MC
4TGs15f5iFs9HKSjUlcIbkj+asQgmY+5BbWxEDqmkpvLC+mQkg2xqafsddd7LXIV
qWLxRpapvPxrym48OmYLz628G9BnvSNdVfTguFckLiTN6ZpXYtZYFyB02r9jthqR
g8VPKDbEPb463DqXuMdRHOVQhAY00vvclAdlmygQKv3xumUH0KokkoTmjM9DT8A/
1Etf66kftRJXlBvuWbvHOi0HxIM3R/hv0gS26SC4T5YK14+B8pLRctrYK2PMg2/V
tIqjT4RsA3lRjIuDVT3/g+os2GBxxfWXpzzQBS2EjytMtQaX2XMhIBSGA+sCZchL
uAnpqmdhebmBpibv6DrVAVlCPh76eGbqy8qsocig4qxK9WqKzuaNNcrQStM11HiW
6LgtawkKbygZGw5U7Ih+zAD/EmppG6vzvkBmIo62nN2cIYHcsN9PT9aSEItgAa4m
+pOwqGak2QFKhCeVhxo7ioHsl0gnGjrUK47Hma/dQsPUaXIFfThs+80Nk66cRq7p
xYkdtu9ngIf4r6SepGfxdF0CiDHgkItdHx0vTlRDG7iJqO92qTPnlzM3E+6rx6YV
jshYRmbECMvXqk53xs+FihRpTzavRPq9/QcgpM2p5Fuh0OD7Yb2rSE0g0Uf7OCuH
jiQ+ilUDwtEHge4u2+GohBccX97XrnxqiNax7gi9ddRnm53BJE2r/kdildJc0Qgg
wsIPCnCiHPVvF+mmjiAGFdWACIIl9aMnAqwVijn1vPXg+4GYjNdE6CTKAcT+1n1n
0HqqkmSD4VhBSI7oPX9ayQUsy8Sc8SCCcCocnsfkLHkyP3YAFVGaQJH9Dcj4Qxsx
dkGiKPq8l1QRSaCUP7/FsPOrn0RWlCnKCo8L/fGqg/4BDVKSoiC6yggxRSTce20I
w7OuOgWtmkeS+gZf3nqFfXzKD22X8VuOq/uH62woer080xGBpEql4abTTwIJgAlg
QmbgKuTKzf1G4xMDupRbD7CG5FL3qTIPQXgqnzyRXvck4X/oYOBbSJFl1gozNQmY
UL4JLbFnXRywTfxwKyZDse+4FbhVEFswzc2/voMAYjklj1tyek2/Aphah4fM8+pK
/hcOTUta1o/E+EGIoZyEDRq0rMhIsV/3cFm5axemE9d+1rtvA1wgmKxqJHTcstYB
h5pD8kWyM5QQ7WpSlHuREKbY2SxPA2k1v1Z+W3eNBhWX7UJ80WfnukfOZGhA9AkW
jBhfH9mddyMSFgDvq7ExJP1EYH8H2sa4sluLc2zqsbzVUH3bq/4CIPJP2fyl51Qt
9Zbe3TQSEkn54RntadwWbv3ExBJWoe6VtapNXKGYvUSLE68YLc25NwRH0jBB+TSu
1ZPAhN6ZJWvD8dTmsO4bGOkUfO+oqzfJqtgKWjhDjQCtGK1hvKByfoGvNdqSx4b7
dGxWVy30JbxoQ0oAUbCBlJqJlZTl86aI9RBHnNVqDSvUVOscj5j/rjrqYn29CtU8
4O4AMdX57pCclyBJuwbQFF2zVUL+/qB71hmiyScxQ0KqIt2MmrnH/QQRV2hLUSmb
7DdT5WIcUSSELDU6me4rBc2NFXVO8it4GquYPgB0+ilqAET4QwqOdVBpsYEE7GpL
VED8JG2Ymho2X/5oUkQpaCIYIK9VmvS6A5Fj/Nk99nFW/lmfqbswFT/cXSjkOKIj
Vj/j7glIuwR69cBQd/pb5CBSoY3am9e0GgQ3j94leF2I55C+hv9Hgl4eSzbpt1tq
9Xiz1jW+JoEyUyaUHmRrPHhzZJ3G3/ca5P9n4itChTOWOQuWXGpFr5g53CztC86i
+x9TGrSAOlYEvkDxZgXOGs0wdSzf24/EhAKgX6nUvFs6WgKjszX7QAis3K3TM/0s
pZl6REDwNGVt/lIgE/J0fKZqrnEibOiHrAOEgPGihflgJsi+Lo+1JCaIVGj96SIG
0m0YO0sovbSeCX/p+TDNpQjE4h2xh1TMY08oqWoMYZjyM/k/scnEz0yHq9PFVue9
YafKWpgt2yHXOhd75l86w1PuVPIW2pCegRhNxSYNRsKAMOKNhkAs67gKGD+KNuS+
+05qqm+m1at+IZ2zO2koFWNdzh4rjbuPMOcIADqZOo732wrlMPPQjKpEs/M/huS3
b4a+Rw7aeZVT89vQG6WbMRCUdAhpVnTRMrHoMcpBG845n6kuNW8b15j21v01QE8u
uj28qhb0eG8YLCaAXgQddZ5hqg9oP23a7sy1jRQBwuuCnAs9iw3Zu5rooqpPwtpW
2CNQXkAe1AEfWj10MLrQQE+CHlF40gY2jCgfv2VDhliGbIHQ8jsH4mkoMZJnVJPT
6vSq/kpIo3kKXoZ5XRzrF876kXojt3KODHk6PjWgalwoBrQAlFg20dcVpfZjUFxE
E1YHgKhcqmA7WjG2FrO0jL0z0cYkoXiZr7KSOrOF50btNTe6jz7nyMClztv1+6zs
UO7fRuKAgQsdhychk+oe7Gxgdky208pL+yDIm3lCWjEcZMXx69nxuLMzKO4F5VfC
0qlT5amUIY2PxJcx66rnQBz8i+F+01uI8H5rvnbxwxiVLAmjXH8LTQDaLyllG1Z3
Q7Z1U6vZ/FkJsNf6LRTwhY8VI09LEgufPQmLz6s9yi7WIp1tsZ0+C3j8kpQUfbHv
HgmRT6BL0u1+yQnSaiWpuTkYxcTdhHDrUe5D0i4u4pp5xzBAiZaHotSP1rrE/mfj
Py/P7/pnHGah9XGe/dYOJNiG/X6cW0UrwWDKpUgCdtxJ7hPPysiaQSfEcjHEFa94
wDUcwhL/FJCKiiaJw3XNM/FPWcPnYZZQq6bfAHRX/niKTxJMwY3TxkugvvuvQ9Sw
177QYp3jpZHdrIViXjazDaxB508ZJua62bS1AooZR+/hPbJSSrH3q9yHl0qm/fKn
OOowq5k0Ggv5UvHKeZk5v3Eoog9BZo+KcVLTR2bv0Z6HRBgRFjCRNDdWPfr3pjR7
feX+86Mgy/uB4jAbrcVq0Wv7Tyl0Esxp1BiaIZI1z0DBYuG+Ts3b6gzvvn3dYdi8
wLK4yhQSljXRbqlD2ziWnepHBJ1QEujGIeRYU46ea3aOTR9Ngg/EG8CCNIeyvFdR
DCeEhksosNzNhM7RjBd7pZNHWCy8Csqopja7G9tq+LS06TnefsUS4jkahHdvC03r
gZ1zLgZlY0l+y4tdeBt17BZNE64dg1w1QAnp/gEgEPWcSFl3/w6/uUSGVS/iWfUy
vXUce0AegfLkrMmIFJ7UVKOtXXlF0pZPpL70mbfJZfsH90MHaQJfXtBy/BKlklrS
b577ywrAtAiBSTPfeZrS+mGPf91KHVUSAo978TyXZdAh6LjEn73TzGYaOIs4Z6+f
Uf3u3um9RKCEXoA7dxNMnptuk60gufSoz8ef4ADx/xFWWiJ02vr/M7csnfKSUcf9
SWqtyEdHEn9RVZXMc1S7lELl++axzNUmak+amBeB4sagSe970g/6M9kf2u2vDSwR
q6BQGZ9inqqosjN4vi/+SRaKijQ4ffpgFawBlBX9+W50ue0pMT4s6Z/tzZg47Rvi
l7icPqNzxq7JfTqv1KlGBGI0EWA6dJYMGzdrIXA985gVvqz7uM9rFE/+ix7XlSLW
vtpyjcevEb4tkx1IZVyjhPf7UfdO3h0XycxGQwm5wFZ8aU8nfE1MV2TDYw5WAiqD
PrQD+C5/LK4tphv25/3bkHBzPCvcI6XC4ONBa6wsiCFiFb+k+WVSe6G9NVbR4rIb
14GDCbhnAF1Vp2wjCT679mGCpbhcJzJuQCevOB18zEkX+93BPAiMMSdjeMDvMXlu
+m/+chrXXL2VaHcxtKgisJqA01wHARPQLZ8sQcqJe/uV1d1fPVIVC8qT8qKt1feO
kHS7RDeF59mmXPYgT1K+/4pArCfPWQat0X38njPmQuRzUmJ+ODwFQniRZFCIfYEM
fMfTrt3dl00IoVqSEhQr9Ojwd5T2ue4FcX2iwKSErim4FnqlwU8Afot0IPalQpi/
pH8DbkSAkG50XIqYP/9IYQpHbKcqZF88LP6LaBpoOsy4BZIGF+N58rD7eonfmnCh
rEHiVwGxtzmoSbuaZJR2lblu7vUpUB0tMlsWswZ3JxPqhZqarTRRukLSF5X/DbLN
jVB6Im3wn5TgT023yUDk/O5Z7/mCTCHBqeGewbTaLP81xA6tHovOqQ6qQ1MLMWJ/
ijgu61/RyZZSvW51uKR+HMT4AQ/wA8JQOl4gygkSA7hq8df621n6/Qdo9HjqEJvB
DZj/c7OTcsYxbnSK6SohCiynIEGwwWrTcq9xkZSO5WfStAz6U7kvJqxyWq6GOS9Y
uRhxaRuc0oqKy9cbxIx2EZRz+IGezjO+/OTQ1CZVMWyrIVZhOrAbuLjKU7r/FISc
Xu/05YwR5BNJS3vLcySCPAT6rDME++nKsBG62PZhWWhDuN/J0PoS+q/nJHj1xO26
f+yzIZOim0tTagprHtCkUdrfFT0a2tUM32zbnX1a+82++EuJdLcnYxbMo2lh/cyu
CxG9PuWvDBlmnGYnzROxtgQGpGsFzyo1CjpXrvE8rFVRXPgMWg1P3IRTGQkErW1E
WEUmxfnRy0NxxkS+wxo0E7IISuDb6ACAgAeHD5yGr6RZRSRbvvxjzudRUBck8jou
mmWUg+PuVS5Jtn11w+7NNcG2euHoUJaSqXTChXRJuT7hMo2ttSsLw03yg4RAroxK
B3BFtrmQzu3PXJvOOjws5MdxOIAuHGKiedLpumkIzyq+3NjFaNQLCv6UzN5OokPA
JORcCYVAho/jkh7h/wjmr3HADEGnvxWIejHj2iyNd+52791xPwkNT+5LXdu8zYYf
OP5xOW6fTw/oakuLUMEFUtrvIoLN4wWbGruGZC60O3pW70if2s3tltO+rQ19LM2o
n3/UGiG9N3Cp/H4ceUx7eYtlHLS5BLNk6R9dgo8cfZ+uYI4Nn8SIx7ls2ztoucKb
HTELxWvzWLsRITORWuDozJMgopKxukTaX0wg1Qzjej6Q7nImoR07asnFisOlyYd7
mMPsu90xdi4nvtL/zrVQ8RTdyQ5plxf3mu97cTiRRfY+dXXm/TMBqqGGeuNf+0BB
Ncum+RYKRl0TqPVEsFYUs2MyibN8ngA2TCwLgwxWuEPptDflJWC+RRzFKKwCgDdv
iXvawI9pGuIoTpsC/U/2OufTRElQlHu8/mcxMZFdF7/RAcZC4D/Hp22CLCocnu9J
yvwPbozWfhvH1G4NcEGGVIxj6lSclzzuguQElCiexdkVawfTMNvdFhTpXdatn5m4
l3aLo2Bhk81rzCEIEAgViLE3RC06i7vsaF+uJfiQLW1DzEcD0EWoEDdG8MOZZe0u
nf+4QioiIf/c8ABfTN+4yjykANZtEy5altsh19xNE7Q7/zv4R2rjVEogod8t3MCD
ZmqyUmTIPbd9m4fwCSlFj/JH8d3+pIXY6bpQjN3hiOSGa9byLTO7j1IL1jHWUK52
hkvq+kMwXVFMaL58274dMVIWXxO9/cbrbIcXVP6ghk2X5z2goLteOPlqkmZaP7bI
4X8PlRSY0Pm/xO7EcaRFBPKjqn0Nbl1tss/ZIZvqhNKDOwLfS+IQe2WEOTh5azUe
ci+BvptWh+5+SHUaaOX/wFylsBF0TZXWG67zCWdcZ8Q3ruDNfUyOd/tKTZApNhOm
YTkLNnI/i2vomHZI1XmjLogzR1fvhZNOAwGhJZmLx3p6H2yRSeNwAn+UvNPl6O6V
PQtuc454YOh7BQmtKaY6aciTtW/O7yoSJwC6vUuaoKD1995RiNJOcBPBup7cNZCU
cGtUDnXLKc2WQJ/M1Iy+cEGQgls2SuJZ7usI8SeleUgluhPkBxqTuosyz0KIjHbj
+rb0csNaeRPvZv35xoTI4eyErS9bc1SxB1OOrbxDgc5d0S9Z4AC0b5qrdxAPQ6B+
Ylz3+gRPkRU6QqWdRwILHSfwgL3kb7kOQGfnVjH5viD/z/xKJLn0KYB+vyXK1eT9
FMpkb5WxVEB4Eqt7T6q56jAtdc/8NIVh1Z1hX2ToEbzx0Gt+ApNMxrcj/JpliXbV
T8qFyAJQljgO936HCOHYeQmwTJ67kCEOvHkZgEt/23EuiT74sJFI9+0+7nY3t43N
e/8vlFuku30I3FbyBNAuQkgzAMfxKAUUx+k2Nh3Im9uJJjJMLz5hMumaQwtJPlnY
ajYb4lTYoLODsuS+eyDKkWQUmaudkrm8XJ4tlFqiLVpeOf4OjX7n6WwUo5mYfxMG
1zWIZBOR1NK9qesJUDPTyREC87RQB98YyPisAMKb6L77hVVYugj2dFI+60RWt2GE
8q+73W8nP6+wjAGa7/hxHIepTqtiNvXXB2H26cISAe1bQDuq7EGYkZL6qnMfUv9e
JrMa/2tQ0l3n/PXtjYQZjJ+Ho9c1+2VyMkfNzS7UaAKSBkCT6wsqiziiQSPX0Jqj
Lo0VbVw0OvJf85KFfcnG+YhcYGjAWxzs3cfRKjh6Pnq/6VHeOj7LCVhAGVzA5g7u
fHM5d3DMfv/Mn8A5M8gNtNNEZVjsJmCxd0rIlPax3+6MvMGIZ4MbNv1ObNaL+/0j
AuBNFA9Ko+YpqVtoERlYSN9qny7aVGOnrdRXC8z5PoDOQ7Xx887pfKJ49QFyJdlP
fi4NumhuxEs6JCR98SK0Q/O7pSIC436QztG6Kth2XNQ8M/VQmRq04ZOcVZcF2EJ1
PLYm1cRB2ws3mmPqgjANrqJLVO5KAKhr1GA75N3+GY71ZANZK00TPEHGELxydRur
aI5nrs+54u/jmS3a+l0Fd97Rxya7HI+r5nxUXlSDOcvzpvtA7LjJi67IsD7U4BSy
fG5r6A0JQjB1YCl2dyliQKWIGIUzLOTVNjR1rWxkwtYoXxSLl18/BDLiHUlMb7XO
UelQoqnLC0vGXtiijJZUSeWb0A0YQGUDfvlAafOjHpnv6jh183X75q6qPGVaYYIT
vYFxC7SnEkOhdbblDZQjhPLmZQv2h50yUoy7ZaMdG+pyVUelVsGkBMo/iEHRnpQH
lwM4MhE3R/+S/HX+0zKq5iscPgXBEbxjrKJTnzxR2EgOt4Hr7DOzCVInaiyZFgHk
5nB9JurW/oJS81aj5YnaLeiK4yChFovwTMom7kYxsWmiW/GjQ5k20U/OLe/ziLvD
p2Cqhw4qcWEtoea86JEK+PiTwIQtXQxGsdbZqxUVu5Y6dom2qV+Shp0Zl6XwRjbW
+Rtb9zeQ79KFu5LmzS4c9GrOjad2ca0nxv7Z8cKPxd9HtE2iS3dn8WvLBI+/JL/A
liq+E1jhULxXCR4A8bTNj0fpycuN2BzQiFaBFAEFGXb4mOvLDW7Kz54j+J9lkSyF
JmQXlooriE8yx7kPdqsNsgRuNKrvFoRDfm6k/wKzCFiQRFKbcQeBQ1PzNDXTa+cW
JrzbHj5zRC2IFNpBPjLjLZBxy/TcrV6EgByfUV2+TOZavjo0XXZ0MnUOO1Rb1SnR
lK7bYSARKINiUgUAYhQzorEe8cUR/1T/W6Ct0cQiEe8UA5wLLPGdBnbCMGy4qNUt
9WpeT2jC6xi6QOUWDoyt07fLkGhP0sFA32UpeLlghgblZ33N/AR9GojkOcLZVjlr
yk+3BAN9SX1I/wTyjKx1w7f8J1mmSxJtyrixAOWOjK21vORGIa42FtGNKcF+VeAv
clIuSQu/snICb8BHTEiaxyxDMDzvQngt/BdiaIU9/3EZIxZHjN6ZnDruRs1EDKmk
lVRSz6Ay+j0UgvemmTha4yoxrm491pJaKI9ZOJIODPuqpUr3KBT0nXxBv3MchfYq
Zluke29RkaSM0FnZ3fu81LCNIY+CyL5Age/LVyF4vOHgT7cEBCrwvfKsdIX3pcHm
fdFpF2CtugWTQpD4eYHIhMGyxL4rFs84Vvkhdw1gmhSU0zn6B3qyzxVoIMF+7pX5
9McnkBx2HjODy1sGDf5CSs2zNcZcjI5ioFDWTuMigl8JfOVV2wbQeKwuyy/h1eum
93D2MihkULh7C78BcxGZCePrRK47hsmY2rem3auh68R/KHRgOIvq7cCgUQfJfnAN
LzZ3dl96KrUvffzTHh7Oe58LAFFrKXN9QNHCnewVdmxvehj3L1OxPUNc7nXMmh1R
RJ/NnJUWUzKk69rZSQRr6KgM7uVHfllveUFk166fwARjZuyJRedajQDlYqbFaNmp
o+HS4yG0+VyGfz0xapQlohXB7PpjdDCUvTrb51N+FlAZMkT4YPddF/qC8RdJ50Ey
+jeC36kt5y/In0anugRcxc0g/OmOemUSULIBWsV/J7TJmB14kCSN++Ijh0ql4Nqg
bxSykAP0G9tOXJ3SOnDuUsQv/uoPtUa31gTvnk19N/kKsOEDxc4/SLeAucw89CPi
TGY3VDEI0LJCqbDRwnVtcRYFdmez4gl+HW4uef1MGbqVFg1hK5Xkxotc/IhBRVKR
csaHxA7juVGCprd7laULux+WsXn6nBA9h2Zz91UeDGCKlv1dkAkavCECBF0SM+MC
9Y7cQIHoFtlTSyJFn0UqJXwu2+ZQx4WfgcRgalR0FV9auOoQ2t6NOwFbOF1uMoRz
A2m1dxISs128bFPzc+SFrDZo2QWGMiq+Eddsvd9iObGX/Oc3ghj63Benuh/0EJM1
6lvqbsH5wGPz8Y3Jm5GNd1THdvXSxtoHOKFWIrJogxTXQtCdWtmRuvtwATTOT8T/
eJT49NJEgnwpBT2jCJRU4Okv8nrvp86iOJEbKpeaU4In9HmzyY/EIGhSJjzKZtPy
4TljAjSUV7bXEPDtOGRx9PvPxQYS/FqptKS1s3MkmYtS7odI9Vqo6Ix6NB3ivO+5
5oPiZ2bDLkmO+Uv9RtVJ7awaX9cnNUVCwmiQR9qarkb/9x4qLS2Urc2hIdfK3kyk
0eoo4hn2R7FGys6jdzHUcF+RXU7XmULBZ0xjT2T4DpoU9KpWHZ+ANgoKs1AyKLhe
DwtFU7Tq37jyxBmwlifqdnTuUlMLLbD0lgVCRYl4LZJjYwfeDJLm1nDR+3Zbg0vn
9dZ35mmOw4GnNy2S4SiKcLuSYK058LTBIoNRmZKPl+wlPfWws382ElRrqWoZoWIP
NH9q7WVnDV/QeysDOU9N9q4tg3loPt8LotAj9i2D52h0UXqzrkbo7e52cqYO3gOD
iS3p0qfW9uOidqX5480hDQXRKIcjzQf8WwJ3q4R68T0Mb4biqDQ2vSE6HtU9MT1Y
xoQbqwInKN1LZ107jocCbmfh6YqD4n9SXq3At612UiB59PzL4YoKFiLt/BYro927
IODT7pU3W/WdcDS9PztcKcU5qtgwZKRqLZTTptp8JgOCg9ox4iMXJ6YMILeT/Nau
g8OajTi1XtTqZficP8oxqy9HW6bReA7Ct6uD+HsPTFgC382crIHWNPoggNKpKnFW
dYU9nr8ieSSDvgybSEt/LFVZ5dO63ij+lcmoQkNWAxrwxgDxGOvA6KSapMXCu8mL
WQ83ZgkS3+nppvh/e3wHRnpfH5WLIErHxXlTwHHYRgxpjmAErLwymGPufJMzKIow
b/l+rX+7sxyf/faNKw48y58tmkeFuVhx6ll57cWcZp7WY9y97qhMAnXd5mpSzNyc
V4dt7VTN0h0TgpgEutfCTAr1OKknW1B2b3fUnBXNHptTiFilSLGBvewoSsuPJNf9
ZZ6Er8+rqx+P2uE2uEI1mbFKzyJ9g0ohBf6rW/Mc82d9T3gHJDD12c4N+eCf14x6
HpEhT4H9Tszmm55UHqkT3y3RTS3JLflCb4H6CxbpteYuG6T5IklSBsVvjqwB6pi7
wkGbci81nKsVk8RkCeF9gDFUD93Cmui1I6LHlr06IPfA8Sw7zE1EtBRrzlqn35pm
UEaLPGb+bDWoysFWa3RiyLP+lFQ4ZYN63cy9iUC0SnUgZ3BN/hz5g8Da6kHDvwqC
35o8VYTYKeBHAbZi/TiVb756imainrmayyTMuByenJXPw0LuNfaOx3HEwwENfd3B
140w6hmwGu+NIgaddKoPbPAbPn2q4A3KoCFtWNcA0Hd1NtJr1W36h9GEoPN6QGzY
uXeItoSMutWk5mcKC5fpxw6c+1x2vYZAu1BHLsFbc80H7k5n8tqYS6+MCYwfX/0S
aoy958EUzF/klxPpXtak2hTmm4JHe4yeOXSa0gLYKHzMLbfoTWaUsQLlikixf8Rb
2LMN7p5bYTR+ap8NamQuDIdpEXp8TV/1i8x6oUntH+UH8F3C4K+L6uVlcqykgFMu
IlrxHgBliZi3pqGBTMK4eBa4WJ7LiC1cO50yckxiiWkuCJTO7GtPzFBWD7jTZfBu
0dI2RCYgGk1R7L154vmbiG+GoL/IdzsErEENdX5ic/e2TnGk30DAJ/A+LtmlqCj4
tsrH4yKlhd8t4FGTwWr9bj+wZXhuVeP3MWcJbrEoit8Uf8cYsGi6lXyxqzc+zNEU
dlnOqObVhBwNl0kIC69Y91XqaBL0TqrUbJ3lWbvm1nbxQLqEbO3i6oCPCF5fY9je
W4MQ4PozSupDpFiUZSdC7B1Zqg5X6sHeLMQoVjY8Iw2gtO3C7qiH5Ip2n2AGT7ga
8Cqj5qxBD9OkBqCH4D4NHSyjVqqsLRWdHgDIlTJKGcmERNOOO6C+gdOZVcvMULLs
mpKgahArLWaRwmdKZVHkyDkkcaMLwWcihcIuTBWQoFYwwncC6T+pyOk+HURlx2nU
Mia04FRO8iK685IpGrg3qcyKej1ENvpDJDkori4gnkErnXXRuu8oPZhj6nWKS1AK
uhT6626HTkum0L9/zuL21flnsyqz9gPEdLXIE4e1WLNMf47b+XvpaOkG1uv6F2C6
m0QwTu03/RS+EvVkQMjhaF9WoTMxOcB7u/GQyINlMdc0Sig3k4WYD/fajzuJsaZd
pg83J0MC7qYbV9rqtPxIwB/yoDKjwmJqsaC9E/s1yrrfBDKLZKCiPU4aTeb6ZxZL
hHyMBPWOpFyOIo0mtuSYpXUkHmAqBtvaagCU3tUJQa6VTmkb7CrikEbEhsicVxzD
HVkkmEOgkia7hQciSLpnM+9OUe4Dpqkfy7V+EWrm4WHbQPwPNqjW/a/EuoYudCcx
OQX/ZF2YVVC61G9bHYJ8b/L3zEWT1oBiTiLf/XdpRV9dG734YOcYYZyKZleO26lJ
j+311XtfWkf9F+Y+yYFbYk/Exj2Uti7Z+pQUtHdv/GBPz3dhBgBCWngwLybQP3Us
TkuI4nZjJgZDhSD88TWc9Bx3JK3gRVkADci1iXr2rdPu/jmkpPDaBaemLCkH3Yym
/FPtZTk9N66777Wi2lvr6kgg0rwf+JHe+zptYC6WskJ8fGN2mB5jsTfuybvE3TSp
o6IOeN/osqxtGox84/QmLyAMtabA6XEfJVVoMJunvjuv/uTnH76+T23F3mONu1Wx
ty2brUiRAVQrjDrqQdtitddZsJIIfRg7BSZ7STrFB3mUOiiteO1y+UmqgHoZYnm+
qS9jgHVeX7+lOVlfa5ONhSXMxTI7fDNQm32eqTnUlaygfttW7rixQZYSEhc53x7K
aAAWj50ffviF+CuW4jj9X6TCN8hUHZdpY4NFYhVUBAWUwp/ZqKhV/i1NXSxh5WAC
2iQ1OTkgVmbSqrJVSHgmA+mJyMU+PSg7V5b61NTwvtNTHXpMuUwCLN4gOXRMz0mG
7YxhAPuVFdIqBFKbus5dOKIk3sOnh8QkINNn4O4DRwoxTA1DVIywmYpRZYO2iTu3
ueDTZzmJ1wwQE9qsAm6fRN3icBbETvbsc6QnQwNFrSiJBEPZOyBsy6OPjs200Eqt
L/d9qQeNwoqdYCEWZ4SGFUUQCqs2/WpptrCWtU5bMvBxZCH/pQ40HedjbIftlH6z
y5NvmBqEcmucLmlDCScjnSSg9vWc4XUIwcz9perpwzxccN4SRuA/fa45yiSbPil/
1VAq7VTqIJZ5HqpXfzluUG6VB9XswH6OOetJuZIt4TR5YqM8CLlaZi7+kQqicrA0
Vg2jZ+now6ZmMpUKMOGBuSsLhjTOKCAaiORmvA5mJOnRJ1SEL/MeHCbFTuTwXTx6
rgTmyC3b6POCuYTbeVsrMqDrxwkWsuMESSfPByNHFWsRVlhu1R+Sa1FUPT5VzEJT
RE1/EPa5UgZltDlfHnftskCeGpufkPnQM/TrklcgwYZ7Pe5gVFh1qBnvXyAzjydq
LQzGAx4mcV+x+gFyat4C9OaWaXcD5oBJGBk3z5J2htDX5wkI6hEc8GEmrK1mjXyq
gV62FkFSad19CEIUwgPB1QA5sKNyEBPxcJuHg6zS1L/QrFjcj++6TVfT1WQlcwRm
DdPBDwTLWNDCxcWPMkTC77NPqGoIddA1JX0nkPODB6NPO8s4LkQRRBNQj61/qRLv
bLXCWfUfqDApvoDyT3cXNtmpOuXHwSbIxUQLN2PFS7MRg3eEipzyYrNakW+jSOub
nK/XnC/BsMSpmdVfDxRrBL90Y3Z3YUSAFzQbvqIL69KsFwhTpCYUpcvnNf4Q8mQI
cONFZO/x3PS1R1B0Zu+9wl7ibkDT4YTxxgMh4qvrJaCN0OcDeqJX17Cbp1M+GQw/
hyichV+x141CC9DLq04j4Ca7yYJy6/18C660+vZeohgSzcxI0dg9+23EDIHilo3/
8wj4y+tIyVN353HcycUAbVyYz1nA4XfV7GuauQzfsLzmYwq7f2Xfdhep8xgxte9w
9BXwhKUVvXoOBm4RLuM+naVaThcNF6wn7Nt4t9qS3Gvt+s3pyneTC6e4zfUO+2Jk
rRBLADksTH6McM94M7Yx4o4G02oQ7asQMLb/l1/JjK0YZTClOQLj480dhLkUvzok
1/NxLpTmlmedMmx8jl6LqKOhnRalnEdlHcv/SAhDTkk=
`pragma protect end_protected
