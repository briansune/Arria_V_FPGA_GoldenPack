// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cpc9VOPEMMBofPYAx4PKMB/otNgWdF99P0IVGW5xYONbuqhD6uYC9VgC7TVDZNY18acrcmWecBIi
VTAxwdzwGPoKwC8080sEyJiXUGXjnh/8KU9sXa6goKigP5J4JBB3tpXDjt3XA9+hfMBzqkv01UVJ
34WYdboEFdqQUStq0BURSNfA9TbttpzwHn2Z1NtZ4ZEc847KimuXv7nyooDfpqODP4BkJK2AA/xG
8vZzGZAIbf5CwA9M6I8rTr77G4q4tLNQrRhr8uGtesi69QGhHvK90Hb0pp1u/gK+8buO5Clwd5rI
/zP27repAAKh4f44hucmHQLtzgJUwlYH4FYgFw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9056)
YtYUYqt+52S29oQ6KeT0LwKU9jI/h+80TY/Nvji0TLA4rns3i45AFoVAtDX7V7jXndSws99q5W14
4b/uzxtez9txT12eRLPh9Pu9Bq/yBIUy+RSqsdBxE0zGF+hda4yr7uByCcltwxq2enfnsT35NkA7
Bw6Dqs84NIn9J5/qmdKkZXvJOpCnAe5agSvLqC4rX8jpfJVmN2AndoUovHn8Nl7q+TR4yT8u3Am2
dcj4XvyGNjM5XeQFowNjr35tn8zs0tsg+VowEKkG8qHq1kO3qlpbThcdYP0VeKV8yhMuEzjxyxU5
IQHlJQOBRIHWPQEAzpBWljO+5pstjp1n+GPDNukEN0W1z4ZKTgrXVbww8RTdXGxom/G5FzQLIkrY
psV6H5S/J3wJGhQ0Re0QrjoLto8otsxjalHMp42MXDZvLYh3+bx/yafZZQwKbtIkQZqvZUpvrBYV
ivVMGYceZ/YITtM6Wdd+jAMYAg3D+OLfMYlyQbFhOAHJ4xfOzKkldjLtp9j0oVlxwT8eQ7ngKuvv
k87ASco+AhTtYVCiqcE1mrnuf82qtMuNwHSQfjWXDVvYIdkcHPcSF8JBKktU9Cx2aYAIM/Vm+tVy
MYUwasUxHqwypn7gSFSWdI1TGFAMznlSBgPiz7vhk8VzVTg5KrpC1XL4nTwV8ZBncPezs8RrSSl1
a1Yloz5OlTPD5ZCnQkDUUna/5QSYmpWSwrZ54WUrAMNCSwsBmdquJTdCwD/3NlhPbY5ms8r+krNs
kwE+sZ2cX9oIzwcugp2CkQ7hjAsOh0jbeA3uhMwDBrw82mvAhXF3H/F2THREb+EKfQBU4tPmWi7L
kUrQhvG1dfHuNSknHxn8GMuvymTIgAiOoDvTosXBteZ1jiG1R0VFSuXSP/7T6fMxvO6pjMW7EACk
OPHBqxlRwXrpR9N0MnFUljAxVy3DT+oXW+zQyppGHBJLism9c1fP3sG/8ZOhf9zoW02+t2UNIYk2
//vH2drq8DTkZBVXrsJV0rXjjzMZ//LYxdhQm1l5b+jM0BIiI/UH+d7wyrGCN6jcGLeVLY2r9bCZ
tSDXM2Qi3Ryc6WVS9/5Rxdd/QPLaJ6rDEDOdUi/2XHB3ohYKY+4NXOfur3SiZj2nm7Hixn3D+jFN
c0pJuwZhmN6hxFiLuvxM6azYt6BPYUb0CNzUB6eKNqsFJcm6rLqfsPXiiyuwMB3OD8HCgQWTqQSA
naya+Jti88LPdzKrnhxrxQLCRqiPfCNuQxgUplZ9eTqHml87jY6rYAKgjCa9neVvNbQWX3Eluvb5
QUjNPWEWwVnvgQq3QZ0GtmvnyjS+hrf7C0w1cfeH4RzlRTkmCfg9JFLBuUfo+uTE5URxtKCqh8KC
+cLbmgD1GqjaH6qLAfPGdCxHKxXqsGSdQMRv70pUBsMCLaZZdJ6SRRkeeDLMiHDnffLgFmLPrEop
fm1J/oYRzjCwpxaM1Sduw/YENIKXZEfqIfo4lcnSOLtMb/cVjei7PXpEF4+S84aiTly2oA2QpGHd
xf4rGsOqPNeAAshTpPzNhVltbOkqHZM+T8wtFbwfKR8hY8SekFhZcwfZ8m+e3NSviTJf6cPX36DO
+Llbwrxj0AhVnmVkdUUwlvUaUPkeSlKgXpGZzc2zdQjplqZLu1iIx3zZQSvENTDpranvpdXjzb3A
afOJ4UefSp704XveUGX6ZVtbMIBscSmqKO7Knj795xUjnPinDYrAIPDzjUHhHW/Tl3roXqdm4ygD
CmdWacNnsQpAs0ETl0cHaSmHzXPzDCGrHGLJR3EzjDyNIWcN/mpJOdHFl5/UnqxcN5/sAB2e4euJ
e9auz7j4pPjwl0MZx44FDnN/g9qsYtGMUXFQe0C1MpGrA536LfuTUBHDg/nEirSnHPX0lSN8jxGr
UdhEAr8QXvN7kvqj3TCsA7tHAfhe8aBxohYVHgpQR5VDSQzFtQEQx5wIjgtJcL1hJi0OKY9o0KFQ
PWi5mYMsLrIXQIhK8vu8yks2GAJvWZFSjaIY1/EPGSbCtR2BzbdyMjjNl7boAKmEIDkc3vWr6L36
NLCyf5Ydn5eIyoWa0Q+USSEj+o9xSIw2QwqCsnoJRNeMnLi3mnRPBEcVwbb43cIKieuTviUOQQ8m
6Tvh4Wm2JXNz2qkM6BU1G+qCAgSgf+Pjew/P6BXitcxnW++oTMiBRbQEgK/KFJ8DkqVDmeDPJh0p
3ofHBqfOOy0a+vfkZnKY97X1atpdsUNcBfXnMCMnWHj3kXDle+Pz2JlQuKii/KzOrQuCwtAqC67w
X03D7ETyQI1Mbq3Cfe0e7IeRlZWCYFQ7bymy2o+A8zJx6F31gQ5/x8+/Uij/owYKsYZIfzoe+rSF
aZIM03vYqyqotUSNKnwk1UR+WUkKBnKvDj6mN67lDBIR7PpAj557U0xklZwd0v5xxiLBihaOxlmX
IsZ+XebwLE31VESGptZUOxoxXMPyjR+hRc+VxQzQhfjIfy6sWyMtfMgbspNu7GmIohW0fKNWm3Pn
R4E/B7IENQ5V4ZydURdpBaD8ap/vJ+1/O2f5rnWD99WuaQTOOEDCP2YV4mNt1Yt73Zof+um7KqgZ
tC52/x695wmu/jcXfnlZMzrMXBdOGO0j18zreR4xQXe4eqlPkvDuikrMXQoLV1DZfzGNXNGsMxQg
V6n2qwzHkBPwxhY3tXVdzFiudy+XbMOAmq5L7PRMuvtYkk6lgupQH5QZ2bRcfagLlBCGWpvGsoTN
Cjr7Vtdbkr2y5OCEw1TXKnGIX7lOkhNP7QcNX7wUDICaPC10xQutDlCV9Assr5tlbDiK5N9oI/L7
U0HDNNvghXdrqfGjZLA/watPQI3HJyzzm7exg8J5/AWWEvr00b9GYJ22/BNDeb/IM2jsGrRfE7qE
IyOV3V9gLuBJDgzJiOWUlsSQjoGntcNiHfXxXtYtDKtZxfmA0wLqketagw0FON5uFdWQ+r80v0rf
3RIAhKjAvHUoec638o6e+TSiiz+lY9Rff5tEnzGeMBmCvkGEa0K9R3pqsaakePJDRmYnbkp67ger
Ss6e6VemLZL+E9koXdPs48MfRDz17pFV0I62EX2/jyP1dcQqZMJ2kB3j1v49+Imm6Yy0A1aAbXyK
VHBAVS6d+Zn6qF56E3DZS7THY2v7fwcUrx3EpV7OOiw9SV9y1ElVk/G/ppjww7MZSszrykWwGteb
T+c+heWca66htClfvw322e1KD5zRJYHLuM7TTzpMM4bV6mTNvzIjm4VUcxOGxYGzc0603ZS7qIoF
Kf8zsygH4uNfDIOH8MwjPRchRwMJL5d7335WcYbqVOm6MEi0p6ZnCLyjVeoXiFuIdacimPMvaf2j
fg7VMH0xDO4Q+QVKvmE/i1DTcTLdwUm7aXF0vp9f6ye9tVlBuQO6RyC0XDksATXwaLbXQjlg7dG9
sPe7gMquwVbDoU+48VEHYDBcpheaCaT1/1onx9/NEaQaxa5ZeC+p6cW9aYZ1lZEMifuQb18hj8Nw
TIyWlYDISeh5IUltbzy6hv+7UTzkU6Y0O637Myg6U5DyXjZ3eHX4zxJLnFft+wlvAEM4bj+g3xot
EVSArqWoHGONvWpPP2GzgDva+MiazSBNoYyzbc7h3I9ZRPdmKDE28tm53OkAxhBZi6LEBIWjdFKG
9yKNk76LP+Igr9G46cSMYKbsNXWc11NUMrkoqNaMsmUzEfK2/aixiO6BJd0+/QTceLTl5W5JfTHx
ZIhwDby937bTGXRNSHkhjzgSOLXXmhJeaohACpAWU1rqrCQDewKSA2xQVATQEgfLCogiQ6iBG8Cd
YtBxoSZU2HUdF1rOECvpnI8pldgceSDDD+/C5pPAAFpbgGp7MwXWMDyzwCN97wY++Tj1858H7pFi
XHeDj1ElOLt4SMh3ACWho9ia9f/VRvpmcT+TdbsoXxJiJL9oBxsZmuo4VaTwcYSB0wFNes/zyhTj
B5dSq7sKW/LCX7cMlYRwh7i2zyiEqrDpwl8FeErf3g7/XVnMwGoJJ/0DCq3gVURNeHDDvdzIg43M
hZWcD3CNWUWCv+5VDtTPC6sclk/JWsMGsq/JVEz7nd7hdk8CAYMkWOxO0ScroN+l3Jutv4Ynnjau
pBb8/9Bx3Xbq7TS59V3wcBRVWF6fZ3fpXsMzgF1gMg+bsBlwahMHO5ZKlxh4nP9XLsuY539Kpoj2
ujBBWaC9MWYbOCaCY0dTIdxqFzySpCNbx6fYaB2HnPvT4pZJFqfP2Yboh/hIUomaRtnu61MQzY06
auvdbiSIxraOoGC8BXuqIKImTVzCQ6EqRjNKqtoObt2VTCtV7pTGHady4UMHmNGcJb0TJ15We5tk
uvrZsIZsTrsdwDn16XHTrrVwWp4oenEkud+lIQ6HGR/dg82raDiAhI57othPKPmhVVwH8LUjWVmN
Lceg2YGum0gEaa9oEgWd92LA6HRJoV6+oomjtkn4H6YS5MIrM1zcI1ivA4RC+yZkoBhiVs0i1reR
wSGohlJc2RdUJOeiDOWPikVYm9wfGLFFDwDWyP10nXycxANPAbwc0Pcg/T9YvUKSsRmvAyebnT6j
ETFZsiubFAWxJV5QnGyW/eQYUYNiwIjQmKgJlRT1CHKGS70h3mJy6ZsSmioG36bKlN6kMgDez4Cw
BV+5UCW1E49dWbfHcadtVm2Hj1871H+OPXqM7y/B7knA0/KakvDJdHH6p1MJd/riQ+sChK1ICjf/
QVxNxsbBHzUrdkAmZGVgqi/uR+so2SsCqGeNB7rg2UThdUsa9fG6FtsC0tf6MfE45HF4pJ7XI0+4
efNLOzmxButEUsSolj3mNA+oAxztTHQnma0rWA+reQ+KUJ/BzQJwtQBZJL0/Nwy1Haabgu0bccZi
wvJUDyT89nxixAN4AxBv4qV1hLz/Gzot0KWGWGLFXDQsYeSsNIPKvGshQbOKgtjFpbjB/pR+lKpe
73piH1ZH9W6hB7J08t9H22w8D2DufJW0NqEgEs9n4MJEkcshh2PyPw7PJG0q8aXUFyfihgCh1EfC
zD2ACZHvOd0Cq2yrVx0o8nvOhGzbMsn0BAoDtbg9SpK8fw/pBbIC1W0fvDXM/B0G/ZDjVN94yP04
isSf7lHvCXg3NYJkF/hf3GSpjIMjLkJs95oFW9A0WjgQk5XdOBiU4+P45OHKj6L3Bglbgvpeuo6E
Fu2+xMwZwBQkzSZNNgFPF11MtO3hGuPBQvw19RPqycuARmzRwljMwiGnzye/sOTC5qfFvCwSmJ+/
NF/Lt/nDJTvYAH9D8gwrpy1t4SwxrAdx5Lc+g5TrcTz9foZotKpDjtpFzcovLReeUrEro+m7CXvJ
K9I3D2mg0gORvslzCmIp55ZIkqzh8tDwc1usXzIH79gZjKEY83TET9/YdiyZ1hMvdmIOe/5hq1nC
CBGwG8RJMdpaQ9WCNM4FChWjuA00wEqnvYp7mXJQGvyi0UHYkhSzVgXOVvkThZ4p51b9dAnDk/I0
Rxhum32Ox5uD19Ze38bnYIt5y8pv6grIg21IkGcsNVaIzrn3C8KEqjFGwPQAWM3fNKnX13Uy5HOz
SlQfsKiYWXnWNCgn9M1BHxlzmMJQc/hBJ2txM9gC3J2FR0MG2+WuyrfSRD4Bh9Pk5A47aJ+6o63i
ExY0FuvSbDuRVXYgK7cShLwceENOSmiBZikt5UEeKfWqjCHvSc3vfbxVeGkjDCJnygiCWVbBKAih
pUdC1786pKgSYPlRulcKGIBBuPMV/DKAg7eB4p2zzz/f896HzAFbHBFVRU+50ATDP9yZj1wTMTPU
Gk/k5mlcb0ZrWDkBnNRdH3dY2ofDjrn4by+LE4G+wS5Mw6sHaPiPY3rXUdTZjA+m/gOY5K8MgpgV
aBWp/X1MNVyON4MEgK52DC0A0OuY+/HGOBGM/mRR/DkiFrUA6PpRNdORToE7Dv2r3gLVFTTPXDrF
kN7lUpIrxoGAzBvnrZad1XL3T4/yNI9GDlD7sI8n9FiLARFr1n8bmJP4OC5rEw7FnlZR/nt/20sZ
iuhnMZUcHkUZPcdQY1sTc+X9rxwChi/25pyhQSHGXwVncVw+UB5eWypXU8E8tq8Ut7pl87WKMDlL
lto/IlzOWVWItu3XzwzlQK3JEZr+S3G6QgsIo7UUdp9ypRCVuQ00DQNMSgSK/UU1YnJdCNC/BvYk
rtmo1WQrM37fo3UH+zydrCSkJMAHzbAlRL6WlgJRITWGyif+gAx0+2gNj9jCAudFZfWVfDS5syEH
/MXco1VapeCddIgucZhGKuvsB5ja1rbe7WKMd4+NW+vNnyqzk2Ep6dyhOgjLDQbN8IqaObDJEwCk
SHKRBe7+SlzTuEHQdgCJJHgZh++5EvP7OvfKyePSJLVC0GetEUcKG/ynFWSVXYnXfML3AK0c1g5H
+deQXFZ2DuE4QPM7e9imS+t5OdLmFlfAMufzE3cXrRB8UcvSS6Mh/poFpASe2fzFOiAE+xBj3d2I
KjDRYir31Eis2GXIInoI84nLS2U5EifWbA4mxAghIGPHthCTEzsVzY1N1HwXKBYgJF/6z17VZ7hv
8IiqNFyec8e7UJOhGaOvUl5A1NfdljWdmuDRrsSj/mniyOGZut5NYbVezkL8/r2Kuwn86/zozzHm
SxSGdAwwZASfrPVpHnRcfd2pArUXDu1SaDZE2igtmXdUorjHpF1oLBu1z1Jj+dG3deGrXu0BDz9K
8A9Q9fkQq/7Jjmk/ARbm0P/zViXK2k0w0yIS11ow+wfAaNJzDTvl9GuUFXH1lV+RAdFW+W6aetU8
BGSRT/cE/Z0FdjTF76k2uX9q/pqQrK6RSpJ0GYPx5Qi+kOmJrfCZ1I+uDd0AffGi0IUIICxe26Zt
H6Kz/TV96cAhdFAuMIWdVhdJM/KtRuQyvIj/4ymWEohCsxO8L1FP6pNEl1mBxUXsQwhSRDazLykO
4FWVcOvS20nTyPJufese+7Qt0Kw6lDizSTMOofytFJ+mWc6+BahnTtLCQKOujuIqMB909MAnR6B+
Nq3MVoLwZEdOkolr1QTbINx358Gz8r14+Uh+7qPmAs0TmTwKsxsoV8Zhk8tW9RU7VVnxOaqxlu/C
67EgNBhHxXVnPMyj0w4VjrbNls0r2sntTU8ocVVW97m4r5b3F6Su2n1ngWsVCVV/WSKAqv2y+oZ1
TQ/lX1Tjc5QuS/QjMi8emD/HDlAi1LvQEd60JmeRu7yp91+G+NiRIy1n17bwzE+HLN/V7WcLcoDp
UJG30cv9rURGGOL08mzvl5JGo9BgjmplwOdZGyq+6jN9jW6+lqBJ+jp+bSwNu3VF6vkbdlETL0YS
pXZjcIdYGvyY8htA5EBQ+ALKrM8OqHfBkNFCMFGZXCPQ/sD+R16JvtXj6xCm1/Ruqw1gs6BviyYx
X4xC2BJw2U4ns7TtsPaQqKq5/H8pdx4oqHwPFPutdJm18H9/cBX3V7VTpEm0W6nUlJ1r+83OEqUZ
7pdrvRFtp5Rp5vp2OCX0w8Ywk/f+mdEVSDcFbj9vjdlZql45H/vRVIEsBvBcszIAcYuEVJVEarJA
y5rGUkPIwNkV936PfhqTkeFX4vcWmV53z4JotvDpUqmDlP9++9lh8sWTik+USeAODXxBwve+p+G4
osTFPViouz33Mea49TweMR6TP/ozVwK+owJul0d2mYOSF6y8U8jiq8rTcIe4tdzz128TpwfFzxVD
ZcNWceff57uduDqa7HsJlEZ0iijJDTUynBJnpwt5PH0Tuy8MlFn+yoZ3aCfOSZBFgJlYbi1Mv0UJ
vlmdav5X8mqMDNACqda0+iIlL7c6apvhAPOs8Fr/YbjuuLvjW6Fswy6yHiKm+hPJftvsBdXibKLn
swgrEX0tRItDrOQs3Inlv+rI7zbk01xi53Wmx5f3DFzQ14AbFPSfin6l5vcOhIL2e4SvGFDwPOlY
Mk71XQYnoFh5awRb4pI6tfKfSROntRwn5E3Z32/nFfoFDTkaKxSxlOaU80tVsuXREXqvsX2RDzKU
y8guP+aAXqmddEcBvEk5ESjhfpufbHHJ9xn9VgA5fSNS/HwfROWn0TCtfSDKLNoCxJlCTPFs1zut
HKCwNy/oqhXEJTC06obVfFEo/tk7H4TlayG4uYMuxTnlnD6ZhT1jqKGn+gP2KeXMbThvOy3iHMtH
g0whAijysQtZa7lRgPSow6jkOAzImlwOh8MEMxJZl9FEKvRKjL6xj+wYSlrpkLUFFv8vXtzZheee
2tfLEyOKT/G7gU1fP9hNWLs/MxOWuF4WpX9pvrdFT75IJfFOL1Hd3lMYbgs4Tl9ULnRejp4D9iJH
tHGrexH6DHI6h3DdKHwCdGJgrmzerMWuZ3owSiOCq0aN4lRrMYLRAYyAkX7xxgCdasWGyfawWxtp
xqLn4ypK4DhAHVGTYc+6UGIvp0j7gUWr9/c+OjVqGoX9WMgV4J3jYmIdVPI4RPdjJTqCkkO1yJ5h
KgFp24P2li7XFTUZ6BHUq70ekKLXIpwVvsYPS+JcqfhUx3D0tuku+V0Mxs93bxHkW2+utQ4AOFVa
AtQF/E2+cxfr+ZOjop5I5tTi40UDNu7kjurA2Tm3xgvjDft+pkCrWiCnYGQO2iArIMk4DKkJIRYD
fq3QG3f/zBPzB7dfjDiU9ZEv9cCQFYUyFmSp3si7mBDCuU4lOa9adOXcupdzCe4rB1HZOHDZsraU
Mj75gBbQWfSesK3uSCiPwa/2WZ5RymWSbRu3ntptjZtj2o4Un/TK4ir6IwzHfXtFM7AaVMqF9qwg
trAyEWlI+SMt0b21wSR/J7/rRmrIQb2Iwykmt6JS9Utt8ZH9z5s/VGY1/2Zy+B7/VScosUze4ciO
8mv/I+QVSXdVFouKuqsREByG2my/2ev/kAdXs6ZP5dts1qVf3VkZjo2B7CNOcANxV1IkvaBGwMp9
lyCP4qzcD1V4hRhuzhklKv3ZVKafr/vifNk05KMm4unZKW0PNag25XyrE26EzQEYdHSUyHnoN9OM
qyx0xOpfydM/eYQ5PxDpNKFPWi+VndI9Fe0U6UN9otZtO0X4bFH1xo94uTCMHwYEqD2BCR3/9vB6
Kuz1p+xTynkDwMcinKt8baWY9CQtPev++h3/O4oa67COCnhFxzNCKD2fNWRIurITkVxbqMEZZo6d
81Ob8oVpnMnGevjz6pkQTv0OsxiURQewZxy4hURkbcxX6ZC8nscy3TFx9+oJ/AseGtZbbJNzty1y
KYwr5hThLusQwgqONBBaiVh1wbdqnvqgjI0KFqMYCXK023vGe6umdas27IMeh27hFIoGNQ1/yXmO
U3C/yi1i/06XXjYjZ8fGB96PDx1GkxzFJBcTcaD+IS4+QNXbs8XPL55TULg9Qa1fo4IKN+cRlXfV
fP0KocF6OU/d3ywYFwSUtc7E1laT0HNTDaPJ+JVN3TXfEExnPcg/i3xj9xmsRoxRx2OkUKfyCcqw
WJEGkTPJDL+wowwNioxlXZa9gxIFaRkzNTKdjzZMYgC82dyz82NIk0dKaxZfbGd2G1f+fz0yJWS+
OPjUbe9OHZtvRO3GfFQ62IRuFtNDS6w5byfHnq7y4i4tyBoSKQSEiI7Nz5QHRVQhUSuN3IoRwXqW
Hd8HtM/2/fAz9zLnxWUkh1xCidRdRhP1UEEoDv8eBLvrhUOPInLTUaMlBg1W98/Mb/f5vOQ9iF5R
qXIqeuzZME97EXDWOKDPf4JGvA5FTeeGWv/mFF4tHObHn7+Ha0A4UB1elaAz108Oqe0d6Kr6pjJX
AHx0dpLFLNuzDD8mDnUhURqsrHxP4ag2oKBi2T3a+D0CWSp51uV/MMd6xhRS0jzNEPPskpFSj5Wd
pCa6iuPmdUaSRKhkoXijuAtkVP8AVQRaXYSnGzXFdC/NqovbrDbUFiBGa4bjQxtgx6Qtbqy+L79e
yooOqPVjp7beTjlFTjDchVX9i/3hz8mDOsjLYIZKnXn5FM0KReS2z0mw9e/5PiBhSRS4kAmVvYD7
WZX00s0UiDNpZBUj3yXAd6ah6ION+IYN0nd9cB4Cxx1BfuAGiPiWW3ISMHaPrdsVvagDv337voLo
BNxUfhycUo3YI5xvEp5uhIMxSwDITX66p0j+McXU7sk80PUBzKcZyXS573l0+fwLuawH5tWPTBIH
ofBXMvUrvQZsoFg76B2TzteShtku8tHqVt4Mp+3pO5T6Mc30C7HXBq6SJSlmTrdTtCw+2EK6sNvO
EvvESAzy+kw0Y+5CRjbcAV6WKBXg9r4h06ZIkvgrDWeEYVdzi9fCOngn4TXW27VDyPtcuelPJ5Xu
JobKXX0AAqSUUb9rCJsLT4VcyxEbXwfWPEwGPDeak+bmDFnOLcxhZTSvk9MAix/ky2ez08Ril85k
G0AcjYJz+Hi+2vi/2twcWnKWHZWEU7FTI5CQ1SHGPGSn0ct5/96e4RyHbhIwUKgqSdCCvxe5F3bd
lynQe+H/rGJCJRkCbNdoexulcoBSEOdF73qvZqekVlYKdgy1ay82DFXHcmQCrpQTKLoRodbzEG36
ujSPYnTpj6Ol/OZqxzukHKUfzUuwTE3OlAFRjtN1gWmbejs7w2Q6HaH0vEJCsrGrAdSh75ELLJoQ
GhChEp0Vot4XPZvwk0r3o8T6C8G4s82lkCO7lQtQc+3vsjwCJn8zl8marZgGgq3gOcJSTzBpxQpe
hzSvoEujVBhzZAQXgpogd3qmlo9Vmuzg9Ns0jIE7q4gEQEwBUpT5pttKCty8Uy8S169OQ5Y4BRzd
s6ROaeLA95Vvy6GsMcgr3oNL8PcQ/2fAV6RGBVS+DEzWLnVmMaWUmS44O9y/M3D0itg/YfMQrxkl
FKdimj4NupuduYePHpzsgyKxqwn6O5WO1UTR6piYwwjnWgEcJgxN3ESFtLiET9+j0BWDhm5rZcP/
VUL6k6pZXPGGiPSHcmW9e15uJ68MEU3HocuGF410DlWljmiIaDwiXiifSownooFKw1OMgnThFw2J
cLNwTZAEWdgWHzmnM11Pab0HGNh90sMdYkXhYsCLyT3vRk0K2bMbI/jPTNKEEGkkPMU61d/ipA/C
O5XIV3wOvh/RrKtp5nFPW75QxMbMY/NYIu1hT4rKdFTuUrlNcTwUEXMW4Wqba1C21BLmMLjUIUnv
yt/eHFXOEQ71agn8qvu57uRZoVG2D62YuWgVyxz8B/oHxymIKv+D0u51pWktCTylI5A6YesHWLdm
v74GwMt0tDWv78fLY2ZMyj2tsm+egXfC39S6T/m3aPfxu8UKM0uTLKdRZecbO4+pk8HuhPgsEovt
2JZJIsHhPVdjomKCnD8qWcJIZyqnP3nLgJu1F8GnsUgeh65QNJP67muNBRfzWKyA7IsdZ4tRLFvg
ChtHztIkQauoJz3pPpQWIIAsrNY5qhEb+2Nc2TCz/YvoHJ1rNN7P73rhxgaT6Mkq6x1my4JsUvyf
A+jmT03bOzsO9ClShH5xyPdxZA+vj/1EAvHFiWaoOpd8BWz1ZyXdrxRt/KGLGRgPEjCHaRaTZ65o
KzwWDr8prQVIQaUTJIaj9lSYM05/F0T2VQFMVfxuZv8OPZXSMunoGeHp15+fmX4tsChhsaVdNogK
xKOOIz9hPZmlaiQ2YgQmXbbDHXLgLknFPSk4hsuhW072EjHtqo31RMKpAtTwujtIworAGJ7nkJC8
EXoeKa6b7BSxnyTEfMtMzlgCHneD8wjdudDnXIYhgrPaSILidxLre+vOSrKv217YcvKxdAeRDMPR
zlJGq0PkPWcblWgF4MDMfC4F6zjdPW/jAqefTTSxlGQsHbqil2VnNhS9JHLVDjZqLVWH8VKlRy/a
sVnh24z+zZU6sdzWe/wtKA3NFXXBPJNhrsjjRRgSlBawra5fEhvytGBfBcxK0s8unZ+6KJgMufXK
akDAAEFxYCbaMKdiD28aXQFdG7LMDynNsiqBDRaichimLfHEdhA05aqsaTS8eg7a9fVdNzyco+gE
3TYJoRfClhA8K7PEgtdg/hQs4iR+LUg5Srz5lGWLckWmlRVpj4bxqwY/LAkuri90UH5jtzDwozql
t4dVub/Ho/0DAKTo8bO3YnppHJ8KUX+qTdo9DAn4KvmHZGuKdm1qHaxL7ARCtS5e+cg=
`pragma protect end_protected
