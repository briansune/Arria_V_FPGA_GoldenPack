// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:20 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V6XDn05atQ/gMqZJ5Gccn2NE6UeVkqRS/QswTkGKoLUrlrltkuM13gCOWGdeVqvp
1xRgEvcdYJjFUBfvPqbsmjrnki8tNAnsM890EO29m1Y0mHzPEInaHHVrZN9bGn2o
QIsOomn24bNRtRSYRj4fxMrt4Gyf+7M1X+0ynN5V66E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5648)
sDzfEOvvFKHihE6Rl5I10Dy3GHGS9bKIy79e4dcGQ5AZIbJsifvmcrViakmb8A3T
QR0ge9e7TgDURaH8IMUeyDiRpfbz0DHqFsMbxI70rlTjjeaIPu4ewYUEwDbs5pxk
dN71MN3L3DgeXILdKq38FJflmrb9n3TcPWTDho+8FZEoHtQaw6E8ACGjnOBSOAiA
PK+jhPh948VrRpdn/b66376qrXmvuQi9I59WbGYMe7VpeedY0Xq5CR6ZFRKuSNrr
zMP57p5Ztiiw/BSdDLNmuPDrzzpHr/fInvvhiehcaUMF54R2FoSW6A04mUtGGZ8o
37WjPxj33cMa/SruUnBXUf+U/GhsPyaT1B1AZX4FQaBtMHcu3W9dcEsX3t5Ckr16
s1/xzcTzLcwurXWacIQ21IBhezZkrtlnx5Bt8JTQW5YfPwueNYSgpRuYg7sohKkW
cVKt5CFzHL9M4xBgrC5gTipfHrdNUCvGL2qRQAfxCSI6Wk5STPY5kFk4Oq2posjg
Pw2ScsSxIxcPc/yVB+QuZgKPTUjKv9jXotyLV4G2SRTuZvUvYO5riX4KKN2A4ndw
IJ9zE2BUsYrKHz3fmkO1kDuGiTStUdiRLmQg/86VfL4v1u3X1O+KNlsgRb3pvyDP
yL4ZbYOWgsX1TjsjuRI1cPo306ye9czG0kcjv9o25oK2BjZmATiD9E15fC2HKaWW
IicqAV8f2dMWNaNTap//XkgYq1wqvfA89bEMepFv5uOQOuDgCQP0nRg0zf6JJfeQ
3HAvklnggU+fjcMvcOBN/hGxug+/Efm55SrxTOVe4ro+fkE5E9LGEt+cA6aAR2QC
DE4raGMtVzYcXgiGVw9ftRHaTmDzI/OP6ciEBhoEE+lvTnB5D2bjAfZEwskmOw4l
Jtkx4awQHGf67DFn1XOqL/4pN0EXCc6lgRdseytXviM4whjQIllBCiGI7i+Grav4
Ly6zd1mxFQkqLNxDJHMpYJeWCA7WYgxfb17saHG9P7MGiH6uX2zBWle8eDAfKt4F
+NbGWpRG/Ww8XwSpp6Uf9fxWXI35Nx3u4BtlSdHhLmwLE0ZrWtH5yLYLa2d9YEWu
aCm8WLP1xwCL8UP3yEIz6p//s9CfFJo8ld0qmyUM9437LsPf4I7oMSN+k5UUJdHU
ZUyRDEEWG1rBWqhuBkNxubrEcy4GlD2fmrjrcnm3y1/V5IbPsFKSyRUpQBgAny88
8LqBBYw6qwx1/1lTj3RfTv0aEnME7B7MhLYU15HgXrZz4FMT//9QXnWVpvAl+jBY
KNmNmhhaAb9W+RyTjrkFqZ6+XLwp46lY0DNmE5LFkAtxkg/2YZzOyS+bTW4N45lc
DhbapRzTNDRIvSns6t8CqQYu2NvIDh/yXXIGrBxEwuiAiMKZ44FhsIPfD1hrPzNc
Pp7VsjMX7EAHX62KOoPYLGXEes/m7snxX6UJPiM0ZsIHidGx1CvE/shgL2e/yDg1
5nOGfHBrMSjezH+4TsPthUuQR6v0v2IUDqR5DpJTP11Qjwv/kvFsWualcr2kBq48
Ix4/nGONEeHXvcAiLlQLL9r0v2y8RSHfvx9PJVlorRU4qikW++ANf3lGJQkS8/kz
tWiXuOEEOjpYtQuQSPDZgHPltSaCLPHhhO9nXKwKLfpmDiqz0zgvU4shQz4xet4n
OWfLXof4VhXLM3cS+jHgPZlyo3+mH2Gb4iN0RDGJVCoLCijXacZhklXSU0K072LI
gqpj94rfDzeki3QRIg4ZPksqfdc1vwemMn6Lh9dDd8OJQxb2+EzZ2YZGkw4tbBsW
5tPgYOg6RXzePGfxIuB/wmj2qs0yiWEaXbLG/BHWiGauYYFdkJTFiFWM+kaChgBz
WuaqNfyV8S6XFgx2BoLQ3X+KXmI2GzuKbBEUKww/rLb53d6JHYxyfK8tM1yIPCFP
J1iXK7L3hDev0sVqxOr8KtfzQ5GSBwehMo5EQ8aBhS8f2HHUmBARY4WYV3Ro7VmJ
CABl72qDvhafaf13lp+l2gRgvD38PRWEivCEbiZCqucYqE6gnaPepeiNCpeqaXqf
DqmyUtjm8o7Um9OyWR8h2gV9qrY3eXiRJFJTWQVivpuIxBE2L18OvtVZzrTvxOtt
0wiIu3kfYNAGAepb40Emfsa9UizpJ5lC6bqouAgHx1nSIBLzUfP6//B7PbEx209a
0wlIKJijDOw1u5Kc8HBFkrI0gpMfO6JZytnDZtApmdHErb1ukc4c2gFFEXZEPNhH
KwelA5bu0xkn9l6WazylQt2SYETNLH96xCL+C3FAWiIEWCi+q8UbTscd4FGhU2l5
WDvrM6L1dYi9YTMHlE2VuIUHGoQJe2cYq7hd81e9L9/oirGzIQInOzVe0MV/ZDkt
vqec6MneLquDLT9jRqKoPP81D+y3VhqSLrTqXX/B5NyOrOqV69le2wrUNE9fipOd
RDw140w3m2ALAsAjRgQ/mHVoy/gywbU2v120/CBMW2iz/4t5qy7yM67x1cKILOtw
xmMFLcWqIF421n4nHPskraiq6tS04hioV8iCCVTE7679yRyTLdTOP12rKzwlx47B
XAPzuLcqJUnfrFF8dhEVAZAHy4Nf8jcyCexGfRTu/CQGx9GECOrMgpZsgOTPq56Z
p0JgM7vfJZkzdRMve+lD4TXexKeJCFMnlHMqIEstyBYX7HvQuuUME79yEVk2WG6r
l6s359EPc+cRGDu9R8uymfdQKbSVbO0ScGQgrhsrJienP4V8+5DFt5hU+8xkvJQ8
H2DGAon0qQnGHwqim7dNjdN6TNmDnV3wPTOMGDl4TIpzl696zsBsdar72JiQU3tz
uE+4GoMoneY7w4uGTboziCy9kZRErQwhgVOa6dSUawW29pdOpNVoS2scPPqs/KTI
039UR9+FbQen7E87Gj8AxNMJn5oD3TSXl472+9etkm/wQH8DAjtfFdP8mHcia5a3
dis3YlP+Z0fkmdomxc2kIU0gpo0a9GMFgHmWckmypgL9Z0Afay8VlT6sJKddEdmR
qokDtrUEj1wZxF0lt7Sg6Sg+5vrSU62pRjhhQjyynpIAN2IflmDSNC4cSG7AfDl1
T6jWjrmFfYCCDmPYzwqdKwiZg0bnJST+ZuJORGBVSeCv9i3hpYCcTAjnI7IrG9iY
cqXV1fIV6X7Vab/850EAg2s9LErUIzKenFHzB+7hrC3F+PbxiHQdyxd0INmekh6N
SoEBnIXxWhbWd/p0HrbIVrkls5+PJbbmDJWMSW5f0Hfgt75JpSPRHaPtCTZumOJQ
numrCsS/HyY6/DDR1fgYcVhy2ADnKb+44lR250SpstmdAIXvH9SOHBEpWjrWziej
fKHtyxHz21LElyyf8uyWupiGCkgHsRYR488LYDvo1+R1QmIHdRepL/hqmzxUyHxp
oTlK9pkIYcqDPB/Mj3ha21gBMhCo5oWBxKYiqX680YAmAyH0KqTMubLvrK1U0wOS
GlEDeBzBUM7htf8P6zRENAUlFLSgY2zvQeQlnV5TMgc/F6Yf3tNHI/OxtPmwIDca
yjjLCgl7Xyolu6MinruerWHYF63Y/GwWMaMN420N33YL994PhEV7KPHNfHRLNjhn
HPkmo4WmIz8c2Nd6Myp53weT2VQVvTaLjQV6C5U0c1wvR2+wErxerFbiH76agZVu
6HL30J/BvM4Qy+4hTTtr1noOSYheIHD08ZPKz+NVKJ2wXxyk0e4C+LdV4RtfnSfs
3W2geK94+IVMgaewW4pL0oaPZ+3d4PFPikDKJBiiEJ4i8B1grA2z8ZFLPfXn+tAc
jg5hH9rD5hxwCEcHFbVNFcZgGru4+LdI+z4oYqkOOvwXlNqVhswgcWm8uMOUPyy/
VUuCogbyNeLUJ11dYc9Wy0NwLTg+qNKu47XdRrt2tuw+jbrxDH8vXUvvre0Ua3Dh
RSQoVSWXPT2BnnkDGt/KGXrSXyPKFT8pvYMw8qd6CLD/DK2n9H1VjXfywUWMj6At
chy2Ep4pwAIZN8IRuycbYAfslv5Utqy3EPTDqW2hWO9OTYoz4ukNLPka5KZzb8Jy
kh8QfnTSPEWTwyzylbExLlGYlfqmzBFPvm8MDKFDw3exiXtFLHAXT9QKOWNb6+S3
4jpu5cJ2C9XGd2U5CPbHG4M9bKrukZRx5//efShDxuvtYhnK9yoTfNv/njzn2CuI
GfDku7PrNVfLz4+CEJgp5nJ5zxOyQUfuBHzzMWt5jyg5le4kCtMVbGxRQ+sHorA6
Z3ND+rfllxOm/nrRrab55RZVVrPSkCHKs+PFDVFYjEuDcG/huIp6vOoGladd7Z0k
8nvhm0nImmnFkEAshY3fPOLYXbQkU1GfBxSlZtPNKofHKRFLAIYPd/5D61g8ij4e
LjZgauf8NWty0OVVVQrqV38uQR3uykVdMY/ZL2fv2CaaS1UFdhDAp6gkrBSlekFW
BMYJQrHXZwRxXnT/gZk6Ea4MCOzl4S1nl2Gh8DBha+hmU2TL/qg/9Z4pnWaDrpTn
Qmn2IreiC126WyUJcgMIq4Rv5UD3EANpKUp31lrpMlEvgtHG3jb7WMeT37FhZj5h
an9umJyQnA4jYvxmCfJMbOuKmMNBQVqU468lc0g4tmfP4XeSlZ5hgTRChZshQNr6
2NVBTfnbGd3ofsG+P7aoRKVG9NOmWLk41y7erbx+A0JFDNLNdCDw4ZQ98fyGc6Ls
kZ/bfMqQ+v1vpC2P/7qEioQxZvIW2e2RNq6EjEW0Oa35BhEEQvS0awWU5NrKLofi
Rr2j8I/RRAjdqObS3n8lEj3wVektl9KqIEfaMk1wnwNSKHDEr+qE1bsF7C7a2pVp
KOdgrviz1l2GBq43D5/gEJ5ePQvIf8ekIBvQJ/Nco4ZIX8M+93oEODwUekNVJsgD
7tqwqqoFDsuzdTP1P9LIQ7PfTyBLQyoAW46WHZj/fH5nGqhbYDpb2aMisI4qcQZf
QK07zCZwzTrLMZlP02IcNC//yBZA6V44vE8dA3TzoBuEItOACIMfywESsuqfb8gg
nMwsC2nZKHmXmgJNnzvvFEEvPp8cuqAHtbZ3YU9N8U3uLVYpShjzeaSCCE2nZgM9
2xLN0B2Du45OKgHmbSZFbinBQGpN+hkXBZRJYN8OL6ZUoaTsV2F0NPPuNTMMtLmX
5o8J3r3PrQ4tmQdbN1DQJziUyRp2R6xiVTAJhqb8we1KMrCtPjm9b7xwq9H69u/1
dQ74sQoehzQxkYdHOAZGIGlcRLGk+IsvUURyb8kCxVbNA5m2OTHo2PglShRCDuQg
NGtBOEGiUh7LVeCRlrGDHNzA+6zNx70Be4Wf4mb0VAKn7G0UXfRUjJqZF/mBpsb0
16DKjuEUKnX0OuoUpf6cN8td9Xw/2GQmf6EyPPwVRYeRWpxE1XZH3tPLxaFuUx0h
GwqAc0j44fJT7LagyslNQqMapXD0m+N5vIHmK5sg87Qjf16MTF1opuR9KCdccwsJ
3BrqJuesZHuKPFDx84kg71s9d3gruIKj46jTtA0h2Tk+FmbB/996gUOklduyyF1u
CjFPTi/iGyPL34aS81dbGI5OE/xNJq90c32O6hevu2vtj8XICV3da3iDK8mEAzlF
RTAFbBU+LJ/Bx79tFRG/18mublsaWGuHW2gRQ/2iZEiReILxocdeKZ0VudFn8xvF
WNppnb6aEsxyxUFoiDvobm8lMp9VaOosAo43EtOCZ9/+opqpSkUNJTI3rCDgG0wc
vmnaHCz3n+VmclGrtNdn5mnWOBJL0iawT8QrP6p89Ptz0DJJOiR5mMPzJ0pEaOWE
jBIJfjMJkCRmcORFGAyQIOXtGwEa3fYcRwqFAijBPAP4k4ENtbXCRpYAa67u+s3J
yC1++e2VZ5aTG12yQzjyKoq21USaf8kR+yauX7WNU1Rfc8BvAME4Um3QFe9YsWOL
RsdHjdYlTuf6rMm1AOkYC5w4g1DsrzSCJWksVSsF9GYIpmK6pSUyamwvaMmvoIxH
W/6wIY4r9CBIpDvU422XlaPOZZlLtFbQwFVH4ClC5DWHCnOBV5LE4cxOhSGqoXjM
8m3py00xMvo6R+bM1NRmD+kRNBEpaph1qw0yH9IUkEk8CxXH0rdUHXV9vjnKUDxt
Uv+70LSuud7XKX237ytEe4lBawoEjeHIpQ0OOknfgPZIYxrsolLpSEisfmZosQIu
iBrqVVUPJV5wcYztaW/+mphL8oHHILR82MOITWMVi/FfTAsFxlVU8mA6cj8+OcY+
0Sx0gVHcw10ps8CWloYrEb7tMTGLfCAsBBFg85mlzMgSX5dtoEu0tO28AEvWyaYE
yJA6vZbK3sDhjFVaXDW3ESqGlQMRdCPRmvP4pE8K9/lu4THU8RosUCFXfYKRK4M5
ZHDT/MDus8m+yJVx7aYTjBiRbRMliFXYYFVQchmLlMDSiTwhbkxK9SLfn0FZ+u3C
CXFBlMdshLgrN0nP+a43gbGOObzY5UJOOIm/dXTy28GQfic6KNS8thq9b9RsO/tk
zat4VGREJZzYGLO161UvVjgWH+MtVfN9KGEqUwEzMVOlKKDu3C3VvWDrPt9J2yP/
Z80+oMQlQGsvH7sHQzB/QnEXXovi5oDjKWtfmfudnLobMlLujlPina1JRm4TxtPb
7sALsl7tLR5wqCa/Vsg2KG/NfVYAc5+ZzbtsO9tP+/Y8Grr8dgW/mkIbqcWil4nd
z+EOuDx970pWZ8Yb8ydgtjEk7VEx9UKpESF2IlUgBkytly7cZckXDUVG46P/ZAc3
xAtFU9RIdevTEoRCvqZNY10ZCm//RItGh+S7sR1MH4KBoPKMP8Ga0hOIYE9hRbZ7
03JXWrxFO3MH6Ue9jTTgpsEL/w7AFZMr/4lYgf6IdMYOaExxKNSQ1ZQ25esiVBQ2
je4yqg57UExBzna8liGaySMXp+dtVv4mcNy8OnMUrB2t8pqqKS4K3lKhbYZoiqBS
do26LRPrA//rnv84kubdOyvGJ2IF8AVj/NGp1yYSVa/iKitGf5ae4wy+L+nq4g3q
478tHKMBLcoW3xia8ifQTD42Blmz7rrTzb2SvnozoTC3fzbhcnU08yKdYIOC8Z1z
kZm6DOWwDDcpinWantsDoFbAjSjcIeZ/BvVKGbXYgq83c059LcyfjT+dADASKl5f
1AmOJSFZhf1ixKVZ0RJVNYzFCi7jOCa9/ORS7bNmIhOmDwSVuavv2JXJSVetTXqe
gNZSrJkGOYN5EftR6rx3EfHfXDe50KhWqKxCWPhvzHlEzHSFGTkAvaRmLSVyeYpu
DSerrSH86YmZNrU+bAzWhPxRTxszeiBvhAo81m4qr6HsM4UlGvlZm+Z9T0dt09Hr
P2vDxlswvoZTuCjYceDZ4EelVcTayWRfC/ntDMlA0TGOI4cgU/hFGbGnqw6tnKjE
bJhawkk6ltD6ig+kr1tuyX7pOxAyv+ubRQf2B+nIPGq65LW4cujoEhhqmLfdHzYW
mSGeHVl5J61X7Ek3Gftl3Of7Uz83oO5J7tf2SLOEFK5mz7ZlBh2u7JuabFM4NJkk
MMS/bFp/8PI8E8MuZTVmubGPFppPAtS6HEHREyR22co=
`pragma protect end_protected
