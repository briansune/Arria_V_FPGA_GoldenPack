// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:28 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XKH++s2po0OYgc9sgXwPSv074IEMQkJUDQEnXFlX0Q4z3Oka22vVVXLpQn92nNAh
0sPo9NiE38vMuM6daMzvx+lXPbd7iYQgQmvSszh5MfnDWO9jezkNuPjdgPEKy9WR
7ELqghdpH61RT6Mj/YMnC3GP35Rf/0P2TaXYryRLZ74=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25648)
6x6V88roVutlQo+RuU0IGgLQJRLYpHRf7WTvj2sBBCbi0CErzqgDOlbF9k66Zlvq
s8K+1uMUwt7mjEHCcUvCNM1G8Ks+WxiZ53If7JO/9fw0xvqFlllLaWFg5SnL0YDm
3mm/FAmNu1rMmUVBNORqrC3m42sK5Cehb5vV7En0zqjSjVr4WyLb4Jc2X5M7BEA9
SPVDifKHT065Y09K6rc8r884wdb9mTEFz0Z5gE1HfVlb6Faa4rcfdK/tjjoVZS9+
PVJZuuHy9KanOv0EBUm2gJhCskHqYaNYylpQFku4zRvJyZQw3Sgu7FVv0fyXvljl
+lnatof3GpcWSSIGZACDDnSKBbtdw4bgZInscUbz6aGITOVJTcuIMqCMx57CouMY
88Wm11nFglLkiPE4UmeqRHZbnAhTZ77RciSQ4nZCO1xWaEB6whDfQ9cZXTpz7xhT
eqkYEuVHBpWOVeV1O9nkJvlWwTNb5/ncRkwCCzanJUCc1nCM5B/gP6zM0PfSVKNs
WEWrh5N8fJcsfACp/JwrD1DkTZ5pR0fcwWQIcEFHZW2WE3DMIw9HV+vt5DNy+bAc
H2oT4L4+yziFkY7bDJrWSmcTnTec+TJoCdbI5m9uYXiGcWADBbV4b2O/cssNuSdq
+RRm+em8vHd/9VjoYQI0XuEJHNXR/h6nCXLtz3Y+GUJUAhx80Iso8/bUdvNTK0yc
P3vH9PqwYYjYV4BUlzLxyBh3WajfU2hKB/vK3otlEmuWR6z21znvF18j+u0ae6Sd
HyIDyUWMOLJVGCw+BqpBBSktZLaqosuHEEteKy5YwH9WhW4M2diLLvjxrCxroAkP
9Yoc6Tr0707c5dq5QMAT1YZoHxxm3YjBYNW5ResN+NPs19rM8FUh+3ga1douCEgh
wOUaYcdxZWyBm3NvbwrpSZmiEsgNJYPsSJoCsQt1V5i6lUrdDV8SU4NSZCo+6XG6
1+GnM6mXRPc5BClywEWTyFdp4ITsPiXFKrOCXkDU37IlRcMfvApweO5bEL0/TyQ4
fSY1XOPOYxwFJHlAm5fXjN+qMtDVuSW0LV70trZrVgEnFhxKbqulgQaNgY58GCYt
LQ7uWBf+pU6ts6GkVhfHwrJg5eVSeu/ZJPmNpMz46FSlw2iNAKR9AUQ7Qqoq8zh2
RhQa60XHLM39NXxMI+/j2pJfSnoMqrn7tzBnBJ+le74G2Lxs68W9HQ69oXF/sgPh
tvllfgvkYpGLeQjDPNXE+DkwP+V0mg4ZP2zQRhgTlQXGHArsyFTHfYk/qUylTlqa
FRTjPBNyBDTlyvWVoDJNWjxf4Ts6NG+uMyzVd3guW7fwrmgTCalHGdBMXQilKJm5
ElyFPf3U9nTbGagPpkMrx/6YBKQ+nQnd6uZe106+1qapTd60gGk1rbORsc0cYWPe
eS+qcptG/ObWvVH3mtTw8NMHcsOya+6YTZVg6WjuudzfYqrvG/fEWLfZA3bSDcPF
dbZYXd//1G4kDp2fiNwSTSkUhDMKioxCaNlHNNMAbcE1fZr/3Uk2ra+w5fUedJ0C
mroQgUBjq7wc/KF1nsokXxU4jZhGJ3oxoY3WL1YFBmm0v9+CZTO4uBUEBvaIvFst
XKnzD5yiGf/5KpJ0UCwCqn7aSmWjwqqDNiyZTZXYeRzyI4c72CVsGGHeMYvuctoL
Ar6GjyO7Cn8Jtmc2vPMhkatK0omyYN/PS9thwusz9hF8hLGWM2HYCF9GukLQucZY
Qp5sLX2bkGvpKoQ5lSOLS+JWVswcwIrsTZwNw6wogfz6TGZBlP6NgRhCLQqJp4A2
j7ivJECEDw9YmK+SVkqQtjyRZUC+LVZMGze1+YZmLPEQ4lcdGx9z7NGp4oKGpiXP
uHlnVipJkmo6DUl0GZCllD4TsALTI+1FPWJNapdmJZJXbaq56MmybRkDS8WViutq
Eb/PHYH/gNX44KTi8CzaIbZcLOn0+T0oXltlCbshgPYwPwLKMQzakSuFFpgnaDC1
242uTzHA+yznx8H15Vi2p7ySdtZCcjVAAVra00Jodjc4wKjOp0PiJQgtXbHjqrJD
CYcDhnQ1QuFNlDlPkfEJUDCaCJpHfqYcHMQFvR1d+FHGjosiC0lEEv9x3Qw6q1a3
9N0m0RXwFUvAJWABjJAcKK4tfqsZMUTIqtUHzkLzdSRRm+WEtTbYRjVDBuWNNHBs
G6GhZrhQgCfdWaKUC19QPicEwmp444M0dOxSksWpnLwpQte4FcG8PN1aRZG0zZ4p
yoYXfI9VrB/UKbKnJXXkj9+fqZmDOzJikW1r2TLymM0C76XgTE08s8JB2h8rzXja
Vh5etkL7EFdV/dPiFxQkDbCszWibHmmQvf21WY9izTkFpjHO42u9pz6q8ODJ82ma
R/r2Wm+Cdihh7gskrM4Day12Q6U0NWnRF+dXhmhWL8OIaRPpJib4BAK7vcF9hXVD
tQDexDsSIbcoIo6wSgsoYNmrENZzL4ghHt46OHXtJS4RFJMQRaxUcsdsDicttCN3
IKG/hy441yhOus+OUOQ9jwRQy3KJ0P84/zSJtXNRBm4C9ia0BAMVnrFg4stxsqNy
2Xjp0qL8YIMchkovtdwK/d4rvrvPkKazyqyPPAOOrILJfOF+GYKZykAKHQBFHMCF
zzohtztF+VIWZ5r0Wah1FGvkwWe6il7/AavMS2RW422mPCR0AZTzxOuz+dLlB1L3
WVmnK6+G1BAZe6/DVdR16CNxzRIV66iGNKvJ8MmgKBEeFk8yKMmRGXWnW15oBTWy
S75/v2yon71Mx3vi1fGim52hVYlSSu3HzUQ0wWnejHXEnoT5GAmXkLo/VOpa27JI
fM5lZczfFLcsorWIUb7pWiqsp4dWiOEMgl4bqJHOY3OSGLMUk77jAsH7vUhORGO9
1QM2hm8ITmaeAwVxzx6jhAUspXvbQ2oC3LDpOpg3TYtArxulKDPg/QbOZ1q5XRaV
RHu9fVh2UJKLpoxecDjUhr1oFETztciaOLUYJ0Gn6BMnOJ2fWsUSb5C9QtE/aA2O
zazeVwfnzWUorFuzdneZpPSpI5Ll2i1Y+ioTtS1K+wj+fvTX1XSox5Rpg3ixw4AH
IBZ9QG0aFypcpclnfYROj5ay827nJfV1AK0io/eCoqNaJ0lH+gHOoWA94MhCueI0
FSig1MzTJSBEOUaUg8cELNeYuVOqdU+m+zDc0lLkZrnDuRsHT1TdLoo22bd6XD1K
PoiH8A6szU2xBcs8f+oOJRyNcblzJuydp8nVWhJJQk3EZtfD1Gx/fxMltR/woAlv
yvjyu/rK4Icb94qH2REUx8N2OF1eJVoVJut9raMIzX/pKP97FOUW0TfSwn2pR6Td
AlUfLodB0UStqse3AeP6WgiW4ynNhI8ApOpMg0ybO8yQ/zRhRVXJeTLEyZr/6o1B
BJjt5VE6OLVK1V1/JowILxUutG/hdChXMQubBZ1Vmadi9bWH5d2HEuWqxWuWo2hf
M516JUTEcW9OzW4oUlbK60y1vBskRMa0kC3PO2XznrP8gxiqWWfwTKmFNYowgLhD
4m/rY1a5oii5J3CeikvCOOcX7HMrmx1aZJiW/XMQbgY2JxPgLS5fXwKCrb034naB
+YxOMq4ogcA3S2/Kdc7cENyFspgtEG7X0phMrxFXqEEHyxALjdL9aS0O+SPTV4CD
Y8EJzcnrWE6H7GgXBVBrt/2ylcoD8Oyx+Dun9P0eb3fpB4Bcl7kMSfyyefxCGCfd
ZOAbwnCVPOhe+aAynxrFn43BpEPxPDLF+4sXH81sMA/1AgWRbjEgks+9iP8rRss8
clig7R9p0/ea4ddP6N4rk33WcZGd/+CY1/Uqz3mvKNXVVtoX+EBii3CfCRUGnCUu
lfaOE0u3ZfK5b4TqATcHEtfCpvygvbeNsWKtyR5xdi9aAshWJJwZstmKi2yHoSWH
+C1WrPedS+S74MtWPj+Ww+xCNs7zC2RzTijLNTdv//RZiRzYu99jfkPUdNWKUhZK
+Z2HDjnMLDVCr9vY352OcC0Rapk2fn+Xwi9YQxIo/fkMPQ5JJ5AtBBq8Ggbbh7g0
FgRn1o5mx5o01CaMdfVSzMVk3FDI8lLXHpF3I8klxMKIuZQ4volT8MYpd93T6Z5M
lw6UhS62RqULoAkjywIw5dROaad1IMP2rOTEgTnPVKEWEYS15dpeMhnvVeeYXW6z
vbZ7NXDWzuwbuCSmNHV/DpVIN5maHaQOFQ8RAJikeQH2LEZkLFIws/HX9/ZESAJ5
qnoL/0NxaqPxBbHekfN2tcIEHvmHypeqeCc7zOAUGHxHfPmoo5wEL81S/HfqPrk8
xZucGhrJvmfHNTrussZJpKkrJNeUg+6puOQvburgawThV6B7bS3526Zz+T6fu4kw
qI6G78hAPC+lzRzrn3YgsOYydFkTCiL6T9NVtwucY/AceForyWZvNKAGiOrVaWP3
kYrm2bxvhldbELpAvAeHLU8v42knutPuPEF/XgihdRgxkkHWQS3TUCt9WMfEc2/V
3AaMG7vLMUGPZBzJ6qjRrjLdz5AazHfgTZs2CNUfOGf0fG920PDK8PmGH949nUXL
JNk9c4Um98CEiF/IGsf2iaoXWkXJYvpgd9pDQs29xCdvQFHgUNF/fkcMFvbeVavE
MRF+JFEu3c34Q1bBIFhVd+mveo6HjZe7MUROaEv/DcRb6NM7EP2C5ITfqF6fD8ZT
5Z1GhavPU62jkRGtt6OMmoAsBqtMCs/WTQkgU1ES+Gw8FMuCo7Sf4pQtj1OsAoLq
sjFdoMmmM6uQMFED2bqwHu8jb0o8wy/DdSj5dnRoJI5m8UyK6Oj6dBMPe03Vl6HV
kDXxsm6jZ5fz5Y+DsuSGzwIuvKUVpfW4zd0uIE+iItiprN+lkdiIvU00FR5fs9jC
CM1Z3lkDTMCZNyYjqdb6hHPLNqNh3ona+Rm3XCaDZ9iOIvgRzFT5E55hJNHpLKiH
dvIZV+HYZVjixKqlxsxovDVSANUfHypMW41MNh6ADAJCZdAi+DcTtfqHHzk1l29Z
FBY1gou9k7F4cNh1SDwUUcsYblxFPjTNlbmch9tRdDERz8EvRPPfgHYi5IgGO7QK
DzlNuS7rpff7QAKa1IfdaisVe8u21JOPLdaZMgGvW3aeGEmlM/i6Pr0F3hniUcHc
EDpObnOuZCbCjkEaobT+kr16n3a7ouauFTngMIRXuc1Ds2MDQCkBGW1LMFaaT+JI
OOVbBL4vJF+9g41J7tLw566yzHAUtIhg++7knnPU8klyG8UKBimqQdoIKah0ZdPR
1kdSnU4UBSk6Ha7pneRwMscfzK6A8YldknGlvQoLS3Wr+At/ph8RAcwYMDuASeJ1
Ye8Y/JcJQb5TJ71LJdImJR35eMpqDxFMq01KTcurrfs9v0LAI3LEts6/n2KM4hQF
gyvBNrpIMA94d08fC9YG6T/dS4UUG3gGg4+7uEp15a3PKQAfCIeN9NfD5aqKfSnV
WdcN0qMbdUj5Itjr9Zb4B5+SGgbFSCM3VX/KH7ZHCOMJG8+0Fahhok5uQ2BgkwFQ
jaozwbKw0QAsrn/uFUfD1ivPhILx7/8T4rvF5ZdBL3vKF2tfdKnj5OWzqXpT8tzc
Km6zwvhdPEDyXnXC0h4uO2HWf/ImDhCfLIddvzqimE3LMlXV0oviS1IlhAOjF2H3
Ajyi4XQhKWmr44usWwySQftNXrD5r5rkfepq9zgrZ8Y+P5Y7q3ENUsOIYPBmWrYa
frYTT47oOqcdRUeVZiqgyHpUlHNfoYcJPUW+Y6fwdpFt1+yU2WSh3STLUtzW0VMv
CTnC1Cip5DY4bsoDuVvbl1Lglz3IjYcGAcqb+yGqcu+HpKsD4NZjPBa26kXrHhGw
j9cMpu4W7jYEMWUXNRJpqTAI4Ug7SzYmt6qQ4W3DqLT0PKYBFZ/NKZOl6dPAG4cn
RJEEtuqVfaka4z6xtlHxmqxEq5ZOnC+e2EGVw5G+kxpQGvu0qWrAGKlgqKSMywos
9d55UcJyYU/LrIKMwF53AKUXshPM2jlqaVREvD22ZU198/YrH5gLf1esv4xRx+KD
8TNFpT6s9L4UvJt+nOEFIVzxoXGSEnSlgIj7lGYxnqdfyosi7XLKLwOQMv6oRa91
lfKHCU0ZfozeCkFHyODx1cBa2tGqpWh3MNlxfI+qkNtqr9wVc4XkpDXRR7YTi4n+
2SMXyM1Z1oVC6xSL+8OAFJEaSF02+haVKiX4zg0MPtJSrUkVOXSAdGWFK/50TCoQ
tG64067axd5+fOPDz5UMjFKsmICyHhuPYe1dH9Ksqce01w7j1K+bsCgiw9kf5Bf2
p1bSDGcxAotcU2ZPgaEZz8R792Y4I9G1iwzmJNmZ4zYf6z6G1zOuvGXC834pBuCz
G8SMWC14MSkhgXfz/gDaE1b38U5ZivOgFR6m7BkaOfSWuwHpwxTKAcPt7+jVyjgJ
hijqMIro9nFhAp7Adtd1CG45cGUjeSxtaDqf5NI/BfmPtRpsUOu7mvNxWxVZwb4k
2OnsNKTk+st7TSPkCXvDxRg/C0U7ScZiTgd+vLKNa+mric+MDiwiHBnOnieHz7kQ
vR4zYhFZgRlFpSH7lY7EvizdkNwXQidFrkITRAEXbCvUU7mMziL3AY9RPtLj0qhA
gLyIQzMgL6f78Fdtjh/Pk/+3f43H3zpc5nF460dRbSc/+Hityx27zlFoOoF2V7OZ
DEzRk82AEvBPP9cp62YfZ+VFM6QuNkR2T20/ElWNnhxx0HLxdwodpaYM15ma0Hcw
gd3oD8Ox7P4NaVLJWXGsPVwTGn55Bki74bQX3k78YK5TRBEGDj818C9AkTDusOrN
FUFtcL3Re3Ptvq7IXF86F5BmhRrCUZPOgNIjeZ0zODVM1TWSPuMREgUjpvv977u/
NUCra4Ua09CBo7M5Ewut+C/6yQbaO8YOhlEfmmfO+Ylqwst7X2SEze4yog5sQl0L
HHGWmBvKHdo1vkjbCaTt7AnTFFHenRjBpkY0r2vKWchnSqKfc9Z8B606AcmS6OHD
uwlbOhz20q6g2ze0MVQNHnu+baYSGEQvwRRgEksVcjGdqsm7aNRuE4bjQ+W/ZngY
VfDmYBG4AnhfUb2X9KW4QBLikfbtI/K+u8UgC9Die2YZLevxsQf2WsXmugAvgWv0
yqZANkhx/NGZtWQoi6QnWC8FOZqbzKOZNtFlnVcFKsELUn7/1AmMc8jfv0A4K7pk
6rGD6pRAKaBOM4T3UFC1EvTKSGEet9vox8u6L75w+ewdeIzjZYyLgBknigrjRXET
55/cDH3sMgg1KLQR/eQbFGDgzRZKHzJrkC6cU81sRWlSFXmzRoBSEL0KLiFIgKiz
ylcqpdhoZVVc7XlbgGHZpeUmEeQn0VsHu52f2uXEsuP8yZjX9z+T1TSHzb7RA8ko
PGK4niQeQ1+TwfRZTCYRmA/+vmV1o4VSMV9xUV07UC2O8Rxt5npME2HzvhebqnNA
iah2MO1H1Bd+LCGm6PIrvRrXlU8U757OeUHey0TAkSsqQdLgTM+JnoEtN9J8bkvR
xLA2ld9uapd+/3OZ55WTxRTX/puwWY86r20YFCnvIWnjqP4jUhm68FloEE85OL7o
VIWSPbg9z1W6x8hfzLbrFVOkzXapRf1KQS9Fep9TZxxQ8/VO4/m75DDqbXsDed9y
ONk2UTc5kovHS48zIybuTTEsZQcfnEQI8c/P0Ux1tn3bdE7g0I78H/2/CMnDq6bF
gNV3umJ/owde8rUf2Knn//55eyJjpvOsKiPn9137Kgu6w2I344fXtjRk/PCZwYFG
7gNuFSa6TzZ9nl0QbwwOPcBztIGvLYI99Ew4pLLwEF+YBThWLbtCeX5m2DECuSBx
VnNWjAUP9iF2LXTgd/Gf3lbM7Bq7Ztb5f62vIDoJoY3A5rYQO7g4iMOba+fuZbxl
07FvJAwF1zANbyI65ECctLeHzXxn7Ah7oVUXkN817kNgKWf5ShRNH80vTKZm4+dR
tXv/vogDHeFoYiVVYulvB9CEwyq3SXUiENq0JmR4l0rEFRMo9yZh7d1SP+oDmx/G
jm0aIquHMXIW5euZowoZHSdXNWjLkgrtDeIwmFSGPjaPMlxtlGER9JfnD3ntUOu1
rQxHigQ1uEt8fOYLfO6rd4tjP0G1CqZnxE+iCTCXYfHF4K89htNnsElvt7KdD4RJ
Hc1l6p5/LyEHOz1T/lDfZMHn2DT2vAxUp0PHgjcvaAqeIG/5CzOOEFstM1azOTab
niupN598CIL5OAiucUpglymPEhybchg4mYFElFDJbRR1ejXaoGU3AeAHzijjH90Z
6U6ZHyDBWz7dBCp4ZxhGywcYbdRE7dqAOnbKXXYWaEmXYKq5iO/3M3tKIIbZqeyQ
cS0Cvm6U+/+m3mgCKHZuoJPaNAU1HlBWkW/EHIA3v041Vf0PDXsiMrKkV6cidI6d
xcsmiJiRNvNtZUNRK28Hfa5Rs5xCvu70jroGwxBhEngdHXLtu+duZgeFQdJKS6ka
QSfKp6WIbG9o6twIZKJcrDi65Oaa0ffeZP4tSYPeE180Ed9FPUjUKWpkWNF1Z73/
oXSwEvXDV0B5DypYO3r3yjfeZ1Wy4lgmUG0621wxx2Al4Y+iHU/vpurXeZcDSq23
lPhJKbpVFz3jxfifSYYMVcPrcqDlgz0tXSSFmB40/DUuyVs4q3h5A2TAsyjEy/cw
f97pjKpfH66wWL4iXWSsrNMn7PKFcxy5Synx7Iu4QVgkmz9dKE+DW5DNJGp/2uRT
5xTGQIUsaZXbeuQtqiLjZYs/mG62U4bEIS44b1mXJApeUQdL34nPzd5KisZ9J3/r
/LMd52QFaLruDply26HgRjSZdkGEswcD212K2J8RIpMGbuFCEblHPAS8rJiTiF+v
b9MfUvIDgrraeuHXplrPs6tDYFcBCNZCOBwezscegePAWpLojdS2k39bUrLdATfH
DOGkvEe6b7cZUm2/vUo/faLkQK3R9SWxiGIMwKJ3pnB3WOXJ+dZN+aBFjZzN/tNj
KdSbQ5o9bs+pQc053NLP7ir0G9N7Ij1GPxPhVIN32Rka97bnDjduPyh2hQ6J1mYJ
y5BJkbUORkHUI7lQWZgD2i3Ffv1ECnF/7ugNmXum14+9RBe8UvMmCkUJE1ScUBHY
mdgb/TixEv/Y2hrNEXhl4FL4ri8cVATJh9CtgglPjF+bjDSp7i/hmZGYZSdGLCgj
rQXOKQ0DH9zJ/PZX6OOEg7rCx1O+LehdZLLaZ4GTZsbKcccN+Dm6K1qa+DYnl88y
8XLUYXnT+QlVXfvc3PkBwEgZWWuSQrpygNwu+Ifpktoq2Kp8UXRPGyrgFhNrQZ8R
O/6TaxzWvXRZ19C7JZsWpQfNOaUJovE3Ls1bXuw4yGMXh90EPYB8QDrPDyCoLfUp
V6BOuG/O6h33clGv2vo8u2MmApAzITSS+tB7i9QhgmbyXKgEsupjj0CAyoRwajM2
jfCL2S7gAC41jF7HFuwbG41lRcAlIAqZNlqSY8kDfNuIZSejXvDfv+74u/HmzaVT
vF9a+9CnTCn1CBI2u+7a1rc/BGvkebtnVxyCfAUzFjCH+OrneaJqL13qa2VUM/Xj
yTv05zHIK5LPaCSi504vM0q2AndK+9BzFPFRJL+TMgPlkH4gmFRo4L/GPZ8RPcYq
xSlMD5tUGVqfjxAmNVh5P+UQhdqqstdo+kBqlZA7hzFfqn8wtiaExn0p3DzXJbtt
k17iVG4em1FGV+2Tpsw9OvGBU6uGQDpPkzXHZDKXEj7aFg9yADGcPeWEf43Yw22x
cdKrbEeRUWOiYZgtp8T2JDg/rbB8cVIE9eyzew6cQl+jz4lKXfuJfq9OuFk/j680
++aV3ZzYN0G7jmxX9ThDJuXxSWxN3Sv6Rb+rhrkWaOgCpKdB3EfLBGnYKbgJ0skM
LoTcaPW0rufi1mGymy6r35SXZjmBvWRcsyjS+MDGzL+gYaj5ICQ9PgMC6aNEU/sz
VWmsrthshrXxzzthXp0toNtUIhm/k4+XcoRPcB6+IkidlJ7nlrXYKABpyo3hegob
3HvG96vkUHrjSbKrNJIleWSb+W1QzYxDZEDusBeFPQEKQHvqPuiO0NzA2/D9SG3h
u9Y0AFyvHKPoARH7GXWCpDNtmBdoLq0X8GpwDNVH24r48MjjROop6MmAEAVitaHc
Hc+2HnvcwfbLqg6gUbpNciaAFwIUGU27FbFhM9CpRbKjnYVehzftYasr9gJfy2ZM
LZWx6t6oKYYf9BZMWw9mRqxCM110NTYDzadErsYRR8PceFw0oXlG+p632iWtHyFm
RDzlNcwBgSYq8oZpu5yFmQsQi15pAoC4mlvN65UYOdLvdo0xBgcDDaZJV1VtC9K7
NN2xWx8CLMiyhr/15uZYfwnCb6AgxlqTs6pW5mLoJCQ+4OxfoakrIjBj0IjORxMj
ks7Pni+Yv4XzGrr/29I+vkDqWyn17CkXSCKa5En7eMNq8qTizMKHESQZOphAwHtV
YRzWOuoZB1Yw/YCZQQUqr2qfFwjPsKBqBDNIfUzXIDZNlljjR7idgEHBiqpJ0mS7
3r1H9KcnUh3CHtKcS48LJJ7CsTt2W54ilk6SXGPHKzC4+FjZxotReffU2NkwhFb2
2hBZkwquTCdy+smAQ/6iYUcFf9TeDaZ/CE1A+UQA11bVbLiVA2yiLuwHkmeEGKBD
vnEJ0zJTJhzz46uGy3EL041sPYGGIhfNeqoqSvSwMq1CYsx6YjDZbtYXZqD6lJDY
kNa5t7Eu07KpB0KK1lx99bPesUOEcflJ1CR9q1275KY5lQqYyrxAi2enXmQHkHQU
ODgXld/hVB1GEpn0HTOQoJV2kf4MYypsQWlvzB2ymEYO1myc1NZPQlKDUtXe7xRg
VmE5mbEGCKGPPRrdOzJCNkUXwLy73xG5zEhTWKWKHxfOq+ltmZ3FMzQjrd2uSTex
pukivU0QdUfGYTKjNy5/MvgG4ba0Z5DFJ9p/e8E9+VL0Nqc7criVZGziqOUphCBb
5Lsdmc7qF8WIB7brt0hOZ2D0+lQek5A8bRIl3OoAMdmMQedHbsljrpqnO268u2qi
h1cSRwIZ2UWLi281v/F5+fo7Jpn4ZCSePrJi4sgp6w0FCGKhWNZMHM6Lw8DGdsYR
pQ/H2fZy44/8UnUlfItPmnkOI+Go67CZlLnXvA/HBYUXTIuYo+BC3Y73bYZLVZ0Y
75n3CspTwE3VRwmF4Zx8XTa6W5fLBErvOiUW1h2mHDMEW+Nywt7i93tpwfM4CqiH
RkEmpxemYcSdHchrRenjfIXvizxxYv8qn0Xu/S+zK+7ON7Tp99qMMsd55frpJHjt
lZxxeEJiuahIZb2Fo/jAxqq30CANJtuLapkSZ7ZLH4pnM2LxQaUz7cnXPNWV06NE
JTcJabYxg9boTmGUiC6cvfglUaj0ac+ThhGohyyC3eWbFe4KgczQX3hcbMqxa+yc
ZDEX1WhvB78W5h93MIINCoeAJIXeEpSSe6drv21zEa371rxXdy67c1WQQ+zavkDP
PbZZ0P5dLd2bDLGYSUXq9dHVcTmhYZLnSJyeZ1KCenw3o1SmcRLHmD1De2D8l22Q
ho9lNkRDhrLTF4rd1w8HL3oAbYAZga4l6CmNyyuYbfICJDvINTgTN56z9TnuWnAx
+1z9oCknsE3qXdblFMT/NGS0LnAlpFHnXWNgxuuFem0oNJORXxV2F1gv3WYwVlR2
64Fus3IUCWgT5e/7jqWFryehscZTWqDadNEFH6melzHkFN+otXgnkpPJ4M04UOrQ
eLDhj0nLCGDySrYiUMV2FuOGnr5tFhDJM38p7DqO5X1isTLbEM74w9K+HvGpsqG6
r07sspASx8s+jGb4PBOHjHo5Cv+WRtJyHbq28p0w4SBlF1YEQE+8NqUr8oCOYUFF
hTfwqWZkqB5gGwCl6+7jle4/3iI2FjM1rEVQz/8C3obw3hov1Xo4GLayb0TreqDe
8T/d1xWLGimvkKePRZtrv9zQ8jO1QHIQNOT9zsCtnRCHChMBBg6hHkXTMxxhv6Hm
2N1OaxA286dfGgL5EHG+KQooLqvJ4zzMmSXWdFblgcDMyl4iNvSFJ/WHZHd+3t1q
dYoGQigIOhSnTQsT5djL50jpLWOxXy2dYWZd0YcWFCluJfkSKoYR2I7NHoDWXne+
rE1CSjSzzuvovowUFnBbtlGdogd+dQfAgWIkiykRURW/+B9sipCWfizdsvnUmyj3
M+SXxCMu8rX1Uug4GgdIqt6BMPK7nf7St6UQVjuBKH0XQl/fcAM2g05bV6g8V8kY
gno0zGRBVqHsu3VqF98PqIGh8KaWS+275EwrhGUG/ctuURDL17eRxVF1qNzw6hKe
h1+dFOjnC8UQI36yKykx4DGTn3okNq4RsVxjWr1ZroS0ITmFRUFIItpW56uryDOq
zSBy1/nX3RP7RMdKQkGb3akTwU/IyeOg40MCnmYljZre43+kNge0QoQ6W27zbYup
5bCP+HHu1U/J1FwJ5yfoBdkwuQ3HcwFEvBIAC6O59SuVxXLTY5VbNhjqyRp1ASIf
EegpmfHRaJurVx/gXCSazdBtFL1tu8X2was/P3Fn1TZo/VT0bJ6cCe5Fk13+qO5S
bh33OCDKRq2DVi6DBvnpmCmZvJuuE3afxfOABGEcHOzkVGC3I6jS3wqO6v14uNyf
QrbYMrT1CEhHUQZw1X/1FP1FK5oTm74cdwkBff/qqYmeHj456Bm64DyPxPKtwJt/
fMMCXCIVmp+jW8B4lzwy030Ku9NKb/Tad22U//Ge0NS5Ofqes/pxnCp+re9DBuNt
6Yz3ZP9MiiyonPp8KS9vDOTvPusTjedHxIPX/9rxoN5GF2R4sg8zCeXOURKscSwB
F2gII4HvclF0CoX/P0IaXi07zfxYIhiiqQ7/HdoEVcveaDnOcsCyYjcajX3nU8ZH
afx2lLYoFI8CNUv1FDXaderrHrF0MEMvskdOlsbAV/XTZoV686WrXhon1DS0SK74
EdOQi0oMX/+RrHIaHhGlGAHq1HRJJqJHDttvM7FPNGlQ/KGCP8dgdOgkLSkZuogP
nA9bnzWO/66XIJEplGBYLHkDkMh17voTF014Z2qWQ0pxCs64KJ3zkz8vytyEGztF
3WRLhVT/maRENozEZgH1vAZWxXxS8h7B3XCtTaGCmLseiR4d1BhiRb4W3l0i08un
SsItcz/TocDll4I/cEDfN7/e3fXyb0tDSB0DQDaDd8vk5FHYl/XVHgkBr8dlC70p
Ddh68T11aGoY2KoHcEgUcRLZaBIhR2fZC+FtGJ+mzf49jiSkYeEnkN5YbjinYjeR
NxxDMjJoITRD4QTcChOjuyLcQWhV9PyeBnL/pQutrpGkEG2foXNtQSP4DOss99BV
RfONMk4o43gvhH0vYKeTAYn44OBobFTLdqgJH6ZjwzwPcdr3A0wjrQiw/C9m1PxW
sJH4PJy9/urGG3o7TsaX93EWdAnqNsSh8C48jCG8ASfuxmVjncq5DYHcRpEPiMPl
wSSL2Wsg94oOwsp5aCwucyS6+S1zNlNR0OCSb2jKO10UJDDknpkn8z9tERQhJvht
jaWx0U0Q5onwDowW+GO89quFY4n0cnbIhAF11flL9Jt/wt+wEr15c8WBvPd92/vt
UGyOzGO7yP8ypf7MWqHOG0n1hU/tCb+yh3i+q1uChiEUYcZCr+yeuC4a3EzSKc2W
AmkxiOixr65D/8n9sAFb/oSPve1xLSw3m8Z0uC4Hhv8yCOLVo7iOSYBwo2GiVlMc
tc5pivyCgBi7Gv5z+qOwemvi33URbDSAOPLUUaOQUzB56MFI8NpPmTau+mxmMpKL
v/CYXxV4AftJAZJAkp/3COHZtTlEmDJ7y+kRT7inj7oivXcpDJGj6ec+BAmQ3kqn
gbbN++VnIvsFAh6ZmsYz35i+zbL+do7x8ZFGrM/ccmeXzcNXK2ylUAkK98dD0bcX
0JjPfz1sb6trar5TpqqPSftur7pbFMuD+yfC/piDt5ootYDcehXoSg5mh0MBaWgZ
c1dtZusmY1POi5HHHrUGc9eVzO88igYjUiqgEx7nI4sT8xXiTK1mIPnCd5DPhshC
5z89l9iTBch6ssNXytHIFwcW0u3HnPXIVGb3agze87gLoWTeZ5XWO89tcGlUaVLI
xGV6e/ELNC/YKl5cw1ldQTd2MdZFryOE0JPB/MuFder+6m7fBIQgN9/J9jwgLVEr
EOA1AfwQ98ogQz92YFIy6duhJ33EH/lrOH7m94bgQwBen2SvCFHNpCFZdWoLj+Hb
L80y7UbTbZIqI64WQBACtlwISB/TBbNakUmddDhesQANwb3pJSXS2d3GkVPoi/G6
Qa4atqY+qXpzdDLzATLs6ECf6Sv02BqRi/CxEWFUWkuGEeq26/ZyZq1Kry0ekxXh
yymhht9DDWuHmIefJ4Vje99eI6vFai8GQdcN+h4vwkDkif0V7YuddNH28FB1vnI8
B+KXZYtRjdV3BZ1upKbN8MofWPO0dxJCdQaHCE5V0tEyaar0UPDmGp1fSGozxl70
MT2mtNgymGsUKPRHHD+HE3Cy3IEG3RDmui5v+Mt3gOd1ciuiZtWZRCITI2u8Pzh/
U5elhnnPandBrn+/btLBFP3ePqxozjcckusoILqXQv9+lLcoksLf0MPiplfGllTE
kSN+NC3BrxsX7L2kmV9ZLQK7oQntIR90zy+kfqzxOB2lnD0WWlSZhKkM3byGjzsv
2+uwpX6b/gPUesJXwIJOI4dkg2RWStDmD4hAuUNTVHdomex8asHRuyoL9uP1kzNJ
5hexF6uH0Z8UmqlFlRD3ec6FmaxoZJKR3h7P0LFrVf+WARjE8eUV7f9XIkcePGml
nCBCLvVHHrNnGvFehYEPDt72kNiX2Z4tzPeowphQkoABv2U/RF9jgB9e8Z4cf+ql
IhkQeQY5fc4Xsk4EIdaEN8LahPIhOpgDAGgo92Wd0trnjDGD4yA8UO145iEpHq/r
3o8sCK3ykFIIolqXggtJSCQWFZaZxQdE6Ik0S1zRu84I6BGOiXevlnlK8ttks86x
irfAUo1nzQxeevQC+/hK9B9XoFqHVI6pr8Mg7q9VZg95bwG7CSKR5iZ27dfYspNC
/YNc7Xc/l4PaZF1IziuQtn5tcG9qkI20zwhT9METFdzUyXiFG0Ec4AaMzgxSZCeR
I7LbBKb5xZdg7TJRlCjR6B1yn8ErlifRdDIo8ob393vNpk1UjYB1rrwXFeHyAkQt
hy0u+RWr2arm5cYlC6kfRLxAidKvyamUAG2G9xGmSv/z9Trw5Q9HWE862g71vUbE
V6Aitr2LZ6taviN2Ht76enCmxpRyNQhanwgASndFTFIsLOxTE8lz/xBTHH3x8RUX
iNOFQVIFoprlNYOG8rqgBxRInViklttXgmr8ma8vZA1VXCmB4zK0LJinVyi9BgJu
8VUAOxfQVNCViuQuSH77+DIm7gKvwaxRbD533MPgB6B+a4rbJprvRZrnz6wViTxm
tYlLc+Tjnupq2AEx8j4OV8U6lKCP5PoOgXwtU+ZKkqHXOp96F2DgaSDkU3HKbhQM
87t4BgOFpQwOmHGg5RyXkAsPgiyVuxtbWDroT/LBVpoZqgCv6w6pxUBtD6vjKMM+
mzcZLR2kmBycSHiJYWzeQjetmU7rU7bYGLOACit+ooq4F7qfiRcLh4B2bgAHaAJZ
QFzrH0UmVAmRHINr3Go3J6zCAfXofVm8pHtD3uh/q7K5fJssmDR9psidPTc2icX5
rnhYQpD95tNS2UHiB4sgKe1r8c0xaA7B8bFpkc1FuPoyporbozQN4Kds8ArYT7k/
/7zqlc1Fp64Q+B3K4N+CblgtCJ4S58+mrtFYdgWmlCrtyHHKnkBQeEJ8JU0PYaVj
24Vkc9RNe+hu2KoqpJeUWupYsstVMM3GeqR86ivLyhelS+OKbGQIph+ZEwOe1Owo
1AMZ2hO4ZqzK/62tATgcnzDDql9xBn5nZMA9eVklpXl8K8B1iWXZTIhfK3pts7Ee
OkTN6Kg3/eyKodKIc3mkZlZ6+SeTCkns45Uq9N/VjSYb84CNcFgf14py/MoqF/BL
Wa3xykjhr7GrsYHmT8c5mJAgaReZFleVri91sQuLdttJ3cGzTNu3b+oPnMZGQ6Cr
20LsBt8re/IA9ZKxc3OoaAVev9tJ6/kefuUYueqT80zOCW/tL0Iofe0bRt/wQx7r
mawBB6Zsjt9TfBietkpTRvkiNXukfBY1+4LEDzMz1PIXjVfjbpwnJp3NCuQwqgD6
/vq5UMkah5ehpa6e64OA1CWZ4otaTfFhdT2DmvhOqVhyaoNDg1tXzVdrA5FU/iSm
Kcyxz1qUS68YUdWP2qSPtMOIRhMlfmOOfsWX/2BhkUBppzTqHFYBrCOh35SbUuY3
qnU1wgGcu5UYjhHPJrGg4917T6BJy+ErWiiPVoLZhCXIH0GX5VnIJA1xXKkf7uZ2
c2cWD++ZwPPrJ47oWMlhO0ZwJG0WPos4LLUqw2QVa7PDnw2ZYCXNuIKsVf97ehk1
r+5+y1wPQngsKwrfA10lCw53P4OR3dmKBvTd200bapfjeUa2pvQMstE451/0yCHL
c2eAoV5Uh8fSn9eVA+07tWV3T63JtkFOE56v9zEZ1nspqLgTX3ghWck86bcjTGB6
7sk/gBAp+F1DMxWaJTcLrYvEZgcTo6YKW0nNLoyh1gVxsHpeDJlLiq6rL3DOz9nJ
imvLfcy2joSrxBaRJrGhHidAoXTMULS1Gf+l0USGJ1zsm5hth9wiQG9pih69+/w7
qWPRd6xpPeoz/MOTDpTyvuv6y5Pwa5UQJnT7dbqFS0qdUtyFerYYs6Kfj7Uk7bsX
Pfp+cuh7bp2UpFGRNVm+Socujpe13yYXK+7qRArD/I/1mQkevPryD7KjvRnAMgXZ
0e7Zpo85F7JABaIiS5KHcivt3wv/OShRIDsCFyyoHS47oaWyw3zgtN4wDGm+GSo2
N0az6IvFNaLZkqQaxaauTWBxhhdKZSWp68jf9KkEsAGSNw1u0dpxUCG+EbehN8NY
7QkxK3jOY5KdRXNZ6SXkktFz+OqQJ2wCxtsYfNSxnl+z0NSobWTpGTbaj0rGVvZM
VZspIe/7vJJeFgnR78PhUmX/IMISiT4oTkx3f3VGc2Pd+uLFZW0dQIIlFPe11bXE
HYLMVUmxHaQFoUIDRq0fluvOgu2tSkKABPbdLdwLmADPZ8wyvmHEAP+PnjSwvaaG
RSSakYwYQRMwhG2/EZE6Iq50lZQIuyjCOwrdzFT8CcetweOCCqnrgXAMEo45BfPI
vVKA2+rL5gifYWxFPgUXDFGFGSCFdbw8ZQbuc9UHJkCeApdmUMK6i6I4uWfXRCGm
Znio9ReQSi1RA+loVsrj3MsZKnzS33GwA6HOH8MZHIrpp3X2pPVP6e9L+MqhOsaz
KPI4AnyWAEArVWbnv8zpqqPo9crfBE6FlCs1nb/AFAD9Z8SD3Myh6NvFEuqWzIxu
zZAOv8LsZO9gPis798s/PXzc1tK9aIKyGwotmzfg01uwVqFtPq9RabAl6CY5UlcE
lpBN1phVqbxusmpmdKZS+1hPd7311/f+Pitslo9AycuhV69p34uPLrxfgttHiXOM
k4coyhRDp5MB/qLjPmf8U7sqbetMWlK9R5vx7E4vpRg07YdqycNtJJELHNICzKe3
rTPbMk/BF9Ve5Jo6+ggyLyBtlNH4DB5yhYnBdQG1QebRDEaI4pMg4mDzuQL3s0+H
acrq9M+WVQ9PM+7KQ5n/RvYBW9WIKR28iHjK33zGUlWJ+e2OZRkVWgKtltAj4bdX
ySzXxUQGWeSkJu0kmgiN+fk0bQLZ7zUn1wKIgWsaG+aeUJvAPKRfJO2UjSmQ49Hp
ANoeR4CCo6uZI/SI3gVYm3jo/V1Y1CQobnA+MuQY29DDxIe0YsxF1OlsthIn8Cr4
Z39Qt1WiSpUqSe+hVSM/qNTUvUynvRNIweFsu7Ufphyuc1W0QeTRs5m9V62oeMhc
8DxAdprSy5x7V7FMt0FhMP3fs/emDBVUR+A98/dxeDiGSeD7c6aEfrknMjfLP9QO
RW8A1gjB4Q1DWllliGQdUiJsOSS+g+duObdjnKm42xqnFT2E6Zkpq1XrnY92ldTD
RML8ssCZao4e4PEcSY2lLWar1Jgz0SzFc5KmsLGQUJ5+UG0yfcPpJVTGRWW3X08k
h5z0sjAi16SUglVRFujYHDAbdjk2PuQVDjZG3U5S056LSEeMXHxgoufypxLzyUln
ZgBbNX8jGMV3cICUmGkbB54LrRkFA5OtSFb8kRqIzGFo8YqaSnjuQElhNdeJOB7a
ntrW1VI2N/rJsup9H37MIi1XxX7vi6ppuzNZV6XbVOoyhXVB+XkBIvE1sGDuyGXh
xT7i87nc/b1gIcVYMOC4QkS4JDjVfb9rRGqw0H/9Xydg5zzrNMh1PPY6Q10LjtNc
+/GoY9ZY72FdDpPj8/wAMjQhMMtsFwYU2bJTN/l4F6OTConN1L9rmHoue8BwvE/J
U+TJgHwKFEzOKVEmxRJQuDWAhDO9nmOdGYD8FtSSLr7MnwEYAbpYePp/WcvdhXZ2
tJhY4jc1aLs9MXTmHlSec/ezyMBQPvXwTMP5IpEHKicFaEtCz5xoSSXmeKSTz+le
zeYEcP+K/fyrhHpEpC7e9kWAYNQ0ePgf5HgGH3v3kVlIKti7/cre7D90+opNiA1J
JrX80VLQ1nD2WS6pxwL3sMFdpYQ6gwuQzz86H0cOjiCL/vDNXIpwx49e77ZNCa5R
//z9jzUaSV7lDm+E4ASeZZlcJQ5jK5JJtERpnap+ESQPNAz6lTSUI4ZfaXG1+RPg
owffz+5xBx/qlfa2PNxVxKccDYSiyT7egs5ekfQ5G4JCU4Nbtb3hfF61h70AsB7S
PckhfZ8PifnysenaCcw1WTMf/Rc8MkBcqiFXcBaj9zaQCSv02omEps+E4nt5yaDI
3TgJ9rQIAA+RlrRedcYWRBw72OYjQIPD6QoabJdLjU3CWSZ/Wt+gROXbj89S97EH
OLsen7zqEe0y+/wWWp3U9AyoqhFOVp7KUhhpz1azL5g3m2vDdRQi7JvQtBaoI4dw
dVFEYxuTGQXmenoXEGWzDvHdYrINWS8fe+x4IGnPRXrdrko0h6fzWIrgQ+etsZoh
pDFrTnmbvywy3ZTNeSioe9yKwHDYvw+k+R21zYleHrMhlyl975wV2Ml+E43siRZ0
OwwByenv4HP9evSpKUIb314cnBIzu+xdQg0ITFcfkCEoPoqkw+pXoLQPxHV3K16r
p1ekkQzQeT8LSuYXwDEazZyO2J78nCbpeQtR/kVg4vNyj1evITPvll2pWnRvVENE
7kTgn0Jk7IVLFLOUQ9mLQvH5qZhQSRdgRLomWFYdhOuXFgstVWOWw1RMtcniUF3c
PcvwY2HaAARTkv/5caIw/5szc1ke7wbXbaNeEAHZN4aTi07m9fltG5S9jO/8EbyN
vmOgcRf8gICBx7omJfbCzZjx7DOiltWE8apqFsXUT0yfVfD4j1gWosQIeKmtdSyf
LDB4T1ZJBuQwjodzYEMg+OXdtJCf8M8iANBrpDlx4UfVZkv+3ZVBqlJ8SVtyPEwU
AK2geVSX/DV+z63Ou1ihAIWQRqC075te1288QsIHxSb3q3lRBo/KZKJUAjEPU6me
p3KZSnxnU/8pAySLrgu5FwhV04ckSqzhs32qTCBnoyRH63fDQE/SEyb9P1MvPemT
DMQYExj5K2Kyq8SETE4E1RZyHC+8wctdPEE80PMnTo/fMCcuP1UDEepg8bzBmFYQ
e1UkFeQxoaHrqMSfAXlRSmIdz8sKdAoF4sOsCZdlkSZmcJPR1jaD8UEGOS8IewLm
zmsKNe9EI11VsnFeieqJfQG5JSsOlLxC6tcAFQxRkf/Q+Jrfw0kDHZ9Wbx8uO+y4
fU7xR/X0d2ROcXTuFawjmUq6pbGyAaP4njDKwFqy+YQseK+/27w3t+EdwZmvAcTM
rYok04B6UaSOaqkh0WXYwY3lCw37hFfYzV6qJ/n4bt4bGpULOyj23V4DKLeDrRwM
fRmDyDp+z/X/85HCoSOVFqPZWjvwFtglSBPlIXHDRnNsPVbv9zMnTcMTtKaZxeu7
qcd/BQb9FQhLAqEwzalwM2UEom6eRuSi6GxRSYgXGwgnQsvEzCTN1H4ww+a3/XhJ
RrutwG++sZczit9Khs+2VIbsISuSh9iEmUI+0c2APpRmp4V4s5MZ9OcXFFtYAuhk
vGe6Hc3qT/rLsmpey4V+K1QdhYvHW8AY+yYl3UPWNP7N8ysZii/wT5uHMsT76kr2
ovzM+yUR5x6r7TuB8HoaZKsJEIIVLkQrcqNQ/wWOBZBRt0nQu4CzLBnXabqEf+Zu
iLeA/4mbrcjoRULSEGBtG3NHvbmjxtHujfMsbg9pfCdqwKFWT0sbH8sjpOzUMfkE
n7n2WDtjd6vdAeeBJvLbnu0UjsmKZYJ3PEwzdI5a4t6fP/iZekfhpfB2WkeT9Ut7
F68dVJp4ZtLcrKj2Sq4JXVz3HtedB+N3pXaso/2Rn0BOkRjr9qO4jFVcJZ2DcrwM
FkUiZAgPrfkLzvhzpK/FJF26Zf38ghWMsKVF+DWAUWS+3lla4+xyQ4VV0vgPrNeQ
Jv28zacD9Y9nQv4MHf4Tfy7vWfE44C1ROatxXKuDErtEi8EUgTVg4Suvi37TZkie
SZQEAPF8YGDrjohzWMJJOhaT+X/dQyGV+Zwtmt4r3Ll89QGUpMfIlySb2zuN1A8x
4zG2zC5C2XHbJdaZFrcwr4UsYnQ4xrEhO5uuLq200tzcWUS4n+Yd3V6VLDX3jbZG
e5whU4gFAczoKXUgjM50kXk6OacUychIvaVqk66hqvXAKvA3aPWr1M34PItDOUiN
cdjvtXsSRKPZiMr6F6ac/0MC0U4SJOZfGEYjvRSRN41Xy0MZNgGnKtf4Yh5Y986C
3ADwebFv1P0BUI1+JI2Fcr4SBgb6PLbhFV+Jkap64xmKzeIcT9MEHczNtHwMLt/2
ESIP2lxZDzPhZCblaYeV0jnepttPWtlmugBbu76pj4w5HDIOUwimpOy5Egx8oE3A
NvRhgOeGWYRR23IVI8R+GI17QlkFOOy40qT8nZ4nOv5ujzLzaL4rIeCP4lr0DMcJ
zl0b1TcvXdIVtbwE7OsPMoy3V7bW0XrenIhbOt+oenM+bv3lGxmgif+vSV8cwrOJ
bEp2wfk25OZaTCNbjYBqDs282oDHFPrnKUlYX23gPuppAA+PKVxI1xGxOgDkOYSA
EZVNbniNDpSyH25G8/9w5DuEW4+3zLU3ZHMiQAG1PSo8bUT8mo6vgrWaNXNzO8xW
mlzA0CImwxyih1wWZuzLTDeoSdbZ/FmoWQv9/VFssIUvVID5ErpEVvAP2Cv4KpCF
xc0hiBuusn4BoNg+GuJDnX/Pvu1CnWrSF1Q1D/AiCk5z2esFkq14q4iljvJe3AAC
izf/Vh6Z3+sODvsizheXsDa78K781gcoP3kOT//q+lb7Ih61Vlku7/6ZxPZUOFwN
95nCmM001ZoxbsivXcPp2v0v1/AW/IpzRjgKi9isegcBitYYZOmMWNzieX4ihGiF
BXro+MVP/pKujn1mayL2emx31shMCHmbTX5OGYMV/iQwZolpARKqb6uiNHTCmPNi
cnWOHc9Tk2mY4NlpEBthr63nePux41omE7D45FW7gbJqw+8CA/3QY9D6CbIkbNPW
7tfE2A1bh7tMQ2Mn3By2jD9VP10YcuN/1Hc3kLujYLckgp6EVgTRtSA+1pPXqlE5
XX//6gkZBJZuSJOPGJtpDO5J3AigPW6phCdm6tlRhAUB9vaW0sStUFFFWuzpjlxe
caGyiSkyeB2aqP50/mb7KC6QThua5TLewdVyL9qb5lFmsE7jZCzCKhgHnGxUCW+3
bUIVoBZrIaXF+Rx56MwwEl/ZN+YoA/jsNSZWLnEMF2H2QCFRAd72gd21UI3c5NDd
G3/wh/2o5bk7QcsTaHKp1NzJ6eofEhxbYdntPQjWkktwSkZWNtksyMC572QmR9zL
28EomvD9DGiiCQtbEuz4jhcAu08FOnbP1OE880uL1jQ0PylHxGKJm7v6aN07MNox
DGMoARHEhgkS8s9N++gzKrJk2QgeWlM5Rlq+J0wTn/AiLp7ueez35M/8x3ih6pxv
xTYe1RT1rLHPr0CufMegivuY/yDvWBmPCwnM12M2b7eE12TTbMhkdHnsuBJaoTjx
/8an77NB/UHehZmeGL/AuRmMr234Cc3CuAefCId0grmTJERZAfwjqJ7ooL8mUrSw
g1KJUooWWIu3qaAB+Ry6ys7Ocm9uRm6VRJU0teJTaMtpMZxJ4EwO4Z7pG7DjP6k7
IFUju5YelsO7Dhx6sdehXHAYViJAfIldUQp0TvxhesJBLlbHGVDRcLWPHuqBizZ4
l7ggQEBMqkXNWSGzuVRY0XnRGC/imxTEVfJAYHSNi2B8mmYePrcyomXNw/8bUMw4
BTa2XldUpizeoZYC/kBDmcUm6rwDGau2CoDHPUML0XmrCevahGi5zd6vbDhNODkP
C/yykTArasXXEvbtvJSzSdZf9WzwESVOi2G5OVnoj8t2NG3PXbsTiF1C34YfTIkI
gkYUe8grJIT3nD3tWPfk8o7kOUANuxX8z3e8gVEvLr6zA5WZ6LKmd6FkSCMlsQzV
u071uvCqBGP3gNKmnGzqnSvxDPGb8Kk6qKzhmYbuFIdnHAGfcEpb7h65LFxFAduy
2m2V3mWAFbMsL8g6S9exYBusqLeJKvn9T5G59Y+Lu5mJ+AP5VVjIAGyngd8fDtZs
+Xql9SoY6Zk5DgbvLRKnmhQWn39D3mSlExVG/4yh4Vp2ErBlg1h8MDDqorHDTjys
RjnkjKMBYCSG7Yrplo6DKafhnF3rJOiprU/AExRb1USv+BNlLxJXKVTznq86NgpT
YI/xsZZDjVUyCD6MOl7vBaQYQ95LzYD2C4k660kY67+Oru8dBzpBhKgQRkZUYMPj
h0Rx/cFYtRByUoxKPejNUM2obE0J4FKUhgKWUr4O0/XNtuhoC38O18AQ6aabClVJ
39JoXJ0XCq/2rKgvSdJhB4Cg2iYgKIf1/A0C6JwxFvnyfovGmR/ARRwLukoEhqOH
maJoDpZAbT0WZWHwb8awmv8jUtcdeQRZ33jxJTLJU+T5ZtqDl6YbkP+EX4a+lYdE
VJEAVuT+ofANe/JO2onW8s78bv1iT1SpJh1SrXjxKH3lfOx1/1JAE0UIFP2JZYPK
9q3OTHoHS8cW5BTItU+FxTzmJnBsYuuFtWeyf4WfzskE4IhCkMd0MaOMt6fz8/xm
VfQ1fx3GSD+rKsmmd0FzKG1Ru9GmTh/QXVr2DU+M1T9ON38uLrnopUVDbAQCjVtX
DtFxCEhb+L/i9SNlZZhkLeX6zwbpCzr4TVMUHRoTqSSvaFbcmr+gRyNjN7eQQV5o
iqL99wGKkzOPSaYTuD8sXfgD6IdG+46GTZyyHjZUxHHVfktEgpGv+esy2CHC1Twd
ystzYyX21qCCN7XlBbA6dL94ZmEqZkKYrx3cBv4Jrh4fGSi+LSB6znHzpuHiWY+4
mHmA+WPJoV0/3uYHvOtF0TbQoMX/cJyzpkDIaQq72E31eUs8ZigkMHlj0v0RJmhi
NJLDkTKP1LDZSngE8rUr62qv/arGNiv/OdDX9p8MF5V6uMD/qrneXf7Y6VElXmFt
5EQ8FFZpLEJpPGSZXlC3GOYDxE1XuTruShELCFGCGfgE2FfRLM5kTyfTOGLd4VI2
gbQm4FCx++MOVDi23lyjXKyrf37TCdEybwFlUNjZwvCZA59wYqvL/Wm/ycna7fLK
Vmfr2E5R6iI5jVk5epb+aQm1ADKqjlUFzFfA3GsWG80zv2FUavk5ZEnJ3xtiq70C
X21wU2Tqy1Hw+FoerHTqFEUPVnFVUkkktDulAwMDnkzK+kxbZU5m2pHnoXW3YesW
cdVmUnEcN9pHsgAF5UsFGmgmneZLvD+E5xCvIQlH/Cml74r9i9dF+LelXMuhVxGq
cn8YMzOP8AlrCFMeIMC7bpyXlq5Sz2AePqx7cTcrYIJAA1ns9WoayU/HjY4+78Ju
U0O9AogbhSulrTMX4ZlrAgBdNoV8rSj7t7qSZljTTYdhGecs60+/Cv9mDX+oNa6r
j05SBbA83YYZ3fP/aSDa63f7QLf1C5lGl2FqyPBscn6WUb+rk1851gJuAzca3QUi
8dnqIgBb4/v/riOEAaAxRHsNKdalBkiJit40BiR0kKYX6Rkusg/d+CN9/kGiavL2
71weTqFOmkU+u51ojhpXzbiGiKgbojBuYXZe5R0n0TazDOisFOtSGiSqFSeYVu0A
lzOKGJzyOPgqi2S5qPX7kfwN3SYBrPcvrKmZkIn9JOz0ZokgHPTrea7aJuDkkjF0
XvX3uDhvBF2QF8Y66T+632apg+jKJs0PCEItFOMsYBnvENWMSU7MkUnOIto+dfSF
sP0I2PueV2/AI8yN+L0BFC0F3pUGcnrifc7lAZ6zkNkseKX6LTNXA0yCJwGzvOye
GcBMaM3FRrKb4sgLPyT7uAh2l3UVsaLuOdiNKxh0EpvZxM+3fwR8S19gD8pV/xOb
LOErjZF3rTPWqElUoEgWGA7vex0QTOcEjRa20SSRt94/hvVNa/yM2trYVcJPI8Qq
iNbgKRqC4T1p5j990FLcnEwE7jb8jcCcHZZ4UEE+VkCwp+EYwbGnBZ17qnuasM8g
Wh8LPiS3NzWGBKiYplAnRKBG/7SG9LuIMJybEZkkYeweeSYXfS+KUQ5uBe15PMNV
C7OAOMA2ZFnfww5gLgkEkI5JmUUCICa4hQI3IAtRY+lsEYvqSB5XHIaxbUT3rW3N
w1wRjHTmWjCGwBhSM62kfmjYmbzgztEKjPzfQU7Rey6o7WGZH+mgmlZNGjxHd4cO
c4D6GXuwL2J7GcXkJVwcmZLc1PH4VYBccoyWR4ChitOIARhKQDDrhOmbHRKkGMaJ
BzxtvHaSwrl4XMsTofitylhgwJZhNJWOH6Upa4Wz1JTJv6gi56QUUYsbLCYJ5IcF
7rhEyfRx1wcqZrEU/DAR+L1mkVlJVcg29XJIIlIto4SFcXUVjtQFDygrIRvJMGwQ
ZyA7FDfu4reRrj2EHAulvmI6WkpmP1aMnEC6XPLoC9s1ihKDxiCPUvj2nuZ25J3g
ntQ1Brb7UHGWGPfPdOkZ6VtFaoLeGfplHWHFNmjqNpI1cVi/kBuItK1ZvoUpJeKO
HWVSS4DsaBh1SI0skbRWEKd+UGmC8/pKSGCfiDbV3X/gCvndLOW5hRyPRQaNE2kw
leAqdVZfHb//7c/kenBHwAMGm6iCTfvjb1iUaAanmLELcmZH7YYwMVuSNXep3pUE
MH861yVCgPXlr12bP0A1RmWxYMHbvsy8mF0Kkeur0Vx6NEgs/JTxEVj3FszjnTUs
gpLhbkBQBQS0fPYdJYDBxfmkrzeqjY+3KkyZM9CBFUsbykBtVyQusAGX6A/CGYSK
/gc3pdRySsKkTguzX3tkBoYWQLBOB6Pu0uqw6qOqjoYpodZ3Q82h6BW1Z6PL8B7J
6aaNvCEUyGZzVAExJtBk9MY+sj8vFz8uCAJ5noixn5ftQ9ZLyRHOx1wqbXasc1Nd
U1IDz5NoJPfEalQRMM6gWPQEOt6/Ruf6RspX50vn0AVntc38anuLSeE/Z3XxHCCU
I1M1HCwe4fvBh3ZfbiBVFlk/dM3q3oZhozk3fWOBj6MLePhHft/NCnjDCRhV+PMB
QGwAaC0NDYxcFtjwZH7VRLk4O8TZITUUhhWzwZyPy7TZ7aclw9q+C9BAtNaRJo76
jb/ZMULLlUtZCa9gJ4Le1RN4oqUSg5h/boTy6o1I77X8c9+2ukpilMAGaMlc8YTN
DFotIR/QJUtO2c/TyGsH8Vsf4ZyTHJNcnqWLJDmU3S8yq3esok4SiBas0nj4xwhg
h5q+gceSRjw+dZeTcXlMAQ4AIQm+E6mfIRi90DYbuxkIsB8klAj/rOb7P5ONV8SU
S+JdN6yJqyKj+93cBylksAMyb1H0lIFuMUumX/5R5xVqfJmSL7sREBDWz91TD9A/
75ptcsyNpRvTI7kB7BzTBH5h2BqRku0in78I8tmNfj5+NM4eamONbRim916MzpEh
0YCz8Xa0tpS3UJDFfQjOF6pAtUJbBUTEtC6OhZ2LO85N/IoVhbUsGzXmXES/Emy0
pn9XXZ+YyHZAYICs4hQU6VDpvFMs0WpG5B5BYOj38/lwG6cURJUlVzMgNy0MS47w
kvtfT4GnM4QdHrr7pI4sHyj/SWau7VMuLe4ukWbQLXqT2P6/99lnb4zQfPMFWrWU
wxvy+O5pCFAGaE+TxfaMynu6828R1FMTpcewddU29mXH5437hKH+Ry6aJB93zl23
TiGQSnhkhw/mrM9JSJ29ul7bqOEOTyj69kUTreDOYqmL7Z2cxfCEmYhmtSQvhvts
JmMBTEJik6cZFYC7oNaNqI8eeGmQBl2HyQ6jBBo9PBnHv+yUv3OCI5kVtmRpsHi3
cm4RSkm9M5h/WKQhn45iAbU+CLBJv3J7u7c9k330PX9UyUz+biV+0PYq7nZYzuO2
3dO2Tb6blMULbCZ4WlPMILnKaAQeYRkioLzUA5lna1NRkAymec9cAW73zTEV9h6R
JVN8VxxSYwL0UZWTbMw+PY/qC5xGdazBpf9Ci9g3u+fYUaN7zu7jG/NZKrooJVlD
BWrYT1lsWsxMrf6GLoXQX+k/C07JwkzZ8paHk0wuWTwR5degWm6ralaUkQiLtN2n
K8G8d2h5umS+dWTR0OD6JfpU+cD0txnfFGzuM/vqY6V5OrqsCboZzlwwYEVxlK3A
S712ih4vK4PL4oAZM70T8ljbHzQyLYnUrpbgOrKbF9XNCQ+UsttIOVJ6CNBhG4QP
CywFz7nY8uv1d2nZiladBJ/KK90MinN/bG5hz24jWAYMobAay90l6UidzYUUoxyL
s/PmOihhj5B7Grxi8bzgT4vqnHv4VrIvdsFlcSaqBzGn43mFZ00RKJVzXw9nU6VY
jwR1AS9TTsfM2NuPeoE0EeLGElApWtmyBWLFbJK5flc2yKo7Uj3Frk49iGh4oGvr
8YAuE7mDF28/GmvSP737wJRcHg8vXXVqinzzM0jaee1/l7ONnnHqiyulflh/2xie
L9YKPdl6Y65V/GI7SbK/ytIosJEJ3oVd96O9Zv3JPylg8iBeb03aFNRYX6P1uRVD
j/dTupo06UGBTSuXUMnAA8Drjq+zwKYz/Lld3rXKt6cbolXca+FuuiYNJxvkmH3k
OeRW5NA6X7lwcCnsMk6nCWm8m5Xcj/wkX3FFClejym5uCoKpPBw97qUAVT8251Zc
LLYHqgSAjfNgrxTNF6kJtC+mNNZ60eufRvS0Ni65fpdScCG63orPUtlKGPHA6uEG
0g/tjSMhPsuHWJ/cBaZP98IIX9tH5BCtGsfVfN2biaI+lX3Ms48X9fjDBERn2aqm
ZblwgDGC9SjOhpATIfRO5P0YRgEte0EA9y1HKNj5DX9K+8kDpzKq4Ro8MIjdu5Eh
LBQaqE0YBazbX8g2d0JEOPFvnBCFYjx5uhbpai+r+2SV5vNaj9D/vW5z1cCtE+k2
vuUzfVw67t6WN2r1EQBD/7x5Su5m0M1tozmm3n/mU47D+GyjjGRmPtKBdlrJgn+9
N6GhCvfrVDFxf5rbAYMuccWeheux/h557Sp94CLo+Aowo+wtQTp2nApjOcdUGTyS
K1QIJyBxEjjd1xc9Vy4Xk6w56DSSyq4HzdJNivC8WDCQnT8komluYsqY05ySVZuP
DTaBGA3x/YqLx6Kp74osBpC57f3Y8k6mOma1Jx8Z8Y4blLvvVpYM3/p3sDqmk53r
77bvBs5//fs2Yyc5sO6BzJT9CMeL7lpvSb2tD9lOvcNK9qYn+oAu7V87USq7bH75
apkI12l/GUJYXnnjS2Rhw0qKteIhDJlN4KdBWcUv1zg7s0dSYcyRRyTbGER6oQ0B
L1AxvIg0JVxuE2E5kWTHPu2Z8kXRhoVZss7GZJohbhAqXWffE5p2u3dRQqOanFo1
xcG4H/5bfVj+R0joU9kOIWHbCmoFr7FDG5qj5VluoorlfTPNyDaSZQhHrjjkkqqs
OU8Ao4N0gzt3oT4YzmHe+cvRAk2PzRvBA5qH9nbpXeh2HnPCyQmnPoSKlFIyoyU2
1qyff92c7RQVzINzbnTOjgjgM/ExZyljtPAICLdIjg5CcIn9hLbK/QwOredjAcyF
/2Lzfqd90tlhe7cpNi7IVuJOPnBg6OLVGLc7p0caDxU+WUZ30AWo5VI8jrPKeBMu
f8yiXoOKPoCQJmJfQf+VQPtjAvyvb0+tzq5/2MNArYtIbmpoVyBTx0hRyCv4IdFi
CrmpLJvKDs4G2St/HspFP04wenEYEtT/dxiUzRYQ1oUe5dSgkaV8U7FzkYASmOsz
Ei8OZ7kaSilX6+/aMc+YTDyG438iXSoN/hehYx0/b9mZ6xBcYmdlOSGY00hc2nvF
KD1pOBTTNdiJ1LyknkL2jEt3W9ngEuCb5IFLG+NiJY+3q1h3X69x5rI8wO5F06Gk
KHHofGRc0b0Y9kvS1RtZByyAWsEjlhFBUF/J/0NHKn6BOenOsTyw0Qfi+P9cpbTu
bw5UjnfOkYF/5zPSn6AtPUWL0nMZ6ec14H1bSUUPqM6SEayVZxUnKey/AYJtrenw
wZSa5S/Of1cIiUQzRsduI685/HnY0PxYvHaHZnwidNXJyF3qnNWfuvoBDc2dYRnE
xQ/VcY2DPaIjpThvaLAM4+eOhB4RR2XewwKnVFsiLKxOvkeLvnfuVTGJswN2ZpBz
j0YT5GaeCJYCUsRtsNT5eyh/CFgBlg9Ha1MLho2+pGgtjABmt2qNpwKJ2Hx5orSa
o/L3qexqdLDAHfEjCGY28u31U4cSRmEkiKLNKPK5qfQTHGc71fLYagQWDOiwYaIQ
0WQE1f3oAWBE+iNSIhYjg/Ng98SjuZI8IftzH8tEInUKXzGGz9cceLwxRL4hJX95
m8mllht2JXoL/UXWGv4xGtPsSQonxPV+IBo8HUcrnlZW/QVLdPNGuPPuycJdzMFF
GfOlNdZbK63Suj00yhGteDpepHpPPmO1WjBJsC3KlWQrrPo4tO9Pkd4PexrvqBew
1uKgvhUDIT06vXKDldqPE6THALrWD9xGBEpHBVvCbwSIIHsWWXvzHXGAfMTCAnel
RdtML2CLlVoQ/v+W9W7lTtzsX2PjwzqPm8KX7kggpkL5ZxMjAgAjvZ9BP7kCwSbf
OJtc4cD/fb2YzGRdVduuYXXm4mUR0KYBT9khRy6aPh+Vl5X3nGtMGY09Yn7z/3m+
HUy/s5B35Dls+2FYhZOgOBEbQSuE5z3iOEdEXMspnIaWLK+u9amJmMMPQzs2xzFt
DVsw7vK8/pS98OJx6Spi3e1tkdv2uGjrrcWoP/1hd4Na/JyjSLDtGXkHxZdOl60O
9RqM21j+AFsvIdVTgcRk6YvrPPS3eTtbNjwOGFyfxK3F0XhcrrHFvo1FQZG8Ong9
1cfJokpZ3xcgk1aaB2ZC1SQueldEhBsmlxuXyej2UoGjtYAZzTmdfy4xmbEPaAuH
lZxp+txdfdLf36qyQY5tz6z5oClCbcC8N+Jx68SqI2iNHDJhpcKXnJeQ5oEWKGVZ
aCRaZoMalJYP1w3zY3zXlvMzlGdAmzcciMDFwGKLP49ffJAo5OfRMAJVTVtDPkxl
pRWPs+kR14Fe/9AJ3hZgsDSw4PT7xHECXOQ3Cgb2kABKSzbA+V/RA5WTAHMbf+pL
ftLe4S3lGJnvVWQeXWck5lmi40px0VgjHwm4Oc73C8Pwhev0vfZg0YCSlcxRTScp
c6jti0uqcJfE2Z3tfn9oAn+oh15/xn6bWmZCR/uxf3iYp6wdcaRnOf0mRTU5Gjbp
Trjbj4q09E4VudPv5+ueSRErpeBez/avcSXjNdCV1EV+P6ZiSWjO7IW+6HUt1BTR
5T8tINpYJpsoSk6y4YBf2ysKtzAZ0C+hbrkG3t/WCmB801hSDiFZtd2oBHlRxENy
f4+T2URAg8DuFwyHozdT2tUWEirkGvYHkCT9IOW6iLlk3keLX8ZAB5xV8TtdJeTn
4ocq0ZlcxEVpjHUiJlcudRV4BWpEuxeU5TI237bmM4wmXRzKQKFSOY1RVApb+qCl
7JVX0TwEEdOsfL6B2IcdRf7c2H6K1jkZTYXO7NK71mlv1yjwmCk+N9v6IU/Zcf5i
8D9cuHscxxuol6Hw1dVbx2VKi9cExrP9050eMpDIgtJfVA2Fc5D71lJX5HAA1QIn
9jTHqQ1oZfS9SX2T78+QXecYnvsqs3k+WI7B49LIlqKYQEei84WsJjYkfeevuMT/
vMqf+dzQLneFGWS1IwO7m8eQaX8AxGo9Y56b4NhQ/rRtHrCsJZr2KCUgPYWGcKUc
EShjKltHpYyBqpOzEY35UY0GV46yYR3zGYGZzdGZOs0sInKaW899ADhccBWRcisl
Zdpz7rYtvo6MZiJYK1g0yyl9IoitOh46hO+qfPN5bl3rCXVuvr6MALrHiwWyYcI5
hpZ0VPavUp8zpouupDOaEpjHFqHT6flFpBirpMN90tw5U6BJUt7mYLdkb3qQPJfD
hamM04oCzokP/NpRkIx0gWX6s1wcyW2WUo48TO9mbrrdJzCAbryeiKV11s6T5FSd
BKHxHTJUPGd02czOYHz6YDzGvuJjjUGRlVOhXSrCRHjd9DnQtqd/5o06aQA07lkE
NDntuyFOFOF18c0f1rCDQ5odf321majrVQsa+TZkfAYpg4OtKJ+joJSzZbTVnL1G
7lv5JXG7oxS9LPMDRotfsHRGQcjoCCaw4UOzIc9anMxp8aj0Q7jJFU7Z6OFPyOx9
9+zJMW3VtF0Vasg2u335GO/eCEp8Y2othjD5+wcg2mcvhCutUVUGSJ5aEnA8p4W1
PApgZWiOyyzHLZ0Ia+fqq2kqdi6klyZHGpDMYqKPPF4YLicTQtK1ag9HVSt5a4YY
KzcbVgK3Sk+d7ZvR6hisvmqzalhmRmdlDT0Hjte3SysKrbuqSLHbgp5CrpqpONOC
Ru5ByvxXcXA5NGtFsGbCvjPcokfKLvMVKedGRT6MSfjA69uUJZpc6OKWGmqa1i2n
pZkPwH39N4ZHRhWiuHD/Vs0siYgjLnodXaOLevdwALgdAsKSuOU0dBehkZHStYb4
ddI2XhsgnzRf0ZzALTsv4ByhT+WJKMulD5/egNEFOLqf3+daVQ+j59d4yiO0neIT
zyOj2m8db8e35o7Rf28EYA7jlJ4xBRz6hAT9JSrdM8KSNOoR3gDcjAVTLMbURMJt
PeHV2VKM5rSuRd2EJ97mGAqGGS3WYvzqVFKvsqcd2JJt5PK86AvLPR95GhQuPggc
ucZkP0+eKhP6mEl3IWRbTsbdB8yi0sA5SfEkaPaI7fxUZiHuZ0PVSuAnPTICB9AD
ZJG9hYW5+mGJojt53p4388SjqqEGLKfpSItAOj75ISPGzlavnfWffEzazf6jRTWa
Y0BAjoJ1DY++edrv4aKRfg1VF94e8Cd2ut3ZNO+oLGebLTXobvxsvbmZr3zqMg4S
Ux0rE6TfdgCBXaxA/FJt9/SA9gnJeO076DWx2VJxG2MPbXcMQv+Ik6lIi+6c3x9C
Tc1enEVIOBb6A2MBGxtwoVUDDXCgZuULgYqq4d3gFkkps6iBv+oeKwh7f0ByvFGu
abU+oDGPAqmaIdmQSlZeJM4gwD8HkOJQ9hC+2EEWTssgloBysHFRZTCSyKB9t9Q5
yEMAhjU7Fr+qwEO/U9KulmES6yKNpMKuZSjmAkrHPcMPaWedL++AT0W1WoFKx5TB
j1iS6wGYNUrfFRXV5serk6niRid0WrBB3UQGguQgK24OhjpUsN3ch09xhUurBJer
wW2A8/So2szeb6IgjnuQj/P4D9iHODCrBqqGWTbWQiKFj3V2nIm8FwdMf/m/RZ8o
10wg+wpQpv8HZ9NDxFvr/bPtKj6WGXjgTqn3gYUMdO6uwYLs93KcZSa4MQXBWjAa
GS5IIYwXW/DuGXHv+evxtSmOoVrq0cCmp4Tgn0EukY5WY4vWoRYfekzftu2W60fA
Whbd60d9UCwvfXVUSGNU3A8U3ylyJ/ZZVIGA//ydJh64Rxjp/Xp2MgDP5jL4rR+C
OcAA+Cc/0NP8DBl5JkYUE+KqjBouaNx9SeVhpwY0A+WcP3jQPCcYzo7YldvI/d0X
Uxk25fe7a3InXyc0PcRxB5Z4CnRzFr5KNAc99qjFX0kEy/lYRlbVbbdAcoAKWSzE
Odjlok0nyWE2heSyRn3sr9XKolsOx9cu/CTTEp4L7AodhIRypTNDGHydTXBMHZZ4
Hjf5E/wxst6eDzaCa4CEOBZtMhC3t1IY55zhYctCdPbCfJ0T+AFzpp7xrd7UUuwW
wg+evLf1oMdNF4QIh9vVxYFTh1d/zZ+7pidQmJTg8qUISkF/RVzhvBB9anBUUUU8
JkNGtveYEYs4WfEaZT0m618PBWaBw+oADhNfoZGzSOFPbI4zcURHwUF6n8Ji8LmK
CcTjuVOaPwT2YNkNA5AgkgzOvXaD6+jZGwX16rm1KqUlX3BmqnKMHvoxO9PoAnuB
3liHpCTG2TyqEkN5A5YPL2DcBgfVOive++Hc6afDL8bqWEOWYUrQ+oOwE6CrjSBL
X38ZShBtXltgU8BvZg5zkvUqGzApUeWsmjzbrThQqwjahTJ7nlSz5+L0nfk/LYtH
EoZICynb5nDjnvjpHEjm6LdQOJ6xMV1iUoeeExk62+SaKPCcx/E49efTaem1hMVM
97e/0xcnZijw1n/uZOkExkDVj8a/WGgDoJBHW4Wmg9nojC8X712Ta30Lxm0XgJ6j
JrHkPmI0ut1/FbSc828q1I6R6+4dk87nO7A33r9m8ISUn492/oaI+AH2UvirrmMp
OqwU2SwFFWUkauq83ClqK5BUBC2TW88z5pBpaxZZositKjEk0xZaQQz+32OkMKVV
2bFnxq/m7m/MTluKUtXQvo3sYT3F12TlB7PMNKWgA5MOXzkSqUy2Ei4qMV2Xfqhr
/XlRJ6QdnuImEptYZ5fOaVDOE7Hgzlow3F+BvnpK7guroRMynDu6DqjkQTz7Lk/I
3rMvx99Mduuz7SNer1pIdSq4ImEBqJRTTg9skvkTKQcQURrkHw7AudfpoA7F7lsV
WgACGRmIehmZNuEXupXU7rcahEQuPXQ49nSDOgXQgIZx/ZBvVhp6zXBRaq63yIn0
oM+Va92zJFJ+dhnRqaXAxJjbQ2tJapfknoivr2k9h+dzGDsCV0pfz25/4K0Wr1is
ZYdY+q/o1Ny2uR1S6s2k0tqWh6oMDz5ltny6t/Ai/gtZBT8rTymbkb+v6Z52MSoD
z57mnUarhh1lNHJf8b+OkL8w33t2fSqBE6WLzKy/ad1ebQ5GjM6J4o+zrJ4eO74H
wbvBny51H9Gypcgyoy1zuIqaji7sZqqc7aln/ten9ewNQMR/AWVK1kDaP2H2Wh48
4en9zNPSBy/wlsO8bu7dgI7fj4QX/DB3G8FAL5Z8hGvHzdk6hcq2GIO5qizzR5sw
fxla/zH/0P0bOcvPlk3NatJvNyRjBX8r4dyvjy5SkM9UJAAuDowGoLZV5/4V8rGn
1pqjvHAtBzcdYpvs6wtyOko0h6poilMI11Z76XHDyb3UM8hh36r0w9eEcYQtI9Qg
7vHBbOFEehhd/veuPZlfReeSUP57PpZDYShu8USjY2rePnnJa6JF2CJr36KfFbcZ
54bzRhlBoYgBQrkVl9ACTzVjiTYCArmBkQNi36eSL5raQQpfv8tKaJhr2IkGtzK0
uEj4eD/uh0GCRSyBxDrRYqwN18uGPtbAZaugFMr94TfcLRLDpUSYV0cbFRgzybHC
dwJRuRysSIW4uAEBJR/be3xe34Ab8XM76jX6uAtVUJ/HSFutPGLx4AUlX8kLESNj
EyhW0gEWxq5m4cFXIG/ISbRIo8JNdawinZV/7sS4GKHHcNSy5KGmHZgi5FEauZo7
qqUaq2aZBCVhmB59c/taCRPwzyCxVNMphCbCBE0UNGmYkra/ukQBxCaafh/XW25M
RTVKai3HhgIKiRyC9kTsQnGbELheINNbXcBKhzvfYazhy8SxNeqOZPhBR5xSohAK
l0NfIscGjlIpLTTfxve43y+dB6ZncI2tUd+fz0okbSWbdHf3JR4K08yXY6MFwpw3
v69TqqqQeJRKwULjGfI/q6hDoc+n7cJtaAfcnL2tH0dvNsLtbzV3tcUrIv04xueF
quTx/PsUHnJWzx4ww+sEpA==
`pragma protect end_protected
