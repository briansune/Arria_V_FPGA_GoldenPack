��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t���g�l���)�eO �v�q��#g�ƵqOl��T����D���f��=i&��+ˬ���sz�M�l���y;���^�W4t$'�T�h2ʀ�[J�Ь�\�����Z�]��O�K�E�9���W�P��3*�-���)-F ����7&z�e��)J����vZ<���|v�:��'��.��ޔ�Ѹ���KL��JD�j�+�$	�3�7�@����^0�|�^�)�+ˈ=J� �W1��b�+�X�-����!�c�N���x>���whse6���{�e��:q����N>�u+� ���=����wyە�՝���V�� z�X^BT�x�Q)r�Z=C��C�A k54�Jd���	�����;{�P��*R��7]I��'��O��S/?�l��!��zs*�����N��<A���|�n�b�5v���7�U��!�E3x�~����j:ؒ�U��S��{(�z�O�/xb�h�pP�&ⴔDT��Q.\Z���!�v�
`>p��8s4�jX�z|+�+� �ӌ��p16�ln!���F�'�(��v/���9�bqp��m���K���ǕHN�FU]�tr���u~w��yuEM�� �z�pjK>�]3:`xk��h<����������klra��Y_�.�Wyd9 ��.��>��b��Kqg����j���В'd|��ʗ���湧�E�b*а�����.	�#y�[.v���1�ǫ�ֳX�q�|$4�#���{ǹ*?C*�ԥ\��$>xҐNa��� M��}pyl�^`%wM��酙���>���x�gR�!����r�88��2Սs�׸�3�ʚʅ�z-A$�464Gð,�6�%I[&���r ��\��T�ؗY�4�"�g�t"���o�<hO�}�+���Q�V�F$�v�����f\����U��g��f�Z�S���s�G./pO�,M�-����f���@
Fe�%�� ���YM��$�~ �@_�'�S��f��o<��aX��R��Z���u���aH�8c �x%�����h�N��$���FX�  �fo��'��͒}Yh�����q�
1:՛�uN��4.6\��$�}R�RG�B�T{�C��Eu%
��nS7}r�>b���_ �8���m�%�aUM�%�ܽ�5�@GG~������R,!@��
��Js�"I�{~�Q����o$5�;M�io@r1f���g#�����K�sW�������kXC�o�6!�rBL�2��3������$nJ�J����yw���$���)���ᄝ)���ңFX[��בZ�_���*X�{A�d<.���<���.ԁ>	�`�e��jy���	�#�F���o�$�@�d�9�a�y7�J�/����V/��8֔џ�)[D�����@�U H�{�������\���)�湸\��j��(S�����v��D+�R}�x������ %b�"�{����e�����@�4u��>��[e70B�J��Do���/�lQA��%��&��ǧ����P�D����$��
��m�\�׹
z�z�ؐ�?��/b<�N�
i����J�	c�KF��>�MG�i@/��u0�q��v��ؖ�C)���w��Z��T+C%^��؋�M��H�u@+��rW���TcI{�CH@�Gkh&m��F�U=�t	�ł��;v�X�%����)�}S�E����ݏ�vY$��s[i/���G����R�C~����'��%����A��B��ntn~q�!He9�2�����sG����@HZִF� 4���O+_���u$(�zd腲�jj*
��*����{Y�"Ǩ��y���)H-�39q���GL�'�������/�K'!��){n4��0��K;qP�B�A�E��a��q�� 9h�]���[$����<ݳ�%�
X�EB��_��R�O -��N�6����s���6)�Z�����h#{	�il�]~�|ŝ�H�}����[!<��������m�<@�1�]�,m�?6C�
tq(�/иSIh{kvw^����{,��PPq�<��L!9z�١�^�EVTY�|A U�2ˣ0�vny���<NV��";O'�l�"�Fr�\�S��|$c�e5��Eٖ�Au�d�.[qK�!�Hr��p!�9g�,74��Y������Yܭ@��i�UQ��w8W����~s��>�Ф$~�\�𛺗0�	D���v�{�E\M���~���Z���������A].]�5�-BM��Gxe��]����N`�O����Hd�V�q�0���()%�s�-;`ra�����oI*l�g|ю�So�%A�*�X��L��1mW���jT?���t���!x;���7ۍr������e���Ǧ�4��Qe��j��s��c�	ߧ���W7�8���E�����×�*+�:�M�,��xĸ���L(�����HG�Jl�@:���������S�FJ-m�9B*@�C.H�T��4|�2(b|��-ݴ�쎛ڨEsǒ��7H0�Q�d5�&ق��=�4��v�Ov9���ml�d���<*��� ª���E�>y�>P/�̑6�,�?7mƣ�q�P��@>�� NX�FA�t�l�����e�=�&E�f�?�7����&՗d�4���0ȡD�':���?(u����pW����t�c/�"�-0��!��+�`&���dH(#��4�cd����?JBPC;-ƞ��7�LDW�pz-dw���m����[�Y��F��)В�9H%�;��@JD��`�cp��~�%pʎ���X��&,ظS�t��\����!��dO
�����M�ͧ���v�+p:�a)�0�a���n������V�3��v	�c�}��qڈ_�jӠF,
�S5��#����ƅ5��	.����ǿnh����帇,�Ȉ��ANȯ1�ݻ�*D+r����;�d��V��vp�W��fkbf��B�k��7[�Z�2*m�ُ�λ���(� �1�{���wv1�λ�d��-�%��
ʼ��F��2]�8c��!:�+!&4�����w���1����:���NKa�z$oȲX:�WnK��1���[����O�\\���l*L]��ڜ�4�>B�#��桭� X��@ ��*�}�3�!�L�^AF��J���ݶ��]��A�Yv(E0{��ܘ�P1xY�9ʏ4�%ww򏋻��ni���U���.k��3�=O�%䲀�R2�͖��F�*6l�)��1�*X9�%��]�v=�7G�|�la;��@���f�z<�+z�/ır�K2��n�r��kӎbI�~���������RX'�3�/�O�v ��f�%�}�+*h��!��S�!ǘ�Z���0�D���xCQ"�F����¾��H������{}�!���5�ߡ�ܹǀ��w%܅��H�Ȇ��
/|��f�D�s�5�/ia��2먖�j>�]�8@mMW�ۣC�	*�su^�T\=o�׫���x��I"Ҕ4�$Q�-���6����빟?�D���֩�b�ɦ�}A�:Cme�;�/�1��sp� ��Bq�8u�N��y[����*19�J�@a���U~���=(�`̌�NZ��Ԉ	J��c�z|�����i�$��z��3�$�9�e��w3߈� hm1�?v,���r��v��uَ\���6���&��:�(����[od�ګ��s�� �܌�u�"��<dUv�0�%�PY�{*���i��?��Y��b�
<K�0�q?�CL�&�S�f7Q�-䵘���NH�	����4���j�V]�j��d)L��CNTp�lE����y(��tu�DP����u#�F"q�#�'�	��9�P-��f�b�7j3(�d��V'��Ė��aڍ�v�v6�{A����Ǥj��)ыz�3�bPA�m.����Y���@�'O�~0�G����t���s(߽�I-�� i7��hh{��8����ah�`)ƣދ͙�9V�T�����gG�_
�GP#)R8d�Ɩu��������I.�N�ج5�cpy;� -7�?n'�Okq�m_��MŮZ_9ɪ!tF��|l�)f�����񃈇�V�5�C���3���
��)]��`U�X����q����d�i����_�}�����QE��1�d�L:Q��2�W4���]�?a�H�uYZd�j��9\���iګn\Ȃk;X��L���g����C�7��=>��+�uGPmI�x,�r�+Uf(��>(kl�{Q��I�FZz�]N�S��XB#^{Z����)�Q))&'
�Ԗ��B��T-`7ti̅^NF"�n���}�O���	v�����"��Ϧ��q��E[�!�TTp���橆1�d�02 ���u��&Wc�E?��5v��PX"^������ۦ�a�I
ǡX�Z>�.*��,�h|���2!	�#@I���#T�	��N��a@�bNZoEj�����@�y�t��ty	���Ȫ�B�j�ÓX�+kS�(@�:��JT�,A^���o�T&�wk����Ų���m&�F�˭��[�7����IZ�'�4��	g
��]�&���#'�+Ů�#G*p��
Y/y	y��RY��6j;��XP.i�ɏ���)����&{��B���AA)C�����er�tY` �)��#ߧ+ܱ�k@]X7�z�r.��c�DnSx|�3�pE$�F�*Ï��>�/�6�s~4���+{���,�驶yvL�ar�H���s�vOk���ZJQ_�;nT,_�}�8�9��O�;�W`���=�{�8�r����8]V�'�
�F�alph�@��̡��n�t�I�G�{��*Ę<G���7�wD��R��E��XV9%k?"���ӌHa^�R�w�8���n��Ʉ�,��ަvL@���b��(�n���
G�k��Y*�@r�ye�����l
�V�рu2f]&Gd1��o�3��?���в�&�������$5�z@�WX4��s�a�LNZ+/��|�S!j4	�U�8�V�v�7v�_�9z*�&u�������m�f#s�$�)[���{sIM����q6o��������e���U�,g�lf~���@W޸����F9�;�?��sfL�C�j'1ྂ��#����{�w?�f�1����V����8	y�s���9����Hٮ���=ۦ�F3ٖ>y^I�K_�B}����c7v�e��+>Y�K����@�}�$A�Y�8)����P�&��b��mIm��nm0G�b��g��a.] ���+��r��I	��x�6�K퐥S���DEQ��p,1. t��O��`�KY�y��95�\RC`�(���5��Di����ߊ��M�Tf3�Abe؜߯i���H6I[��L�[��!�^"q$(�
y�NN ��A����F�����11H=��s�����v�I��RJ��Z�_��v2�~�~	R�0�d��.I�4�Z��!\[�:3Aa��ri�&�e��`Fl��X��Q`�j.i���T�Isb�/3LV�v� �M^��v#3�Wv��F�^y�KlBX����+J��� Q?��[Y���U�(2����Jq������I��0��d����5�t��紟<:�c9��j��f��� P:����b�ɺ4Bv�Uq���e��sB�*����a�L�8{K{�k	�.��?R��#��rh�S�΍�Ѐ8�}��T�S��ĸ�z�B�����\�As��X��d�X�m��k��5a��w2�DW'�SGL�$ˣ/�_�Vh�U)ͺ��A�����I�����~�
��!�57��&
-���]���а�}�2g�^^;�5�nq׀f�yk�