// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:23:29 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZF6AYuyCFl7MRR3rN8BcGkToQfbSqho62ZqsMGzldAY68biBTrSg+pW7uYQds3qy
6GFaW7kCdPpSbIayiWUrw3Gz0stH4fDyxwHypx+QuKGik36KcjDNMqXotnXnURyV
uE5srErvFB4BcFMWt5iK8h+t8Or+CsJ3fDbHd2lobjk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12560)
LnsEFnaclJvnUvBakM4eed9sm0w4iRXOloNjj2jUuq5my2B2kX4cfiq9YTnHN8WE
Y+SFMZeeZWaNr3YL8PRIpeORJQrzvXCl1Vf7CmZBXgB3PgN08MpC/m73XtXTo+uI
ILLWGWnqbzbo1ruupHq2w6ogTVidHLwJDYOO0iI2kQ2gFnD3dMR2f+FdtfxlPKIB
BudnkxIlQTuHyiZJwwFCUY1AQ3YqQdR9WxGuKeKr6XhNOTha8lRpwyYl06EbK7MH
o8q/RgvXj6UWwmdrLj75cCV9qI02fFsvkYGJfqpOdKAEYfOdyTsMQD2oJcpPEVw7
T2U/vTIB2eXdeyRGw53sMMxGXohjdd89BvsHJAjU6q+GDA6/W19p8PbN/Utbmsj9
sHeDjLrUmOKbEah0R9wTPcY2V56GtkE04zq4inMXP59WR0S0vBknZEO5uKLzpZ0p
TPMf4wqsqyYk0Zamlmd7gBMQglkuK4FnQ3UMcR7FKY2ZcHJ1f9Gxnq7VzqUmzfFm
7ZHXLqn8iZ0d8OVgD2FmaDo64/rViKRpzn8uUup0mAd1G/wq7eBETMeJ7r0tW7xL
l1kIKaovU9hG++dQ9SX/by+oy0QpqG37duOPTTztGsM5RUDt7YMGarLF7tllYZ1z
qn/GM6lasF8qumluQPBpscrFwP0wbtUoYw5EBSPWt/vN2sQd2ci41VMXGmT35gw0
7eBrk2T6j+JWo3Jux97H2veKRE8WDCICcXKsQkLip9DcCB4LByb1jhRNBPYNBGxb
RKTvxz1xUe/hEuf/c7N5Hdf2HOqTa2g1GS3PBekZUzS9SNFerDPLsihn7zd4Br7A
OHIxhX/3LsgrfUiR+Q7Ent5HUr39QLzZKyEy4L18GOXFsQM+aBRZumDvrQQUZ1UI
9IntQ4kYx5Pjq6oSJovBx3/Ob8EKKWm9mgD86w1PwgluRilS4XE6V2nk6d11klX3
MWDp/I8IjDZiz5sKwCSSaMEBvzvabt5buhYA6tQUnyCEc0WPW+g0vtch9P8uE1ht
+2cZlD3JX8Ygpa6QxqPOBTmutuv1Akpcsbd5FLW9YaS+iayZHslToqg7EDW5mvbw
7dQvXmCxZ+BVOkasPve4kAi7gZaj0GudVhmDvJcjitr7QpVNSq4dZFZ6ErcBTrGi
gGdcxdY2HAqClXoRp6MmrH8zT9+l1bhZx2T2SViPXO9IkFUnd/Z8wHWL6m9bcjgc
8kmfE9VL047IDk8mzwX+y9fl+1GWIaPNxpsfWal3X/RsPanW5f2iZ4I/0fj8f72A
T0Yv12DwD2GwsxPSb3CRKORXfoUF+sSa8N8nA9dUGBH0trjThlORKbsPB3bHZj96
R+vHy7b7orzyGmTuQ1k22Q7rkBVtnJEhZ2XBNJGIfuUVeVIbe0Owu3x9P60abKty
7dH3IId/J0OGH3+8Uhfw00IMX4k3uqmnvRHBmvsj5CIUMQsINS5ipqQdKeREzjgh
fTMMMENIcWDULTVnmwE+a7PCUklgVp1TZfzbew7ouvhGZL8O4H1fRBqmPvM0xJlZ
zfMuI2w9DDChLMYSavdi+iDp0xWAyJfUtAvuXK4Ov8k5SjjKo9Qt4kjlM+61thor
2ze2/UmVJcRYUROhyKwowjjH05dEddTWq+4ilgUqOwOMw4mNJRATX8Idoew6vRqX
PEs3DChaZCYbV4e2535xHymnl7tWRJd9DDelu7ar2DAlN+bPb0tm7kq4hcfa3xoh
FMz1aUWq2bD4LKsiinfOrqvGCV/L6yWBOJ/4FSX9ShbwKIDXAjJ1Zu/vj/s+PJNe
FE+vtbQhFmUqZEv64GtFzD8vTli2EdFx/egbSBXty+AI9Mz6BJoQva0omP+SyKmM
gIvxlzqSPZe7+Be9DTQIjACGIj3wK0S9GumXnHRXxXlkbrDc6nITwAG9JtzhPeXx
RSTtbz/jc7JbJjXFUMmphM9LWngUEOgTMt9oVrScy6QtO8jeTZZVa2Xo3Au4NgmE
MvJdJXmHANLjm1n192t4RnG+5Thij+6H7/4f4Y8Api1XUFSnoe8EHTsqJ90I4BYH
LaI2aTkxdRkIN2Qv7A8j18U4S4JeAPYd7gtldvgy57Y+VKh48QPR0VmrV16DyMSo
BcJOFKLbNwA0LfL4rVmnjdAp/Icw9PpkcEvtHn3jN+vF9UU8bSv/LRwimA76N9rc
8HQBsYGu91UB0rJjnNCGu/Dgg9N9y3JSaUaAKYmL5RVhVUg1BhT34URXZuH2y2Pj
CR/FcYqS765VXZjdC22KnUtRd3W1/DoQw+iJgNJVOOq1+7oNpPAAX4hSdLT7Q/sg
laxsyZs1QGOw4xkPOvJgvExCLL8hSQd/TICL5ucoKgNBLQUYjlaWgJGtNQCU7uF4
ml+xAUWqLuXMNMVkxfhJ8UeZRGNWk0kbhrFDoVGDYnJa0Y1Xwp8wmQDwxgwPrBo7
OBg2gSloSYHd8GH9oivKW+yYX8wQZSeSylD1v2Mf0Xk+gNhA+BLNR9Hyvl7N1fFa
SMBGbC2ctzmrmzfOuBVSAXczS9mq32pFAcZ150jxZOLxm6akzykQnsQPuqrdmXE9
IZZPRntJxWm89ELDjXiWu5QxLlGQjWM2XQP6WA7h0YcVywzWOnlKWvOjURcYpZzn
AoLXqNb5msU77rUZRRodYZgguhwjDaSrfNGP13wBexl0Y/zAR3Eja5EKda0kwI3+
uClWEjM3N/rY2nSUDIJbnK6+47c282+ts0Z0H2AsC3o3L5rJ7iC/SFkgyEUyteke
spilfcqM97qAuVlyMnksA7yjKvTVOzp1OI3htOxhoEVEUmG+pipOJnZOkLMmKdfT
5qJ2beCzCdIY1wczUj3fXzUy3dpzSKe8PiZBnLddsznhkaXDWlm59HJM3hK7UU3T
i9K+bCLDOM3IAhRPs7yGs6oA3nEB7MmPnDlhMID7q1eb14wJnoWf7KNcVhUBkl/F
blUhAA01ZShYMbnHH+j7Y9TmdiyIIvNTPLZ+lloa8ND+KXeh92SEjiNpiKA/3a9c
LZrjCmlOpnwDnXzWuIjeYN67TvhwrN/X/aDYqzvN2MzGvji5nqATgIfatmdIEzhI
S0hVL5OXlCOLa/Wv134hiBDZCeGiYwRbycwZPLLShwJ7GCytepgjcTynVpWiOWkv
0VXcS3g9mVasdoENmq776gfWWdyYcRbYudy5wrD1G/IljcoE4FtgSusqcXLLKVlf
aEhuKDpJmUCiB5glYstP8wr4YmV5xnwLuJmF8UQ7P7aFoC3UXP/k6NEKOi4CnLVA
NCDFd5w5KH+1SRtHomYBdlYSRnSL8AwpoVnZ2S0RTItKH6tw9DKmk/iEQhzgnZ8o
gJdbkix1u7dCCMP0YhphTfFbtDye0xMlKRKjU6yBT7MWLOfIwEc6lwqBEsWf3sxO
/OoIb0G43hv2DU74uDioN6e0WZ7Uxm7ZyOxjSM+jSkZFByjNtzXi5JnUnrBBD4CD
vhtWEtNnY6Hz6hqEWB0fPM7UiRKeONfWeQj2quOvLdj3TpIF/06CFJ3q4E/likP/
OyGBP8ALmWk4A38N20CNKY6D9yQzvnY+W3tYmDWSJXlJG4pUJTpI6Syq65s7lh2L
HAX/Bu7NXG2sUIFOfJEz87iHs1TLMb6Yfsih2ZVIz9omPcnld6kawR54f/d2+buQ
VtC5EabNvhyuktSvGotx3nTA8JJXwXJXsRtxIpKkSApRiTNqfeuD8d4vu/eWVdPV
FaMwqjTtMH9tFKPD1Pw4WhOZcsZcjXwQTq5PohViHji1YfqGvPyxmsp2sFOCk2cG
De6jcEOasHr31LrpNBncc9n9m4MTWLveweczF7a7YOm9JIv5plNuuEa2YF6qxvKv
f14iYr1mpY9aL2CkDMujLkwZOwwIGkm6vruSxFedIDyJUMplb3KCpwO5t2q2M9Nd
noNHAuSyh8/lVLK9P4+DDfWRQ7z/aXc3hWptstKhjER1Jjwwzkt4JRLBu+X/qPKu
JHgEGqjhwno5ZLyTigjlXtaBlUXsc+8dbCIxPzA97WhDjXwXQYknT78V6zHLV31F
qR+gGhJtxnAdqWSGcbzzRrLwossKreXn6Bz7DzPcSsZthIbdcGXzSGSWfTAYqK3l
nBXJdufJi5k0FzREQaNivOEUZlmI90lfd3g5S3ogtZ7L2sTZ0Iz5FV8w8qS65At5
ZVN8EVMfuRPPj6gSM4h22rWA2dcrcFoo/MNTF/82OYkt03YIwdCx+b3vouvIgr/a
myJHbwn7Nt91x6e28Y5g/zZajGpIO1NiFNmQid2TbVls0YPB0wMazZhWModOVCV3
9pGLM2OHZitV7ESgcn4oyOgUlgF74V8el6hOfPS9E7mBVwJuAM4Ode1n1HZ46unW
taV1m01KjVbfKaxIZBHLIyzoN3jzygwRR1Ya1r+9vkpU6+HWRxdIksGe7cEvXHwo
WKhPPojdaeQlAffDwYeRxr3nGaN32re6hgEQOvZECDpZUakxvSqPFembS2grDvF+
uP6cSON1u0D+6R21KxkcCi0SJUhHb6GvyegcOK3hPLth8Z+nbA0YCLqUbifcPA3K
NXj9jwSM9URF/FuBJOcynLicLzIDp6gbsmhHXtaBiJ08SHqt/Wzk5tlO+gD5RIFe
y/uqLCZwMN8W2ccMNruybkmKDoNKzJKj88YNLNKOb2cLS9JQRswgiXQ1Xlpax/mB
WZfT/XQFziR404soztznBUuQSHMAohjt5ZA9YOUZM/rCT5xGp7k6HTpJn7kJ0ERX
YEGvVZW2vauEjhwZq1/y+/bMiXibl+SSDQoR82RVLmgH6+/QdFC5bRPPm4WCy1F/
iFYAQokukqsQep7OJ9lQurulDg4QPRGIkX4M+Cu8UegzCyljNdIeScTyzvnf1Sxw
IfK4mGrvay1ZDbJEvKpzxfEaFEn2kDS1NlH7+gQX8iR6wgIYafmtkfHfoC8K+FDH
RhTKG/01Ly4ws5qpNeOjP5dpmHJLWys48CllNgBPj9Xc0XV2jKjewkDoMEEWY6w6
az3ZNfuFqQEKZgk06k1EDQH3sBNQYnnwpddwt0fACmrpHhjyk/oLOFibNiO3+7Uw
ynaOODWnBsPsRiNd250G0yBqvtDC1U9EShvvs020mEqC/GnpazZX7FkkRr6FrdER
0BgT4D1J3EhnZwS/710ZsbW2KFOb0lAmrmHxBQWq9BOYrzvyKkPy4nS5+mo3qnZL
fqaLYSoiYqct8ZaRVVdI6tvvG/slpsBxsVkk38tRRKSxwEZJEOKWC3Hd6pj4sfAS
grMmZmqF8wdutRWKnIRNST8vKeJSYdtgiRQ48MEOtfQjLKglywC+Hju6kgbI29xj
gEd77VABwdf9j3jPUV84IhcBsl8pB09pXAcZaMkgrUL7Kmca7JlePqwoGm686Im2
beZL90dA1eHO51hBuzM1CPk0bNs2ex8Yernk1/Lp57ISgFmqPCqWhpfhPs2PgVSV
ZEPSRwIrPft0ME4UvF0Rg76Jvb4APf8VDj8YZ6UDJVL7pwErhSin0pgSGsTqwb9w
iQpj2QYQpDdOwYvIYpMBB3ssed+N6V4DJiYRQPjnKr0zjde2UByiltjcWjiIg6nv
wM5k15BDov8a5VFhtsDJ5e7y4sW1wOG+k4Nxxup/7x19kFU/2iIYlxDLIguU6by1
IBy0IClWrgMvZS/BRSjjTM3g+JQtBYIxn/es7JU69fEdOUtFOCFJ+/Vr6TQBmmjS
Kl3ep2jIe2lcQSVJ0kGctXIjxGFERNY8EebDhnUBHsas/xTlTQiF3ZL2ThyTV8eB
Jxoce2vZJZSW5LYPEx7B7B2G2tik2W/zkTT9GQZmQ5TMtNfIKjSgPMh6iJEdACwR
fkMsIg7VD8AAk23kastE8B5YRAlAqbzGNKPqzpHwY9GBVfuTO9O5mFHso29bVB6p
KMOWUQhJqY1R9FypVqS24yeMNAVJYOSa6ogfosozpjQUVIX+u5S8Hv1o+ceJ4Ywu
d10c/XTa82XA6HuN+wTdfZlPu11aeDkvTNTdSnKSOoXRxCpJOqUD7gmofXD+JNoF
BqkZnOZjn34ssinpF1Mtx7YR6j7fifwbqAqssofcN6dRKcp+Cdonw3RXejM7re1n
0vxdQQ9MEbbU6sXbq52ZiXGNoqbjjYAarzWG5+TI8cRZWBw0CWpM/nNVV0ycfhd9
yZDIS/KnRnlQEOGA/c8Qht/vpadoH9hd1z3ZIGOBoHZBlnYhif6+R7iGcRIvzxZU
OiDMoyCenAj4KpCpEytaf9Zl4XiWu0Y052Bsbq+s0YurJDGJjMbiEVlurZBQ30IT
w/lV+G9D683fOhHtdwri2C9iKUs5mTLHCHDEv67MdKzEs8R0TcQuKOFhnQYBDtHP
VQkVmhWQdWUpyT7mZvJhplOgoKEOy4xMbJcSdoGw8JAY+CdgziX7JGIFOrAYMdpi
1KHn8rqKildvHvxu8M9Xp1EKEkmh9q0jxdYJi10dkvRQoevy+1mZsX7lenXS84cI
Lr1fWc2GvLMymjG3nSEqA8X/sCIlm2FdDAiAlK0UCkgiT2e/fnX2xC28iRcI/aLA
QBKk2UWbiZb0zSJRL40Bj7wauEJLt+FqiN6jLzqQ9qIi164j/tknWxw2MkoIy03I
05V1/oIFu2E4wE34x86Xl4IEym77YxRs83LExLlDVPyDy7RuN7K1EgfE4HhuZVWE
S0oDsiA9LltPex10P7vLbU+MblLZ+TZ8Q1vjuo8wXX9K3reZoUrOmMvkg2SVketV
Q7UQPJEz8eRhFAn99JNQGhEXQBMB/hqF8G3LhPn0Ie7kfs8jnGbhFenpW2A67sPZ
y0ldlGwBa16sDO1EKrmtdEEglsvgi6Cya/0Q/JRUzkpI+McGG/O0JBs4BdloIko9
w9f/FA5+FXZqL8akZc3jS9chYiQgAyn0IYW446KiCq5KTgpobHx+zNs6K+JuhM3Y
KTLeX/oiN1qPeHTISwK3BE/C3YeEwIriVFqJ4zUjeijMVNWAORByMg7hFpHwDQFm
2PruWUvuMAIFLg/mJW4iF4Z13mgAcFL3Kwr/n9+lWkpjR6Za2R489U74HXii3LO+
KWfeEHiypbVS3DNuqAtaQ6jrRgg0/8asCSYgW+2bcMxOlPmbhhBRJlYEEVNxKwvy
KAKO3LzeENV2cj/oXkTQWscGsjXwapTehF5Xv8AbbtT0rr0VelWpurQO0ZSODnDB
zBEHFu+CqkuWHwYnXnJWy+VIt7cubYb7jECvUYT5qljfjLVJJR9M7qIFhE34kqXG
QRyMAarYqiSYAmrMakhkjuF4EutQTy3bfvefWUs7rOwm94Yd7jy6Rq2ZzNL2vpTO
OuIKGqLTwGo+n8CcgIVx6TlqAlIk5fofCOankMovUj7CBDDb5apOlRAzmXaoIHVh
RXrOh/5JrU92gOKZDtVPULpROwsnEjfbu9tadMnOVhuQ7tdSYRHEs47GoTTESZqp
1AK/MF8g6gOD2CcfeNXHItQQ+OTxOsZdBOCnC1yT5lWePFnjX/fX3iWtsJsUNDoB
qf16J6avN4jcbYP9MyWzFIiQy711SAU22bWiFEXGMVxJW8REu+mcvv1vIX5NxzPe
9p/fMhRUyhBn98nGXdeWsIsPKY6Ia0Tufdf5peD1MCwo9JvSF/6DBKAx/UmdjoNa
5Sg95V8Qyxu26nQLc+BmzYV0c05xxCfVTxOtzS2z+fdVHHOzArM8JhNwmnkZSCDy
PAu3oZS56kSTHTOBMPXbvWaqR7lgooS/9F2dy9MbPC/ed4QEc9m8kUxeNrdrtODW
9kJO4bZXBB0gK/f4QUegISAC4Ll3CftfifkJYO+qgH5zOjqU25MJ03KCmwSSlh7y
FbmWpQZfcwGEryrgtji0c04JMbNTMNt4XqnuXqy6OYqV9n6vwcqbMBQjMCgRo7nU
RHu5GNZ/4WecrVq+jQU+L6s/Vxs6hP58b6LU6me+b5nMxFthooIZTP0nOR0MEpmN
o75re9VjeBtrZTL9tH+x8mHe7YABnHvRc7TAf6vd8nTQDehXWp25fdl5rA+yFT5c
RpgydyVbe760qawJc10v2+PUU223UaFfXWPDYDJqJYRlNxxYPr/Dhlg9LMraCv5k
YwICIG7WDWoySvyGOt402haHuYaW2RZwlAZkYak5SvRmJoSAol46zvfwHDSsMwjb
d69W5TwPjFNldj7ixyPvoMkJj4arhTVNYZhxvCNnQA3qvso9n6G8CqnVtDyOmD3Z
GSNK9JH0V/Oj20XOunW3Esg/56ZnqBFCx/wMLHV0uNmh3y9YliSP4tVwg97SF8N4
aOe7aHvG0Rblz2lisBC+mEBNWLW/hqKExJSomT1MTv4WXR/JT76g7/U0Y1N895D+
gffE72E7UN3+CEkSdOMx3yxQv2qSw+kFu+uG4pxZgzszqjg4mTvINYAur9H+RyIM
nxl3qAiw3vQtpbTsySAtEpk14E8Nu3nMFBHF/FK9N0QiiWc1H0hjwI4iXAdB/+D5
N/hZLaqzlZr1qAIqievbA1O2mf5VhCKfQo1uvHCeu8PzAwq8+ucNyGPMd8pzrclO
1vG5afM95AVES1AWGfFsgP78jmJ1/Xr+iCXlVyBsh6HUQXQQccjWWhUu5ktYCXxp
r7GOq27ttj6OXOXXtphegDesEN5g3fEMOpbu2KEk8bAmzbHDF3dABh3mGJF7GmBh
pIwxDaT184ZdCtECx1ou92KRtpMhDmYZAZkRnVivA/9s6GFjhDjYei1M51G2kNWm
MhD177AnEuQ550UuV4HVtdaxw/5gRoRI08mGaTT6ejyuzGaZLy+Cy7mSqaChO9ac
cB0rQ37M4RQaZeHUtFi2pLogR29hgmqZ9Go0lJIWMFfRn7sxyQ/NZYEF8Bm2bX0H
/d9yl43b7snVK4kCBHfR3/r80uFCa0QBnVlzM6pLazZ+kEmaDbQprvxnv3t0CU4g
tPJnIFVzH5QYr1rZUV9Yp/o1jot62Q9aEE4By6PhwrMA6TumqKfxiO+/ufLR4V6u
yz7E1oysD0PIC9dNjvGrxBSDU6YJ5VqlXZOt3ZLxm2malCol61oEPccCQpFOxmgN
1ZAKrAFOKU7Ny488U2E2ixLlUYM/G6vFmrLprpJFHcW2/KhMjUSl29BGgBf5s0D8
suWP/yPraXoQEPpTPtcfupLz3YwOyQB7zp5rISfzZQZx3ucFLFSFMADbaO02B1w9
TNOql7kRj3wA9QMjw8o5hTxK07Mr02KUIrhGp6Jf2zA4CItRt1n7vjuBzmDbot8y
5QQ4U0nN88XS0kmkCe9MIsVquGMrReBQMCj0WlDENLDqw+bc14IlZ9gVapjC+kw5
CZ5VdDDh3yi7/cuwD3HJkbB8VKBqAfz0eCEXJ59qtW+JH4C//gCh1QU/cRIr9EGZ
BQK43YctdZJUi+Qx8LPX6L9hhbNzjfiEZ1CNcLVK/XjTDbADcg06pwztozY6IHY3
32mv+fLHdBGUWe+kYoK/IGYnTwHg4y2YTtiPF94DukP3FyAE+KXCwbwxp28RE8j0
08j31O3wK187TWTWex/NlOJJ+wra7IpjgqfEnZEFXGSPQD1GfYRWLtCsihW+1uqA
StnOTIziYUV65j7O2wNv7geLyTjGpA6SQLJ77BlTNFokyepPFYooCIPe+4GlxYYN
Ojf/oIXGJtKg2i9uunuvGI7uthUbDMLQigb56NbTvS9ddXP/cqcwuTFj4gzfO5oD
YKGUjxcaWB8reLplVjpR0goTfVRiV2x7n51YC1iczRGvYN8DeaMYVQ8O2u51hXru
cgt9tg7LjB3eYh1QCc5MBWFobQdQl1X5ZGXyb837jAO0N60t5xjhotQRbhWGyI6E
Ug9N64fvwk5dL5JruG26zq82SQgIxWusIgcEXm3gLxFdN2cTejXcGGF3R0682Tr2
xDB0RbkVdFhkZmE+0g8KYKyta1Fk33p28u2iXmCbYSE+yNYH10RjaLmJARF1et1C
tLA7MSZxmgD+HepQsS3JyGSI+827P1IcA60nD46pbZPBejKFkSsAzpzxnlGC9VQk
QGmwdRNyrd+S1U+omdY6CKAoTsl6UUAgB8oO3BfFw9FgXWJ6op1zrtQ17sN64xxf
iLcG0YNHZnua0YUU6mV7R+264GFmZZsdPBDP6YfnngC6Ke00uaAzMIcGgm/iwZA4
kpz9ks94Zvtl7iJVijhjL3PpZE4OgdJPaLjdTce6iT/5MpP7Vv0auBzPefQORJEf
w58a0364pM87gq6vbj0FApU5CRHNoxLWo0WG+Hv0Q7U4tYFsPJ5ZA50rM7Mta/5r
OfvhoEsZRiH2QvhGnYrvmS7VusECUqtHU1edRAM46ZEoPZ9u8WX2953N3EajjbAL
Fo/C0952w04KANNCQfYJCJGWvLW214ouK7wa2RO9W2j7TvVqASLEbwh9F2zZdDt2
QfibgG73BVeWZdQ8SpRJ+V1wsnw4unkrSm0olX1tnhbPhJbjwEBjt2oB9lmMpY8Z
J7G55JsFXRqXd02uqxcIwRN/6OMf8PYCw9D04mDXoL9/vOj1/+iOt/UheKpqshKA
3tqyRW7H5lJV5QLm8Z9t/mbVaEfq9FskGcKHlJuSg8BrR92TFw8sbyRG21PkW9a6
y0aFIrQVBUuxZPJEnCS/R/dUpeNiQn3T+lFKaUPjszp1MtZntRWimLN3T0PKQtAN
Vunxzy/sQCR3VKeqHppc2cf5U1J0xhxw8BtAS1pvyYenKT7K8lmypCJWT+h/fgpd
vIka9y4FpAV2W2vv/wZwRHrKKhC83j54Jz+PniZJJqmqoJs0vYi3iiPRFWUz6y+o
23oGl86XHzwKq9+a2kwi+dSEpVKzwh0iNpEVVwhkCTUzlIL4DALe3Jc+TJgVBvqy
CdLpGyw2fxvESa8epMTFAcnKqnYwSdUJjrHj75+fuINERiq2RiVVSBU0/9SnsuqD
5KhnqUWF4JLSdQxpivdrWyKn5WnoPWsk002NluRCZsbIBDFEjujNF7NHxXPBOsca
tkqKHcQy+IAElh5qnUjdgpTr339uBTw3KzNlkGWJDkol+kYggb93mEiC2aqno7WI
AkmfqRVnmC/hGnggabLy7fWdGWgJJKBk3IfgjZ7U5RXYvbGTs6hxS4L/kysn3PAi
eMBykwApr8Rs+k8YDPMqt2S505aLLqXNO7F97yqMHqIA9aQ5KBMVP0yH/tFlCUDi
zmkHlxT44h8TSlfJlfFMWR0SO9wyQLZk+EfZi68/NKsVNOxQAzWzOmk3SfCl2QFq
ZFldMzsRXSm3ukd6Ldpp42MzEch+u6ciXtvUPUVbf+BRjJW+Ie58A2wdXZ8cyxpa
CVRrB+mKxYxMMLItR8H0a4TdUlwAmM3NzwuBrEnH1E2Xmz4u2zTK/Oyi8eoq6Uuj
E3pAd7fllZyF3uwfr1KUP7Hs/eJ9Y+r/HvjPqcCh7JFUgDeJEVlbYhBzP5xcXDbG
vS6Rt8TRQ98LR5nyHLwhv/8Zsch98HFETy84M8178SmL51ptV3PlO//EU6k3LhVl
iw+LiskLqtC3Tu2yCcQ9XzdlH6M0jbN3EYTVwUWc1ltRBXN7y6PnFHzjD5FFIVUr
6DtBfCoQ6Y5OiAgk73djwfIXxPW5ImjczzZgG0pC6MmOZLdEwsjLPgB88kNm7cBO
Zvqo5VfeAcv0If+qJALqu4AQDHGB1PKm2Wq8kw27Ox/DaabTZ5+J1vCKErvJV1Iy
4pwOIlUXeX/cgA9Z2qz1vo9Bdjrl3emW+CF9IMw1dc3wbTiDRDsZxr4o8aicaGwI
LEMt4VRxl46ZT5+7LDRw9VmNiByfQkiHJXSWH1DCkFlLEa5ZDQZYHbQ6ufqRGyQM
HYBi3Iq1lKZKyeWDtCcv3JSNX5VawDTreC+AsjGj47amOQZYeGIaEjOD0LMJDZBR
yAfSEdmuugQ6CLQ3+sEMi+JtPfrefLmMjNXEi0bWiE5OYHEJFkvFxQh+bEn9Gw3R
m6rdYAsrKcBVOb6yRc5n2iACiH8Myy0DcmYOb81ES6mrJ5Lg8zonZIDnW5xMLV85
NzO1RasFzWzKk+qhx63SnC7wksmuS84Q5pUYA6Me3ldZK8YnYeAS6TyK4tMND9DF
kl85dXn4QGw9pfSO5RO2dUEV1T0oECmPN+agXQkz7Xq+NRAOIt9WxvzaUen3nk8J
6TfUioP2tJoLlreOUnhU6IadFBcoCvICR29OvpFMP3Yk9JG2Ht6VbCCW1xxsWJdM
BBdSpjs2A1D7XOMaOOzWbNL4GHp3rNQf0Ixv+OuqfJYyUQKU+nqLfO3pyZdf4dYh
ImNIwWj6i6J82gxGIfMARmoa58nR6fLBpByuZMT0zn4ODDIg2egCm9qsUIsPzM4U
2F2lRBYyn3qn2AUCW1HM+KCHD+on5ahQ/34SttYBi85eXtgNdxjijme+R4sO5weR
Iruplsr913lEqqtvAqsfQrbMQVYOxlRci5Ue5CTWF3pUQ+wUBH2A5/2xe1wjtlKD
JEKKXxIIZn48QgOfhIvtn5ZbdfyGgc4NJyvRGU9UFuOb0AxEJOvqxmkrOdCv7R4/
5Ntdrw055m0l5ARn0tUY73t5C7Z1hXIo/hoIuvYkh727XCcJaMl9865vpSYYhjf+
bVBSMKD9bua0gG1jxEeRZ5yVJe98I0Wv4tYM4jyl4cvsEZm+orulhEKz/t1Hnqrl
FRjEhcBDofu6rgQtMb5EORbXCSptv43HozSw8FdT+VFML5tjyUpPdGqNFcB49LYz
AY6AhIvYjcyaebpU4RCohh639D5Ute5JCusPMwB3wiUj3gR0ARFfFnT5WrFBaUcx
PhgBzFZst93MuTryc6Jw2c4Q1Mo7U9KDlA/M1+LowwTfsIEVig0RbjwnMLG8NwE6
wRxYcwhJ2N9e1h0XxtEsp96OOeXYjx1dHK85vcVutXZUPN9IeMSnWTQH/WvdHn2X
VHebxsuv80s2z8buXnk0OSd+CHFRrsTiFiMOpj5hQcBp5UCqwPEVD3ArmGgc6jMy
6xe7LSX2jm9PQyLAN617WLY2FOwvydUNdIu2r+VLoyLYAjf0Qby5/Cz6NvQBCcaL
VexFAdYcbwUo80c8tw/HT9QJEsbwL3rRL7vTiE3S/7/FYy1E6+QPoAVWi+ipO+j6
gT18dO+8F9B59gnqIyPLMex4DYecGGG7fVuIs+rMMkhcwfIDv54eB4xCq9LBxFix
+ttkLZFdS9i10BBkuPBLujPZQfKdDoh4jLSjZMSFxczm6tLdpcaSW4Y5vQlt1tEU
ziLtTqOOptxawK26EmEHy+kH20uFqbmLkAVHyz7tufL1egzaY5/tlnaVRl2ZVYZV
2GSln37GD5tmyWd6Y2m9IOdyDJ6P2oGwkdrjOoGX/HVsTIeWSuNnmklDo4NIWvhg
bVpxxzEFyQLf0B3fSrWH6GT/582TUztboU1kx5Q2KXPIR/Jy+xjyEsTaoiJ4F2rR
y3kz7Bfw7LKM8UCeaU+X0zuTUQzHkMWMG4I05rzqaIh8a/DpQmHE9MVbejBiIIsc
VWWkBGvdRkDxDb04XPJucKs5DTfI+P5aQFGvVYTusAAeGfc0VDGEtnU117gLVYO5
QXS4OAcCrOKsD9Qr77cy/Ft7fF9CDpBIM3XlTwPn+/pFPEKwlvyHxEuFczd93NHo
cIIdqydktQVDx+Z8ICLe46Kh6NQxZZg9gB1lEUrn+vQ+LRjgPLd6EhdALhfqv7c4
XS7qS4q8m3Z8j92stL5wC1+TkfTYUM/jcwpor+vnxu7DvVM8NWPTySWk1KQQRK2i
8XzU+sSGXAwLB9gj7HLRYLJ/8oNgHhDKi42dlzfP9tsQbz989I+y4TaM7gPsvL/A
x4kKA05a/0sYzj9ObhRyFoFw0QaIN5IWpPJxzSquGr5rWcOlvA9FvKoJ0MKyzI4z
tVHlWxTDbAB3A5BZRkz2Zj266c8T4ZLL1wCBMs4Z8nXT5ZDyLlPRZX6RuC4SOhtZ
jlNQKoUCdl7+IkOohcQzrdnQcssYuKomTLy6ujWCsEbiP+IG0WmkyqEOmpx8GGKJ
pM9pMT8JX7BeRL8fIsKEwAB88hSeKBGy+7gHxNPxZ815uMlS7VNGTQNnLrr+UmSE
d2XPKUhgWCMK/JRKCuBUY6YwK4ns9eeROZKzCxMSHltl8KljWpXvGo4RunI70gXX
QZFA8dH0R2GEMh065cqkurTEzoDXWqlEXGjzDYDEBCfJdTUVI1utVwmYBr9MDIvr
S2BSNydLEFoKVMaGsGD5XsXt9x2lXPS8d/nDeN1854FIxfFfoerYNMq81R8NUhZo
T9hEmXyu9V51IX8ryMqlYLo4geBTRJgiuYBogrVApF3qrheMlD4cvIo+1FDs+c6h
BEVnCorV4d5kAV2MCJfMYBvidfQXX6nQGOqBNLY/8W8dQdxJNV0OCCEqqZRAyteN
zTHgXal/nyEIJUtICsceIRtaoaiMkkFwiWRp71jgbR3Qn3WiPTQzHjlA9LEChCGh
i40LQgKYUksCiafmR/AJO7m+5olQK2VH5jxf2tW4jZ1Maz+nhVNBrmYmvNOfFwv9
gmRU6+JROS7i0TQ94dmJGWPtuMLagYin3/axowgR/xqyBF2Lf1QJeMQ/yPPiB60B
86pW3L4CUARAQzG0YviJwkBRXyGIPVse0PANEgvgj1MnqY0z74BYMmgixv7tIR1d
f4oGzmPMBpZOpPst+zJZJIBhPH4sb2IEVE76SbXhZAf9CX/fYqxDHRn0eSUXGdFb
5VzGAUMQboWfFVmluQkUF2XLyAHVe54Mlgz8DrcvNUvdCiVsu7+ysAQMvamzmr/R
R3G2OBtMD66S/pf4yJA0AeO2Zg0HwC9C+MMLhSLWV8HSKA4EHvklpJNjVnMjcOYR
B+iOORVXDI6GkE7UTaM/IMsBcvmD4lCOADyx0Z5IStiwcgXJfpJ8uy/6mjvmwBeG
hiq3g4Em8RXrwQhogrz2JfNmL6J9WCvz9dlWsRZGm8oSKQ1cBMD6XCKEcfnOT1dy
HlHWIrSB18ZrrcOttD01+IC1z40YVSzIlZIn3nwPa0lNI+AaBzNfP08a/we4Qf6T
i5dnO3jrHmqRyyMprm7x50XvxdK8yzZmW3bV66+L8ktOISEVpe1oNrKyX9yVzBLN
KU+CyPYLQy93LNPc3u7iFqndBlR68iInLMgK659QJRKPJzoCoYfNhCgkrOwGMNYj
EeIFH4LhSyrz5he3AfP8WmwHB1Eo5OyOsmqrqk31QMEb/e99lGUVhpInsiwZeoUC
vhxb0vuf/4sS6S2AR1Iq6AoITZ606pmlR+90XjPzu29cYqi69NMMNNOA8xEd8AfY
0yaxJGrs5YJlAB+9+m7315S3XoLlobxDG/6rTtK0mQu9xEEk9/OXBbmbqBlIipJV
RIAHdnY+KXwmmnFlbaPWN8sLkwMNWFslZdE30vYLZvUwO6K5uJ26EzCeKsoNdw6W
448W/yXSJzyjYrs/nZHGMG69fN7RvETmKc6HB1TtB+STsndHIiv48RgftY6RmTa+
ukhvAreX6fVv2zcnrG3+N4FRuk2kSJk7dHir9usMC5Bw/vcc9vCdXyHCK246OJCI
LYPaox4UcheZFeRG84x4/oUyXQ9SZavwD4sI+OESEWH2dRMPA/VQTucS41xM3ma5
2aOw61yldBeJCS2lEyAsln3ORM8TsujeE9kdWTc8M8x35koQmqX58zPRiWnM6gy+
BQdE3PCUGM8i+A4T5Iw+gu4WMM5r9rNaI2GlITz7WJvmkBdH657hSIyizt7vwgXW
ccTcqtKkY0VEH5+MXJ5pm/tXBaZCVSDxxDqq0teqdGJqvKwWE9lHiPBJkQmw1nzJ
JnyptHm9hMzUBrNUh3+jb9sHAa+uWtxryMqCHopmupA+MLIro4sjZQUCoishTitA
++z3TA8mLVNqCqCffs9FvverrrIMqWq54yiRmgCXWvOxFdpCFH6UJb7GdGOIhIMj
lSvafIhAEgdAp5g9+oB6YpKLnFgho/SbC5bthSDnp+kvyfW2KBynr/udmO0dPnUh
PlYuo0TIzOFmEYf410CgmbiJhixQTR1FOtZRDLGgwedcSfrwYQo5L2Cq3AP7gqQa
0Q7XnHzn3nItwnYFdteqGOyl/7WpAB5IStFpoB0WnUI16ikJuwq2VFrhGAIk/PdB
6CgZCFkT7d6VQvwksUYXVIjblOVx7KpTOEkBr7shsd3qhnj/QJ1qMRgMMPy/ih83
nIR6sE6IMU4CZmCJhRfjKdN1CmRxBWAeYZRqZphtA/0bw5RkPhh49drxRb25hMFb
ZttRfn1+7NtcKUTanT06SobFYzK2WbUXe/wAKGpC4HLc1DhjqUqj5h6gEqgeHuRo
hEnq7KgOGlFv6nc428F+7gLJL6YRPxRZLzpwUvNLIT+Efb2ssXhxNeHSEfzwXOez
wIjSMlx5U/Y6pq5grglP9Ozy27DR4WnLcAxiqfATMkq15Yp8BQor4Lx2bYtC54PP
8o8bqFnDof4a8e+ZGgnAk4d3SwArz9x+pf75HYcgzVcU1G9CXGLaoTlcrGHiNA8Q
Wwap6ivOcA+IHPT/jHCbD7FFB+tdlswKFDHZQAqi7y7fLwvv1CgHwzk5TqaUDEft
ZDSW4Udzp37sSDJvpQaPqQKzeojDXDQdf/2ZIuqPumKyZApY4TLL3Ez4kL+QBuDY
6HHAaBDykQZpDYDFfIOyjYSATdayVdthxOLCKvC0Ts7AfGXQu47yrEEfu9gds2wj
3GtsiE2jycSwbzv5NRAmknCBhlo4t4hbekR9c81OwyaSWyArzAprr9LwaK5cBd+n
rBfolB8w/Or6RJI6UMEHdom72uirR+jJ2qQsojEp9pM=
`pragma protect end_protected
