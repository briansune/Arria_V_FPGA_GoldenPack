// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:19 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pEIx50xwZDjpfUlLKRDoSU0abNCbwAL/zYmdh8+nmp70hnoirvJizXMmtUIZgRWQ
vekVKW+kx/g7Y8nvb3XLr13DhKlGG36Ms6zzlINljwPAiwNfOu6kEolSPh4D7nil
9QIHIB08Lfyib4CU6rfWxJ1DWvfUSrHLey6MlfpqchI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
oVXGgYfSsr8NuLvXFOf9JoGqXlTtUcq1kXg9DXvmjepuJbdDrfOlmLH3Q9wFmCuW
4uplhByt51VOJrPFk9E4j0CBGCV+FUHEi31XkCVEq/UYTYh9foR2+RFAJlx2Db7/
o0V5mXH3Mj1/gHzvRmvmljZLhyiTNvRwwDhmEyC95KYHFBxr1qVKg5XCc9s/pMQq
wqEnL7nY0ncf1DQl0RFIQ1P0hY/u1Mq6PeC86Fw5wkisJYx6HzPNJV10zYWyn1BJ
glyam09cGSDqTxpdcSQbLvyxrHvnnMifr0TRa/1b83xfzpeEw0aNW99mezssPU9V
xNxnZ2jZVKonS1ES87mpFO6Q7ceit2IpH3OU7QwcjQhatspRwaERA8Ie7tSN+i4i
txSFi4OdD/+/RZSCubCahdSHmbt+v+xbx+D8ZP9AIHOJ1Bb2BW44lCqwx4HbSDsc
xncIbOABd2pZtJ5BJDIUIxJI4ZitMtObnUnDxQ+m0DnRT5PLsPMesBhJz2D8rXsT
06RnSOJIRedzR8QRf41tBO8iu4OP5UKW71EqnOYeBYQccKYFNomM1a+o7mLPZ89n
Y2uiW+ULGcf0pzkJNSA2uYBgE48+Ksbk9mmkacIl+SfB/na9OBS5NCBAIm/l19gF
v+Wy+V2KQuw7iqNrdm/72Eagqmu8qj/L7BV9O4ihUj4X7q4yNmfXL7ML7VtYl+n/
8zPXh4SrBRWVd7cYLj2HxaE2Jjg59NWpSWyIDj3URN/vkXeLIv6eUnPN8QBa5gw9
Fa7UKsgM0cr/9AeDvT1UZW+J/TPC3m8pBVQaV6n3VEfWJe2MH00rWkQ+l9xJfwx5
k3+n8p/VSlYT5wYFlFE6GpvxXG3QB6sSTZa+89NUQiZRgjgzYWGKWmPnhHredqQP
JGs3RGRdiWtSPoWQ5xrVlbIPvT3LaRA6yQPtpdshsjU3HDtarfxe2aYYrSDnSBGS
D7KfjE2u2bteRUN9FMDMi7isjLtssYEaIPMMo3RidDsv61GtdqCWL1jadmcsXW8z
JGuS/cn2qESmnZmBtnBmFzOqGXgAXymwDLHE5jiWVw9AuCxN+vMEdXDc/xKPsYTU
zg8HlL1yD09/efTkntMFHhyFF1s77Hzdym+gRXFT6FsnRgupyy3Rd96iDDrv2pkU
YTFoXI/g6DWyIb+fq5cPmh9VgunvmEoavDQrF1fCQ49bWVDsexCSpuzgri0mUSma
eqKhmgKE4WePq2gK8yp2RUE8gTKImKgCZwNf1gCpQFEVGhilR4LH+8+VGrhwUhWZ
ab2EClOpXiiMyqDB3bnGbpO62KNW5teOWNLUP5HNSAuv7K+XqY8JKFkp23s+FzwM
ZpB+o+ffe+zse2WlR1XjMLMZcl/XoWgMrG/LMEQI+VXS7zEIH4P6i+wGsdDrL5pu
lHoMQo89E1UEzXmi/df3m33XS59WIfyp8bb/6WSzewfMDM4s9pq20rU+3+r3eqse
EyGwJr0626rYs7HC62tUbJ64eDGtTvp/ktIyRxQq01fkU6Vb5A/FI9Ti6yop+2xx
4XeMy80Dtu/91+cshxUd2F5rxjHvLmwCgO4IKkW6vYuVGoGafTMM5qKsl5QZhwdz
CJmy8vyyePVRN/RUAaY3aa8x+As12PodnMmTqKXWGlR1cyP4ubHxOn6+CHDUO/Zg
xxzDJMWzLiJVwud13fujHGPUnOJPVRiqz6IGnGA+6IP2FsN7OPr4zQP1+i9G4rik
Z4ppZgXnBcrk8Ktr6i163VrjS3OyhB9cZAB4oyc7GE4Svpi7p+prHhD6S+7pxR3E
h4QsUaycVmcEl4CNx6cvpUkmXarC6mTeH2dGQtOXBNz7ZG6PxBeT3v3D9A10L5Xa
pCNUXrURB4EEX5faKVKBX0IJAjksHXauO9CZ/tnIJFcJHSvY1yT/TqtBLeyyysNk
uef+nuSMPyDmAMz9aPC2u1ia/i0pK2Rym0ZeFpV+xY9721WJlulnZ1ylFlzb1um9
9PYtKjMCCxM1llAvVJaj5KPG3aAeyIXBmv+IT3A6bOSawsAnYjn51/AYt7LQ82yj
okHKDgNahSGr6AuqGihHbJcg0T4jNK9tqj5UQZCO7HVF4sDDiXBnjLSxTwS0PFTI
sdJoNmKZG8I/J7Fyad0A1QPGHMWWA7O63IPHNdNRuB0KYyfEU6402cYyLjifUl+a
sY+cT7evOtOsChmz+2hJ7uimX4tgolOhWkyDR8+quOXlxa6gqZAnmC8qpSoiewUE
cCC/Gg0KTZX1TMqvg0ezp9gG2U3RB3TxG0Lc1uJrNuvC4P6YVF1tUBaj8BzC9P0Z
neDGd/x8AOz0RXN1uFWEJQNfUjUQIsGcOJdKFvYlwHIcrIIIYoLRv9QW6ZGPe5Vs
5ZS2Hdl6sSEKM+ndZtX1nYjDPfFoPyUyG4hjiSie12PZ0BLDz77l4daLKpMNlB67
N05JeoxkDGFV59wXIxu2hprlxah3yd4W+hgQXATFDuzgRAWqk1UnQ0f64HWETMLO
uT6ZF1zAahT06TWJ4uqz2hh0U2UWo67CGXQpGOLzQeJaxD3us/RU0IhuWpAhGlxL
nFl30AjjagVm+m1QskggGOuoOYXw7DayXr+VHJuINP+fhJKooPXUx8ryPXr6hFvI
REHRGJQRa9DKwq3nf6Mp1C4WuvQYWR79I2iUeE2ERg0l4PRz9rwI1KTFBIWlyScC
NouFFFtpPln10ZvbXpzQ3E4bQ37PfhnRWQMT2BwiOD79mzeneAQ8n+L/bfeYJzY1
34fk7tOJZzETvcCQHGlSfxf9lIDaOGub9ecBMlt8Va1FaTEP9QyxPgk8tSWrRaTi
D6TQMAxfAyICZgKTjqDd9ePK0n7rSu16MZI1oiPt9ubqQ6GW8bjkJ6uCxR5V0cee
L3N5dzgJA6D0vGd/Y6YEXrpHsjZ/cl8cEuISpmmc6EANVi4DN2RddwLv3cZ/RkmY
cz1z5puQpHZwgHoAUJM2lT6o7ztLtBMLTrWCNQkTuumIhBd8nbdXQqR6DvOTeVrV
ElZrpqoaUgLQh2MUdmpNW9tPwgkWfHQareZwzk9uK1LPK6CyPpnF2/CP3y5piZ5n
15TwKfRd+9is48qVCOvnpZpWKRZ5CEk7ePcy2YtzZj5AH7A3WSli7L9NYjgcVsSh
TbO2aGZPk1hblZf5qGLKQq9WO/6SXLNYG3WzcLr1kaio+dam/h70JB611rJcV4py
AiGX7aBESwNvH99k2Wr101YT+g9OhNJmCoE+BCJNGnAHPqEHs/A6gWs82ISCtPb2
P+rWTstmk2eWT3tBgBTGkMDGMuCfIiQsikLT5kwjqhIryyFwW9PqUluZev+Y9Y5M
wU3/1mP8S2r4hsLTDtJ1K97Ty5faBcb31YlSdSX64RfgHWNDn7Eg+xgZsHd4HKm0
sKOVUFcJ0bjGAX1yPKmadmR7aGhd99e6bp2beourL153WRCOJPcyswrEbMtSIKQs
U3yRUBS808qLB212OHWU7z6kWVT+zfTf/eFCvgeXtBCy5hc2dUs/T5byUdJrqTIo
4cUMNqgRW11wSxK9vwObxK+h9MA9HJ2oGwm6u9amrWlIBcrrDPvmFq24zw6inrUT
YUbua42+edE2qsWksmLwjssITBS+deDN3As6HqVPLl8bqm2YcfQl4gYjjmQyph2O
lmLMXr6/Qv8zJL4nw/K9MSPXXV/S7CS02WzLelq8nAZF8RjHPvUjq5U715gb5kB9
d2gBH/Xc74EDIgZ4azobkfICKni9pNZVOlPVA2r67HgHz44Z96ZnudxGiOtjm23v
ihyMC0iWe9RawtyKEP1aXqoT3baTpMTq8LUgHIFbCV7vgGtOrkZTFa65OLWPXzvW
QQUsBFmn1rBHleXUcKrMiUJ5YCfcHI47YmiNFq5Hqrf9FhwByw9+SUBGdLIjrfE5
oDaycrZw0ZQjGOGWuU2JluyNpVBXM2mbxLJliHMzU8i6/LB1VXAukTRaXlDYjYLx
BvCsGV7ryu/pV5WrfQqZ+e4QN7QS+rQICQKUvrHE15YELItDlSgOwC2dZpyaN+eS
wF5yEF22bBAXNNDRmFV02SggntZhe9/zdD1/Cun9yq+YsvvG8W3ILTGNE9hXAsqP
Hr34Ne3YPAUtH52/qeFgctecSJMQqfb4Rl8SQ3OFWPMSyWcianoiSoo5Y2N+oLEP
OTOpR85GHX/vxAU5ceKwaZR4ai/A2JsARiXz1fQKnvpmSRFCZeeIhwWUJjL7VKJ1
4jJpprXj/9Hz7PEkKjHUEFOKhLsVG+LFChzsEnIba7XTKd1NiO1YD/5szho0nA5T
89gf2fgDdycCTXtgRFsuDJS77ht9xsyHpizSWL0iz/oW/6UiaMqGtrC0ZhOGA7MB
f4TX2BEbjXA2xx6t62jkUM8z4KLLMHWld3GdZxYWUJnZgqp+vfPpCGVUby1dXrHW
BqQXFUEJZiqVqWZcCDmBv4478DZqrdXRUT+RUka/a9r4jk0RyU0+x14XLYT6YEO4
H4Ewd1UcL/ReYSzcsrS1UilVsuiGl+Qs2jR2ID8IMQcCRJSbgmyjCPaT7FLFRbJI
obFPXds0EYpsLHHHs/hBH3iiRnJE7wkOoVeJtnY/A+Dn9XNHAf+maM8zBCPkO7nL
0z5aAwWkWBnxDqOKkH784bQtCUt+FaSJIWtcEggqiibRv/dnF7bDDrXj0S8XaXAP
2uBgUKirf78T8zQebhX9RQcNQU5yTAXWSQ6snptNbzLBW6NAZ+SCSnODCYKYMmKZ
fMcr70jldsnzhcvDcnoS1Dj0I6jMX19y/HEA2ESvth5rTmX/i5HLjVHYqbgcBs2P
Py5KWK9yhwAxtMS8liWeqc0NHqlR/SLmf685vpQuYry2LZHP949OSFXrOjW6U6Cr
GGyYZfRGfutZMhQtmPTAVLZCvgivYIlGgsxxYj0f5NU2bWlL4JYeP8d38hEMQNN5
ZxvQfkro8JkjKrzbSL7WJaTwyKc2NgGelgQI9DGpoeHS81sRFn66FX6P9jO1avAo
y/UmuPsgSaf2+1NzpowvSv39twvbGub0QDmCwngUODpra5HrLHxpzFOA6peU5R3n
5g+UfKp2rWeuilwsmPnJj5zf4RjjShcNmCO83Igs0ielPeGp0Y9nFb4Oxugt49ps
/TiFLCPcqwUClfl9pHH3D+deiryUL8NKodx0okZJ+PVOEEuY1szy1u+LqIOauy2y
gSWYnBJ0ZrEekiQtWkNHuF3GZnluDxS1HL20XZQ7JB+H/cjvORf/wEZgzXRIfENR
P83yqKlJ1fRriC93CIHj88cMoSh/7naAR2XYQ/KJKnGbl5G2B2XNCypUmx36fjdE
Arr4ebzOWRlJnqTnOb2SCC3lHVvfuaIee7rIbhc0OuRqAR7oLmcUcGm66NZ9vPvf
OoBlBrsZsB9kRojFitUXuTqijtflbENFl8QOQ70OQ/ZIDff6RmhgaOf/YgW4F9+3
TuXoHak8POrOaR1Gr8ANUncu3k7u8V6cRHIp1jCSQJ0JGyYeDhgAsBzcFzbhutDN
GPzKwGA3EMsJ1FA6LJmAtgwGsE8QLJSA1wx30Z7ZtX1hEv886fJAJ1b1xrdlsnix
dLZUFkkKvkAbDStnE+6vOsV3n7IJijw6CN5m5KdqjMvdPHd0riVm6jsYj/fq8LgL
9tqg36mCrNArA1/WERJZyCbI+igFhBkweYetlPJBEcvzQMSgVHmZa77OwAtrGmKq
Qy97MdZ4TbzSXkx9TdG2dFco4/311bAeaWWylP87evaMirl9FrYOQwga/bp7S9tJ
eQyPQpu0FsXRl2uuId5OqDCTezDLVq4Uiz2SJ6wW8IIKG55sxz6aT1KfS4Mgx95R
pscYKVwgTRhvnPxpt29o1fr61UPMOLTKzAMwrAq21Ys8l9QvHPXiX27wr9wfDEtB
KRo2c72ikWvBb6vO5nwePAtUrrLC6gk3z9OXs+rDp1DOVeLsy+xq2S1L1SHN0/Yv
eQZsAkwLEnt9hytPma1WSoPTcvhTOUGVvqVrSlfhNo79qbhOyCs8lZ8mFk2bO5/6
UjtTKpPc8D6IiCRWk+RgavEXgsZ5GTk7XuaIgTElsirvroueKEs/V6mvb6jAHeNZ
kkgVGm4LNq3MdWwvDsR1sXbfS2i/jSegJSzQ/kqf62no42X2B7FmsEZBpCAFBz/9
pTGYDD3XpQYKvEKzIhMOKZNZGyrNnqOVYPZsa45JnsHSE8U0QVr3rRFGWAj89d4g
AKGFkiLyl8HWHSpnujl0uw9WsMIRKWE/bheVVHNf6kpCFZbNiaeWLrEv+DXjNs1w
IyQDJSNhONUDeCZnW+fKKkavkuooE71VogWvRIMltpWMME7hSK2pz59qx3OrIGLx
OnC7jAQKd/nYCDgabGQBl+jAmYeKmdFaJjItCsmOAJ3nNWBgPigrUob2CjJ6rtle
csqkmTgv2KU9UUTXvNEMwofPAzMe8K6nrXYoXev1oUx21hEoJ4h1xK2ywWtKpLUW
B798vCY1PtIfDg6kozKq5XOXaeiuHZ6e/6nFIDDHSJ+9spG2niGzAJe6wGImhnru
gqDJ8deP9eP8pU2YNLMeruNj5EV/Lhvxd9P85DWzx+UB1pXIWedkorb6+XgdP6EV
1trr/vJXFUPvd0HZcEw2gjIu0MAoP0O6fEh/dS97ZGxXPKN6/7pHpDIFqRGmy8UO
sxyIqBHzGPnOonvGV7LCyyPBX+07LD0pu2YUiwUBCdVQx1drcytINTxHljjuk5Qc
l5XwZrZaVbv1bszMms5isxQKbrcZ3y7OcbuL6ry509v7orHJg/14rHeE0ErPFW/r
eiWFXM4DyopARK43Ki1/aVaHNySkhzVTZttUPXkeN6PxgZeqkivNEfOeEkkCx0Pq
CN4AuKqwBjEvRJ37HkUHqcBNmmyLeTUOndZeEb+riiQlbGRv/fWn+hrnR78t8xwC
meM7aXlP1KWJ6DzLJNZRiwuqDBBG31Z7xkd1c52wGBEsxk5neDmc8712Brk3QE7D
Nq0XrKU9gL/0g3eVILNlAM0duEIcaIGUy/1kh8UhrRTQlJpU2tujnUSpDmYPWd+N
WEb7xwhKKBDURs5G1lWhTS+Uh+AJsBKaaO8WdstYRxsNzh5agHAwp6xrGS9+Fc3M
LuThN1mX05xebY2xCzXz59B5CdBUTkrkQ3lM8F2IbkPWpPZl50Oi7irNg8WM7LrF
Q+wTpfi2WdMXhU4qujYrXvy8G927XpqnvodrRUNN8XwD2qNxgk/DVBx/yrkYo3cQ
W5maGklDEHG3poQODzm/98Aaa96VbFQKr7STPjUTwl4kAFj6cGWECnTFe5p8QLqr
Uj3OQK/9qvG8TIhoBWVSqqiF/aStwKgb+Z4J/qoknShXCgHd0DFPuRFwTMbvDzcA
tdCZLUq/U49G7xCXFiuQjBlKffIK6Mw+WH/Q6nURwsosgr+UVL15ItiBXpp/QSlV
3TYffp4GzdHlrWcAfwFkFg==
`pragma protect end_protected
