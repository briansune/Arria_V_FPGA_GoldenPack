// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:42 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fqvfDkwaKHgyuN0EgnhBX59WFylVJdNKd5OV9R3bprK8LvkrfgDJpkghTam/g1Fk
2aTrr0RuhiLS+Eq7LfD6SBFahB+uBSq0B2d/rVDkIlsPSZSOUkJh49Zggv5Ybs8Q
PEFv9e2h+X0/rxCxkT3cW85q4l75pi+9WerC/opRdLo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
ud/qTWq5BHCC0rahrSHt9JFoSu9+2n10bL3MPdSz1U1+ymebI27gxkxncSbGSwbV
75Wyw0vQtrEJh8fQ/HuxrZuKlnPTFtXknFP/W7NFzN6iaJ09mMgCO8k7UvFKuexU
rOfOUbhuh9eILCjsO+YflvEV0CQY8zRN20wXsjIG+lLBUVcucU0ZFsP740pkNAwe
Q2ykTf3EdDFSRksKI+ULRg43iMImsGg04RG76GUQxnLZAqTLK5hITZ8fCZHC5gaq
xC8FX58px1hrUBLsQyibAash3lcF7fye2t6ogfgOih5LZ07a3wqICkJEjFww5dFm
X+Jd1l70suqYMzTyC903U1rVfWo+/KdSGM9or+JuxZuWBFNfW6/wcSM0tj19QHQo
P/Du90h0gS5SBPV+aU0x0hEOqol/qDR+gzSlWm92G/uuoVWgBkTT9W0AiufHnAvK
skSH9bx8iXugEd/KAAefUSgRLnn0o20kHG0UODuWtzTVTxU6vksKR8lYMtkuG1NI
l2nXCnMzTUEiMZy7PLLiyIcel6Y61CHPoxFFIsxjLNhn3tVzVtDigch9FOKAIPIh
khzgfknCARXFkIYmb0/jVSAXPSpgz10eGeZ+NIbdkGDcXNXoRC9ufh5eIXAiJ6FB
fvo8FnV24QyJK6jKekPPPMmqwCChyMACiJab8dmaV4ll5MRpWbB10GiUAUgNosrX
X1r6GYMuyTd8gwE9WvdEy9hxExR+d/vOOXk8DsIoTU/v96PAE8LlTdLpxYfAksqO
34QXLVyz1N3l9Zjt6kquXx+2L1LyQG8kfnQwgPSscQoCkYXQYMlzVoQrHHOIuubc
uvkbzB1Fb+A0oRIl1dNPbq5HPFTs52mGDcmRo4sLKHS39gKb3sIToo0A1SuuhzrR
FaOgM1NvxhCE0myZiysA1FYlBqZLdOX5Hz4w0XbryywVtRWQoHJDZtCdUUgIbMIP
QZpBXxWe+t6biWpOfY5zlJ/B7Q1jG5JYVjTMJT5qSAkOY+ldDCKyeAaClvPJ68Io
NxbXz4WnR6XK3BphCXBuCBxQahp60sDyE2OFpCRi6/Ebd+ACq3Y1b/yk+c6eBo8o
WOGmtA+XRphvjcEmybTYgly/WREzybXIYlDVfHsj+jMpnbufejsbXBWDINmHu3sB
eDSxxShvfRdOpKxif1eNgw3H8633IOTvdqNKH0FMVGNQfNBjbfJqrFbGaI0NkfZQ
qGVeOxH7zt2HTvO7gCVlVstqCaEFgBjMgybJ9LIae01Ead7Gjr6HAKRnhySepe10
wRdskY+uGDpa9nVofpNmICDHSoZiVqWRHgWKu11r9+0zy8rtR9VEA4+SFsoGdFsK
NOWrPQeLg1JgWxELrRCIpXVW4iLieFtAUXBf9LTajJPb8VLNvo9LxeIT7x76Ky+2
Q5U8uQvWbRpBmcQn6JpcBE++pYVyplj0KGpsBByK8nJ9sNI+ahkaS1CEQ04TZSS3
k7/cArfm1Im4tukwpblecKHbPvBkyP8wsItEmpjKoGPQekaeTKGxERS8G+x/x8fE
IKkf0PYmeh7k+ZNjTds/08JRciXG2ezvDn2+tHDu/Ri8fuX1XoNeAr+wshrkqDWB
fps4a7RNgaQIBaG4lQ5WJBt8tmvsNA9K3EPZa/9luCpg7NjAA5wEC3LekftGb2UV
yl0joMAaf8oLIfjnopSInLtr9Ff64w3tB3h/b+g39mX36+UvRx2xRIh82BV2O+ww
7YzeWsGnhm62eKYeAgCZswr28aaaz3T6Aov6AY83udddTQeL7cWCMolYNZOXS8Al
FAd0varoNJi1dFivXlHulN7e9DzQgzA6BibU2lnrMgVYnePFewEFWr3ZP0NvpTPH
gWiTnsA6jSP4pqYTs1COSbb5yuPr/E+5OBhsKxA+D25opPSH9TaCxmeWEuTp5sF7
WFS4BmoHgenH2FqHp4KGvfXPr7DEJPBxPDluz3KhSBtjhXoQoMVKFxghMMVP0PP2
o3cRF6a8ege1riyTSMcZzK44lfoIR+4XJRRjnTQzk0TP4/SSFGb+C/hgJltHT9Xy
zn4Ggy0nGJMjesXWYfoBuOtBVQTQA28RA+NNuh+lCAHScwD3Ux7Vq9qFqajBkAas
ms4pOaxOxuOAEksmMajbyxCYebrRAmO5cdhxvaXavjno+hBKFVhRWnGGAp9YXtLW
oPc3NI6tazMXo474HBSb1XFIzLI6X1lgcrzvbtd00BgqX1kjNrJAGHI9eGc5Vlyf
DxymnK3pMNE8StFLN9tIpU1JLFQ7eW+0qn9Oftg38dmVwtUNdOg+TWr5jG+6rjIZ
t00G4z/jhtVBgoujhTm/Dl5Yx57Eq3ApEYdb6UDx+DH4Ez2zP+gDtO8S9ys/5vv6
1LRtt7Ow05DVU59yBaXCEGUKc/lZ9Q/UXAKcH/WMQuBG4sj8welrvaNiLuw0j8ZG
o5b+bva513yd2a/+5Ki2xVjT+sDWsLm9zBPxa/JCMe7jK0uo5aTrtgeyGDQsDoho
Fpyvromqb1jpkQ1+2V4PeAVikK2DDLqJWSngNlhAMi4wPEXtcYatxN92QHOV3GwW
Cma9N6SZsdNTn+2TBDebj2UJketYz/k93QPucHxKX9A3HUMmBGiK6EkDh/6T6VEP
7ZK2nuuacGQQ0EiIXkeMhhu+JDQTsM6DSR6qEOuGdpzlBSu+RRJuQRCHUoBM/ZNy
l+hhECA7jfwHR0iCF3W7a7RViyUtqpcfk7+MIZxeSdKsqg9nGBPIiFAzYTE4ALsO
5JpArGYKjOL4tKXPvKc5O07Izq7AjUNgBs8KaXtDd4Ffg2PqaSjLWywldKktaIBA
3KUnMo+P0p/ke9bQVL3kcusEvcWG9mBJ7ciJSfa1ZxUlBQhhD8737NPK42efSrqy
kzuciXjxIsuqqDq0rDlGTJvZCC0hGjEHgEhzrxXDRliqbN3aG2i6XZNXnwE3Ohvo
0jzUMfbhRdHDNqpkJnBwujt53VHE0X4Ht4x8gaw8ztNpkw+CZC5zDKJIpFg1c7eb
9M5Ao8QBFR45hXOvEK3mo1YAV9opFRu8wirUu9Crmqa5OfqRoRqCP/+se6qXnpJF
wRDCQOFvhaNqwGuxJF6yQLi2Jd/ijyAcjulpZn4xflsx5cDbEZddNoRNDzUiuPdA
oUiP2RB1+s/vjdslIvDvcBmostzYhSyzRohdW5+bI/4zQTS2riYAC5KYyt1KCfFx
wmP8pkNZnKebkSm6FWKDsaKj7ySK/wXyF+6hqM1Sf9jAku4JeoiQhyTK/skMFlIn
IcvRhiGeYDGjuN9CpaB9RWaUZoqbxECDZfMMSfEuRf/lfC4dpf9BJFXGTifU9jcd
PWHvZ342SYC8TlRgLi9ytty8pExH55b62uiI2iB0L30UDdY7MH0Roe7cbNErF/v8
LUtS+SOQZNs6714leFr3CwVOzKGZ5JtDLStcwLCcl/Z8aw5GqwNaX+XPLEKR6tj7
yJdWnMtjLWSIWphDwClkc5tvpNiQ9RFBe9sRxVS0niWaUEtpriiK4AKA9Fok8Y74
PndUoCm4QjJY6fYrexjQiX80DfmueCi6nzhzV9Z1jMUHYtJaqj9kor0UllgcGC/M
p30mjwM3iILg+y4MgvEE3UTItpRsNldznHNtvGUR9auaY6a+GAxbNsxd2fVdfbe2
9k/f+prmYfeP2wwr9hl7ywpqliMcZG0JQrI9bwJwnnVjw0PihRqR1OOYrujbuV3D
+lKu79k0B+34Jm6MvsyB8NsPR0U+XGHwgex4riGOVcTqlsktxgNBnmNw6pZ5ACQD
GqRGUICsaMD7+VSwGsmoAfXONlzux8fNrpX6EkavbuqE5o5ZBao0MXQ5DwxLKHUx
eqKZLerjKILPjzEx4ZbJEQ+6XOu1agH6lCDB77qQXLb2xO5vG3sTpcUaH5yEZKrH
mYLpxNUK2aFHyScBWUqA+pjOyuBmR9jT7Y1+Hl2fig02Z2UY2vCPYN2kFT7bOXlS
qUMZBd+PDr6a9EiuA7wTZwwI+LvAjcDCklcCJbaTtPrAdheD7KhxWUXG+b4L2q6p
mcu3DyqQNEoVJoZYRgWIpuqZuu9DFoxZ7v2W15Hz22iRfRwE7VqTfw3SAB64FtLZ
Kg0MMosFQ5Y202JyOtNpMm2XcODLxOAAfTSgUP2qVQNZQu8GECZ5GfPCV3X0ppTr
5kY1q9l2q//8I8DN0aqg90JpbKu9LY+zLzXH1BaSMI1nAskjT4Ui9W/K+/kPDRel
1aFQpaq1TCuldH5gNt5R9dyaReY3aCPS4In8qsEUj4Cs81Q7po/Oljo5GuMcgoWq
4IdItwUrJZZTq6hAmrEBaakgPouEQTW4lcOda1URITtZqzgytTEch9JsIAEC2bcm
v+lyGXFIMujCwRpsbLmCKcVr0eY5WlIajrShobClQZo4Fry3kH/QaMsZ7dtSYQco
gH8mHmr/hOCliTopW+VNAKhpCTpR8MLklx4Sh0R2Dmy0wT75evwVjDbI6Bs6ZPoc
xW9ASYSAtxo16Uhn7Okj0aAYMJkC44xLzuve9cZ2QtyczjEQFbOhzZzYo4JuVXQw
M8wfDZ8CO+2YV5pQTtbSsvJhPQRPAinGbRSHNH1KhAKw31V6ht/no7XMiRQEBy46
DqiiqcWhKQPyXPL+z1w/5BFfA17rrXhu34dH2R0klFsHWO79jPCvfG6Rh1DL4NwK
J0IHbwQg+aCVQD9CNYg6Q7hxP9TRHMFR02Yc7D/n17K/LhUzoHOa+XDPJpllePNF
BOf8AZSVCJah8KNHy/dDNe1AsupWb2sO7QzH2wvXAa0rfUrRcEG6Tjjfm0s/M4tc
YHKYBClIzzEWs6eyHuCqPErOs48Y/HfyN2dCyGk/rwF590C56WmEMkJ5SVmy9NVR
T0GIX9my2K6+ZLeqHzk0WPNJnATnMksoP4GNtPqng5G+fXfsrLcLTl282pe14Zfs
ghZbsnbmTBlSBDzi4iJbYFQUVnSmsC63wPtK+POmZGY+Q+xPA7RTf7BAVtFlTbHv
JabKQO/pWA50epvIis4oO4KhOBH2v8YtWS+ETaZbvwIJh9YoLpdQjQqBag3F5LBV
mKgMo8soPCZHVzSpBEW7kGE07WTDgx0mnN2K6MI7BAs/EEpfxuzzXLy11SipwdRg
ll+iQu0ZS1HYN2wN2Nz0DWrOIJ6iHMn37VsDUsCNVikQ4c0KnRl42Ic4CN/1awmY
vKRAykPZnz5IoFrZ4QDVcsuZn+KFm6KaO9/4s/bOjk0ynaNHR2V4tucvU9FLP4UH
yjeh25EGVyKJTsIbSoRAwKGrdyBhMPsvG0P//rJP9SxMHxvvXKT8Nl5HFrcpH3Ab
bTPY12/PPXKkJlWjZz+zAI+BZKid1TbXrXVSFBZaAOHiy7s7fk629hHLSyYmbkPn
tXnrmaXpO1KxyOeqnRU0WVJ37FlE7xOYyrBbY5TJpv15Qy8tiX1tEvWiPK2W4HbE
qvMYG/cI9zNPheApyb5cvAF51Pq9tA3QXPNm50D0qjg1Gwzhk9cIi6wSZ2f267AX
Ah3EwLyA2nX2/4S1O9KXHYuTrmIjnY3k9w5GVcyZWHEJyh9pnDEf5NGVDM7pcBA1
/iuZL83eYhgJ25aBnzVbTtLD4B4CR3kqyEddnHlZKDnLsfGBZAUeuwgbq/10MwJq
O1dsj/5OXzE+reG00kIrDM4PMB9YScB8z/Ab7JBSN3oSirtKwWUl7NXCY745ovSh
FyLP8iuSoJnt/T1Xbw8q+bBnn3ZSQU1kgXrH7Vslke6S++twXOGZKNO6xPpumOuM
t9HFPeXrkxu1T61OFHcvRYuLK0nCN8q3jUBVr8nakQTHzKakk8UG3m3K9PyNaO8M
YOLH3qspc5+yBKMQoe5K+9awreOlo2e/7fO8feYTiggHkiCAP7IkMZR+OncHDbc4
7amH8JmoFiHN0MOYiVSB8DM45FG6qNyE7eMrzC5awqy6djXRyxRpg8GpJlIy4tri
tWknBpkxx2+BYmo5N1FA9+12LkCVwPptziAh5WReSo5x6o0FW7IHuHD1lkNurqll
HasMQtyZLOVDr68REoqpJM4XC6aeW4W+HCkro2QGvmcVVRre/L2YiyThlocKTpzP
B04W9cdlAgf468aO6ZmLrwRVoTUTUO18QXe0rBwTcGJOgZCz+W/wnl+P4emUkvBt
9YfcV/UJQIkZdhprD0hFzZNng9y3qZFu3z6dwjYUAS9gP6RMPaUyBLyuXE7Zkvbr
MFuSsoORFIBcv2v9B0XGn9GNu/x3RfcEphW/KYJeOWURdr3QDWcHb7nuwul3EB5t
Sbq1FZN+5oy+N24Q9U76Ye5usxnlpJ85FNTNPpzZBbKLswGmm9hYFViWbZb/uv2l
CkKNQUMtlySQIfGILbrsv/rjw/TGXrKRdJIV1js/meKO405mVGSGWKms/GRd/H66
TttUtL4CWA57dSDcGx3LshCd9rFOMqxKm2kOkQzwSmrdspR35t9Sy5ZdQ17wznua
qVUbft+bqlmW8rCLYRUSbgEaMRwszLMK/yagUlUtbOIbVq+t4cMEPM4zaFviqHAs
OVTSfnuo3ZtVst/ev6sUD5E1oeOrABYR9I/EUyUDtlsX4h5PLjZBStWkuf/djS5Q
CF9Ea1/A+joVZ5kZFMnqyQAHfm1bCVH2hoq3d/WK2eCKFnHSjBjjc0tENt0+xI9P
Ku0BUyTaKdCC4VR3FRgJ9l8wOTM1HAZfmDWDle/rB8AX7xlrv/NIF6qR0WGkp4AF
snHkV3Dh3X6plJld5KD9cG8+ol+ryLrjP9ZKFUMytW7Sytl7EGUYjo0c9JbEQ1oO
1Y0Jlcl0TRGQLfiAaq6w4iL5Td2cmhpiIVg0WYRo/XjeztU4Q1Q6kTB5xCKDpe2s
kiHveR19qPw/WlXTIhaBfbM8DrozJMhmJDM1z6lgiHG5672bIyFrWGsfkgHY3omH
wdf+NQae0wborc1IlqpgzrM4NILlrLcalwPcz8O0Viuavjo5zgsksU7gDqbqoH3Q
TLJ6l2oVjMCRWwF5AUxIIZWUb0eKGi95Q3RzIzNHhdEmsISphWbeIbFpIvlAtHCI
ui634UWo2Rbkj3Vi6o0k6uQTbK/Pu6491fMrM4ceNUOmOKQMh1zadMquNFdnFZzs
QxIQwHZfzJsGO3oMwCwpLST9XdJ7NP/08t5zkCrvEi/BTKh043WX3B1MQ5xc4IVw
YOlYpzxVpJ/NOdV5reP9RXKKqnHzoAYMEJCurhmwAtOneLOdgtn6GQC0XxRl9W3K
IVrVdbMBnymj2yZixvgh9onuy5b+HwsfXLqqGimiTwoptZks00CrTr6DRgkMeHsE
BBqJzymVjwMthqPFmHRpivQY30k28Xjg7YT8QGBlX18iRSWg7Bx5fQbL0W/5UchC
0a8AoV4E/a8WyYQfn5NNvM0LY3slXHcjs1nlgxYMTRkXWs8vpdVCnlWh7FNg9pd3
rpHrOnd4P1Ok72O0W9/QF3/mfupUESJND2BRFMRCk38Ft/YXMHBQg5nRRHwBDzqi
O7AYFRMehcmSImc4eD8ermJ/tV6qQML5BVyYsQxWYtXD4z+7XA0wdbFuXZwhl/VY
gN1zrUWkjZolPe+KFXO86+hqLutq/OOBvYbyjFH8md7VBX3ZmIfByvBB8hHcrFFW
54F3yPoEk7U+9gk1U/HkY9jrr7l+AZgsS5gtqWyUETf1OrAq3pQ1NeHtmdSt6L0Z
Gejv4/NgKfsAnInsKl5E1sSoDHXjgX20LQUG60enkj75Jxmg/fepZtwHJTLk9z56
BlZA4t2G61i24kck51wo7Y4nbl0Fl3wMbw881kB1KGZkpDhqWdVBe8Vu3DtiJToE
laxwi2Bde0LscXCXpR+MzcqyrFcL2Ak6yjA8QMQ5q5FCE5AGBII1Dor1yQXhij6V
Z04FMpZUNTODC0jmKz+LZ9uCIT6pt9PIIMJFomTSanjNqvzvJLf58R28eAxsks6C
XJRlG7cMEueOJ4B4gMlUt4+H4vwtorTIWXoJt2jcVACRiC3yjHz+Zq9OgBl83wsR
FYhBIMbsSUeYx02xfsxk6yYgZ68ufZV96xLZpkIKMBemC7voEIbKku8Gjh1qbrp6
3Vxen23voqiZXAmY6/ZFtCxTn3415Ix2LrwvsgxdE7wAVdOGxbzpIQIA+HbYl/TP
8s8w7o9fsKiPtyX5NlMlHf4Pr35caJUE8i7BTtXRv8dPQlwCIx/vj4aUGnwB4dxH
bWK4BoVynYuv4n5+ifz5eMUxwRmQJtfh9w8pGZIspGev3CQuZIbN4Y0sl8eWiej4
P5/uwJyhyAz36jo9cMwvRGJpzmlBWGzkGw7B//ulmsxkqc/eSIWg+Tm+5EcNVUDi
S4UZhCUypXgiBYBVGDAJ74qhScOThyZ0B4/I0zHbjOuYdYh7peO0bcujOfSJaZb6
OPfNBPcirzEtFe8cPLprQmN4NkRv4QODTCwfH9DHFKrwlaFYWKcujSLhPRD1wnqu
5cBEt7Qh8iDTYWN4hp95U9YmUW1A/07MWajXrdU1xa9xXCrMpKFZEzImzffB9V8M
hsN6fUM4sinmmTzFxi6xlw==
`pragma protect end_protected
