// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:25:48 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EoAYAW1TT8XVGD0Bb3QEkjqdqwASwhrgYrdOHTIOco8ki6o0+VNetbLSAMgHDxBS
MeZVb3B+GsbqfCaIgktlDaZBU5EnKOYrCdqEln1fBMq9V9I45eWdJ6X/SfcBwYUd
PWeyH91ew9gQKcTA/8d/IP/kzBDoeW0fh+/5ijyVOic=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24960)
J2wY9OuPBY99Nwl/w4fZZZZq1bt4PtScJ8cjsQqlzkFBxIx6z7dJjw/btMt0J1jX
JzFznCa+ywqZjAp0TMCFU7dQXjnssAr6GatQc+pQUhXZIrin+H2YxDzEBpRw3x5m
0KhYmCeMiXZ38MhtBKs7rRNvlhgvB1dAmjwRQgB9GlTuOrqKv/MbQ+m6P7+kk1dU
tFW8Q/IPxp5ff7k+1UEPceVUJsMdMHGUjUS8EKkIjj8t+3CS3dSzpsUIk/jREDD/
H3QzOD71VxLhVwscKWrbFutxC+wvEoFAD7WApsIKeB6WiYbafniMousu0CrW04p9
JQyF3m9QZlnfHTbWEHHnKB/kjlKJxI/ZLglJMiooi4ifLPaW79CRn/DA+ZINuEu9
RPqtu6xbCkyL07tGkHSYks7HCVtVR7XetgW7Bu4psK6nKvQa1vjqpcg2l+QFRd5l
X1V+2c0eysro6dPxjkwaDe/cRbnxgYQYMQGb7w1WcDIR8E/GD3xRCPvp+098vWz+
+LyATrIPAahDt1BdTtTGFvzyhhi46Y3hpfmWp6ggaxkqAyHoJ9tJEUglhYna1RUj
OSEpWPd56N9NjMyh5pSXxCGsc3lrFwXfZJ66n0OzSy7lDnHPHhg0vrDpJG1Qqzga
Zvb/1Zmh3XP6L8TN7H4HIVGgKpINqRk5EIiTItqpty8vD0FXPw3rDoIKQ4LHom6D
hiwP3Jj1/1V8Y3lJSbRf6MtAJ2D0cxTIxvuHjrELme9r87R7H+vbLerrwioafbye
TiBaZ6MkwmXdlBepcBqqChNjFnXmiYRfQ7eNhcQG7/aP38IyxN9f96/BBNKZLTYH
2ZajA2i3hp1UADLbln9WNkGH0t2FFGxyhcpGZ6NcjRoPGgYYoy7+9MTwb0Vos24l
R0iLnJG5IUIwyp/kskF+FiYkoDjcqRbYXs4NU+yu5aPt4nopyfHNQJ16aH88buQR
RqSPYdKuGqvzBzc7U3kPRX/bO8XMbUFB5/wLs+VhNs/0RMJPoI54IN9n7aaINv01
42l8YmHBvErzYTW2M5KNgUXfbrrg5UPJKGkybXp+Y9Q4zVjGydonXo3IN9cx/Va6
S6TRbPsQVZTOCh08+Cgitw1rTZrE972wQt/Yd+5f7qX0SYukjILcWoOzmQyR5Nlc
byr1dj1fELpsPiQpZj0xibo4901po6b+GtT7c748OEk+7QPrnfcPbW9StGL7xblT
HPbx6ttQq2Ywsm5nWAg1bG3NwMUxHWihcm+IeOLx9fmCtv37O3j5nluBRCdFGA9L
aO+YFYzc/11+EB7FqsThamAbcFvvLiVhLCCOwIsZoP2c0RKAW3b7EABCIoKK8M/R
5aN7MWyBS/B8wqqRB3708rmQT0efWym9n9Md1FbErRqZlAFdid5EleYJL/dbXPDM
xn803IVsFfaVyIDN1iRKCU+A7pP3HNerMpA6k5PlqNPERISosxgypHMooj6ZhdeM
Zve6Ur9QZ8futQagVxKeRqPXGQ6RFabT6qZJX2D2HrnQTcPds5ZKAjsR7Yu93W0v
Z4WJ6kPlbDS8cb1xFAxqY8ylzXI8OISFOTRghs2/r81VG+0syNFU8+wBRXxAPWoY
TS3L0cKzfgE+AW+89voBKW1D25DO/MULKSHPs+KL8C8FDhHXBsWGZooNCV97Qt9p
U0HRBsXaaRXYnV0vdiiQuyf9BKAO9cHTq7o5esIekzrcN1n1gVRQL23fVUBJy+u0
reRDjhV1AoULGkDiMA/d5oFhDNx/oED9R6obOuJcGyCXiygYN32SRwFa/cTZfhGo
asmS1sX0yAEh2xC0/e542SItEUOvP958WYVqZfRheJI8m/dPgkZu76nxbsTbIOL5
IZ9lkxdcyOQcawDk0ZUC/RijoH1cC0Qt0YuE5S335L4DchfQ/Hz8Sni9cSL6Y5ii
8QhGk7uBWo7cwxxjX1NwpAXgnzBN+yO71KpUs60M8NZwvtiL39VkrEcYojIl0raA
FSMQjXLYCeg36VFuJz/p2UUfkKYaKozN59eg+Qc9nhSxGBMZ6SkjYOb2cFsjqWcQ
RPfhdODpUzKFyN/gjEEKqqDcLqnYuzw0CRllJN8JVhUTXvdrKN1D+v3I4O4a90aU
+CQs4p0EidW66cqLTni5nN5Ui+Qmd/eZRTHenAez2vw1Z6XjaQ+00gi1qWhxcoCO
7MarRHAElaCF+fqANNIzOPnZmje08NbQIJmn0uFwF2dFGyVikkVYZqqhdY1LFnyO
A0Rx1sGH8hkU3TOxWGHnvDij7/NMUzs9Neuq6FhTFc0E/MFjWdA5xyxSPxQXN8hU
XM5TXQd3YWzEFASK+Fu7QUKISqOyzaaWkbX8X8CKYlnKDP7O0XumvtUdvDE4qkDT
DkJf5jNUvWH/xZiU4z3GGq1bGyr9nQqwIoy16hQjT67D9DzyFaCFYkiva+KaUgeS
UwytiOkxGMSoVyX1Zczzfzi2cGgPvxtUx0jmTO+vAw76PNwkHfiheB/+pZdN0T9x
5Z6ufaPCTK31n2k0xZ32iIV7KcP7SlN2MbC5Wpe9y8Ez+hHitU6bmbDLhb1yyAQZ
aS1qJ06hQj/HXjX0fvifkxfsu26ef8EQU1Gq4P6HcUP+eV+3J1wsGOaTw8WVI+Ad
bbkqlPqunBAMaEGIkAoNW1D4YJR5PwR3bTIVfsQF6hYAwwzwfOiJVPCY4yqgT2kw
hoWO81dyop1ZgJxQjntvvl1NhJMmtPziqRxBh4ay9ULbDJz/0sA+Gbv5FISa5vZW
KF0HrKtPAR1KxQua8rO4i+OHtdkXFQFHbSmjKso0Gh1uFuKJun2xB1wB8uhS32HI
tssl6yzk6PLEn8DJ6Isvib3Jf6qB6DFldNK65uFktzQKdE2bjC7kKAslIryI1m7v
n8KmNdfUON+i4PFUSSJHoWE8C9jBHJqhTsWfj2FoGRRf/5eIamFoqz4IsTaHqOu5
IQXLVSsCsFWxgFZtuNX9K82M24Ia5VwKb44zdY7MfYNyX4kahfqumgN3VSr7xwRz
UhoOcBM/T9ee14lvs1vws5khzq3Y2tqOCw7Q/q1wQmvi9tUoZED+JSfVNvIvBXDW
UdjaZ51iGPI35pk03kIVqmw7A+8a8gGqmWi1Zb6Zn33jqqWoVzj7YXdm/HhK1xff
4p3UhgVj3Rk5AMlF/bbqt9K2nUGUMfGe/yGbL+m2ydTt6jf57AqyFW6R/hvVcpOR
gojqttNH5AaOKCmCr7Lu+e2YTlRd4GF8Q0XXo3NqPU6O9LETqljtclKstVYFDoMO
esUjDwwPhVT5uH2/sQO+KR/1vgBGeoZ/IP+L+H5RMvc/ATyQXUfHQy8EMRGfeF8W
MKu2Tcfc75jPgmuvb1n0f6ZY/B3frgJFFgxd47OcxF3MoM5PdeHR7MKd3+utE1MU
155JC+jOMG6ecGxJVYqLmkjxfKNouOCt6NkHA5Rjh6UZ33mcRpqYvAdZ1T8xBrCg
cuYpofxJpteIzas6z+OkRokfBw9QJvM1tyuaPbiqg9wVnp6m7D4tgKZbdl+yVydg
STjFHepUH45bmFc3FzqN2D2eGKrMt26tB231f9sOlrvflJrN5qg+sh3nrFgGjdgd
vMqiigl4o0m6Jd2w/3iMmoVTRsQOJ+y5EpT0pZAkcIXX7JFvgiRdV85nJOrWup6u
/R0/OG1JaZSGyImy+mN/lHL6IkFvVZoPfBSEClr/oA3BWSYgZ8Xv8Wg++X85Ennk
/F+Rux7B00tvhhDgxNZbvnkV3pxxNS64LSs0B12E4FQggt4hdYiNVvSXA5mOpIt/
PaBWvxq0lZRBEh/y2EBCoZPkb1gwFidB7qmbxZ2l4qkrdnMJLxym3RcjHLdGCfyC
XkFx0bXfz8hHW1An+DmKHerepeylr5m8kNkH/QDAos3gO3G7CsJnnsNF5b1H170u
Qin+ZwACbodNHhcacJEy+u74R9KGjJknCfoUyU5GOV0/x+hcLs4EdQDNjmz4S0HW
6kyvCKsZJ/aGzOGjTQMThbQ+d+bQc1HD7hpV93H0Qh801NB3UzkZYH2oXsz0Savh
C/DrXL6o5khNhzSY01ngicAMM44sTaxD92iB5o1WKyYLmxhJBU+Kp213Gb7VZVMg
HwR7TYPV+EEy5xBww5xgbht9YZQw5lYKTstf07toijzE0MMgScA4s1YmtfyAO8F0
lHyevzQsbEQDXYWJN9/8OPcj9VDdsBEfPad4hT7bNYIAJBTG9CuPqmf4o/IjSR0w
nhsexJni6U3JZgJSEAZsbvnITz5KkwMDUVvllSswTv4o1RIepHqkAYs8ZeKcNUSd
6NHnDKEUafKmlTBBEXSsLCS2iZe5wlayl5Nr4nsU5yESzvkhEK5p0B4XSaf6WYTw
CBFuhdUmGmMLxetG6QqNw7gRpJ4ODWCcRW0i4jPlceDxuppDx0uVypA4wF8rcWw4
eInPNzf6dbbO0L8v0MFGvD9gIkMX/6bSqrpXbbT35ZepS9nSIt3cTSo7GyAAIwst
tT6RROWoJacP4AmjaduwNSslv/WJjEETpS0LsEiN/AoIW0I+qSydQpm4BFNkSjUF
BVuGpJ0YfP9Chglr3lTxGhtklQAiWz8JitXW7USKXgeQY8ncX3QQZqrMsLOZrkF4
jVZlqHuJcUW/xNPPxD06DayleqMgzxlRb5B330UYT1hzwTJ9jebnmvqaRftadNsx
C13B7UsJdX3Y3zRqt/woCrQjyzZ64X4KJbt9vYqnoymNtBHU+yMaWnLkwPrFJ9qz
UgR2ZWviY8fYb0R+nx83ATgvOrm3kOLy8Ijvz/ABVBeHnakThUKHR6i2i2QxRh7R
75Vxeer0TZaP+dLWBF4ibLf+66F3DTMOCcu450HYNnh3BrPlmdTtk6v0b6Znyo2p
4j0pKOJQmkIgxqzti2FIDN7vudSsT0jiwsoKzXjoUA0+miUxpSWDoNhoi0en49Bc
cIHSIEpbM+Hs12Hd+m+gZrM7QIsv89mYIe+YZQk04ToppazlhbYfjlvp8Yo8WrfU
5NSdfyEf6UK0WvxJjjbE1TCtOObtas77Bpzr3Yz06D1NmtH7uqKIbRFybXn04ScJ
rpFO4QLaiUEqz6GWg/dM7VMzxhEe2IOV56S7ndax4LgwdMg9UfmxhYY9sdH5dii9
5qDXcQ5hNsymFs/IAVehoOmWHM4BMkycX9c0qcbRI/r5LhYuoYOvY7r1UeSzjlyP
K/Gvg3B2EcvYCvBBr6T0QW2J4jhlD87aZz5338Gi+BgrqRzTBXjtBc/nKlt8Dl4h
SBaLLrypEoa82gdMAgZIlam5TD6mk1QoKAQd31R+vYvfsAr7AaKxpl9ZF3U3clzr
bbsQYI5nLWcNY2WFzYc3szvLnJocTSfYht/RSs+ZkXNJBMX1Aql3LIgKd6R9Zezw
vQJ5mTrfpU1+onIyp1jRaPKA4UAkSxkmkR5bU1vs1F2ILYD81PFbLm7JNPdNSak4
+ixugzkIum9ej0smkWfUzF9eQA7ogKm9EO04pP5vJh+hvbQ45EvSkceddsOHOxiJ
CKhHWCtuQjdXawkQp8Hl09xZfxv3rOylIz9RewntoE9/aMut1VOelKNcum8PsGZO
7gS6poFKzWxrhPtPk5wub6gD7mkasdCg16ZvFqjl1ggB0untkPQCE7MiwQG7RIXX
z4v0dEhQuXSr+A1858P8Y0Bs2zgqxPapDupkgjXdSh7Y8//yucksVnz/cjlr7sHT
HAis2HwD6hd8iPbAwAIg210s5p8xK184fOgZIoSEYmbOVpblMa5gJDkCz5u8z4BS
Tv0hzJHQwL39G+qSUc0q7PvwnMyyIgmK1FsJSJb2ak3+fYFBhCuJnZPKovqHFf3o
XwY4uqoIO932NZ63SFHoXTmc2wTDNBA5inJskA5GNxfnBm9uSb0+TyxmZdsSZZEv
3K2EVd2OsHUh1BZf64livW1ucvqVW2Hbg6aUM2RZ+WjfYFIDdjoerOpqSoXRsvTV
18XPFNK4r+sT54LB8hrHQ4XPpOIUIEm+xQkV3DNa2uFPI1Kbz687JtfftwEVDlpc
gwl58L+S8YXYRakwg9aARmK+FAAEtPBRsAWYCKtTYOe9CGBPQhGg4lH8eDboUPF3
zZ6xhlQX7t88VoJo31zZn/BFx2Z8B+KlLRNHfvaNzxGESfdaT5I4fpIApI2HDBBf
b0Nn0HFLUuBgqTe+S0DEGd5vhQw7xq2bUNPEPDJp7iNF/BV9gH8DOWx8RjNKlP7X
8BfCh4VThpxkqdyTzwhGhxzNbQYJTn/rBIWqmFJYhfxEjTGW2jmdY9qYvxxVGNHZ
1kkVPGSu4zdB2CQ8x9XZkP0ZOu+e56f9k5gs6GyPHsDT6ySBDfdlbjcOnmKUc48B
1HcHvGCrHfk0Roniy1t8suu5dyZP9bB5R8k02HTY80Wgs0f50lJOMaqPi7ZsKcvl
EOzRIukq2C4ZqV8sfbg5W0Bp3Qwm/C2ZQc3yDLz+e6pJAQwsIWd39peaYa5dHZF2
BxfhzQZFPGMAjIkcS1J7iKFrTlEf6m1gHeBxE82BOUW0robNCDBTWEga2GFSmzhc
dfvObSn8jzzT49PZGpwrOn/N7m+cJ6cF4h0Yf/a74RPJUeNU45aVYDgS8q4BpLaJ
k3h84kqoVf2nj432NvM9xpIOTatNn37gS4fPyi7QNPCcibT65/m5Zk4DhB8y63EE
w7+hJMQfe8Tr26Jv77D7V37rlGshd9xPwxQuM0aKWU2e/oKMo8LnMntlKod7p/6P
SFFUcxT2iaUdnKKHLXp2tDN/RbeC8vvdScsxXadovrAytqHFMtaCTajq70VIY+zW
2voCKlku1Ei9YcUwzH0StpT4DHjswBFfkN95q85BmRz9t1Gvp3eBDeCy0NR2mypz
GvlEbvQAMVyL6KMlp1v6YbGFOpgVhMEECMsGJZYJdz6LPSG+7E19SpPh4qxTNJEh
niqZBl3pMukUICSgYf1GK6EDWCgV3HNVl03XDnSyjF1IscEJAIJERH/rsh3NbUnI
k8n41d04+xegiN7OXqwoEcEYFl+CpMsgIzFNjKz6RKjNGtqezILWivVdR2P6+5r5
q/NqpYn8QWjtSEUNubUd9vuW25n2/LTIqBJqi8TaQfcglDeAgS55xhGdLG5IOprW
A91xcujhQGIe2liu0wzJ3p2YOffwFhCtAROlvnCbq1LoiJz9f1vsRf7OKHjeJgD3
7FwdXY6ZJ+kz2AXl8fPCGKHp+nay04QdPkJFsw6nDxER48S1rdgAlkm6sksaiR/B
GqFIPafhKGIQAECEKmHn5MixPBGHx8jQ87j8lP0tT+DD2nv1pN+rZorX3yx3sb0m
Qywr2N3y4oAovUBMn9oAE92kvhHfXE7VZsYn6ZUMt0GcZvxFcB9mZ0Sg0qRIa4OZ
EJ7thhCcZu7ycIEUsgE33iAGFmX2tXHJgMKLsK3nlHAsO7KZNJpHPJW2oUHS0NRv
CkBji6J7SvGAR8+71o10g+t4iJ4/tqa4m0Jk2EUl9iGnEZSibbj7L1iiK2pXom7Z
4s3qPei9IuvsffJrG3hkXYX1smrrMsumVm5nUqy0+Ekl2tT+eVfI695bP4BDmeQN
mmxsDykPkjngkv6V/jLBHTkWEBwVim/2m2qsmmHUMuJ5xF9b+Z1U29G/pyTbiNOO
8tX+6wTWpPrtwjG3Hdo3dl8KzJ0PRJFdkIAleUnLG97sSLM5HwxLkI3AACWIWPAk
g9t+5ZRVM1FR38vZhgFWHzQgf14bw9/Rz8kbm8YPdUd57DPPAHc4aN2l0Y4aKOKY
oI/oN4FhxEh22B2qHwU4r3FyUkFJZrApesptwtR4rf6BD6bhCkzdj1gwV6yWqkV1
LUJQX0Cw/sGVn5TRgYAgU+j+WSLftByaQ7ZH1KM4mvNf4UnC1Q9JcPcJ1iaK3XMf
Kz5NPMar7HeJfKO6Z2MyopN5HnpbjlcaI1WBt0lxAM3lxoSRSsLDkFfl6+wF/kSO
BYVxHHQUPI+reV67hUrCRMWd+tmckg6LaN4gUoEbb0PLJ4aGXiHjA5/DdxbYoDYk
8G690j0OgteAqTiT2WEyB69jRneUE/SY3rF8HltX1gIuHZJjD68ZCzDNqNnbr1sb
QIbwJ+nhac8FFk+QoVsTD5dloFKnSp/G6M/1pJ+F4DOzVtr/nCWY9i0SJ9swmAEi
nsFGnlnqSeGy42rXw9STcqxtmExJ2Q7gFGGxQmTeM1d05o8+7Uiv+auNM4e1fGmW
f0syP33Q9RU83vsae285lhukkYY++LCBdbBLXeZiu9C36yfKGa/xYEhMbamDM1zq
Sgwt9ME3RTDXJyCZPZi5sZspqR6leiwUbB88nY+vb3cIJpR0MoGihou69YJZrXOP
fbFOD1a8QITtY6q5AFppbuKa3lz/yMljSLwQh2su3bQ6eMNglsTUOsCHROKcyN83
Vx2zhHiHiydigdZHdY5E8QJkFAB2H5Zw5GQg/YzKVL5JDU/ZjbuAZ+beMSv0GI+n
KmGeP3EERa4/R0XCDVJrXvsHb27//KeTQr20DWu0fLWW8KY0ohxX12pR7zZSeRSl
8YGYXoolWpo8QQqZzMNSO/sfePphfHeM97fAOSDgcHTuBNmlFdUSxQOxRZuwzw1R
dt3tTRPYRKr5Z7AJgYGHBjhYb5JgA7+jnCNtFLA8L+5HBtJpb8n0juPUy24QF38s
j9oluC8I2OYEqs0L/GyMFn1v/p8zH3XmumUmRudrwylTv0z4/fI81TPNPKmgeCSO
r2Qy9/4EmQ3v44grIoJQHHS7DecAVe1YAXbKHVy5WTZqrFLtDq3t9Uu6zwk4Csfc
UDHil9N9KZpK5Uwb1GjdDm2RtOm6YzJYEF/8Ktka8LKPJ0LkrNCrXjxuWbGHcAoA
04hhT03/5XbrIy6hRqJyebQp45V+2j/A1UHszUdM8KUb/V8jNmVCkMhcn1MHFpvg
htiefkGYFtylbTqJyWEts7sHEwH1MLeg4kWQsZ0ngUH30YrCX01cuqBpiOSS+9fM
0FxKu8VKOOAocL7TnwvTuD3zbDf7wrXvY+urJNrYraAjrbbhYkbhSsNQnfrBM10i
HpcFacmjtgdyBiAcrcUavnlGVvVyrQu4ORqxqMk3QPKuyngHYQdmtqOw22WgWOio
2TpuJLbbMGfcL/oERv3AQV3HMZ1X3y8ydbsyqi0iIcVMiNR2I3uy5uASdBeTdLN0
LXryD2fAm1yINqSULvBFdYqfhyTqQHoEHuuTBy6urY/FCQr7jaR10o40Nb6XI6A5
29C7b3Co2gZt+eB24/TQcptfRDXdAY9QMdqaMr5ziH99oo6ez1CRB0aZqAaz53o8
/HZGE3hWNP3WXjVdQ2LwSz8/MTOyBOK/s89onVYSWht/UITxXZhB4D/1xsTr4xrv
ZatXINxzf9XESjd9ne6xAaWqfOXGdgJi4vdZLMo/q37as5rgdaZKfLWsEtQTAQAf
eoMbti6QYMIgzNZXWbX1z7RqyUb3dX7HSiHXrUsAU8gspgvWfS/jpV9g2FF1Gllc
Ay4KN6t92auZxNS22x9DLXqOzltT0U5wGnYknQSAauWEtwQm5nMhcj6h86E1mEIC
brylTmw+1rYAdVaZqkp3yabh41YGRv+gBtU3RZ5iCqBTAoFmblL9fKN4WBty6VRf
nQYMa7vhxTcgsLsj6TIrMbinp6sbqZB+IaYc1honuyGifaMrpA9DTRgnxxGqUCpU
nPOJP/2k+fiJ39aB6AvpLuiaQIU+1iwmM5tyZpOpsgMgB1WDycQ98TLSmb5pvYZB
lUWFjgnkyICyaRazpxtzNOo8Mnej5QOEapKtrFMju0rUve5ymEY5qqT0TQ8+/kye
OIXIF8nODYiYaVeBsM61KZTPPadNIW74UFaodrufB3fqbPTZxOo6uJgCSrLZj9HY
Dc7l/U7T9VSZS9/8h/yt2xsbkc9wQbBwuC7lZ6yDb6pH5zDAe0XmKXhvyETfF+1C
OQl73y1QLKkZC78AC91hA0ISfiU6EBD5ddhVaVnsO/1uYKzCX33K5wXlkPEI9tLY
9rVMN3nYsY+yoRPMMtiMWsUy3/za4WlETMqVqJ8ox6v2uS9uPLiaPJdiMKaOYwZE
7ASpzz9E28lO4lPjZJ7I3y3QyhKi2ut+6EEGF7CeSL9x6I++yh/Q+Ab6f+qwu+ff
qHPY2safPMo4oLN4mlKvm0H9PckW11Bmu0GtjVbMuO+IC7lBZetuYKG1BvPmTdhZ
Q/vUqfRlFY6NkCCqg13r77/6EJBRpzD/KPRL0CcktjXDDR2tIv1xqgD8a5qH2/AN
qGdP/fDziMmQAPFeqaXueY4wXak8FHFqmBnG8jj3c+vk1uEiZYSwA+Xuzx+0XIss
TjhXY/AFEoqcqCtlWZOhiLvRpKJRZYoq1lxAyhNL23vOtf2ttY6AsIbyAzgZjawv
xMHRtlzeozauHPI/G/WTtNqp9BRvxjnD+2ZweKg54hstO7HQlgo21NUt6LEw4RwJ
bha17bnN3Fvao3AdsZhLA4VjUi2eqis2J910JzTDMi+kU1+3NXCSnd5uyzMpHgcI
5I9k5Yfh4kEQDRIVbXu+X32sGTdx7NXZtoXIpAW0dBCgWJQ3QSkPgr828NBgvCG4
Gp1iwd6Ti/E1O6pTHUeYvpG4ASz5LOROjZIdI7K2PCbH0WIT94XyCUiJ5zdqSD/n
TP55BL5aUvBl5HUyqdizXc7bx9CZHFd2jRE3drt4392Fy1Lck2UKNBVkUxTm3NIf
S6SNIQsT+NKOv8T65MUu0F4AKuOgyTxjIlOcqhNefS4x7ESd1XOT2kWN0eAWIYTh
qdapr6u2SAqTEGwLN/NZUMBijeqEhqkg4SupEiGOyQggz66cuZ3fe8z8nE4wtP4X
XkwaP+PuZWe+rDkiyPGJdDPluyoLKvyopvvnDO9u3/C/D6NS4qs51wrwZVObcWbC
4O3n6rdnYYkXEyPrYJAoLnBgGf7jiRBRUy6TtkpsvvLWrMrIzOCstOA1co7wqgKk
Vgkf/5rE4p/GO8H144arwOzrSCyw3d9ynXLzluQrR64A3m8U36Jbd/iGDi6gotjw
ohG0dQZk1KtqB04MrNQGUaeL7kZGh6DqjoaeVWBqxd2z6DtLko82FtUeidhRIbx1
8RG1E32zxvz+WtEIV0YIts46I5LRfDU84tTzqTTZ2HkOEVPFbp6KfupiAwiv6Oz9
duH8/4faafNKRxpCpQ9J0Yap+uPSR04uKj5ccEMvaSbpXG4hoP3NiIQ26dO7ymMB
A8G5V6dbEAcTHiUqWESCEEp54gYnqjTigBM+3cZPGw2EXsdDSJF6NhXw8daKxFxn
HEuS0+57sGtmcdD4IyQdUKEuejA8D7m2hQx/5fEhQnYoD+2nzMh37LEsRt4nBs6x
FRo1XICyaE1Ah+OX6AyLiNcWkyDWWHfrOR/T4ZZZ+n6VwkeGZ0xyLqR1Jc5LIH0O
IJ+zr1AWqP3otoKdR8MxGTNPXs+Fo+YrsfiICtG2jJsBSj/I/yxzOfs2cS+0TZ3m
keIRKBKaf4y6VkDPuZxi9Vn+cKVN8FSXI4/BuN0DdbP24ApCxJE6FiYrsbuqjiJX
5/ahRckNr7I54EwzB66O2A/Yr0xrzv6/9z3H3AVvUT1hd86bH3TSfvzAsvzAw/+Q
foviuUB5nNcJtDPCqIq7680gAZKe6GhOsceysI0TgKjSX1/PQO/jSqI5G+MsEIbT
+Eh+bRG3M058QzHJSB6hbvhobIFTs48yy8jxUA01+qOWAD4PAd8i6AH0a+YSUm6Q
QxjW0o6ZovU/63vEA396atxDJuiLmNxFhE+KTLglnQKXIolm2y3mnPQJoCN7L/eC
D735wBoRof4qCIz+c/bStfDa29ojpxeO3Lv7kEl20S9IuKYQFZTmRMSDKoEIPvbY
kIL9d4tUu0rMdC49oi7hjc0UtM4iW66hhofClXxXuO70wUTX0vJFkoXWzKPAd7r0
njTCUbThGOlYgLTqz8adkZgPCRf2YEoJJjaAxmMCLuy3+bJXPn72cQB6jvx14SQ0
xZXjVvRRd3gn4PSahyKUS9bv/BGd65oi2xOt24lb6sI5spLbAuSAqlhlLk/j4lB6
gny3KZOWXWTrRu/4YW/D5Mw5vL6RZR85wB7XG7DK33Upx/li4SSnAdgwz35Q9kLG
PA4jW13Nrgpw8lFMwWUv4Ea/7pi3G7b/U7SsBn8n/plL6r5SNHykYL8zirkBpzpq
y3vFgYLHBXXVBdF4cN+dla6DDs7EC/Amjscw8Zye4rIx7vl+srxtBduhbiZj+vdA
sP1xn2tKt0rEX7XfabI3oV+RO9QmfybUWdlXa/UFP9z9z0g+lHDIt+EjCqY8wj+v
FQTIqPOyb3m7OR/UrCJiFKk2A6S2qAI3dxuAt36enXGABYyChFN8vyOx8DfjZGh7
Y8jaDKCaXL6dIcSGP8q2nyM5XSDQkOtDWSLRBY2e4hnSKZaYS+QeXReBhHPOxNU4
rrqgxs5d32gX63zAPAWeA9R2Kp0E5EgaWQrpv6r8aEUCPspy4BWT43Av2mIM8HEw
oI14ajNK8lHTn3oWkRseh1AAKt+jPMvV6BTzYg44yhBykNWHf6E9lXWfTjFDjije
DoiicS0Y5tFpGOWWY+2MDqrSVNAU59yWsPnsW2evI+82neNkf3SYUTgKO9KVyl2w
5/th+FLzBRmzYGMqT7P62PnS5c3xhq1AJvU1clu8dI82VvxOz45Gzi2xY4t8lYEU
zi2WQ1AYlJ3vDvS3QD2EDJ1fdLvyb+U5g6RS/HIa5dczf8Garb9/Gf3PSvBH+Ot9
DFPlv1u0hJSmRVyz7If+M8QcP7uB+dQDlxlhsD276CVCU4Sly9M7kaEywl3uDVZP
CBJNyiFtbs05V5R+VGjJL1AW28OJHA1gEGZDHwqV+1Wfa7MqqRanI5d8+OcM2ZFl
B3NhzaowDLFKaTwhFRdKhKicy7Ml5vO3vx8wdHd7uaMPEXwbE5/lgDafOteaffdO
aIOo0ItoynaCnkN+hTU8qM9D7WY1cmB/pUEI2UvfP+OKeZZEFIkKaqZmDmGj1Q8+
nU3qxQQbYUZRqs18rCU6jcnYPN0+Rc/EE2QEEJ4D2ZRN6F9Xw+swURWK2fHYUes/
1jDNYpFvJMVA0+RGmQhnUPOVOBo4LUNZfleIQi1tlhXDB2EGz80fPVzRFgv2BwEZ
6rRJD3koOFr/V9SPXOKP3Q4EfatUh/NLcHVyKINYt8FTI/Iz8ZeevjIoLAtNNGro
1PTqB7ecjQO9hA14hckeqMcOLxeHe9QrXvnE4K9imqHtf2KoWfp1yt3YLyjAYyTV
mQkhvr3zEhFEXyoBOA6T0EBE4TsHSwrKFAkJOFSHzdJU4aiBi1s+H0eNQU10MDTL
/LStaoSN9ZzXPIaZuR8CGukL2M+xoF7+oIkOKtWf1+6zJuMs7yWXW8w4QxOhiXhk
GGP6kzh0cqrYqo82G/XZH3ExNgh2Xw04sXj9wwFvhB9qmdh4mFHGYYD0Jg8aIRb9
s93asMu8prTj/kHhGjlmW+w0mIE5u8tdBvGmFQ348MSMSDi/8sdc8Ke5CTamAr/Q
/9o63a0OdhTiu00vguGL7+psnBBYnk8Zi3amBWkoKCtiFJtjqHOtMSSnOvTv85Tf
roR5DwBQO0VGBJYMP+zw6T8skLgTPJaeRrpo/dq5nONzgfZkvqoki3I8ZOx0t0Xd
uVgr7zVBh+HZR7xaDwTNTy0TXwBAfgiedV6QMdB+cuAoDQdc26+UQtkX5H7WzZpi
6D/eBMrSGtu6HOlQTtYw/FCsAhVCscjy2vxGtc7qPmtfoUZI8QUL2m23CR+4fmBC
kgQgBF8Zo6ddTy1+R97qsGBr341/VtaLnE5dSSqZVtbyc04bArOio6DAEglE5CMP
+34qdWHaWXoHnpHdWhNpdz3LMumfuHdcveVss8wrsgdJm4nvEkI81ksLwdEeBsoN
SAZkAIM9Yp+o+/Cah0fdmWq7UyWqSW4L48pDLfxXQPJgd1EsGo0F3tNIGPD/ckNH
L1gZ3KjGcPxUGTcKnAhwsxI5/5P0cLWFdMBY5hBrsQBThPyrdpZ8Djc90kPzfUJe
yrqxpBAbDd1c+1X5DGMi1M4sX85qvjap0I3Q9rVNX3/NCo1H4evEpjFtAQkMl9A0
gtBJjlX3SdrhUq67LuyL8S74emCIZIh7/pZ3N33I0/YdxHxInqq7pi55ZM8ksVhL
XpO7YPM4UdYlljIObhbXu83uAAKpE5Lrs0MdRQp9rXOpNta120ZSZOj+ujULC5/y
UQG+g+E7bZg2ie9Wpsk7fcXGWnZDp8uQyM0VRtQTCbfi2U54SJjp21GEtael4mB8
Bqs4f3Ya2Ns8SqU1BqsFrSUDeei15n1jHv95CaD80gqbXmG5U+tJk0lmkTHJzS6Y
I5aw+9Lj307orFe3bDds+xdlo/+UBZO2i1ylzp90i+tyJ3L2VP4hF8OYWzXcJsCw
WAEJn662bJeBxM18NexuGronXJascDyMtb+tbppUPCxM9unO63kt7XGHpMPZVETV
dq0Utg62NMC4IO+K5A1Mb7TA4hFrt2BAlZDTb5vfoNRpMQP9ypkYWmmYXHyHJZZG
dHZAfy44DFhIDlMVt1xDNSL8MCK1ht3RYt1IDbbhlaLQkrkaDBo1dvGdN6zJNNNH
xoMNx9Y2aTmM3LuE3IIOgji+Ne9SRlNJdlhj9yHRKb26c346icRoXPo9VPGkso/O
r5uX8wB2CvsMAWQLep3gPv2O7W8yWlqlqC9U8gtA5VssqModKS8v03iD+e4PSzsl
Katfzv2bcK0xu3jTxMncV1nWoBGsHC86U3nD9/AAaoPp1/AIvCu+UrW99O2wiRno
Okd+t/SnGkxlY9lSKI904uKQbexOpJ5yJzoK45F0dguQcgODEIFZqcVAKS0gSDjn
QXG5ImJCVfykZL2/9RZGMbFySovWHbXVx3IdnZI1qqaGkYq2TbkNCOiBTA6eWcju
CwYQOibhIC0omjv7Vv9IHrj8RGHvhcEYsBsw9wvU7PhqKMNeJu+81Fz7XNXJ/b+J
azl/qviY2gXjq5RzK9Xh0gNfAyw+0h4YNxwWww8Q6K6U9JwqHIBBW1pnEI/XXVlw
ltqu50Lhv9uPn4TQflxsQZpIMJcJFbD2Y3p/ADslSL96vpk3avx3hbONQUxYw+Mh
6qIi56vjM0ZH/xIMKp0zpB24TFNlIMGKd0H/ECSWLYTuD5EJEmsDbAF3BTdUOeCe
6h9OTatvmtlXiDp1C6tAZTAY1Vk80/ILxXb0XorB8u2wyXAusCPFZiWOpNy/9gTV
1tZNDzxpBJXxmHu9GLgtaS4L9aaP3teaNcmg6tbrN7dLIbnOqIYQ0BYsa+ANLa8Y
ZEZG8AjzksZKLcjrkgFNUGoE5wBdvjFDV9mIDqpmMzepb697HWApKdqKPyMkTX7T
KCMlVvT25euoD8WNtOTn3cvxr7D8hOq+9y9nqfPllGFfTPAjfkrshRmtjTvMdN59
TyxANztppPAOnuhSTDjpyCxD+UdFfZ3FLKNPD0n7IEa9PBJWIqtGErnW+osAYjoE
3qkhYZ6b8MgoxGySQw2xGv4pCSusPeQObFYmr3N0WXWVWJx3LcsH07QQwZzpVg+F
msdN9HSMmHc9fAKcwcOssdjk3BJlZYN1tIdxQmatYctAY2Z8bzMzQvFN6ojgA0LH
PubW1hXzwQfvZa5mEiZ0fD3bx1MhwucTie1WwQG/HrQztTLzLaMLSy5SFNYC9X4w
C3Fi9UDa+y7lQUWAvdqjnhCG7rHR22HjYgMR2txd0YHVtadsL1kdYmjcUVagCPdB
gObnD15B+hiul9ns5be+vftc4zL9HLvTYCuPU5iepWjx35PI8fFmTf+QzrZS4m17
wdUbrGs2zrSlwH3amFTdqoY3q/o2useNKZT1nnTkbE7HR4loSgpt+wfR7PIvCWeC
MtmKUHW7C7xBtO2j97zdwMDqWzeM+dmwjrWCJ0XtFykZTW8+yRWMCGwH485v5pyM
2d0AAiQVTnsvh1zXlofbzzjAb7kU8KJYJIBBS0vi8V630iU3gzUyEtBCV4jckpgz
A+5gCBInRaQ3mlsfjE6l6+5S/LwfcPH4oJh1sjssccP0riPK2fq4YwdHfsrd8ODW
2VGI2bToUl/SkNh3Pbc5bKsGDyoeN5yLD1o0p7fBKkRMTTIpKtimOsgpS0/ZvQfu
YV+BVjK8m4CVgE1a0I/ZdWtvlFcZq+lC/72B19HFgPaAYlPT3VmbmOqGh7nx0Xtk
4uwgE6KE2211J8/ECM6FYFvd5kuMyCFTXD22GP3lzHdEOP8bZ7IAXGhmPO3O3DnW
RVYkenmlRsKnrCmA3NnGnoUOuN8Abxhnp0ZmuCcFkO4QJq1AzPE0SevuVVft6FPw
FtZJg40tj+HxcsFPy6jC/JoXjck/iguPn27U3Ssp1yW0l5fTRa8ulo/lJvLiOUCh
IhUXQ17xMonkQEk1Ja3fsl+PguFjnnIXq2xHsl4JzFo2+hQuLlIuNEMc2TezbptO
YbKD0VbAH/tUxSyy4BBxJDjFlR1chLhKHo8EoSQur1TJJ7YXbh2ijpeqMpcMYYgN
jv4Z6Mm9iPJAh1n9+ln6d+j9RNMaUzIqniPmq5FMRs9Tpqn3xFfZRRhr5rebe7es
Ypf+cD6JRAHBdnlzcR/SlKqyYD8MzrnFnxVHidWOAMJssKUsRAk7puGEL1Oxvr9E
1IHJqG9/iUBMlETs5wizZDVdjuPBwNxQWcZBOZMyGBxq8HVvLXlh6oLMtk77o9op
OLElyI7USX3WWsPgCoB0UixlpwB8BjDCS7HM7LXq9T1P6PeeRDquUhWVqaMynsCd
mxFwDB9yzZIH+VD+YQo56zQL3HrjRSL9IaOa+jvZ2D55SGTxV5CoRoajlws5wKmU
RuAt6d8QFX0xBmaBpiPWyQj3jnSfMTNQi2Z2XcSnF2UwiEMt8R1TYQ/Ud6AkqZ1L
YlNUv8TR1hEBptOlP/dacu5eYvXlMgkTadDIf23sRAPfnKXe59q3IO0fyGxl2gcE
l6/8mwvw9yq2E8LL1emVzpjVH1f1Nqeb7b+OwITblDdVRjXT9yh0vd/4Dps7wZIV
yR0f0R+2ZCdGVGdsE9suaWdBZ1k2keL+mm1DUlUzc1adXg2WhZHNPoLFJUDkbc9/
dE7UnbyvC2Oi6yiMAqotsSzLD3kQ9VqFUGBLJ4+L3JM9McSvACVRu4h2lw5DiQ+2
+qtPvprBaXoWZ2oel9Vlmm7dPGZVnrsBvmi1+11fBybQns2+CpkgaIFHyTjqLNZ+
mlUkiogx+fkA1ixgBfoTQsXf+F8TZ3M/VaXtyb9bMxC3dxMR71LmdkJ5joQV3c8V
sn0MoTPLxciJo3PuSNxXfPYj9980Ma7IiiV9XFc1MwD4HJmAb/Kh9MRg7EKAjDKq
EnU2Ah4KPz+KQzFuVmq6/JLWtYIy9WjpjB1oI39sUnAaACMRd17oRJ/0PNSaU723
HPb4cPzfqBlx/gi4XfNFCgLQF3W691FikbwESKZZN6VZzsPaKizkx5bO0hDJrZ2X
a6iiYl9tnCZrySZFvisxlzEesMgxQEcYT3zAjhN5rknX5dsUEShYF7TuviZ4hNKV
/XbKcCeW12aZWGNR5KyyxAYz7mv/ESx++mGX4D5G2Jyo/WjIpYJ21/vW36J/cBBV
2uvUeqRVZsXsHvxfJ3/3RwBjC+KVMa9RPZyOtawNZOu3sTNDlIxJPOrvsRXrGoHp
opgSVlEgMFzKJJYzZV6sUR+lYopVEEpTJ6ZbDqhrCHWQYirNGXlG7Tokgcnqyvwg
7D+Wc94O3yC6GYH9Am0u5O4rBHyAkTbEPpGPC/ja32cdyabFlGDzOUF9s38i9WR+
EfBNMA28auAwN935IH1tEUf/5GbaJ1FTuI1ApU2nhEExatp64qQQqp/ommw44crL
NZ8MPF17c8JYktRoV7KeFOAl1iCUEY6dHqiunxA+/Fjw1od1MJOFGHM4cODPqTcu
z5CUJ8iZAE9baCfqXwvF7nm0q69jPKpbEpMhDoW8niKAOR7nz1Weu1e8Dv4LiSb/
6JI5VZmX5T82qsu3etIevG676Qxr6op35ha9Ui30hdPs1tCVebnEB1V66Sfd7meY
9PCveMuTk1Ep+2E7zTNSAWl7uS/Fuuo44OjPNbw8xRCRM+GsRBFdRCCCEv53UXKw
17zCosXslhG/f4nf2vMo62GbJlNNSxu7uRvnXNe7gEa8O+KyeNvrspXtTSLdKAua
aqAL9gBeqjVNAhrMlXeWliDAmyfAOGMlWa2fg9F+MAMVFCwQaHFlgN1OoXUIDBww
fam0cXxpwtsKJs9fmhlYOeOo/a8dhyjB/ontMQdRBJ9iyXMcThxQDnZu1R+iR3h3
0Cy4Y/aBvi9qSahv+f8ACto8mYhe0tpdWNV2ycjcYTbnFu/h5uhmsevhDH40XP0N
6Ho0yz5NpoZWmZT7PkUAxZvDiHSio4V54lZQ6sYVTXfpKDbUv7+QXnJxKbC9rdTD
L0B5u6eOhLUbhJG3i/YU9A8peYLkkm7GxJCywhttEIukcwWAj1HFfLKGwXYq7wvc
oAYVovVYvteSXht3/HSvGNTql4b0Pk10G5DBQz1jeTo7fqwev6he8nmGSFu4hj/+
Neii9lf3h/UPldDWXB405NUvxdj7k4hrQQNnETHXawuxBtp+73+pyjbwbrV7QRpA
kwICg2UyZj06GgLOHISzMEWLPRF19u0E75DeIcVGFOA5Pg8Vj1/roDqwG4TzbwlE
S4UGXAgLo20f5Pp+fT0E6TQ27qO1Txn6F5+mFlQjgefIzn9kP/0wzxZjzdv9hRpX
BBQF47afh2T7GOGcFnRA0qBysu1jcozYlJm5ZRRXTs8ZPseGaONaw5AJgrvZXgyp
L9JdbhL2/Pwnjg3YH+6/YsXVHHkcR7m+52qREW875ZCwQo3DKEo3OdUofTI/zPrX
webQOwGPE2bmFM2LY7UBcR3x16vnaNi9k6zeklXrIAwD2YLOcl6da7C4RmsNmA35
i5NVY0ORCwh+CqY+OycVK4EUIJdv3Havb/cxR1bRQlyj38NxNPr6g3YqomMWGF7C
Lk/RsRgpjo1gdCEo4W9i+uag2dUywr1o2PDbo+4GITIGcNdqzjHEC8mSi9JQX6NF
20L3w/wGJpL5znzAsrSg+TvHLITmpFtRZ1zitf4/nPnn4Tvth936JxvhzD4D3Nd1
2lPzdzShbp5zfQhIZqPt73k38s6uW7nr+pg0t5r30pzpjRpqMceHA9txbv1fk4/6
ONRRIn918yH/Oes7yv7ZU7NSzTBUH+TY3YGibwhGxsE/FeMNoneBwDLweSCXBm9v
ZHaN9Ol7FIoqF0ZaW6CeyVc0R6zvZiyqPU6wBqsUaG1IpRXS9A5ygfQBQ1Epkw4y
rSNOLeIHJq/LijYC84LY/a35xU/bUYIoUQoqv+xaNWpD5EtFAmTbSclD20whiLu6
GQjZSTPMKmCmlTcxlL7GxWYzL26O00kDrS8366m+J5EjxwgSKYCkwQZiFYligGto
K2ZZ0IRZPHYFrsM++293hPJ61DIlTiCJePKG1j5Af6S1GGAPNpt3ZGpZBh11CpJF
Ok7DkJeGILiwHy2607mk2HrrDlrfqxqOwLOuAwmUmAGnmHykLh+43hlV3QK2D0II
OkuPfq9AdAUfKMqBWFmqEGcdlivLhq8B+5GSaTAp4HoI/wuEq00UOadcTmXKm5re
t9PHk8ZHhqSPUOu29Zkw6U1s0ccMn1IpPp+35zbLrhA4Cr4+Gdk/um9cw0+xpGXP
mDzClt3LT2QAm1ajU3gnaOzHAYNFANLa/ddmNsZSlVznxsQBVTT0M9lJvXhOiq/W
Xt9j/9wsHOdp+JeVX03t5jHL8aDzccHhHrhOeiCavaNAmILXjKZ1+I2f8Co2xhvt
bo62YK3LK6hTsOIN0eQPUlMXW4BT18ymxzVt4aM+rLkTs64Fw5h+28h6AyZ5ki8O
5ZyVgGMlIGyg3jJvxSV/7Kgku/CeeRyWW9IrKQx/AMWXv05Vw0i7x1trV3TH/CUr
QUvhCAaCK0bv0JvC/2Vecj5DNy4Gzg0Hoawd1A/2D2rwnqKq2EmiNSTDQK8zoWEm
AWARkHva9afQ4I78xL3dXCZLGkiig4XymAYbiG7MUAPIyPJAsa5GXI0dVzHanzFG
6d9+VUk8X6wVC4tiTrNvDJv8pUaSmjsC9L5hr1DLmcdI5e/c9s5IxSQxeubZzbkQ
c+Mv83vSpraNgPuJ+CTaeI+Pjf7nXhxjWmT8K6WoOiOT1ZIq2exahEnn6dwA0NR6
7aQCvrM+ZTHEI67nV//tn4XigxhuACE+GVCs5nkyi6IJF0dh0lgcXsB6yuFD2ulm
0WOle3qbU6npWgVqV5Pd5k+HL85Ar/CeZfuhEQG5fAOu+q/OcuZZYMy/BTmI0beY
gcAMT0QNcgkvxoCd9KVB/G/SImcC7MMRkH6F3rEFiDawbfsf21hntTWJJYDhIvIC
easeeAGgJrrMhWcU0haX1hZYANABaDbmdxRvLR4qyhRyby7EbKFMwHdo9WKZ4g5N
UhN5whkgyIrcjD8A29Wrd3hm7YIqCmegWv5y+4gVHxjbwqAAFE0q1Q6nxQr5mMvr
WnwAsXBFIImt58UBd3UChIDvNCea1Ro4hwrt0ncWxxBQ6c9/ispvDCSoxpoufDvN
XWc413/iw7UZcAYhbg9BOAPh5kLkkSn8ZDpfdpvTRcv7vJa4CpiSiQaw59I4g7SP
W7+iD+Ae5RAq1NAuHDpbStZxZqLu5EMZwty9xkgyf3rYcuiGNTi66Sneo52uo3Dh
oNFAQarEjQCSsu5zZE3ssat5IUa09pbp1TlCcOkz9yuI+0RpaE3KzaeOez9UOq7u
u9aKLia56abBWoQolwgueVDr1Nli6L6Fr+HNn5rRigdCykcrhiy5I5g4jejfGE2h
nkj33OtmqaigD0PA6FttJarXRNdZy40NReVBUvj1ClNgwW9VX93j3VNlBUOCeYA6
3JGpqePzI8cOcdBUcwC1ngvXSL6UktKTziVNS+bLWy6K86aE5fHEBEGJbPDtYPPZ
KgV3kS9MD7MZv2WDOAoZuoXVGOLA0syweO5erWfu1zJusoS1obargphDsR8gyyyA
J+TH10soUG13QTvcQH9XnhXO6t8W4l7cgvGOxtOt0gVrHNPd9gx+PdwiTrFEITfY
K/hVfvEXGQHVUODrBiUhHsK4fL6XQYB/5kqZ80WXUxWfIjEnbv4AvSbekApli/8Q
2VNmM0GJMPD+2UZI2IO/rAv97r2n2AbnmElc3ofMF7IxAj0l164kmlnwjaA3cg+P
RQGXFzZ6eVAS12SD6JWi5xhys/DtNfmNgIoO2/GqmahWHROyqRTkijoNwcq/rBU1
glk7ejPQXiLL2Z0NNS5sV/vYB0ZcnzejxC+U7cSeNr5lQa+sSRRx4/Yq6KzUsoRd
HLr1k+jQzOwdCLBcHelQCZ8nDVS/E1Za1oYdxJVe301atN1W4K/wr0QUQBoVZ3Gb
kNRTpH551zNS05P3YRZ9TZx5Y+dPVwuzvCxc+IC/wytKwoR375fpR7qd//cv0Pl+
MnSCaQa0yh0ZUN6WopIfbI0dmHulzAlbMTexpUbQNE3xV7MnmAqWNsnDEZ7wEtgL
vzTmbw0ULujkxle+RLx65eeYdw3Mf+nVU23ZZb6kXLbwpjYS1CM1Z4aUhWAJtqB8
bX8D6YQgznHbpQ+8pHwdBF0VFMWPMSpb0x4ztI/jHk4R5DX9MiV7LmVZhebzuekV
3Znc71XT5IJFyvcbqR6BoD40R3PGNcgsvmhOQsyXxyPlne+TA+liMACDn6r2cDSl
sinSarUOKHJFDenyAnsAm8JYuN+/LiMc+r0YBDeDFwNSRjeAFkbTBY6YFmQGY/Ce
J503oYXle7Y1mtX7KYNCr8Z0nYAwOouf8Y8YuGoussQ902gIUAZV3xGuuznq7F2M
u46v5pTVj2+qCDsMfaT/O1+2q/N2YGEWonGD6YjorWHeaQeNyGnm7zNb6MFcHMcQ
SnfEHMVlbStkx/m/mqPtTgHleYkEgGg54G+VWQBrnLzPK/BcE/B/Humv9cAeBs1A
gT+pIl0XSZwjCXCqM3pQ73ID1y9mO5z+9pk03z7mZndXn0+syj81ZHiJlUyg6XwS
fJw5oVisfx3By+uZv5SA1JShPcIuXBoZcDvNTqyZdytj1ndevnXdqVGxXrUX47yA
QvQCBu8R7giimw9zRlpZUspvM3PyKzrBgeMSyDa1l3des4Y8GZ8mj3nsA3b1nHpQ
uoHh8rkrwsC3ke8KaxNxTXGdbDm2r6K/2BqOEQjtlWhLuDtgqpTuo5QOhrKO+dqR
JiDlVWRJjHscxEQiICAprZ1xpFrxD7wExqZD2ufw1EN/hV0mhvbOTiQjAeuZn24K
WZoRSrl/aUKeaGVEJNprvp9x+chhJy25UOO0QMW3LmR53+xJTpJV02PRF6YSisZ3
5LGMGCxYSALBM00VGBYEhlm90LLPMTiiKoRdFUDnwmUgO7KAAy455eZDJE9HSefq
YQwot/O2VUADzYiKTUQ7KYoHhtdMp8mGLvnNuB6ux0MSyPYxJyLwgrDeDojolbil
71/IWHg5bTvCsyzGvZPck7H93BNFZuNdTPfLG6mkNm61gAg5G0P/i4gKZbfTsVcy
liZAZWVUZO0UNbSKqm1sFvsztuwWJS6X429AN3crqmS24T3Yij3Twt1q1q/GO1E0
fKLMovk8vpLtUNbuCeuk++tkCmdcEYVtrQlrx06LeKGXTaC6md5Q5vDe5z6zvuFU
M869xE+aiVK1RAUUcaammnU67MWdYrXfuex06fFUwMXmESSk9DDdRizie3qicNNs
iT7d/PWnljPYY1iTiw+wCKIsZlNy5OLVothUK3avX9AX4hSoYQIlIKD+p4NWNusj
KgCbSuguoUTvBwf7oIcb/st434Ohnuy5IXGiLcGWWENlK58CS5AYB7aHfhN1HK1M
YgGcRqePsyzIsTxeKKTA2MuSfhNfhGyOZVfnfFRcuP6YPkkj5VZ9ug7L5yiBeaIT
6HZDjQNxVBokcli/Pcfdgyo4USyd7QT74pIDGUd5c7hrgDO5J1Fq79h8mRdmlIXY
giSLDIX0EY+rNkfJVRwgS7MtFfQr4oeXpFeqmikq8neF8M1WhTsJpXDd6UBD3+/M
OwEs7gBU6xthjS0ZqiRedmFpTzDasxtb+4Fan6FNXC05csWma9s5AtmoXS2xbYQQ
ntyUTYFlhwZvB+15cNOKU5ZENGIHi0yEsY7v9QrmUo/nsTeJnRXGLoOEAE1+Ko3n
kUD1FFQgJ5Dmt6W1ECkwAxcyl313GylP6g/i4jgII7PGvNlbN0lmjfGk4Fv7pZQ8
QiB80ZKDkf43DjNZ/UVCZ+SKeVlSUT6PAhLonZkm0bfBo0gaobl56GAjVSktPwjC
UarV+5LZdhuRUdaAJry8LUO4FQ7G94VPfEASQ9INHGJ/DqUILVzBIWLoq7cxCf6e
QS7w/MlFFMLfejy6alYBaKGOgBp+n394djo6+nub0/SLDBhPQKIhB92nGKycp9Dt
RcYvUyi5CfURxPjW2r+lxfWzgUUo3GqgKP3rPHXoR5wHC//VwZLyLSbdBSXpP6TH
fGimQi+w/VbNP0+5FVVLsm4Cqlka6S0S2g82RY6JSo8IZNyAYRBDmLL096KCHRz0
8qN8gyyP9Hewh+jIQUS7ZI/N9XT3OsHvtAA3McsldwsuP1+yr/hfpy9zLA1i5yyA
yfNPX91bIgBqOmdW2A4jjBf/lvznzpcNeSyrn4sv/Nhx0IqbHpmTlURwHlzH6IMZ
KXqExHf7ICqo1wPFVt6OOoODl8Eiqcr8+PMBoL6qrfDYRGR3kc+lh8e9win9klq2
8r+DVI26vcrl8oYcZsUECekuwfWrbZw6NabrvtZ15yfcOtNx18F6kED7HWaPZmuL
GYJ46h0gvPR/8OHqLLNM8Hc/IMsPwUj4aqJ+c7Tm7rwNixBJdHdZSMhlNrWMP/7o
Lq7YThDK5xkYwUt4yVeJP/qkjcbbp23JxhzmmGajMVgO1wwiFicT13uOBdvUgj05
tuYR8Gy4RTFViq+5lGn3759GtbIZT3VPnEcCtFwLdRMpO95r1FcRSbZn6Y/Z8Mbr
FRV3pBxqSSZzMw/kRBIEBrJFFTCZZHz8SBbhQ2I9E19sbETGvuijR297HL8hi9z4
NSAZKJqUxyZ4mnL1Qwz4zsb4r5oOcwW1MB9ekYS7QvNk2jOBOXvBUjQNRxugZr1V
lHURB6n8D9pe8gJSao1aLQlRALQIhilVBjq+k2AQ/DBHWovwOeLg1AnCZ0CJ0/fQ
K6C9Tw4+4NmWH07+eUu5fmYJGYklcBnHZUyHGPRK4tXwt0w3BeFgTd2mu6ehvbY0
t8VFwIyAFMVJnibl4P/LJ1HyB25+YWQlr6h3lov5lMWJCqxbDWva35VnkwFXbTHg
WuhjjteSt6TeiFPCarwLIfLT05dGKDTfHoYeV5uCc1Cv4DOv21uvqfA3VJ/qB/1B
uLY80ULVNVkq4/0IdBWWRX5aHMBjCayFhZXKPR9mGwQfxPbUykGCV6/qhctq7OnJ
2geIzvoA2jjBOz++E+H4lGndTozdCQri/tVbnCtl/86fB0iSRNs+7wyxJDSAp7L9
vUvCVJXRPDJfnstwnqoFiF2fNog4aHL6nJa53e3OvB67PvVrBMbJh12VdrJPInBN
LNCu92hOBpZU4+HSPSF4huMfpaoJda0wpVi2xDR8OApPrD7ma/+gVWDoskFhQskK
KlL/2SB+PmYlDVPOuMSVhagpLOd8YleQQuY/dcxJyv6RamCsFpF04lYRFWVSkBTn
ltO0iIJSBLHjk+axwVMNb8Zlbx/4eCSh3kdbgds/ynqE4LmQutCDO560xI6AOOvd
efNIh4ZsPiEpIRyE2BHTLNYzTecH/LJ8QsBU32ilMbKdqIrUcaP//+Urln8IhNhJ
olTbDyvCkkuCCbaEtKqOrL2SN4Q7FIUCAc5e8aGRO3TtpijVqsg5nFz06TJ7NSwm
kjwjdktZRTs28Jy4MyIdXorNRp18bDMlZCUnvFV50lrMePr7R8ibf8mqkQJ1LdOx
FVjqG7mnhn5o9u2nZaU9+qHM4/MCDrXy4BrS5DJ8TFlGwhzgnI1bqB7fJajDhkIV
4Ljum1aTp2TcGaQrcc5A5yCEhf+nuzT8qreEtqLsyAh83RwjzZ94j4vsUgSnLu1i
aGTF8c4/VzTDZgmhMcQO6tz/ktLBgt6HSyt5kSA55cbkv/QtCn5bnLSA1QnlWGFA
uZz3sccrfrCULriW412TFb08dCXPckvXTTBcZW6N/UNaLrjxADLfE7rbmCnjqDUi
skHOMVqeuddVIoF9ddDmrgDPC0kgJ4A483OYFdoHujmo6YvJc2Q63QOi4cSQOKFS
EWEemzeei+KdARoKDmHTN4opr9s6Ml6EyUQPFMYrRPRKHGt6zl0in+/e4kBQVABs
YqxRdGLFxqtdOZVUsZsHHkQGqf/KTpNeR2hnqsN+eGaqKE9RkDzR0+LMOmWsvWIh
6U7rW1+4CGe9Qtw5S6mdoM+Q1Sd7VYeJ8OMC+8LQW+b5BmmsxWJubUjL1/+qg4yU
3h/Qq6TCmh4v8qtUsE7LvZyk34jg3awpVC7xhaRHjGsTFrjd1jLro07xOBueKGBS
sxRY+6Zkdaxp/x42Kp3Y8N+5yXXNbr6SF6w88g2lTA09sf6AIyplwS5k7TyH+B0Z
WGEp21rgc8rMr+qfzw4ewI1NezX5Wc1Rxva1+jy6Qy5yOfG+jZywbZGUpIFZmpQd
skbLk00zt/TH8bvYXyu4T5O9ExIyVB9UX1MiwI0KivSes3lxKF89YGtRG7Q0BodK
UNNl9OtzaZa1QNwZ+hcQOrDnlpSUwwVLwJIE8nL8Q2M4lH/hqH60mHG4MfPkOFy1
uF5OXJs2jRtJo3Rtzks4cwlSAkK2xKX0WTV7eULqVnG67S4u1SN/FBxxNvS4bcH+
3tgk8BAZn83bENLDGbP8xGifhLAaxtzTFoyneX/ufHkymiGB7BX9lksFVRQI4hhP
6GYbs3pm/bKgb5he3s3XbnacCJH96BoPVhHDZB47ZFn14mbX3TkXgUWDkWi961LD
DAGWUpvyRyL16+1+OTsZ9YVuVJnpTFhkRSxBZm6+NxCaPP+ZTOkcLgZQf0ZCh2bJ
1zGllPP4XPGVeKhrTpqxAzKj+c4mwONxLC8+s3CKRNLVfuGySpvGXUplAMeSOEbp
2ydRSXKfFhqGlGoedi3BG98/ub/eFg4AHSRSUQ832FN8QBZT3MsUrKLB/gjwl7q1
IuUhhm3Oc4U1MkDRZG4Ch8N0I560zYB7IlQToMfwH2GQN05szFt8LFypCJJGe8wA
YIkcS1Zs4rTO/CmkKtwWSfz1ROwJDPRKcLfT2+iRD9ZdlK2BA/rlTaExaLMDYc8a
ZDyOtyZWH2cKGmqBWSDQw97yVAr8fnh2g1keXFWNFXOHJE1oVDFsoyk5SyTql0/i
98b1WwEzV6H+oe1W9VUHl9z+TAkPBoQIBtPp+Ig5hC70lxuEIxSswkjNQpkTMaX2
lBbZKVFbqCwYdu9/Sx/uBD16wNvrKdnVjhOGJrPPWxAQwBJ+ZE5t1ve3+M+Q5t/K
f7CB28WwVwh5pPW/RShopo+/t6SvBNdlhFbRxfVxTtTAotBTVSLswqRZbuMHHYyn
NK358U33QioMKZVIiib7nYtM57FUNBxkrgQJeiTHyoj81kT7pdhg8QDECtDazUd2
+6olNezXSfMwKSjnGfkxCIhD8zrKn3r+1fjHFSStvBAzIBmMzyEFwwLjtPfCPfpc
d5MuWZ85BnEsq8qDpMzJolH8Ft9q8IlV4Q2FrAzG0SYBC2iKn4HXhca6UILLXZt3
7fwTiFqvToHVXv+ZN5sR5Bug5r6/qDCcHX3zZyThz2W/W8cE6xbX3JPuMXMuUlUI
foPunFHj1hsDj8dkEPcf3ZF4nOEz7hqHRfGZlZSHm6fK+Rdesk3fd0xXgw6UaHoB
h9QKC2iRkNkPEP9xc/FXG7lA7Jtirp3bKN3kzhwrMFNiM4HIQW3REXSwis1sJ/k3
4E3dh/Hlp34dEAPHEsJoRGbS61LT0uPavQa0TNFsyiHBgbCEdET/+1pQ7NCyGJpi
MJrLqZJ4AvhyvVG4Iy9U21bVYz8c2+ZrDY/gWfspLDtR+D8brSt3b67muArTf5fq
f0Dm8qA1cK5z0qFWs0CM7TyhdNtZl8SRd86LSWKz0QljGGPxUKJ3HKw+bo/jE6b4
ToPqmyLreLQuBF3qLUCeOqkSFCCfgDM58qIcvyaucGec3/O1Bk0f36hOGvz+X5CG
zXxtClAvCJzw5xVEpuknRRM4+J/9QsvP+X5U9UdTS266RKUtLkferSRDvEMYGyuu
YFnKb+MFD4dsqk8MF9YYwoeFGjo1MB/nczPmCU4tbdkznJkhZVRA53IqnT2Qpnrm
plV/GZYkvpjZm6Ll4/AZtQsrXhToYY9F2dkIdSkMle3XQezQ90gPQIV2Rq66w3AC
AjuWkrF1KbpDt6g7zKs0OfjReOYKuGfOwS0tzEnC6rv/0Se1uxiFraPGJhB+uNsS
wITdbfT0MFTu1qfgfsVDYJORm4LpMQSo2JEhSG7BedtIzzjZ1vPB12RMBdYERyt8
OW1x4ihEHNm038CmPzjPMKBnSDbtbt8vZK438QCMNOvHVWst+uqI2a6l8d1RRMSe
Nw/p+z2/Q16kLMxvuma2GZUUvNquJka66gm/LUIkWhYHv4Y9oCPDaAMAGDPsw9nI
ftU3cLIFz1Oe4r/rF1Kh6PMzxPRm52GrwKoHurfBEwbWp+G0KGVDw7VYCQ/S9qEn
5uBhkn/u4OIihe/1XTlM0uh801bXSTpAQLNk5+GsnE7KZu9FYtMUcuIKo5xro0lC
N1kSYEIfU/YzgFlJXUXtI3gknbDBVXKEFl5yKz5dDRtbbu7JIFKtvDiIFB7AlnqR
Xa+do5WnOSuruteH9Xc3eLZ5IexiYal0F+f+Lk0eDAEGqzizjSP5fCSQJZ8cGc7c
Isw6hUN3C3b5NE2yQGUgzIBlhVgMk/vxEdINTX5Bf+EZIhdOs2JtOVLAkQkw5dqQ
Y3vrkM5uBRR2XPRhYgfawAeys6jK52m+UMFrdUlrqdLTrTiDwuyjzq1UksjOTW9L
w6CFdOmzHCjmwLRAvMksCqcyYqt8eIVWr2SZtFf2TekZau3/khi2n+Fk0+hOJrjy
lwYLZuHkwSyBPs3m8JA9W8q9ofINAtCtsqZSDwDvtVxknA/xGerehfLivAHNzSSn
D5it9x+SMCSOP5mSjufn4qxtiwXFNu1We/6vt9d0KYGqK+5rShUetRSYuxEDvvAW
0fcEtUDAdwRT80e/muppdpsrskNIvEeagxs3i3p2bfdamH4xEj3lI/9oERVNgvF1
XrjZ9LhSVRy12vRn62ldHQqw7HeTFcq5iMTjnmPex0iDuUrmg6fIpMRWmIWNn7IO
3qQQaTSxezbBhTEt0FxZJz2RwTiIVKsH26UVW3snBoMn1cngRY2OcHp6/5Uiksmo
JTV56mjuQNY/L8Ot8/ezHkP7NWT90YtSTH0DhxrbUY7dfzrDmDLPGPZNZ+RDma8g
Lsl9EUVQlwedtQ9EYG4qnOrr6EtysBmsch6HkElDPNQv9BKF8RPes2ACdpsbBny8
I4BpACeVOlPStCg4P1g3GxyoMv+g/NT/vRL2OvsmcW40qHPHRFSclPz/cLkeX2yb
DdRxL5eRla26RtJQBNq/Y2Na7iTB6mafFQctVRGaqDJl39k/FGHLJIyF8/YmgDOt
iywc/Crx0NzIX27PIXihlVEeA3+X6L7NnodGiOSq9C7aKEQ9okdJYXUqj4Jva/uU
p/xo6EIzQ+wCIc+QvSzfG39Ma6E7A2t4Ju1o4CzI/VQAo0gpXq/iIHsuNMnB8GcH
uC9kEMzn1J19MB4tSl/wldw4Er1Wd4XxvXrwznHXBj6sva+cbws5YvOOXqgWWQvB
sJ86bezkFLBO305hwNkGEJY5ssVfQi+jfOhl2MSP37uUMOEFWAEJLJzxOHHApYoY
4CQaIje0Zd0+BBO3ym2/ngYxhDFVCHerioUFs1H8ixQCTCblCroXnlSFXFIbTBbk
2JV+BYKKqguye1NibmhMYI64MvepWTX+tpIYs5OOUXq+7XT+bqSa55/AFLkcM/Qa
RWFJcgFjTxp7TApsjLbXHSAMsy4jTpDmDRqs747tzZj4yvJIvYOqSYuTdFN/DxsZ
GjXXRn+Qaruej9rCq3mvJtohPPXuoCJd50lGJxCPB5UfnTA1nouq6nmtwzvNJ6b8
CJfuJQrCxdy8JCVVmJ8UzeV2e78Dv4KGmwJHmy2GdRqhuboO3OtiX7mAneK2i8ju
MuFbUzKvV7v1PH88D5lp1MTuJ+Y7sNA+31VwR1JJuxS1PHLrKs/jeZ0NQBErM/jU
OygMkGaCgxd78S7mC5KuEn0Rn3kmY/5itF9CYqQtNxeYLINzP4GXWi9no3lPURXo
jt7OBQcPfbI3T3gNg839IcDKZCiyuEq+2yPNv6iHO8Jp5iPrnEChzPjovv5x15iY
pC5B623sckfpwDglxM7ufBtYTkyZcziGzDJGP4qmrmg54sH64JHSsYL+EJeutdyu
BVOPHeSoKX8aGeZe4/aSV1lAKc6HjHoUzJKx15t3ujChH5XKI+Uzltt4Crs2JTMH
ZgHaGQgbnoHfmx4YNGnKPjfDWX50ojr7RS2sDCwFyWl9Dy7RCtrWF2AdXlsA0HnT
T0NtT+r6lC6UYqHvfliqNRc7ysvQlfoLd6RnNeI3P5be4bUgvkNFWlK+O6SsopEn
VG+pqm8zd0PUTzQ5u0syaN2I/oz289Ejf0f4HtgIMV+e1X3V/UbGofgk+vDZW+sB
N0r6lqif57BLje8ROg3SumtGa+vc0DOoTtBYfmAl7L3Je9N7RjuN8WMKG1wORDi+
hkEoK0mwTYKzxTRxDvEovbbHz6d00hIlOsmGJzEOwuYl+i8qMR2vuUV58AMhcY4z
98ygphjrswnz2zjsybRL7PXBozLSGsS5ZFg84NgOZKqA+IZG+CScyZpEtUov/nIZ
u3L9xM5gBvLUQICI2aZvxuKO+7xb+iRLfhyjxYszMYp98NzoV+9uFGNjIlto+f6h
2MXFwZfjJlRLfCQaaLeZQe4SC42qfoKsMiufa0jCKoF3S+kRO437DwRwhyHKnzfd
YCidmNoWEQelCoVdpC4nqpsQ4TF99raMdCUEuTPliowV+UaPB2R3MXju2WiOiQE0
MIe8uQF6ESE6fClKIzNirw4a5NzkBywaK50VUI9d/oZo0uG3jr6+8LPKdcqYIfVn
bDa0EXiFgpuy0Y1YXofxUzN7uhy8M4je1Ves0MeCKX4ZlVex0Wsnde75ZdK1Pypg
BKMWxfzcyVZlihF4ggQJMIUygy7Pvip2nEW/0UFG2kyZAqg6kMkDIsP4rTBqgajq
23CS7cezklA3LqPQGD2/T6CrC+rO8teHoYpVEMRJqA37vMddnimBObovd2RrL0Sd
gDcOgnQyz9mH2+MkJzvAfBfEXA8EMWiGwiltUF3fcxmwF4gY+apZzjD3n5bbAG6n
zMn17uR+Aj6xLe+vxx0qmBzIZvUqvOTsWZjeipB7LFoNtAz7flEkxbYdJJ6A8bCj
j5N3tioCZgQn5AjdXvAF57TbYexCrqX35rTqZbrqX6GCZ13v8Co407A/yD9Gn3TR
l5m2F5MsSjW6MiStosIkv591s38mfXFZ2CiSyDxvQtUcev5n+nnNnTXwFDI8kgk3
k7Idy10EvtiNupI3cXyAIYjezwXD5PqAoFr2ghAA27AbNZS7qufjbs00UN/ucolX
WSp9RVe3j0gB7eNQ5kqrvJHwMNH/ZlphnDlh1HDUiGx1wBPH8BTvWo20UChSftYe
e9uD4E0BSBWZheOJ9dRdOW4TsqPzDH219tdeG9voRSlBVA9aUVqqwtD3iP3WLAnI
GWiUf4wFmMgwmU54mhoZLNFmlLors5AjgJqyoYGl7PxJKOHByLwdHs2io5sohRjY
dzTha3TiuCEaRWbl25a96wavnc/oIyM/C2tXZLtxySd3c55Xs984DphMwxdiiMNd
/xAfwxyPBNTosmtbXquPYnmzSPYR6I/jH/TeLmP+YTbgkI9NjvooDqckHe7izhpC
7VD3bSJGI7IASwH0XvRv+1lpGKevJVAQr+tzXdes/tT0N/sTDqgya4HR/VmRsFMN
N+jEfn1wEe44gS+TczjqFOlcs2BUuPPgSBN0NKwA46icsbZVe58fkgmYxf3MEow2
zvW/oTnQUI8ey2p6Y44WD0VKkm6wLsxKSvTk+WPjBxtuyID9SHmkdE96kv9JSFtz
IoAVvQPWTjygYMJzR1r8Kqs01w7PPOoIjN3ik+j8iCLyzOn4taFIiGCxGMV52zOs
ipeff9SMD7cx2blhzv1neCyQMthJ5EmmvfeSMqt19wxXW7OzwrqgSCeqEa6jdm+J
wDD01kP3tnq+sGY+ZFZuGUxrSbpgrAWbXi2ECtmElnH3GV3Eh0zpMiwoOCtCe482
qi2Mki+7cQPbILSnIVpaqwlr7LX4XLZJG03oa0vmtc02l50qH73e06y1yv2uBK6o
ej+O/mUrf1vRZgaubEXNiYJhoy+Iv8Po6XdM6g0zs1fqSPdc6MeHEsgvU5tSxQlk
mdVoPZOGG1pjP6K5Gkj7+g4gNGwlgNJCTAmojgMfb0LOvj/yd4QnFijjHNmezoog
w5FxXc4UbmH0GAccjykN4Xyk1vHXFeamMp3ZUHeBnuob4B10PPph/AUekRUFmoa4
sNrbJwFeGFmkGtrQ6cM0+tDMY8NYMLtQiak708XxTwdXYn31wcYHpuk7JQig2WSd
TIuDVa6Jg1kHZj4G+Xx1d6/ohrQdKru4FQ+uCg+J6ksaV7aPWIcRdiVzpAujIcRU
GKDqx0fPZstE0LJnxbIq6UiLOKWhCXkpGlQ7gs2y8b29c6ii7lWFQGszXrE0NGM2
CdPRs1yi/MUDBfgQmS8iGEw/iVsbpe8A7xf2dfadO1e7xmisvNTLFrUO+ScoTfnx
E/reYswxu9eq76BAVnZF4SvefcBOxFDHWXZUXuVB975eeyekM1W7E3o7aRecWANC
evJ1E0aWTxEj2Pkk+ayA0o8989/PD+WT7XX5VvnzbeiiJpK352m9grrnDXc6De4u
B1J2+TIQELBQK/Q7YYCaHFPoB23fjOaMk7ev4xxwhWPJzuXRRhPwI5PAmIAhJTW2
zadgQVPfK99l72gWgJ2Dt3E/DYnoaDcGpI6HK5ELy3jI597XZiEwas5C3rSRpy7r
Px3Yz0o/ouU/i4UzkaxiSqF3rOJYyWWR4SXpUtXBajL8Me9EqBDTISq7BDSgugKL
pMruuRTdZePuj4k/PaFHyB320wE+XjAsjR9sxTG73mD86xncBACGaEhMgUdW4xZ6
SksShq+IIIPDku9/Gh6WGmmHSZdlIyTrZ3CufOftNXSYQPMMYVVvT2nDoFDE0yo7
nq7JFousSN8EmcbBcTWWMAh0DnWXd0bs0R6eXJxIC/M5u4GEbUNUROqu5Pn2IFvc
mEUe2dkBLbhBP0k/LI6CZCuoPq4kjHT+xs/vLWb82is5kSyhuee+iSys/hncVp90
Db7vBHNSoS1F9J2Dshu3qfHLtBkwceq4goW/Fh3r5xzkrcEqFD0DHtAk4QO3+skT
rBV7pEk5R9KTf7E8adhID8UsTKAOFaeCr4o3RPlJ7QhWXOB9M51fxSKys614MO2x
ZxbG9kEAhXVXtQulNAXbnIevWa4GcjLqsEPmb8qg9eRZtdes4Z8pXPldJWvDJtos
iE5ZOurimDLJcuAKwobD2eexL6mXw8YpDa95FemdXfBpDH/dtxtLZo+ZfGdnqlgr
xpCoHGVsaV9XwbUeq5aOuKNNZrNvqYyikh65A1CsOM5Uieu+at3oStRHr/wqxH+z
xIKHl21Z6RjqZojq0sx2yZWmAjxotRgjVHqoZaKvMxZabuMm2j4AsuK0965WuO6c
n0K7AsPMqWqxzVdR8DnXBRZy/ixcytXxzuMsvUUKevwRZ4J2T+EGb9ybrIiEsMdv
ph7p1lIs4Uu3Jkw+vnEQGsrZETXx0oCcz5DW1RAURriOZ90nXmzA+5khAc1lfmyW
1Cbf3geZIjDYoxT1agO2Gpi1RBDNNd2VBWXAIYP9i+G/CV67vqyooDxUcXHbVNjW
kpVoxxdo9McNIPp/tf4XSFpe1uON5PZfDLpl0S0BKZ2t06NUfP6u0P9+BgJVxYp2
ieKQlEbAy+KIuRd4R4YqPk52JUU8Gb00VDGvR0HMPgFvSf/c/iegUK/JGbcLeqoy
`pragma protect end_protected
