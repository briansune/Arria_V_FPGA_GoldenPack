// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:22 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bUT1TAfQgBhiUxyPn26laZ6cEwKio1Obb8rMW4SpMKO9VUFa/EW2s4oMfnr8NdUQ
2HUttGJ444vOgVgVeu6Fp7t+TYD6iMz7rTtV7KKtjnrlovsjh7y86YYh2wUtN8s0
G7/0QFgHrVjFvo44yb5YtfTe1G62SAAGSt/zezf4ztI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9184)
RvKn4euDDmxGnFl5mcR4G4Rmvl464w1ha1DSIFpORmlk/mmG8C3bGdMufDrzgVe5
Op9+wGAoVi8BroGRJngUBzGZo7mnJTI77uBR7A7YGzosQPcSz7YX7UqbkccOVUBT
WwBpUAYYSKiE+RhVpDhfSkB0E38f3aZ5mAavKy3GXznFf1q4JGCjGmQBmBatuuvR
nilY6lJTjXE2zHJgIKCX7VRb0k8flGgR3ZRPgX5pJ1rVsM2ZDBBmWZsljWyO7VNr
QnfBaM8Nt8u7ANicGT0DzNcIJJUvrOzcN9z+QoWwSltNDcccd4E0889gCnJGeP5u
ZUnNWI8pOGatR+XLfep39lsIlmen4ol7y4Q8sU32g5LO8yv1tgWLSEiBev+6OEAg
umG8r7qcuV8paswCbxYQY7y/xSTLYBAxsL/aEn7j6PLaJHGj8QeBCrLfMT+Tqact
F3FpJYzU/mdrKWFdbTWVw806PgvNzmEu8L+K/WVfUfVFqOjwAEbDi5sZVCAIYYkP
MMfO346DneJ1wC5vRnICJJzFRsrZMWsLaXI0u5ygPz/AFjAsw16rZGrhpdYVNiOo
q2LbgQRkuNwB4Exerfxbt2dD4mBiJRgJP60BsXnnked1awnUwUsg5CgiRDaANg43
gdo7AFN9m4QNmc3DncDnuZlxsvW6J8JJQrrdvxaIzsnELKYITNNJ/e/IX/9EzAAu
XT2oSy6Y6FCfQykYTU870c0vqgFTLTc1qMD8/hc/fy9yKathHSv4a9RO4Akci+O2
rROBgzTccqFEsF4OLBLKaQnad//cY6hnyYGM69gcP085fuQw/FHgAvSns+lmDNhO
6+wAkMJuMdvrHGo5uYF3H6yHD5lz4M9HSNvhh/InkkAPGe+FHIYQwUhhbXkSTCH9
l702kWA1A0nufqevAcJJUD+T6XnXQxZyYP/3xJl36l4mLIYcXYfoPTcuWPedf8P9
8TPun7VtrQIj+q72xZ9/udcF2OBQia6WleKFrxtMlLkJ2x4MBqaj4WKVyfPLYFgg
2HetRevjRqZ36FzhZ7m1S+ADM2MojYv2aCHO86UR/JOdxAaICKF3MT1Wt/hDEtq+
uSMsq/plpBogmODcBFINmeQgauTLtyBSnbw/YuPrEXnAGFe9XOiAVZ5EXd4/8tpt
TEvLSLF/ioKlegYfKDGLNxe8ACPNPiO/jYorQgM+va/LxNr6h/2Q3cfaK9bU2Fwh
TDZLQJ3MIygvPa7aIwmBdscAUSD+Vbfut2HVkRB1rnGppwiBabv+RPxcZZtizqdf
cmBX2JLd4D+Ezi++trWBAO4Wq8+eGU+oc4UqfkXsVbOTmftw7mqfEE5h3oWOcxJU
eFx5YP3WwbDG/gsuWKEFnmj7A8wUWJwdert+xTXjY4t5ZeqpZ32fBqPEuXfW9Esh
LWkM20rVeU5JusyLAcCSl2l13srMN4cJaSNNpLGFJd0ywnXgYD9V6fsh0VG/XXIF
+/BA8LFhIuFVVjM5J5KHH7X+YjhodpY59J9HDZ+A1XABYpteEou2FZp15Kr+vamw
MckkvuSe+ZwvnsEUzr+1WC2LiDTXVJFbXmB36U53q/JTvzW7XSM3X7oB9BC3uCDj
OrM+eLTuFdcK0qtYUA/vNXv5kG81N4OwCl+LeuGDMknTKZrsi2YeyGeoxkqhPf6s
wXKSCEqXYJdNhE9ak64wwoAIUgWiUzcAZspnKaZiy1wZct5n4FJBAdbfPMGskADv
3K3B+aua9gRfuyIpcajDsEKl3yXUgMyAui3TtJeS+FsfeeFS8mLZwFCWcVZNyrLi
/UHWn29edYJFNB0UzYhWUyjLJzScdNDSDqdbH/Q7BvFI2nBNZf6Z1BToCGjNu02y
9K6PusJ1TCm6DEYrGVa1UvnnExjlnLcmNodAdMKe1ZUskVK8Nxdpg0wUmtKI+ffh
xXgeN4MwaY5cZOY5tlB2TeEOFr0Asn7gxHcrv3Yc13s/WTV0rDjXZi9Hd2shb4UF
KpHdiuUMryPTzk5wqn2DGutbdGp0DL1SZcEeg8j/to74ze1+NwqxhOQlIo645fCX
u7bEW6gVSMe1uQMOmHGUEb8nudGLzF9pDtnzcl9Ej+mztpT1jyNxRtezildLZJwH
W7EXJflU9xP4wzbkUNsS01er0/iESNM4MV/Vkk+gw9n2c70tA1ul/X9ZqQdXxuHc
JGhXSH0xg76dCfMuwZaPW6VgJwAoWqq2EQlKybQXZm4OQH+oFKkNow0gspVqZ739
L9zbZaGIvNPcjs4K2K8HzKltZiHLYGGRW97ARILp8pBofwwUqBBuEzUVNXOPQP7b
m3Js686hCWU32PhDr0UpTQzMaplQ9AAGXuvgMPhIGJiW4tejHDqAyY/lH7pRN3Fh
dc+GSM2QNo14kRG03VX79XhE7UayZ+Zl2aZIt9BVQ/MTftd26bJlmrdsm1M37jQd
2PnJYKm944w8OIUeSEkkH+xKHGSZi387NurPKfr5sFgPBuDKwmQ+HrKc2Yf4O5iX
9BahkXJYVUWcn0SH9LNpnDNOrgl0tStWOy7aFIHIc/t8ftaiYejv7vKvAHYuSu7V
U/Wv9xiC7s0vPssqSt5udGDdLIYfzUQN1O4rJ0Lx+syOpIzxJsTwMXEiUG/6b4HM
9YAn5S1PTD9uNbZNHO8OfHf7mUdg/NpaeQxqMQCGF5y1n1YHqTsM8hXs3w/qi7tF
+IUptO6iq+qrjinIXnvoTnxiplrwG7Fl29091ttm8ayIhpz+ol0AYktjqeKttyfD
DKwmIxF2tSZv63lImFrav5fVQkwJDHs/Q+nnXOIOxwyLbm4VICGmcXJ/YcRMKBTh
rAuSxVC2jf2OrThHHVqxcWGFIUWNQ6Sj+UNIhPZp/JT8p8eSgjG3ZcPw9XnDHA1e
1GESCiPsS6k8VgUziPB3KLtG4/MMqI0yhSRMwEU1fYD5ZznPtFZTkK9RaGnog7pX
PfQgs5KvWb68aA4kR7exg3k3ijFlRzWHEFXrJZ4T/QeUtfbnyo50kukSSHLcWn4N
FVQbTQPXollXbMB1KxtZUFMWJdXAmPUoBOmzCvnJxdcH3cnsDxzY3obGmpAaZq78
ZaPjdoG4ydd8QNKaKY9cq4Q5F4gqlt4ERzKNT04VAaAOa2V6iHKLwrqkMgbxRolA
AEaP0Swb3KZK/iIhXR/ouyfi7DghgYWaywmByBp6DL3NidfOdBSaXmOt8f+yWiQ3
7Ld7yarDTJLBrKWvM6CJ7B8ybhgpA/UoyUhkAXPC5qJsB7eGXWswztAd+rwnPAHW
OL8qSlOKm23z8HLQTVGLv3QVOFrHnUZQTmLYs9NRQbR9JDAqLKJ4qsFTWdfaiuNX
uDlZdGjJE/4csP0VWf3O+V0lhizJdo51PofPd4qXqXLkt1htrjw5ifm5MVOTDiez
NLzpIVZwaz3SnondgB4wm1xMTY9W8KKbw3npk1OPbPz3suhIFFgANuwCGFrwX2yb
PPvycyMp7jzXYQXDIUQtiOeawzFvS6rR1tw6qMT0/E98XoPd81Dtk4QOvIM1n1Iy
Bum7DlSKjRYATeu7iAOBiZYzm7Kjyma/X6HC+tHSmE5ip9lt9QzHNiOReOHnIHYl
/kCzExl1Xx82WvP3wVYIqWfBBdiaSqxZhqJOmAWGZa9diy2bnAcTULDsTpiUEGfO
v2A8tryO++s3uwJfkCy9gfwu9i2mUCpsrlHO795yVgKkgO/QngF48tkxry9VluWC
ur8n9xnOHUfQ1DW4jvEDj0X3JHrbOYpcuPPKHhoPC4P0NmdcGc9YsL5NHQuyS8rU
gUMA60sejixXAiNg4crzfYbtVSUTZprl8rzJ8B93g4K7rxTa/wmQQMVHwma+bgd8
Fu1L2HF+vwdQmwUq3IwLM5+BgMzPU5Ekgt00T8gxA2+TeiKd058tTzhr7tSnOcBd
WyTDXhf0lEvn1BVe27SabVfF9mSgKYdr3kI7oBZWwIfRU6WvFeLOjAyOfM93uccv
SEFcEpOUlCodsoBqQhmYQjqRVRQQaMAF1Tgq1WTMc6+CdMJcC7y+pxA2gTdz9gb+
mSatWOkzkadenT2kZHdqRIFwWXBo8vXrCjc9Tpq+yYMWyMbqsT6F5IfaIUmaPjtx
7vKGJlmu5hZuc9l+JMippNmAJi61rr3W3Fu0fPPrQJWKlv4honRQaJYCWMSAudc+
KEah4fB3Stqm2QJNnfjdvlFWBwF9cKmBe6ACcz87xKxSx7w+P5/g/sdxUbuRu4Sc
G1DgYUVMWLRwgMYUYck6CvkXVz0+0WbnuaUIS6eddDVUDj6Gfem2oSTE8ubYh+t3
N/gQ4/PtBMg0I85xSlaYOKjeq8JmRKCcfX+6di1gR/hpeE3+5VOMKiBcPLC6eJN1
C6V/mTVqahs1yJTqNsNGJPrfP6Hf0SynB80axh+ozWjZCwBP4xWUgXjNCZrHLrok
2w2IETAeUqcufImBvjpEznK1IMoaMOYwjs6Xy0LpuveAVujd8PIfYEOO75lhOpka
0XhzxC6uSgrgpgpvjk8R+9TBJzsjwtBgwPG1aCwBBbASoDo5KpjH2cqZmAaHUoJ9
sSl03vVNNBNhEi96yVPrjla8XBwry+SgoN+xF+4q6fNWBkKJSLPlBbSjsJSLmrbi
bHIDssP4+mJFoLniy6bRcjxehzvVNrTt4mHe4MGmVMklEWPQtTOITPESwHcbEx6E
w+GxpWbpkHXxvNWPkN1NCuuFUrXcXYwln+sfjB9Ya8MAc5f8O6T7TICHchyEs0LN
Mh7jVb9JYxH6oDsBukEi+mcfr4vgXKOrO8vlgNgpmPIT9FpVU6aLD9HG1xuqoKXx
wFHlYq4sQyLy/nNji14XnfErO0EGcfvIOVsackWhK69cCmdrnoxpIc85aBQh7XUw
tSjqNAPm5/Mx5F27Tgc1s0Y7GFGNu7dFRWeaoQfy/ND16+oKb7g9o2WN+kuQDbWe
XZ+14Rwk/L94V35dhO1HlY8yT/LyvP7GjzefaphVvaz9Rq3H1jUF9g+aIOsUEyuB
t1uns5W3dedhveE/Xm1ADblJ5WLnv81WlQ0BVdSGg6c0YnwGmAqZcs1Hz4jZE+F6
2zQ8MYSGPkR16DxWKRuf11byOptSpuDNRa5M6UQBkuVJTErMXMd1kETgPoa+Yzye
eNhWeaFZ5qzSGL8Ee7vmyqnzrW+UFsAz8BPlk+A+huwfmft0GpTdBYkwcRLJ5v/C
oblKK3C3pqnCvaPKvjoNQXAvDf21+lGebN6i2ET+0vkYjaGxP7H4us5HuCzXtsz9
hrfInEpRqgKHurKiNDv8chH4fQmO3FSpb+VQPI1bL7/HHPNlVntWBGrE9Mur7T1A
7nVROZ5y1+g8sTynbo53crfqkeEL1GHWokePRkM14HDnd8QMVzZB+DBi+IIPjccp
JKl7M7VwaSQ9y9Z5LXjIO2qWxLa4BbkN6nqTNZKIa5qNCLKLvNhht0lyISWewQ7N
6uQY+7+ethlZ0qzBgI/f+J3HTh5uRUeQXEvl47h9CvJ7AdXuuxhbmcaV+jVSUVIL
pXSqP3o+smFK4nvcUg2dBYcoE7H1bOV83g3p2I/e74pcI6fTWsMLlQc6f0rk7jXS
5ZHLzJelsMj5qtk3bdUBd2nNTLKmclzjUuabULOhGzScaaKz6byAZ/fAFI95/QHM
dBtIqOmInYuMedGUvLvhNJ0+KpfdFqXbQq3CyYIJYr6Uu2iWkoKbFvc8wLaHRcTH
JsQAfmdZyCd599l++7FmpKsWaxIKlZrkA/n7wH7PHG4EaVeDwWB32lINhYgWJ1f6
k5HA58lwOWoE1At/sq/Tizw/aTk7PWdFePdivBtOF1ctF/loyE906WTasyXVT4sT
1jVhrpk5fjNLDovrH3RZbp662/9y5rn4unJB2TU6s+WGD1PXoO+2x363PECXklRX
QoF9gXtsKQKhbSQn9Onkx9RAz29wIeB+VDqg5PjqPsqDYg7fLEou+cP4JGoBFqEN
1XqQ67kcWnbmtQRfkV4aWZY+25tHDB/cxtNIWslI7Oo3mYyxdj4fFFnZAbrxF7Fs
kGduxyDO4aQqfsyNxpirWBeqUqJ/rzqoGTG7gQ4/ymYvgDDMeVHscYUQ9fKX9zO3
rPaePjF5s/bh+462O8OvRpIqPXQluPDH/KPD06e6W+sCpI1Vtvckq0NlYGzvzY/2
lJuveFfCKcGoXPcB6Nsza2sNlhEvCc20+PIlqbsBlW8U1y74xZpfc6hiIe/3Z/hD
OLUY7kP3PKFr1UZCe9gL+G0yIoWW8YSOc5JVcAFnp8DXo70kl6gcL/VVCWdVV14/
Rw5FCf0Z6S5ksFVj4xDeqSmqLjvGvF6Q7Q27s8fLfqIUxR8u5RzwQ3KOWZbimTlf
d8QnmXwcsP0so/ixkE37mBkvCjbl1wxmnkgF6moxzl3pPUz4b4hn7gN7JRl0xfJS
kFaEmv02139qtpZB+fUbxLwU34jICHoIPDM3IV9zaBdDctJDlIRyiCLJhwixK/n9
TPgmpU/jA6Wl3kc2c11q+ReQN7mxhnorq+0dJSCvLwCzBOWgCjsAnQE2bVJ+jPGK
uHFrOPWhaV6qkCBTIQvv1CbWz2QdFowoVq7CI7DKG9IOnEvcq8alW1j8PbWIpUVc
050LWFfloj11/s9qoi7wmdDZR2MT/Jf8Agq46/HgdWnCoCJMEDLuGUc1OhFGpLIC
Qlbr2rM4moN4EtEsM1W3SJ/B7vJ9xKrt+knBuiFz7Xv/sLyLZVhCjClp9nEeTkHc
sfY3F8MI5Cg3yH9e5Zb3d9flr9btI7HZS7wAwh6krnLk+RmMm5cAeEY4YazWtjax
fKPpg1IM89ZmeIBCbjDWOEkjyu/M0TlLgxsjfhRxB2XBY8Lkss3rfWwH1kNhObF6
TfZ2QoaD29tKvD5PlcULdA9+NYxBcDErYDf0EGnhhcwV9sTrzn3KGMTJGpf3r6Yu
gXWs0iVnyk7fRQnmh8EqV3PUQiyrNMV5MpWWO0QF+mxfTibSFAmj+7OauO3GRkPT
dPFRbIH5AP7lx4/1j5Sn4O69Gm4NoOYeYAvhKQqb6yxjzeMUInrXzx0u00VDv2nV
v1UHxNKpWMoa/qtbPTKedOja/pnyEH+EgjkMi5ZrzM6l21tYABa+F9OOZNNkCPqF
M4/Ov+l0ssvxTc4qUCyJVe6GB9Da3JJJG+QQW8g7LwECfj8UZg2ezzEJkhy6Xb3Q
jx6LyM3iwY4pmWXxO9WwGme4TzYxWOWwL1zVaCgRuuvHYAlAxpA8KqPWRJN4ffTU
ePxzZouCEcilwZK/fF9v7M93tZVUlD86Vj1y/tSAW47eQ4BI+KcDeg88ZGB8uemR
YgLw9shfZmj1rCj645pzEkyR6tPKwXRJkpwCM4c6DykHey/+5VoiEMFocdyXDtZ4
2ZzyAD2ect7ZCHyXMyd1G2197NKKOTThSRx7QhYHW3ICmhUxNW0vMPZszeGOtTjJ
Br/OdGdXK13kB0soHCPAQA2lAHw/4oM04ibnRxSTbbqIs0da0UGcSQRKcwPSHPGK
BEURrysCyvF7uFPy5OPiQOH5go/KbYj+/O2XeiBhCH+wIDOK5EzaauS3hKkbhWpC
LdKefL+D5xCOxPxlnPo0EWb9JvGrDJOxsgVTBaQT42UUT/AmpgrTELZx56+rYsIt
5fLsJOm4FrmjaZGjIolfeuKLg/JAU61ZhyreSAIa0TF3THBU5/0CqFHNGMJt4t0z
wRF0oKQ1twzie2hxU6nCCfDTUJt1AoXf8Q1rJn6/aTyCV0vz71HbEas9fHbWFTU4
21e5VujizojY8bKRDBhlbr5G2jx2PW28MAlknViIYp8jsI2bRgvmbyC0Zoq1fWYQ
9IAWxM/ktWu9R/YmvIQaf21sAd5SVBn0nL8b92j0eYnAPT4fPGpH/vBFDtYo/lwP
Nke9BBh4VDRL7Lt11SpEDrov2Klpr75+FlP9dZONkNYHm9edT9qcl9qQj51LnoE/
b7Wi+qIS/WYcTYfZZzIU72IaO6JazVkB30OgSe+aa2FBZFTG+Ol5/5vtrLV//4NZ
SZzQXcucwmPVR/UuGHkavByOFQiUsDg1nqqtj3L7kBsLpWjDzJx9hfp0sKW1K1lp
oTdoJrEwlwRMqiXtE+LLZUqSxXUsiFeJdlzMujYbN0IaCiEaFeQ+JKjhKgmj0iub
wD+nicmamtE5u7KVCuAPWBpCX7vbKS5tZ1EzpgNLFjgirehTH91OeaRBggcLaCDT
ZDiezcGkCquqsD23Y3QjUNgA9b1z8e3G3r/g6zdm26fptLPdbngcraA1Uy+GAV+Q
D4PaWzb+INDMnfIX0lVxqBHyhkpKS3nuVf51dkD0emEot4BTVORuQHU6zaWMBvZJ
tRCVdXVik1KQXuPI6god3rKkeXA13j1+hXunRBR1R1GsWJWPpRK5MBRPtogvO9Z5
SFhu+k2Fmtg7c+E599Wo7WwHPRX+hKk1ImNr2h92AVgNpzU7mMgFOI8OktnJ15eZ
zE8/WoMA7sTCGOM9C4La9UgbJerpvjPJXNICsm+SVpjG4kK+nIMCmH5TykYgkaJr
nYeeSM/yqdQnKh+wAW4141PZkWaes9YVrYbinuqO7lNMpCM0vngQE/yopW0Ktz0U
8W4V1IIC6Ncq+8LLkMnAg87SRNHKdriTCcgtLZgyNdvXx0c+800lbteV2BpmyEfl
1EsZSYK15LtWB7f7x4hzCkx8vZSzJGZ1MlgVUZXLnfUcMUETNJImOXAza6RDpfON
nmmrjFDwDZeF25NXE/nY9c34s38ObWFKQBijHFqV7zFIcDmV8V07q1EkX5QESMa4
+AbqCWDzMByAdVrzh91OpCnR3Q3DXkJwByri64DGB97gfvKCy3J6xAw9nVibd7Xx
Y86Z2g+2OQA+MCkC6HlzG/4iM3+SIfQdI2UyEGKbCYa0kzdvVfqHTHmkJm20Y4VY
HUcH30jP1Yf+MJ1TJzwknLzAWoa7r6MjSvaa99S67WeB46mTnnh27itQJ3zlQIKq
crrls1EmRwEdZEfJpwQ2dur0HN5n7aWiTUnZ2acBlDWc79lenlwCKvCoZ0TQDAIO
TQv9IGfXjmNThbYdHt/BdW91WWRjA2+pQFX+ptpCWi2fUVFadWjHAFU1E95HPEP/
omJbXyvxeRyk+wYEKBOFXQQWtSOiT++8hDAm6XJL+x+k/KYm3TtwRlP7Z4oMzPNQ
KUEQG4kgDeUW2trv8xONeILXjjcJSzY67NJ+fJBZu1xIU4422xc0jtqlML4mRXgA
i9nMlWFelZv/IUJOfUgVGzgfa6purNdpGpAMtRa7lZ4Cof4f7loJCp9fu1j8Hy6r
wdx/HfcK3/q8N3CGpMr3/yu4ZAIrZ08feWC+yV2PJHhUOmtOHzjebdQtomWR0PAf
8E1cqWMrigYzHmO6muBhxApRUbc/sRH9bCyOpc2oWhX53JOiH0q0UNYS1ly0N2P9
o/ewBqq6EjzIwXRK6v9iD5nWP4dJItuSCI6n02O8BPt8PmEi59FxmlFmG+Nxgt0w
adv+APN7qamIUDi+46+z4mdKDOgdaXriw/QkppS92yoYcovq/8FpN2yufNGEnNMW
IeWovA9IGMGcYgPofFqsAH4gPfBbScHzRXvPFW2Q0LxDPdfZ/MCHYLCueQZR4z/Q
/sxGJ4KvkP8Ic0PVodUoN5ba8PbVEYacjwhpwkUxocK5+AbFnUAZswZ5zwj3o3hI
/B2oMkCHFd/DYvERdGBX2P30diaEpH6NUSPDP05NvlkAEacoTSLBa1REgvt5XW8f
0nawF73lipQGe4T7kHtQC8quhbjckJcLVfngRYz3m0XzldqVmA0QAg4KmapRxIXA
Svl3r0adtDTZVsANwdWI9Z4ULtJ29MopO3O14fkesdlXHn6T2x8dlZbRwugh59oG
UWNq5xJnoVLEEw4wBmi9PzuZqDYnDFegVDG9ZgmpqT/7U8oDJQhpNDlldS6L/TXp
M4pFqNaIboO9Hjn4Tj8gmTTd1UkkG+KItFHp2OWwnxhIhDGurzw60wwlL2PYLv8a
mrmaP1t9QcOL6x6PngX0mz98Z04A0r6JCoefLvqDGVZllAjoD7ytVU487JnTYdJP
mDCLkMhAFX4o3Hj4TECrBi9tUFozeyEDIdiAz7Qfe+gbFlf0lqivnmM+taWT6syO
Ap/5BIAX7vsBvsFDB1hRHxC4P+R/4/K+zv0QqBovhRXPYQHB3ywzi/SVoa+26YJb
9ugQn17Iv9Wy5CbgbwqInzWOBqAhkLPIig9YGzplkZDeM3GLvFo5jS0Tt+yCdg/l
S8bfHwJ3ybs8StIf0cIXQuOkXIvmYlr+hfE0uXTjYoYJU+4VyEMqWyzXg9c7dBE5
ZTwhIVrUJOoWwPk9RMBh2XWOFu+3IcPs8b83qX8wm7rSfc2TiYKO2U9yI8Hs5tCC
jdj+G7WA37vo4UW+0fSrYuK/tBR0HqpZ3xjGppC/aMNtHCmwzRWXoA64Dfz/9+/v
juOEOjykAERld1W02dT+/XVLIw32BUezQmns/zEgR4rPv+Ly/C2Oe+XDUYCgzuI2
aFU38UfJtpG0maqQa5yE9VGYC0Whcl6nnU2xGIlI05rEIz4gMdLAVP6jfDb8/Qb2
p/J/eLepR6SNGP4Qu8JzJWgsjlMQRKwBJTxWSPK52M3MJScwbaBM1mBPpNLu3f3+
6O3/zpm/e+1+EUu+ISlmrOwTbpFZryJwQc7jqXlYs6kbInMO16s8rPzkREPVjbGa
LEwGOjaTcPAKPO1vDL1RxO0xdTTtz0Y0kZD4k4bcm9wVNpP7x+Dj1aVa10jg3opn
jmpTfGPkzF14gYSDzkjC7TgvmYnd2ZTqV0VQUz0QqRpwkC4QftSFnDgvE/9y5Elq
IYaVH7+tHlb8GiF2Uv/5ZR7p7Iu9JHTD1csMTzwk3tTCmczp7WvMDnJW+DElPa90
vTv0b7F7gzyusnhXqXIEgehnlHIFAadUNlzLiGq12ECMi4PapnivQfqn6MxJWaKb
8b3lD6QY69DJGLdHb7Zz9rGnQWzG3dRmRBd30vEDWRVbXzLTBYqCKvPB11UOidpd
/Vuh8aVZFoj2QtSKDudqfoLa1vDx3oW29Gb/H/xnTcyv5buEbbaySJqmKfkHfcoG
MIdpr1s3uK/xkKumwjWX/FPFX5dzLA2CWufVyI6sRarJoRLWQMQsHdrQOkD3Rbvz
0BIUgOu8ckvnEbl0MkaUm79wX59QjseCG5/zpkcwWNZstVujM4nDu4/KV10c/qLs
IIpMCJq6hPkd/BPFMExD3L9fcb/OgwMZPxbJL8+iDXXIJldjOtpwm/MO3uohPhD7
bvD705sknpGJzVPVpEHjNfcIGsG0syJlvDol32Zw6NcG6cqLX2tw+ReR0pNazESk
FAvYNrUeDvdZ4HB8uj0Vy+cNw6e7MHR8da5w9E/k2NfsFxu2fqmRTGl7Svnepv2D
+sv4Q3o8y4z+tFKBnIzF1taGUDaYJzZle+VmwQ7KlfEKxXyBeQIyRWa/zFhTalki
MXtdIx4/IihHRyRG3PNJY9uGrqzeT0PaXbutvyvQnZBT8HKxRmnAF5DNU6jrpruN
PC8UzviiIz5O/TlM5YeDpZW/ktBr9xvW3ob+IlINp86kdfGR9bAY6jXOSiOJGtYz
EEDTmKqUJW4/U+m9FIXj4D5+5nW39IkYlazcAKzKsd2n69VcI6pT0SuG1bbaib2u
Ml3NtA5LrN+ZMcLV++mJa0uUslEuJTSGeXfIWv1xLx8OC1J+3BmDQeaF6Gx4f7lC
zBbfyXEk6tRZHJvePuS3s+UTiWI8MJizG6ABTDUlT2/vye5XIUslSYCNybf5TLie
KZQ0Gf2MUTGmyQBa/HRw/r50B2rGdkW2ZcPihG3veA8Y8h/CMO+5Bjn1cbZfjkBS
OdK4vMlSh9kBaMVXNR3jjzGzC18b9e97mYyg1uTahHdLooC+dWflF0oB7fdYd6E/
lXbrC4I0mpNpQkGJ+UyLroSijNEJgqaPdJtbSaW5oqcMA3M7ErlAxjwLVhF622I9
aDTwpRdExuezQH4j0OWtFe6Wm52xP1x829zntTIOOnPjRwmRrNzaQzvhx6fzaNDY
sFOxrvr0Z+w0zMJ/mvrTA+QoqmpyC2hmTcCxQypEVU0/A2WHyFH7DR+/jyx47+bv
FRaRtCxZdPP1s6yotjvxGTkJbXIplRp054MqomQCSTGeNIpHHx5ZEGKNAb+j47cY
dSCe6QpMJ/j/JARUmbT81XSVGuHiv47USfKw+4s0+lY4guzVYBk7fonoSBbaqi3H
l6aPUrbUWyf5Bs9ExCe7Ew==
`pragma protect end_protected
