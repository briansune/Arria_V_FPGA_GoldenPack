// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:17 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kD6/he2NsDx4PC/JEGX/fsv+xvj0ZD7FaRKx5lRw8PbOprPziaUiW8dXGu5nMSbd
pizT+mQ/5dHw84rtP2GbPlAo0lwv4+a979lDJmRQjzW6N3V4c+gER+cCQndHVl0u
o3xGLXc4PLYfzt/nk59LxGlbULaSWmqNHwzg2LqdWO8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
LGvC5g1t06HW/njaRmGjiG2mzRCsEiVW+txNbSPas7iG7ioJqBay47pnjsfpMME7
kYDtua7XyiptKhbmEHxT6Cmn8OeZswoqH6OVIWV7MPRm33sq1b76TR/ixF/fXHob
rOzjkx6ALfhwbJyqepg+wBsX0Wm6KTWKSWq0jutQRpsQXr6uNSCEoNXJWJ3/aKco
RHH7+PeaLyiekBvPRRKlMqszCrsEmrQAi0TYr1INWSTbrjLdDSxtt92SHSJDr9Y0
la5vEgVi08riUlsHwjRWW/TbO+tz0FhnxGrD/UxccO0sv8E6yHiHdue+J6AFnE5p
5ukMSsLL+xBbUImINFMiL0mb8LtHIl65hqwQ0tN5aDcgFLdRR6Wr8gL+RR79t1ic
H5bK1IlvGI9+6MUz4Qel7kcI4EbdJ1NkBLXogECmKW7Eqw0bI0bmlhHTHAMBjNAZ
hlprAmtdg/fwXA8bzWBRa3uu9RrdSTxfMRjl8ytqGxn+nIWEmzuisJo3nKcKp4lJ
G34eJqqAZoziXo6D5/D5D1f0zflpd1FwL9ouIZup5IAL284KPQjyx2UWwoadmBIc
IPgNJzq3m5aXPxH5cGR7eBq6XAP3rPZbPNIPcrs2nOcO5Ygg9PRJXY613tq2cqGK
0OAv3nTTjpXeISv67rZ9qA+pHnCsh+w6hJy40BuEGYe6qwGV1xaWVANQARfbL6ED
Pn7LG781FYeyGZIFhbDED0p/jUN6Zm3wDZkFYwAmy959YRgSU0BdTN2DuEYCGCD4
8HLz3CPxzchLnpVUPtVafVBnJdfIWdmqzhu6B5gI9+eOFcHcwQJm35OKdcneNBZx
i1HFgCJnG4AY4noN6eKZg/2UHNIIuJMerUEW4mMhs7hmMBe91iEBqGOjDgzKktvK
Xzq311uDW+C/A7GYhtQcEuzGphhLYsFV9dhM4cEMuCMHKw4yoLYNSFI/kcZdqkA2
PElZp5eaV/uOMaakp9s7cJIeZWNGgNACwzCWeZRXMnB9YFkmy0nZeNbcB8K5RnEC
C6FSFeS7vdC9WJbRs0lMwIbdtDLJWGqWb2GS/16c9EWtm3VgQ1QLkkO6AUk8KRtZ
tU8ZfOPb0CGwZoipElqH8Y1Vl9AlskRNLkZjhP8JfiKEsgE9d0oSbl8Pc23jQ5wh
uD03bObKXZxjRurQiBi0amKewb/U6o+aeoL74f0tJjpDNjZpdJMi1B3xu3ynv5kz
+mTiT+rKEUd0Pk3lrkuq8VGOyA8wJdGyGlI4M9xX8Wfi7lmXRCKC9Ww66XtHqrKL
lP0mVU28k2jsah/QBtfFN+7apYuozaFykjiPMaND2xLBcGeg8d8NdMLwwH6VjVKm
Zqd+DLR2oaGdcdLfh2cdwt7q7Ivmnps3wWfd0WJ9vPiyjdQGEPEhi9YmqE2rYxCr
j5S7qJGvjZmyUyL/1r4xVz5IZabuAbFOmZrC/1GsUTxnqXpHEmqczC1cDysQUF2O
UZPFeKX2YR1XYO3I+k44zXnh6sxKp7UBwRjH2HZ9enX/4DVkawZt7oKHE8mRvtpD
Uws8TQdkwxWCpwT2zDwRbh8wyBvypQbWLPRrLWI5GbrWnkEDbeYKbAqcFaD4QWYl
zmqZMkNlXGRzYj5DngZ9SAAHvaQ2gVa5huS2vTnKXxopZIjrJMRZpXiqUPcGMA/N
mAXDID42GSXlcrvYAKGOHWn2mC5iEtqYelMBc4LsgwjK7/t+wATlHEU5otIQnmUs
ZkUz988YROqdvdLJotVae/4+93HurEejm+zEH+Q/qi/TX0V9g4Ybz+hKrviuuxtL
OSI+mPSbe9XB/PLyTIBbczpYcSYbkrwSAiRgLXLaaQ9GzjB8FRzZetPDVV9WWTWC
AYcx/BR47Dg9LX3RUEZU221tQR8ouzEpxtkqKv8t0uEJLWHNBhs+adiICl+ySo3E
5ofqL5L3n7M/3k03Fi9aCK6cqVxccyGX5TYZ/QVbmWRVKdpY2RYjfdBV/L8Kq+SX
8CuKaW8gyGfADHSbg/DgYpQBy8LEV6+nhjlojP/8cm7zjPfWneCCZNBmfWs7qn3U
oUbg3bO54K9BaQNN6KesF/sA3gLIUbemrXu1lv5MUChsbgabiezPr1KT4EDLBMjp
Zum/ko/JO8Uc0PCCitkoOOqt8o+UPwezaEoEzY1WDQqBhlaHJosW4ZGOt4gN1Kwx
Mkiihzbn5rECi9rufumKjpxKFLEEstiEVF+Ekm/o53GXb1YmBnJS0ptPfJp/7Isl
+0vaHVoxzXla3nfcIVoew4TIxiK+ckxDsEqDxa+bU8hu9XcGBGgOqlUFd99hqf/Z
WwinqYhqVr7wg2vKcXB5IS0CcRmNo0WJQ8pbClxCjX6B4eTa0Pj3NLyDdjhU29wh
vppTWSSoTz4uoJw0AWuhbOzhXRqFneeBERlLkaGY3TVbXFWXwGDLk1N3Zr7Nak+o
0LBGdU6TbJqeJf8xfZSij8rEtMEOGPm91iiVTZ5WmIxvrfqzrxWqM62nH6GQIn8A
a5M/eukM3YNj5O3HTHfHoRyIbJ/ZhuXjJSRMm6essTm+jq+fg1RdCAdye6R4iz8t
nXMDAGD5jBvYoWW3+EzsifSGvbccmKxspM7beq69mrJ0h2HpqEUyQtWsQgDxHZ39
iYLyH4ZBQ1SIDk8n8whSzhsLOiBVjJc48X2Z/924LvTCZP6/iBbW86LMikmeR3hU
82MZBy/9ro3sY9hwFGIOpXmyBUj/eUgtkeNX4hmvyMJFTbTDkyHWoLSZvbZvdery
7UAWYsk/ubTvnAFXzt+l+Bu5cu79CM3FKtmD1hsdvbiadxDKl9jYsr23o2O69SLI
g4F/47kadIwOIylLVFgp8J/jITSYOi7uhkMxDSLEqqQT4tWb1DInLOEr3ExBefh+
GQNnbEMKjT6xzqfZpLn5wfTjBIIYBfgrLheAj3h5V0+CTa2afQ2hW/VQK5vRhfHx
Vh1qKnAjwkzh8VGAW0vyxfiH96iirZYYHAL0UTE3jvq+14hR86xE0U7NIQrybITE
xMmvdyqLMCS8SyfzIcxsznP9DtuEmyecBZihv2BgOaXGVMqkXTfZgrLIBHrT6PjI
xjGONimazMrArPCsaA8f838sQjvqZ2IQjgf2vjfxy/PYesQ5LUY0VDe9pSDYj7fN
eeI93+cbaDzJZ4RI2rnNAQNd8On7mQQmQ78inzX3WszgW6/YI9wrJFSfmxYXraGA
g+l5ah794EMkzQFYwylNgd1LOJtsJ2gi2CI5OlPLmV+UQd3SMaMXhNT+gickbex1
NtGgLzPHagxGM7YC8Hy9Z0aAixfQlWa4w0iCabAzRVl/w5oKTbsZ3naNiG3781N5
/VbSUYHZ0YkCqSX0p0MlS/NPTLXKgQhzqKVBOM2l+++VbWod7GwVpaDtbzv99zXo
3MG0/+Go6SNgOMmaYlM566Nw3MaiboLbY//owCqK4AE/xtHTSblhBdXOXSHwXrjx
TjRtzwebH6CyRoXcbYU3XGrjPQG8OuI1SeqxpL6EvFMthaEV+MehI7XvQWo2h8o/
ZJ6TaFi/OQZqETuPG9I/2jpj2+GOGBNQ5ImgZY40KGkgU4lRgGAOWUglY9YZ8QM2
q6bGubkB1Z4Lk7gVgfWUfgM4gM3linWhwlZntnO184WQfkarSS2wKBomlgLA0cdF
exRCQAXXuI7lso1SgCvCzqOecdpCgT5+PhB5i0+E+4Hv5YPK2y/qCxMOaXFXIlRc
tTiNig+txmUONqMYa316Pyvkq/Ggo+zif4XzbtXv6pAwKMx3ZAlNr147qHJ1TJfJ
+8i50aMXUThNRns7X1Pz626EZ5rBCc8pnpJexp5mYpl3BeuQcNy8okMMQTBmbdzw
E71qtExbCH4C0OHSdyIJlztOuJm2S6qz6rIL8Wm8A4nv265iNJhjcNQq8DgndIsv
wTJfzJbLQ+MXrTYJF1YW+Q6NEWkL8REgJQfK1ygDUc2XQxojKGmZnxDCszHZkWc9
4sLutSYHTYszrpIEOOd3VK2vx/XwX5WfZ8tRD8D0BMv83minZgjm3qbk6JAn1vpb
sRCNG9MlKoquRT/DjbJzTun+o8cl0zAsHf74hY5SgH11zTVNcf/k0aqvWmZtEAeV
+yRtg1uYgPNgOazNFU2xTxL8Q+Wwm06TBwDUWsM4Ur4updX9ua+uw3Qsb6BJBdyM
TJdOLUpFJ7pEzk6J/Id2eNnrIM+Jhh0fHztUmp/CsUbGNSTDi86I3C8mkAfmjUZ3
1zwKWjxErUGfDOWLbKhqziplt5QF28KihxxLMR7DFYhEcS/IO2i9l2Mi70XjZfym
s50uFykB7b5WY7lY3E67rYiYNxIKVnudsNOODilupXE8nUyVMjfc9x45X+a4shpG
D+vKGVHtfNrLQYfVKGmyAxwZY2kF6mwW81SOp+YW1nl0va8dHMpiVryv0wxOJ7jo
d3JXUeT926/LZKoF0ZTc+ALTCf65ai9ziHhVU9HxoStS27ZWRGILqVpZFYykH735
zL2UMOiwnivk121AeStRv78G4C9h8zbX8/kykuWtazbYrAsuUg/d0LPQU7C47t2V
wd893jDkl1xPyk2Mz7gbeC2utMnssdHQdeaUz5L+OHmsGklCD19ZeTvIEoDOsy6E
EjObRK9fYPyyZi5+MQuDGWxkWz8LIOwL5tv4ha5yvJnK+I7+o+0nvfGKel6dwRaz
y9rvd4v3o80REbMGJMP0RVwyVBOb/uQ+Aw8BA4qAzvv8s+GjjSvRbAEwfHlJUahw
sf7jLsBWxW0p/7VHW4I4Z04BtEaBv+5mzls6CGIVxjyiztB/+NISDQQwpdtKDPjO
qVq6rVEno9V5LMZ35lhgLFT7f4VzhiU2sNHLDBe026vDgGtocPHhcZoTNNl5LAdk
xtrJ6qe35s1dgiJFp1X5xXf1reQNbopZmhi4SUatZtPfxgB+kEDbPZ/BmQMm+gFT
b87BbSUzBmOiWzyX3fzjsPgGCgxmjB0AWDECTeZ9YQuPrCN99nGf5Q+qFJ5beA7e
HZG3Siha8/LsSaz4THGFeJHsKSLCMoJW+GPEPtZFl73oRzvWH3ULa0XtqBLjFxzB
P5nCCITdrO9Ev1F4/xGeivZAbChoFYRjLkeO6skEptTgk/+a79moxG0ilPCcWb7k
n/P9AfoDUZ1pC2JD64clhqUPckKYnDaEfjSDBWeCpWLL14sFP7N705nQ2O0M9L6F
vwzkBE3eD7AJJ+bk6aNJdXa79Mb/LjyHKaWt1N3t2kMDPsXQrPG3Pf6gSJYFzwKv
RC+wjn+LWgts8Boj1VdryqL+UG6c8/TkajpH2Ps1/O/7srBUEaDJ3iRMY90pN/uX
wU0+yVj4+jYoo7I3uaCAW4TATgbX5RnAD6WJekkwYxAwvbOEJCrrODwf22g3Pc4B
dzgQ1R/x7hxQ5c4ZqErtKio28/hA3vqX2sm6JAI8QAbCCK8eXXv/B8u8iO2ldiw5
qeFFSM8BusNr7jerf4hlAzl2NpuVECrzFUZNSZY9OQH+ZIsoN8lx7iIACJihxMVw
dqolrfybAVwAR+RqVPO2EEF2Uqhg/MKTxOGbmMyCImebFe8BejRsReSwaaH8S02E
OvIH1AtgxqGgu46WwVIv4jRnSqDAavcH+pUqTxe8+gqA0p5IT4w++D6g4nuut6mj
i4LI0vDJjjv93coxIdCl332wjSCBPSD0TCmneYr1+lfknXMSJ9G6b2UQBrDAja0z
Sm35m/dtZiKPtsigT4gter+uXw/rs33P2X1LgN5LHshnLWfpOEKoYcqGhTb+I4KD
tY27vKASJ0m70C98ovL6A9YtFp4vvXPN99Ft+ajlzI/KEn9AuTGx/n+tr82+GA5b
tuc9KnwGfJ3hA0HPK3tCu+FS6ApQjTG1ksgkjTS+6xqRVDXndxy99v4HY14l5S56
3dHIBiz50rBUNDCzvf7vKHNQAwuuuSJsh1CrQ54q06AmZ/Bq1mwaChRlP5y14CwW
2tty2vO/l56SwfK6J3aho7UTWF+5s1CBBkSSAi1hWtTfPCp9W5lCUIywpkMGPO00
78qofSKfgTcvY5h5LNJbZMj9IUAMuCosrgj4T+miCUah4atNZ2tMCpN9NcXKAs1W
0l9sivDFzUHRqVSN3bue2VhFi4vC5z14F71iMfZfazDVVBxbey1nUt98cbxFFGar
0vYhqN8QY8BzgMr4j82gypaYeL+92aQgTrAkYQ6HQwTkOC5liYFp1Nf7Ap5AfgJZ
IyhAj2IC1JeVBlbMH1jqQAu+MOS3q8jWVr5zaxtD1aocO3nC6yXHWtxZ+vLPSYrp
6ghpDxHG+QriXgnYtcb+mAv+b71wXEZyQN1F+Agrbx5EB4+1aYo5nNR+tbHPfW1i
ovXzIm+j+0p3yqjWl8n63zzZo3ymFbqW8ZSDE2npUZY+Yk8GmL+BixLxpEwSKuC0
BxL3J0qKglqoqS+gYdoPMpyZFY/L2nSEGZQD57lO38trsN1ZJVnGv5cJZAbsIEIB
Qu8561qs5wt6Ed5jEQVhWVnR5BQ+tbETPjA1M6iEUkrkOERttcVwXMCirX7SGI/z
CTYNZQpvMnd25ivENjmNh29LeTpWwcupm3ePtvmFZO8byhuikMRzcOe2URYBlj5U
kCn3B9b5hphh22CXrR6kOQZyxFAH1DCZ8rqzO9h2PlqEMRXzG6OQzUwHDOAJ2zRT
tWT+YhoBiA9ie3Llvm+qCdw4JBxNz4UIyLVWuVModekGnZAPZoXTHpypf6ZraM8+
7n0oGZKOoqOjfEYqwFzqqUn9AFdIk0/xTVGKigHtgH5pJO85LnndP9IJUjEd63h2
CWXY9LT2NpD24eg+7tCfUQt6rVy5ZZfXg6hyIyw6DAWZphBpRUicKbUzxrwkYkZA
ATXiH8R1Eis+LMhpkKOIiKYNVY9YtNfW3lLBx4U94uzvneHCzvCy+zsX8zByPbOr
GM859RNQWY97wQz+T9qbGpBcp+RDVweO8/CrJtvea+0H+PwXz2PoXzPp6ghFST/W
S+NYmFTqaZL2rBvxyaecwKMzTuamL/VBsoce3BcQ03OCGgL8sWyrFxs98te0ydx6
tsUzKEOXaLLPCvA3vmq9vavfyp5JOGjU85VAalucH9rLdZkgfdtb5Bg55pKjweuV
GWpVNyiM0SxoLb4LrQOk/L5X5BobN8J9YWve4oneKspu4lkzEvMuznsJjIOQBx+q
g5G/E1lEuCluDKH5RML1D7IihwVoiqZukxWh+dFrYwP/wPyWu0Gs3OKLYqxYDIFX
WdclnStJaNfCH1X/i4R0K9+rmiFX1EyIX185lM06MSw4IzY4owHh6EILmnXbWZrv
//vuqW9JnLSdifW0Ltsg5fSJwKMcVDGU/GsOTonK8Hcu6/UFKx2h4vovrYzthxgN
nW9wBCyjvM4HMw9Z1u+l+ezxoCNxQ6Q1WNSjfqg6xciKmQJJJqhyszS1K6RmuiFZ
XYgCdUxDT/e876ve1XNgRUA0QN0EveA4nCMqkT6FNNlgL153uopG9lihUoIU3aob
XmqdDkbPgRGVdDLcf3G2VQA5CMk8W5/y4WEqs+8zHibxQoDrTO5ad9xBlJV3FSXP
Jzkl3UKOuC7QO9E5RxK+RaUe1NdQLBsP5oR0GlD3KfqyXwkvSosPyCZT3AUdWlni
D4RBXrj4Xh6ieyMh71gzN0YNnhqxxC8YclZXCAur7h7GKftkIQ4wvcKg3Sx/SZu6
mwP6cGtGYsrvdIjqo5NM+St41ijfj12r70WUmNnH+6hTa7xyP09OzALHhYfM6WZ+
GEjZIE6KCcOARJvsfcqYZ1dZ2rraiLya7g6HoT3ybhfIQR8nko+VKJCIABVoDsVH
hG7kqGtY/ENr/CiQ89upPsn4/YhYMmDYJhMuDo+7cr1pQXiZBY7WZhCB/z2OVYD0
CuuH31/+mUyLB/+D99qlpofJXJ5PO88n5yNBrwE/aP0x3JpWRb48UG6nzCFHej59
RbqOOCwX2GNJLYM6JsEUAAeMWV3EQEthacWUQzHC2pSUl5J583rUJIEOvElgBrKJ
xxMl4I32EwEIOCnftZsY2RxdZyDdyXpnNM9mKIoaV4/mAj63gHkv6j9gh/VljZ4n
2XN1yJYEBBjYps1I4C2m4+Jn+V+OQ7CP6N9KhtVVCwS6GQT8F32B38Y5ilKZe8yg
sE/vTa1c/CoTbP2E7jCj2e/bFw1sLgE118xarPqgv+rpnK4qcfRN2vOPhUrLe+U6
wiMlNZyuaxjDzCjkbmWMr2OihDpbpc9mnIwtKbBPaRLKjETLr6Ca/QE3Z8kGLihq
l9IffQylZad0sJHX7d5UaAbjffb0CPqYZkQOK9zhYUkYm/03guIEKxpnV2a8PnnM
TFYiKgOXxU3WMrXNdGtqkgTv+DokfoXtuDEn0SA+i1Jzu+Bwasqx0THxTLUIRHz0
6REvlpPIMsDqHFXpR0Nm2UMmuJPMQW611RQ0y8AY+wJTbvDrd+TBj0AxRGXLtc8k
DUsJY3kSEP9P8KL2lftHf/VzJLYvcWuBpK2ZVlMeljY6Lpzdh8mQfQ4A8ARZ00Qs
slI+K2w3hY75PmbPRpZpZM2fi5/RtE2mC9xtMHRU4ZU3I73lVpya/GZUv+AYEAov
MWHT+OWTVNriAwP7Fbc7B61gFaglMedfu7MGdOgrKDOpK4vUYueZqGmiOvbKdlt2
LMUBJW/BmIJ5CJQe4oHj5VHe77o3+DiHHDd18t4TjI4ndTb/6ufMwE87ckLD9z+q
H3IHJ2My9hQv+wEfpxdh4pkIlGBBkVWRR7ll+pf90WQUuMxLr593XNNUxiCYpZ+x
OB8+XF4ga7oKkKSfhe6lbnMJ2LKj1dZNcpVeiNJJn+Shde5VydgR3JagLI8NoWvG
yygbpKn33f2bKe8gIyhWEz6FeB9T+a0TYbyamwqeHfIsKQdllRd3kf15Hj8i703w
9JAL36dcdTDdCl+wfa3Phvd8+lub0BiV8AybBDSz16s2wgb0AC02YM5JTJyM/fAV
NYO/gYMYbTKSBk+O3Bj82bxWcvRjJUkR9ZtBxJeg8rTvWkGXXA9b4PTv41tmRt9A
y/rjIgQxKgsAEu3XUL/I/CeM/gn+PLmckDMkTn4wx4U0azvKCzHNFtN6vuvIjMDM
nbSk+DzWNEFrQiCBiAk9i1gd/8jsaYKP2TZfTgwS2qixnlsmM/fPZTEylECuZDSB
5JszsHEahcoec4C8QUqHUdIMl2vrqU4AXmBwil9qlIpj1E/zgarvn9i8fMuAmNPC
+XfRqn+EsEcJj+Zqy2xM5jw68bS2ktSl4MGgvdL108WUTfCYszpy+Hh0gnq1LHAC
yVwpckCw+WvgPe4phFFerYi0Eq1X3djzZXGZonW+1qWtKgDu/yUqgx7OQGoQASYI
9mLh2kQdaCd7koyYETYe5Lq5WGtDyqBVp4ZEmDSHszhvcS9JM2KJIZDy+lgfAKmT
717IEghCEoUXJbadL0WsJBzM2u3o0qfvm49J6JBpcRVrX9pFVH8XzStmzW5xJQiJ
5MqQTvKyNzPcW/FOjdud4BXbnpQ0F4ne+QHG2ZRLRClNUfrYrZI/LI924I1raCob
5JrBHo9tQVgp9KiPK4lm3oxXWiPtzfeZ5sDke1Uy6yrvKN8fBK+jgs28/hGdHcy1
uzkHiZ8UghcfuGhWYrT5y5bhdFv6C3qgunLk4/IC8s4yuFdUTrIyuymnqh6jfRzo
dIr9S0361JXaOKkmfSC5MtEei4kAOPPY13Rbjy5yVIPh1ATWPWQHh3K0tn1oKBLk
6i9KFM+Vu1UuR8jEmALOWok5Co3N8DpGRyY1CDkXfuwWG+FTgt+jhXzeSTH/P4Hx
RyUK5I8MNZPbswgi7buB0HBvC3h8ndFpdkAw+2dJpeocAPgB5jMiaaPP/Y6IX+PO
WWQA+KxWlccEYfzEakeQu8uxgjZMyT2swzY0iEYh0as0EjDayA1FU4Nh2Kb4ZYYA
XoxgWTCv6wdMkCwQrG7akPSK0fzMIyFTAHcJRwDOJt3j2K93NCdVb/Myf68mLTTq
FCRvU4h3B9GAohOviQCQy7NR3JlchzF6gDOxd5XyUJhOdZigGhyzzSPeNU90g4up
8r1ojkEHoCneo9NcHc5tJWOM4pCWRaJe8YnnupvHrOBYlCEOgLItgerLcfQDCtIu
HAByNB3n1fx8AlsUIU9UtmLAbWL7gEl4msfuow/7E6F3Hfb0iKPWRa5rfZ3WF6l8
0JRI+uiIdXQG5l6u2vqWXHfHkwebbhbf1CuCLFGsCZi02BbMXIWLMJMukVxsbhNT
F3WECQGgKW+0GerlIIFxXsrUn/xojUm+65UWAWmcI5g80Lkmk7Jw61sWdBCfPZ4Y
RCcbCea2H1nKlsY9HR84lIJrpFdriyonwFjU612rC/hluxBwTmBt+s1CINAO1ut1
2CtVfzMdRvN2KOU1Frh30U3crCzNWjrEYpwjRRZMXOMLFVQ32j0AqU8ck/2IWdw0
5hxcAdgcdNWeKNonkY330mdXor7xSkUoYimYVtYIz99u7E1pu2zfHjBSZwCx3CnU
XyhbfGIngG6QiPKOBN9pKY/q2M0sij6EtI5cgUpQg2aM+qBSXTsULIZwIwuofk2a
bo4NqRaABNLFxAnbhvXy4FivIF83qSG8J0maIFuLsNoPOHxwvTnmMnJr4cHXrN4t
xRRAiXLp3c5a+vEvOV+ZtBTWAHhvB+ZcaqC6Kq38jlo9cOTs0cGyTMJrYuSOYOr0
AC3zIwzMTVwDmZF08jKUc6He7YO4jQE6EqtkNBM9WUoeLg2m3m1dQj2S7HUI9tq3
MBNGN5Ii4H1otahMIvy7UTlE6t+tnnecaf2UM5kIrjFHwaeIo7/PqTMJqJx1umTL
DaoprKj4R8OpLMNbiQGVduYDhKVH9sE89Av9LJP64G2Ew6a6Tn4U8wN+JxMc8h8G
J/Ci8JrtQhispSrJkQZi9bZe6TeMlaqUAXYgDkA7RCdMcVJTqLUZlqc5DRCpj3y2
RDCV9IG/mbfbnoqJ4kdtI3LVx0a4aOZoU3aqpFTmbIABQmHw+EJz41NaJFzErPK4
iRSZM5qnmay/bEz5TN3lB2Vbpo8ZE43g4sz1qzBqzkpoNalh4AIzcJPFWOUP1Mfe
fAW7XQm9n/i1r1Kb6MiuwbDDZQWV+w9siaYmweUkh8fhqrNY3OY9GJQzEB/XYcCg
1cdsp30fligOOxEXI7/a04T5flI18NuD6/HKqvJw15Lfad1XRtyPUpxsZg78mJCI
unvZlp8BTI0NV9AKbKCpfxyTXwwT8Y3X3xM9I525nSDeoh6i/6m2zzH+DGpJK4CW
mkr9Lks7iz7NysbR3snfpYO4vqyrRNtQUjV7wKPgJeDyxhqBEVfp5dJjTp3KGCG+
kM7A1k/h+IX836/DEzYohcbUSawmw9/XAJf2xjvVfpAVGHujbCGh6NsV+BhfPeC2
tGKvnL8NhrbmTOCwR2oh1I3+jLQYhpkcAI/2EVjt3eMQ225SqCSOkCzpFstP6dW+
jcuZXwcQxNsixYxvcYRqL3i0V0dv1C5+HdJEG89DYGj66nldn7zbMAPJ7pTII5bJ
sgzMHgQU+ULDPyraKyzmOHDcHCumyVGRE6Y1BwfGuGbuIfvF50bwf5Kude0l5u/a
0Z1Uq0px95B64blMLHrzK4uT681HIp5e55qOS4kpZmyJ7im7EG86uVHoUsE4zS74
Hd+EB8zoY8vxhKAknth3LDOb/Scvav3goJzzV8j6vw5oqHKD88Qvs0yYTCdszJKm
A+8eN5pJwv07A9J/fLJjSByXLXYLWs8+UlE8+GMfj52Pim1bOxYq1j4b5YsSN+sQ
jxY0t7PIO3EFvmvx6Y23iU7eT2CklDfja8SrF+txnPBMO8EnsbhYMmhjmjkhJKPU
9/gbQ0i5D2tCty4IvQKBx1SNftqsLJuQxUYBKryMuDBKeJxOqlXIUFgLfOk+yqIb
/UPa07HKs/EhT+GhlekBQkATuXJV8+Uq1Pvqks6SF37ctwiejxAJATNNypqOsWyw
jKU0m71UZcStmnBxfNCH426TyN3pUYEmUAMy+Xnuv5w89U29W7pIdgRe8FxLonRy
nf8M3h3/KQGf4CW9FIODTE2PZHwqDBZxz4neq4apMEgsXphr5kq4ozCimh2Q7voJ
NM8xOW0KCZ891Lws+6fYOc+TBsSjo90tdZ7PGDxQBU5XCRG2Pt/VcP0GMsz980aY
/tdfNg3DnlX/ppUDQeeDOILZShl79XTOM0I+gq1XOT5Nr7s9R5R+lhto6crDa3du
iv0B7cbPx1wFJ/n6eqIqOFDtG6FKwCArTRAwYLyrxmaEK4AHd4jb3URsdg8mTLsl
wgS544Uj4kvirk6uiPrafh6pXp7sroF54s/6sDml639lc+FJx3Qjfn/M9lleUGne
1TwcpTmgJU97O+EH+VzN0WKpc/YdRx7dIebiOTkF5LM1VWLhZo7Nf+BFi6OswoLW
rzqoRgGHl89Ea7KDXSFuz3lnAL3Rj5LN6/FAkSkidbJTzqhfOSrKl5eHUF4fqLCm
F1QW9ucYNsPT/eh6p4IDWpJO8A3wmQfQrtT5ZUW9NRBSJ8tFp3WvFQqJh3yCUOyJ
ulAQiuiNwHFO/N0YCR3Uvijp2AJwCDrttPbgcYQS081ftAmMUb7rNhqWo8i6fLOK
WskSwkdOjM2f/7tcvaJrFrzquxVqNaROiPMbScB7oGpbnqz+oLkdxNycGNT1C4H+
/jS5Eb5j/1/tgjHxggjkBp+LqRGuHGkBhidO82y50ve9l4XMt00S0PzqEA6oOYuC
aY3LVUJ1GlRmeJI3moqXePu0W4tqosu7KsBdhTT1W+u5hVRpoao3KgbluxeGYKj9
LLO45TtLVp32lciT52Oc3VlvYQm/MVxDc2oXD71xgjuiNyIrdpAS5UyBQ8V9aW6Y
5ROzpYJNp3nDGDGimFn5pvPrWCtDGGB2Brnoa8uTmMTqzxxa30TM/QnwIbAo57GV
BX3JY0jffQtP5Rj9RBDlSHgyqixfuVQTXyo/Mlks3dz86KQJwEOelWTyHuGcUE1R
xAuCsVk2zXg0IiTgCkz0qze2c1GYU+J52TDnFEIoiBWubDiHpRDXJX+rHckDlfa/
7bvRzwtsWDvAkuZtaS3f5xZYcgBbV946XfTQzFj+J+ydZlLj3aAY57/XxyTaICYt
uJQY9BwSBfsTBIbMVsjyJGngM7Opt1OX/Sq1rhEDMhNeVzT6vLb98RFbGvOUB4Ww
8ineApujn53N52ZpSFdHFcF7747Ao0+WKwcAaccEXNuvadUnoEj4i658E6WgS0cm
LhBa7FVCuguIeD7ECfkPb773YJchL7ps4vb56zEMoOOoWhjo9KU256gciccEKhzO
2KjRoRxTJAVrIOy9us2aC0KU7Hhj/MXvxHeTWQuK8tip8XOziyHjTQEV5ZzooQWO
S4ckjwM6IscWFkiaKVRUpoXA0HhQOPFXJ+CAbT5EGyaoIwiZC3xihbZjBnC1vISS
DQpaJ+OoTPhmm0yJDYcjXlz9pTEgngqYTe/PF/RtvBxvcHyXslB6ffQT8Q9UTgXy
6SrbGb40p/DNyNx97zJ462HYtEc7IEYKUyMe1MlGh3SDLR/F12kl2fD8PqRdYjRI
WJihaX/8iOwtrLd5Lvoa2u2oaGGJ94gOniFFK90qR2E9jcR21pGTUO660M0qmq7Y
jfT1nEj5uYE6OOdj4yTW3mEo0mvMq8su3BoVn1mEA5Omj8tUHHD2AWhZJwarBn+F
CIr07D4CCcyDAIvXE3ptl15dVUBpOApS0ldARlAhgcfMURDWYZKg0qo+kdWLxYD4
4alhzB9dli1PlnFs/oHcBf766vWVzjxJx2vCtRBmWg1pxZVhRgxeIw6iTO1qL/vX
mFXPvbWPn5x4+OXbaxNyTcZdbBAZsZoB/d00sr2O05yePckFwoXxs4/W16gkBK3z
oUHzNsxXjQclfyloRmTZXIw0tBacMMwLamCX4bumoKgWj/4eoWYDwWK5T2VzON9q
vZksMd+etYa0wemFGto2c/ZNbJjkQyKWcFfts54jrAUIypIC2IBx1T2U5sAu52Yl
0WWqHOkEJYPg2RugqBtrWy/XyHlC/r82g/+bsS87p/z1uiZ5A0pXqa8JU3rLkmD1
0S0iCECiKAUzH4FMOJLOowDsx5aBmEcp13tctXkeCPr0PEr3Y/h3iveHWl6ckwWS
OU+qoU+BSI9Pbg2FOx3d7OtI0ZApCnqdYo3NxtZ7RDXUkftZH5O/w0tCMU5rM5aq
fBCOU8GLkjw4aDwd+5nTgFe/cN35hZFK4+EXnmxsV1eI2TutiiI/8048Ce436eMq
sop3zK5vYJ2PY1y5+a9zC3eg50di4ve2l4RzCiY6VR6C5INji8v4+HfkpSvFsThI
Nj0W+sne7gikpvXzeLuybHl5PQkdzlaghVrcHzIsuyT1XlX/R/HmyB+w8AM0xmEP
OkvfPTem+e4IPXmt2SiK9kGQwtjU84WjpT8Cy6/0d2WThYMxd/a+d/nPRc7Sz3iW
XHraEoR7cmsFbCvjXs8APsp3u3iOTDB++d7CM9t4P3qlYJLjVj9dmfbQaK7LMeMg
2Z5NJKLfxLuAlbuUwOovxV0F5gf5KSQx6e7/ZVpslD+lugw+bi2Iz9lhpGCTay1o
dwtKTxa7DlpOkvIOMBsmlC7mIWjZdPqHd91F5+5cC0wcjqx4Qwzposka71Eo0K+2
JPvUgOTrRjj5kVRnruaCSAFt3ndvi2AC4m0PJDTJE1Ta6hXCYTaUJk4ck8IggcLR
3wgyIut/1Qg/9zCVIVenwP4LZMtoYgxQigk7lmPurgRsm0Gg4q7p6bqSSeo14zt2
HJXgmC22GX7UOHP+8llewjId3VfXhtzDTJmMuKeVEIz4pQ8dwxVu2YRxNfPBQHuz
MNouffBSPUTWs8HoJFngu7Qi4u8QIaU54HJ9IHjLLlOX1RcxrqgrEF1Vn8T95Yuz
Qq1jGtxnO4vMRkB+U96XvM5VyeGiyxs072gx3Hv7HaNn0gA4KMP6g2FTkFuRkDyI
u4T7pHncUfV6hNGeBQUIgc+5I1KOu91pLfoa3T4TiJRllmPnp85G/eIr6YEZ+O+G
HPqo7gSdBMz92rIMkEg0XJaj8Ig+jQwrLvMOSwV7JvUMc1R1Ri9kG6AB7Arl2MUz
S6e7VoJiryJz5sJIeovj6KV41bHtMMxWHwE5SOzqnVYH6b4v0zgJIU4FVSwR1/T6
l39AaSclvy8hsmiGkpejNMfncFLH6kq2Dz5zw6UkCtI8V58cI2BW3nPkWyVWTV6/
5jGzBDCTHhhVuifdKBzNGMXJgOXGGpQaugtuqfOXT1d2AVLJRrZHHd9njWMy/cMd
1b7Mqp8dbWR5Xs5qIMJibskfjHFCqP3Id5CF5WSk7LnUUpKXRfN50XfgMW5kzB3O
hvTX5TalJKXGn1e+N0ZR4dUcR9RlIDHircuWVi291i4bOfxzyh9ZTkl05wSkpsWD
5UwwTbYnLIOGfoVK/3p6eSh26eR9hp//i1UeH52N1wuHAStTT27fg0zZoLDTNTHY
qA5G5hH2W6/P+Umbuv8Myvsl2D+z6hzGKom5E24/4PU9yJOhMFdTkdeNVPOPt/xl
U0G1wqRtXfNglTLwDt9dM1xfxPzxeb2XvKxvmNiilFQXoe1OpAOaRd3NyObbG51x
qs/FeTIDmQ81TmA3sBXxJ7QLfE81BaD9spsEIAB4e5+sOHOB2A9zAouR2abpqIW0
BRbOfY+322XPymsGx2OMayj+rigtm58mH2sKYA0YxE1mAv13CNz7nSCZvA4pXpKa
wjyhpYwI7KZlf+DhcWYBaMJmOXiJX3iXiEnnCGFApBeirpR0GwU6AgA0my3+a0uo
cqSHc+E3ousOZk8t7ksUGQ9uN8cTfHMUEeJunQR1L91NLsMJZ+DgsgGbqeaR2JQa
UER8ZmZiMtdRsA/df/suzzltBmXN9cdCWHYLcMattCM6kvWbjWfhxw1fjG2OJrOU
S/ieTfNvEztDkmaSFOMgRE/GxBbvIAf4Fig9UxIUyEbtKCUxWdgDPKy/TbR3tLIi
PJ0A3fAr8sfBEUxRJHHVb9EHxqHRZE7YOaZfbjCce79d4u3K7OdhvsUEJWKZsl/X
bF6ontsI/CK0/9nQ7bnYGcx7FBDURvA2QKTVapf4CADysl81ugJRu7lxnWmc9GFn
/JPkX5cValY7YpYlM5ycL13coH961fXuLPhR5g2bWAjZGRi0sQbA6XqrjquovgxA
S1akb09cZRDDuRng51JP4czUuD+a04Sgsap5rgOTFLNB0O65RD/ngCd+SdZdM9lk
FMqJqOh2nZbY3z1HhgWv7kEWxI2Yn8QsnwN+siF8HpBhXauHjA30BTU6XbQI5Ps/
vumONrOANDB1cTmm7twy3pi+qEWLBVKPMzq8PeEEjK8VBOGvW7HbCiOXIVyrjZuJ
69le2irKNhWoJao16rg1ju2DLPl2gYjI/B7QpihI2eXB22ZvHCTUUgASDNR2A8eu
6msrSvJ8LrpulpbfLLUqpPQl+w0xA6SMFcEQihoqMPcZZvkZjfnpgMN34g+BfbzM
b2TQPfn9HeD9kT/yiHIo9L1QFXU227HujIAr5NRnMkJypmMd8ITAyfbrTIoSokWn
xnzsHOIlVoBSWdMAOnoTQuWyLtkDH98UDk6rYu4bT4i7MnHAooiYTIH65gss6MsX
nrG9trR2jK824hgrHKKIdCoNGssfh9roxUbDK62nRJEDnrSzNyjy79NzcIbuRTP5
pHMFFGTtE+oH0NUPHuZlmaPqGXf9v1ORziNXQvf5HqHho/IsFoX/biIEeRcPFyTf
eKjKapLTSDEGiCQs6v48qw+Iwd2+uc+5aJ8SFStA1z6/RYA8/mp6ysfO8ktits9e
ja4ypVz9UwkiIc6t8wxWw5ruoAef/f06tTCfGtzi+loAeaIvqxBrwuQIIcVXQO+w
oE1dGfKUk2mnX04ho8FOlrMqbJpUbHOxRBZ7HIbW8Tz6ZiziSo2RB/iMjWLjsNas
MySL4zSaaasv+EsJs3EkDnOEs9Bade+T6u81oQiIfs7yl8PVQp7DQg6uN3CB46LV
Se+U2ZsIxeNoOrpppDjYOqeazr8nHyMdINu3dmLphgx/pEhDG+rra6M4Sb+eAIPd
JaCSH/DwM7u6ReG+Kr0JoNeZSv/zlnK3seoofHNZKqAknoOErQSrxCq/tVwQb7YC
E/68kB8Mjikd15pZrpLOpD3ekXkMKkVlvTAHWT/j3vl0tylSZF/frjgjHrQ4W8B8
kqJ82noVPTTN1TqlMBGg8zV/yMg5BRk6wGCPRuS/vCC/jcF+1oLFZ2BIvdSA7YZY
3zmcxLvE0DMU2I5zzBT6An4rwAyQjVpYXVVnHwz8Y40extKpAvQNnvbiF6MJU1kP
9VvH6mfs9ALW2xT0Pc4m7hs6Kl8bhaiCF0Blds/uY89y/J9r7Q9nD/IAXej/USQa
AqelT0M+mFOnBhhmPxQvVUrVKty/DnOAR4aDN9pyAkY8VEpgjzj8/zb5mADv3/+3
5StXouoSiNNMY4T/3C49bVap35GYpeSeS9FQJUrc9JQVzzIlkuNSmWufdBak0YoM
0puEdQdUqMvoGVSYXBE1QPW7UWN7nr1Zt1ODSt2qxZHQOVOu1kdZ8c9HJIorf6yk
WNf9a+UziF4++5g0mnTSymmOwOcimQWRLmgXao7vq/BnkwsytglT+45DRitFIBMw
B28TZKiU8MZdN53lWQ9JIRedTPUSAE7Htm4r8g46sqBq6aX9WPX3JL6h4NUsnKvG
b/A1nFadznR/NrMnAd3NEIi8LfV5NC93KsdyO0HqDvTwLuWcltM7Knj9KrCNoWs3
262zQeeU6HZp77t849ZSWgzZkK1D2CRfalJdeL7Hj4I5tgeaqnblcCtj2A+o37VC
nWdBy2LAly7gXnTc9VwaJjBRVXiQV2lpBnqoNfmUOvCrl+Zzo7soujsUyjqtjrkG
TRNF6eDncWkXcDsEUVPRhJ/xPa8i4Q0liHFp8lIvvAgxWUNkxM6/fhfDBPwvaXai
5U9fkWhgZQW+VtOcij1ACQo+A5lMkKnLp1g8vqB4s6bWjsEkaEhAUFp/e5V/FDG+
MTLk8RjGETVw4w/7R0pU0LWd42aa7E9JWhQmDWpSj0w498Am9ZyeZGu5VFtyzDJh
SOgcZeHE+g1nc0egQnP/Pus37UhmH1ni/TkrLTQkUW3CT3F5f8gRkyf2bzRWVNE8
TQsibRkyPp77kIwwujzNLxKIY/Xap1h6BANmIG6mIpiQDUE1HX/5SdDaCQMvs2//
vI1BcqByFWLcg8OQINP9HpVC/VQjnLXTkyrOv4d+M2f4ZC3bNFolwHRB9LdR1GLp
A/CwW72cxxKM5yPRh/BFJemlDPAViBaWsBSZ+ozxNu7IQKjHc8oDZPREWSdlw1Xh
YomtlY2gtuguvjl6vGm+HdQM35Kz+1VIZGdjlKrBJrIQVWhvU5ks0pwvkFilUmlI
896dmen6gj/8PjjPbon/L17hbO12hXPktiXVXQ8waCqZ8Hqv6R7b7Mpm7Qmp6YWI
q6/FBu0gEgLGtpB+2F9InN6JusBLxQ/2Q80/Lk1G3RRUG/6n2mkYCf4XLbyQ+wi5
1xemIKMj9Epj2OizpI0CqlF93sWY/patg1e9dgfpsNwMzx+yK96dD/kZG+kHr8GV
50KG7mpf+MbVIo9yCLBsx5wbCXuEAojBwXzZR9azusgaeB8iOIzXmWjkdtJ3g1Xq
Ucr3zevX8YQRME52zbPXoS9oSTF+d7PnqxkDj/Hna2Xp1JW3fwmD5z183P+Eu/SY
9PpNo4F2wxLB7JNJ4EkpjRDyqHqgBAGwrdbg4ZXk0Vm1fe8S/bUb/LpgK0/Ly+P1
ntzEG3PlzKRxJDew2/SecWQKSk9hAoYyC9UnEpWIwwkhChv/OFcsP3076MVEPDF/
sxqLDq7Eoa5HFuhrK0uAASe6TNCaKXWDmtvAN69VOMKxQILuoPVtuvDb6rI9KG7w
Z3yFUMmY/EHbK42uJf6oA3uwgdrNB93LtG3BR4NbC6Grj3OnhhpnvKV7Pb4ctICP
vCVciC6BTUMGI0Uxop1mWHEO9EARgby4uSp5fTr5sZu0tfBYIBD3HlQ8GA7iaA6j
RL22qpq4iBwMOBOZ7f9nmrO7wGCAKibIZD+Op4q+9Ug+EFmHqOmowWsyvpBjJrZm
/MxZEukAE1oagx6rp9VLLs0qOX8SLA+TBPf0gvrZPwr0xzHd3YYbjlEJHioH4o88
8b+EwBFEtQ20aQ+VPJF7OwI5FKWcrv3m4S7QodkW0hIPvVDQCOR/R7J2P/p8xqEn
dfO6N0gXgyYEsLzzWjCV7GIEnim6ToaSquKMto4ARJ33UBO9cZQmL7Fg/0KODIDc
MPt46HBue0YCygDugXgkPZdYA7ViWrd0Wie/AVhUJjGfybllNDJ3KZspzaecWBCU
xnzrjyvNzDNIf+mbRFb1vJ16iO0JlBW+HXxj04en5A5iEAzLuFdXRlhAdKa8+kPa
Zc2xh41Ia9fiorXuh3IHiBaBmIKv2OLMTyOwhEZyXU6GlXkAjMu99QY0RBEodqkY
h2uapqnmi7/O3TdlJE4Z7eeGrkTiyBT65mRPqigAspCDq8lDSUmaIZ0MX0Ovz2+4
cCrQKSevrCAlRnAm2GKCOur33eS6PrzRPmGyLSuEXO2HxyuhAcEv4vIBaIIW7QCi
x/aBbkKJr/KqL8qiTVppa5TDgrTzcNfixgHmKsVOLPmTuJ9ySUFRluNpunscXS2d
LS7rP42Nm6SYN5LBnZZRnrWXqaCZpJ0vEwT1UQyUVp/71hl9c/PcP1dAlm4Hhn2v
C80YGNeLbZmzMo7g2AXgm2a9y/32pqXH2lthHr0T7ILp/vwk6o+s39XJiXuQFPs6
l709HVJld8uCyRZYiOgLPl1EOKDekA4vrd3tdLPh/w0eugqKYxy9qdL7QhfoV6Vm
xMHXcklmaDSWEPR9ZYn/yd4Pvh2Q8ipbi1/jo6nD99Z4qzqaEA1mhCHbQraQ/T+w
QeD3uwhXNT4kbxylFpPqat3+1dxcrOGzwClpEMeOaEsGx2aZnkJ6xjcpm3eyeJgs
pilkcWp9HQPZQ4qqdDP4OM8g2GSkEklJsbTCdZbBVCdFgN6K+PKdGZELwaDnJ6QO
fquGUnDwFFqLJnAUVDiC7VDnDLdru/nhVKLtzkZ46ojriRlun7xuiG4/tgpGV6tG
bYqples36TclFTFCNaHyQ9gtk8SjxjehxxW/5OE1BU8sl1Cw8cgkKBGgV+88w007
JWdcX/k8Mg3oMrNyzqVr9I0AkgKgvwMdPgfoRAWmI1kssiLdzpo2zMAqgx6T2sZi
l4DuGypaW++HYZj7koNmi1j23LAHTMlcLdTXdJZFTbybBG38QcEh3lr2tmQPFGg8
FWLV+YfQeqPqtCwPez94lKcy0oxuvQf57tv1gqLSjxHZd2wbjznonaryORXlqWbI
INXH3oIA1UOir9IZ9GJ1icwcY+i2OVX3RtZLmMvDQPwoaQaDEu8dvdcErnMQ4GEc
S2jBlfAMpq+epwaLaKtBndk5N0imNb3jErkoOmOe7/YqAoFTyJFErtvRnIFMA5J+
cOSgVCgl+jRZo+9v2HADTXmp1xk8kf1ME3W+ZrQzBdSPjdKjmZt3iJTMSsx/yUkY
FpXmZz3Ax8fa4uuDAgu8QMffKOnYoYRytQ4UZ3AXAf+R+SsHV4Ac0Gwfepn3bAKB
WbFSOhGmCkUEdVfrAxVbPi+YU6Un6ai/Dsvd9itw4rKjuoalvj8c7wabQcEwOmC3
nmHE4e/PpEaeqylyoh81ri1xkAS20kEMwgw4qo5rqkqKJCocdpQV8TJaaLHpgYmV
eJ66qCRK6ZntDjkEGv0nJQX/NFbzsf0DFYKmQJtV2PFOqBYhmVjP5iLt6ukAPgoL
b7f/HRc/R/VwjZHChUO1Suk2S47OdlG8etKfRW3B6SxDaz2xerOfdfZOV1nL2qQg
v3AjAUiG2G/CC8Txd5qlurq0jrc1KxjcZ/k0hDpqZoIUa+L7k016ANec1Rhhc1j0
njlF5JLRohdzRFKRe1IM/eM/2q1ThCcxHl4tyhpiijp/WnOs3npxrpPVJFbU/42g
zkem0mG/n3vnplamV0LluN2eECMYyoBVxt+E+0L1idkbEO+upyTa2xxjXXRjR5zJ
ViFm+lna3LNlwJtYAxndiZQlUFxgI6/OW8ORkvCovm6wCUUVFnLmFAuCNmOaiUJX
dotlo1TScAtG1N2bdkJHVe+ZNHFAGqMutCzoRr20g0jLWltaZc4A5hAf0UrSjV5y
t2zueUqPjFBCztWtWTeUImAosf/edZ5kA/9OjFmaChkHAIxzJnzBj7t7dqfY9p6q
MwRiju8VG9VzkssJKTe5Ni1EUblw97lBYhgNgvFgDrai9U4Npk2NZtbGtFxUgynK
LV3E+szKLZ6h+JifhcudIss+X4B5w0bLO4AtEzTXIgmceesIobX+M33UOQDRLCyq
BJDdN54h9Mzg9AEoDKCDpGaIwxhnWMu1YS93aC/q1su23MSBQncsJj8X5SOCzD7b
k6+wQfN+M6EfMX1oWbJ2xKqyGjgtU1jZXc9buf76PgRaBsdG5THdTX+sEROTg/o2
b04qNkY38BllQsnzdMXyJ/r9OUvWfuuRql76nXRVcXA2Qdom/YQwTuI1Z/AqK0ue
zB/ObXRi57+5KjcyeN4bvJkXo5nNM/KtNjOu64c5NfZzusZeeNxkzwdELJ8KEVWd
kVuEsNPfXiFYMPM+9V7O4s+xx59CDXK4/v0vmq8huFNVu1DMn+9HY4AkcD3YqCbw
tbUbJmhmoiCdiwVLCIypHM4TYgDvlU4MUmKSaTUuh6av25zj9MJtSD1BQrEdx37k
NU9fkEkGE7rZKnnGCFcQqh42ilOOFgy1fSNIMTyqm7ulZRhniutzzr00w/OnJSj8
zQ+dNXzJLEN6/nkjgzd06m4nYQw/B6GywmyF09oHVCMO+KARWzcmfkoRP2ZVqe9Z
lHJhC92aDA/aKn+mtOGmObDssFYj77kOzpaMuGK2Kj00bibR18Sn5KHTwVK+BXjE
wsnPWXVfgxa+sbV5MEckUFI12j6dH5cdtftbRK6j2ZI1mMDXpRvhdW1pw/gsc/u5
te8MLcm3rorHs9CPEY6J32q2j2dsRiX+s2syiln/Z7VmkFRrOX8g6iHk4g4QGX8o
aNo22kSYo+YNVjBIXOfYTRvX3toloZbGfgzuEYmwekbdWG3XbzovGDEVKxDQaMe9
kSk7Dwr/Vwqqui3F26nchh4JzHTN+VV7A7FnT6D2TcO2Gt5JAtVDzIuqyyKbPEvL
mx0QMiT4R/5fsJoZ4NA3WI/CY4UcV/Y1SgejOCMbwQxzhJlPGAdlXOQrxCHxWGTb
oHASRz6boGgm4TdBhkSvt6JDoyTwO1fX3LfYHIvyhVPbZ0kye6HP3npw+c2nokf9
HmNCPa8zOflb1N2yreY1R+LLm30DSguHB2qTHNp7YnlxipIQG1UGBpF4mH0v+o5F
6zy+YO7SjfYSQC5TNpo1vjlaeNqAUdUouuyIBBKU3NGu6eBlJjzKVjsWbSBPd8Bp
XpAuDd8G2cFwDyp45kM06ECOng9sIbPNZ+5+JV51RRWn0tN4JPJxzKB29OUrJTUa
0IwEOcDvTvTU8nWCd2aWKGZWm8oyrpEG/fuwkMr3PRCShHwLqjue9EByzqieyjvB
bf6zjVxHmHFXWt7t0knYbI65gSPlwHD/D54JU6S5VwPhCQG/O1cxUmPc9XF/FVlx
19vaaB8GCnRYlMyGjjnBy4l7qcG14G6Ala10WnUBZHIXSTPsOQCWS46f8LcaWOCP
4OPhDCtFntc1XIBoLoNZThSO+lMDLHRYjvMMJHTzo9EhTy5MRsJYJGfne5o1Ljy1
2mB8TgjAe8im/FQmQUvsMo2IrCH/h/GZWyv7ekIojgfEH6dFZeDYR+2SuBepe77C
ry32Cv9v8p2vgVQ8I9oB2+YLArhga1jecJtYOuaWxaS31dsDkzt5xQXGLNixQ6Gc
k2j5k+u+5UZgy0IqsagEoQK2YciNUDNSJuG7fZpxMIkUuUKwGv1uq9Ri8Idyf9YA
KF8EgaV12hoOIhChblGKxzectK17o8Q5CTkPSwxTLn8KiSGDCwikw2KOmsJVU6f0
Ncv0w166vqPyZyxS4UitoHu7x6c/hcdB46YRHq9rZoglmMG5oAtnW6M01X4Y7Rtg
s1j94bJhz3bHkJP9LWi/g2nKzAK/M1SChDidms8zdfmLc+ED2Sf5If6wQsO6DhD3
uMGLx3JC/QONWxOCwMkStgHFp3FQJTsmf+Ik1TciiZEj6byn/ivPnXvMNU15iCaF
6+G7T9ZqLg8Ypn2TUWzOix2CVBYs/M0wgkSwqiUxnn54LpPxnfMl7vKYkAFpKv9Z
OjQizRj+EH3qylYSABJKfT7wuVcCjQDxLK+BX4vFD870eQlh47WRoj6um6v8i4Wo
Ud5ydfU87UaXOHOSkinFik95B/70cysG71h15MwH27MDeGrNgsjdnkjduZk9JJIj
WqyxFkzYzYKrE6qD4t68Zg15lTy38RPVTSwnsgnFjOGjK5lEfnNFmq7T2vteY91E
XEPFQJx72DZED6XFEzpElbgd4GCnloJUSw0FRwYv28ULVAB32Ln2kvZq8XtaSiU7
M14ClKa1mu7yXR1aqxAeIveh9SC6nSYrEh54uHSnYpLXxaBrkrkCJUYiaYunLVGk
jIHQXihAZ5TA+T0TME7VZfoGYeczn63YBypywLAkUDKQC7sQKAJyfYslCgGWoAm0
98epO4xTDlLrcQwQO1des89gW83bNG3dTq2feDFZPODUvH/VMv9AB/CpBwhhTMIa
CzkYaKWgNjMM+3zlQ8pDQJ5oThweyVKASZ/xN+bR6zNioTir3fsWSzgW/EYeze4L
r77gvuXfLAVyn1fIrzS+u0mSIS42ofn8Dj/Xwjqt/0uIwfP8A9PlDh3weF4Tfd+j
cIFWcWzssFlxj0PIrVa6uk6/XxNajO6mgPk0ZbnOD3r12WcJ4nVgex547PfLgyGi
G3+145az0P25kaWjMxJHKd57ut1lvhMDPSL4GH+s171qtMj05UAZU/xH6AzFktLw
mzQfN6HxfFGLwVfoCTtWzNI2HVHluDGz6d+IeaFlySKcMqABZ5mxIjCaRdWWgtgi
CYHTsCv/3hQHa9f6iMYjBrQN309JciPQ6VfleewCbaJwT396SkfJRXpS7gTkom/T
bWYNad7L0Bn4t6wkWP+rWnRcMKWRcYiLotcL5lt5Cwej5bMj0o//5eEQwOfpw4Cr
2ObJkaHqa4XrvDRXWtxsBArgJRuZQ2M5wKdUhAsN8RGK5RUwCwaoGvr0m960QSrX
c+KcjmMyG+X1nxJyBKXqX70lQhx2e0a2x50RKb3HdLmmK7Dg34VvQ2kiRpdYUkV5
FJJ3mg+weT8pVG4YXWnKSm5shLGW6kjes1IGR0e0QOlzUufDH37MxfS3xoFN3urq
mtOxoQxu663FnKTVHpOnU7Prl6iVK5peuyBlXz0iuOSuZAIMGpk3FAhPA+sqN12/
Q6uT0+KlRTwHvY8Biw6vD1XPvh2w1ADy/m4rByy1YWZbi5/6041Ek7czfQt/q74c
EBn4qftbCzHWBtzILzmf+MFNarLycsoXhbV9WFaJm9K55EZZ0Cu5pI83Dcq2YalB
c06apk2C4tYidJsd/mTNIxJCAKjRCckywGZy6cwsrcOjgk7KNajEvQsjA5/BEIx2
TMU4nBgHec07ZTbc+5SOBX2cFDXL0fC5QSyQbzwBeeLTQ3TKjfEjYhaA5BTYViQb
mnv/KUcZOvRROO9mOaaH9JeajljtDU2bjL9WMCbNq7h+rlodAwexQ05Jv3AyBjo3
8hVa6WM3P5UIU96wVsVMpPVkHcY2/xeySbXXkXr3uzDv1lkPsn0I1yqphxQCv4kr
U24+PX871ROTmZXJ0ZUPM7KBk+b/tMHWSk0JN7qInhUtgatVO4ICnqXbD3l9XBfw
Bf6wnpAjcbR1Y1Xz3c9Lz8FSwdgl4IlubHq4lCrWxHg9PiILOKOSJGDTdpM4Uzf4
LSxyirfbeWjmSzOLq9Rqwc06LMA32so6iWazBvefufBqJPLfPa5pfBitfx1OSgdc
vTC5rRd+4+cYgaTsADD0ac/S6yqzUXYsaIDaAYp0KgDpE8q5TvnysDDVKxl4c6ho
IgqAOI2KQtdZJII9TAi/BdpszpOW0S+MsT5RwR09Vjf5QSvEOtNtIRryb1r8IxeO
2VMyRUQE7o4ofRY7TTCgCPej/5dnl2zg2ziucoUdrP5CxOYY9kE1o0vl/XclM8BE
s2fPQzGvoE2M8Bvo98X3OI0GbvCjh+BGh9lZKf5fukW37x4xUazsgoA32aXyDR4b
TkrRwiDn1+Il/3K5L8purzK5WQRI1t4XHnZRocXhsQl3JYPEp8nrLMzZVZRA1y65
Kz+vwL7KND9AWAwrUzbuJ++I1v00L5nKi6f/IB+ov9xOh3H6NUSxKkjnyuqzul1+
s7+wdaISsgfROdunhtjmTa/6C8/jOCrlvb4MUzSl96eSQgNIDHJ7GmQqKNLmd918
0GCIIKgHaw904mj+hZldcBpMDOqKCAt0i5cTCuqJWkdmhnx4wS8TvpVL/SMOlzjv
y2D6HaQI4Cv31toSlxbH/0o9gKBluVjGwWrA8VEV3IxZhlURyoc//VAPLQn++kVF
kBesqnWmzISDduz49ixjpG2PnYaYs7DWsvyFQIDHVDIBvegQrMsJ6HwCfbW3RdD9
Bqtm2izHwLJUyjjFW59hyE0Sx9hZ7gAKNEOQhFXCoTb3nDSRFwr19EfHijnDYPsy
IOHpeqwMeNTbjQT5kc0oFXOKe59LNYOT/NTbxv5/9ynkpL8xeXtNBKK1bZgBWD/p
4c0j7vWbKQ4xeYShFWi9s5eMQmbJJYReVyq0TMdVxCDJnrK30Z0dJOHscJIHjelr
N7XDoIhOL6dDnxARp6cqvMMoihECPyVAHRUBLDhzDetPYfGSVDo5v248o1xNaO9V
p7ixVNO3K0GAuyfOxB2SjW0Vm4ATEd21vQjHEM4gzX6YVfNAazYfzkzmyKUGMDIU
tnritgGtsvH1w/YE1RNDpToRlI7YlgKRkPrhz6YYGa1HuUXG4vykI9nmS1NTWZik
mDF+wsWLrE+UFEftU5+6nHrQnujkDM1ol4d3F/ng1CQ5yd25UAIwWqnfpTrDCcFQ
4oBIT2VlDtjy++O2CtMMeXirtcbYs47xpPuC1EshvtkYqIBlzPUxifNIPEXqL4vU
91XsS5vaSwcXswDvDkJufRe4IqwW4XniDBHEoOaYU3GOCCm8p+PGvMG/U65UeiTt
dLyMMPo2iHWCqnCYf1bd5yF7AWT7P2DDzbegyW7yTXlDuBHrtSqo6V5hEKojmc3A
ltJJ+qFJ0sB+Ys+BtFs5d1i2HDM5Qb8DaP+GkkELn7L0iwPtMomVf8bMqPikRwcE
HPSqfdQ9KxMnlY13ajH/OwnA+1/8d/By5j7VbEeagksmeHn89MqRcNgnP0DN2bI0
zKPa+uM6hfn7QMPqbjYhMThPrfhR9ffiwrssYFHbcuybUQlkgCQOfTtwLICGaiIy
xb/hdfggQrEH+PYw8Uz1CzHK07pZxfsM3wOmVlTZQ00gAgOcS96L4L+Igo7PsiG/
U9kYfoI09iNr/d4iWqVoSO/egN5gXKnsx9aK5+fLKRDAwPXxAg8pSFc/qEkLphsi
Jl6QtyNgjXkXR+ViE+/HfAzNPLWQjuBe6dDzVMR+wsUUC/Sy59gTxtEqP5I8OvMv
YiAsnkAf8fm4ysacWljrALQpeLZ2TfHGevByjHSxpKz/feetjZXGowFmjNuBN9GN
jvjWcR4bfDrox4+oqeYVPsiSzYuJOlhhk9+9OkLqVA4jLYj0FOimHP9sLVjcYTej
9bsdNXyGU9Rr26b0d5Iyb4rBGTLEepdGtGOMHMrjnw5e5nuwbtijc7aNrVPpT7pB
YVRe16F+vE+fke9EQdXi7j7EO2LTCbOMxxMsKqaJWlkeS/eJ1XRX8Vbl7J/whDR7
1axc0PWPwyfr3OH2Uy3MvzLdF9J8nSmHrKOe1dZEwA6UC0jBWRcywfro4VruKmI2
lCTucpvfk22DSUuIZKS773BVlR/qmbLzb4cLzH8Gl/jfAplSa3SKhCtpqfV+2X93
NZuoH3A1Jew5v+oMYIk12c855SrtVmKu5LnA0BCMtqSH5DhhiivyqlhSAhGpf6pO
HDsevP3wE3x2A5J73TMqVgCIPa4UzIc96a5zA06x4nikdve0RHRnhYAPeOCICRig
Y5wUwobmu60xcBZ+omDeSBV2gpT+O1iHDLkk9KTW+aFu6kwfzEOeyObducjUDakT
iirGGAp4WecRNGOHpAG16TYa7wlTNKkt0OyqVpWwv6Bae7n+dgAd8OcSGb1f/z0B
ZpRGy7ZAqJ++O8ZM862fAWGiNo+GjtzBNpvACCuHNNpPJ8A7dyAQR4vNqMQe/tPG
YSg+hN7y83FP7CNhi1l9UogUky3xoBVzec2UB8HHguAR+EnI0S8h4Ouw88X+giYT
izJ1igKe2N9xG6cBp845XR5JE396HBVmZU9M6l+SJzJOxUoVTu3p72y1kyQlAVKR
+NiWM7TkriGh2Da3rSu0OruPj6aLrSVn496cMQGzY61uZpDDS+CbWP26ZeqpMouo
3m6kS1bFDweNvKZgKAKZ03MujE3rK99JKZzHluzwSfcV/O/0XlAcOvBYS1obDUtp
tHh8c3TETVoDnA5fnhl9cSACA1Kqw1oF8AwMe/84I/Il/I97A8igImemgMfHweyR
MJB9xUeiMYQCtJrH0yQY6XIDG9nfCt/Oi4UHUXQXRBL0ZeaNnrRIPJzvZ7m089/q
wwZpFTo3H/suNUqFCNJBu04rcKo19SapI2p65ATVZTWnUWSjZoV3CpTigqhuT+Pc
iXzFHknlxi/m9sMqRZBQwFqQGrz0GMELRd1DT8LlEtwOQbKsUyCQ5go4ev9HWEjI
jfb+B9eQhXbLrMpwhiRYNDZpBSjb3WjMTzkhVgxSFsQE9Fu5p+roXj6OlxtbHX4U
YjUCEv/Ue9B05eFhRwEiax7bj6lXvzFJWRzSgrfnyh/1eW5S0mAp1XB5ORnm0uhI
r+GgD7ZDKVjtHoUtX0VDjHKqMtTavLv9ZohTzIWa1DJPVhKr0XTFEs48+ru9FHre
+WJcnvyJo+XHr+Nsqw34WS3hrYLiSFhtUoK1dkcAxGitdaigfvdUW1InoksHfpki
HMw09g4QLJaR2hhmfGN5VYTVv1/40qw1p8cd7JJ+zw1syTU+fZ/aP0i/GqUWAoIX
tFR3VUAbID6o+7Pyegq03AJZoD/0Ef0KrEybrifyozkkRU20ZYdpV8zB8Pgbza8u
y/UDHO08MWpNs5BNlRIePzqtEe72EOopJ3KZnGi+imddZ5manci3iPpvArwBPcD6
uAaaFx44oGimw6DIuJjuDXKApLCTEdrlJPpaVz7H8yRqppk1Zzo0cdkWkyTuu/+q
ZYAgn87kTikWlNzP0X0XhqGZN/+rlgIEAuarUobVBp4+KmlGAtHKmRXN3nk47eT1
ZgSBaS0vQHHyASRpn8zeIFtNtv370OXAFZrMUoavrHUE7Y6rMJ3+SVdoWnYT0wdA
/K20QborBr2wTRZpYxNJ6efmKmV6wxYX4FyzxL0lXgufe605jaWhA1lnvIm5Aijz
i+Af2GnM+uD0rFe8jM3woWGu7349e5KQsApH8pNqqj0V44qysU5DetrnpdnWQEdB
46wlNUsLthQcR3kMluX1uIhcZIdakjxjSvGwam8jUJ4ezmaQA+W1/whPW/rN17Ve
jnKlQDipNUIl1PUPmLV8/o00k9bm4gNsa/DRkv2sAga1u0S4kdJg9dp2yRJvNReq
HOgUeKt4bnInjGHsRtEoSVJv7oLbmZ2hbIjE9TQeRE7aSHw8sVP36uAQqOsdD65I
BgtTQgL9kW74cKDHOLI2mh8tSH78zAdYQxf1GP/LrBxrBQ2m/ktHYKWErpsYmN51
Rn7vNQoA7c8TQ2E6zMdZJEbfp1lqfMCuZD509RiBNvUy+B+nUp9VHmZdy2KQSSVs
OdPg367ggYWbq9W2rOP8vhQSQopVj/9ggYbkfMrJsvgMTKpMMpCHhaN6p/+IFyJ5
phuGldnNAID+/AUEFKI/g4MaGAA+AxWzhQ2Z8WGRqOFMA+7nOutCSe4Id+pIMHCh
siOdH4Ye0HO0PkSUK0WzXvFsvd+AHsSACD/WUBGav1OJKvzSxXTXGl23ovBfxl0O
wAJa+QXik9U9yMeiZ7922j0qiEaHU7vUl6Z0KbvN4TgrFAWWs1Ql/QkJoPKKA7Ki
qlBif5Y/9AIjFmCLuhkMoQweVmTs46Kqmqn3ehoYnpTAp3lcki1brmAuf1gr02p4
eFKUaiwzxJj4FbdDuJ7yq82xidpJ0HMFEeris1XVH5PcHKA0skmCvLVocIDRwTO7
KcE6ccsqaMyoUdq8bvxMOc6RLMPEs4keA6eI+V5kt9RG44EhFoY2UTT55qMG7Gun
GwdHq/pvJbfR3fvb9ansqrIA79ol2alYUPKFhz0dUXnBYwpY8uJItbm7XTczNFKD
vHky5716Yu+wejXSAtRL/p+9bh/cSJPYSv7qe/4nuMRYJ7Yz//6DDVTOEaIHyaLf
6XQyAKWhmqfUfb5XhoiECQIYA1xhiB5UOkRti7+jDMCQfmy2zFyAjiggDSgRWG2L
wyqoxr/3fC9bvJ/y8p21DWCV+YIzg+PD/55N2evQMa12guv1nx0Md/XK34uRrv/A
8RZqA8g4abz9D2bboo/EyKFtpGy6nyzmI/QMXVRG/xjF+JuAeVMFfnx4FRkD25zz
X6inzLPaIhe4DRddF8wB+x1Y1gE0YTUIa7t0lExgCOQkRY0LazNT8X6fV7FzhCco
ijw6FjPNMVGaHw+/ZTTt51yu+bA/rUz1YDWaaEmKCXLUutdKcimCNvloNInuWzeM
wjoTZPIRmscrbcKJEei8njd/ZKJ5rEV+Nj61eIjnB4QVeswVr4WKHVn57mV/hG6C
kz34MOgW/qlBGKj85lO0D160uI67RjZUagA23wcz7uUeSe6KyJDgXvjrhvBH319l
dNuldEMKZcCT+Gv8HTgfL3oYD8qKYgXMfQmFVbThHFbtT6xi+7ZyE+S3H0/tUI2v
/2HYFguH8bgOKnr+d+AjAAa5sg/ZukyTol4k1sTxcfK+v5pIlQHezmFD7A1EOlBc
3aUV4d2xnxZBV1jE25e56YWkSXM6FOvnXyZ9IczjZtpruZoarKN/9T2/sBfUGMRd
YN6NUTC0bWEQxgb8UroJYwKxZEAZC/Af4gSGNfK8w90vBu96mqSv+052JbhzXWOz
i3401LXazH6GK74114DxyLHbcG5hAP3Kp0bSxcn8LLbNU/pHIBJcqbzjVcVjFRAV
/YcI2vxK1CoYtg674+hMmKz2MvSsVhzHHn9ZrtiU7utOAaEaBS/CCmWIGbpJ8v2k
/JEit+f81C4GxP3mLyv7hU+r4/Ibs6KWKQH1wqzpVam1o7tlnuWmOyXFxf3qQsdT
deaR0kdYBKVVUezzUYqZq52g47+Qs3uFRbncZTtrKMghlHFq3sbrTFR/MdsH/z5H
oTD3vjGhG4DA/JgUVZgEY/2e/Wrpg8pk/vA/mzlN0BaSDl35ZUYd7DsrbZCdW3EB
KP1NBuAWFCDbBROw9hhx4/AdflEcEPbRWfwsjxwYUXSZw8BSnIYIdUht+qq5/8sF
DxPl2mcX3029G+FakSZD+LZ+lIDcE/EUUhQk8e65px8Nc+God6p/g/SPrXz3lcas
ggwbQOaghXfHRaq2TTg+/9K0AMddi1+9SeqBtXNq1dTqm2r8ozQl+kgScQGv47go
s6noyc+CKz6v8W2LwrYAuwsU2cJGajhBlv1jX6Go71SlgssWm1Zc8FNk44QNs1Ap
eOggVOJhHf8fXubwehW6FptCCTkOfMHX9C601hXFLEBbPUTH09Ze2UxUoxVX22LA
ZUoAeafufB4VdYpeQnrR7TzIyoaCNEmLzSg13xAIVI2AfvC+scdzNdJmQvJVhpR4
tBHYgXIfk6nqJBfMSMZE0DNRxEiGTEb/J8mDicSEYnYTwrvXYzvHxXmtLwBBjrPk
6EepOa1w8G4ldG3AA2C/SgrrG9iwzMpAi4tmB1JCv0BJVbYz9AvZ22Uy5ZG8Dysb
1ptjVMgk3yQ2HIQfpSVoSFXGBpnx2Js3aI457Vf5O614VTPs9fBHNuVU9EeCEdOU
wqigRSgiWSQdvCcwwMNyUejHCpk+c0D+PnQJ5iToSyvVjGX07jkFXwmQ+xNs0RrF
ItVE8pfsjFyOKEUIbjYzANZfXyiZg2VfzlxbER1l11mXjiGKz/4Ivm5nrnLrUcw/
dLFE32wiMaadgnY7CdC0f0wY6tSS5PrGuYTolGc5oKor/ODsQ3BO9MMOaYgncPit
KtHl59kioGfVOzDJ0Us5gW09+Xg7umkWwdIGt51G5bKuQBQshbcelPnh0ZBjD8IK
MRuoSjSxfT0mmaEhRmRzYyonr6q0aGLpuzNIsWepiHoTFCuHWQSfONXWxwshE1DI
pr2Sh69V0DF9Voqm2BLSw+vzek+jDyGdsjIQ05Ut35BRt1CtGOL9S06Hn2AbuoU1
xIwf037B/KngVirbcsEXIBr7eb+MWWQSSjnTmzD88NXrPfCZhfhClqvCaTCg4de1
5skCqW+izbjBymAMFjcl2Mwegpgb58uGAbcAScJ5n3PdOYAHrrVTwcnNCDPKaQTJ
ayXNj+9alqzSYRo/B/HmnUUVqo6rHFpHbyMfM2j8gzQXrkHL/PEregwZOgwjSOMZ
By97ERU9B9xL1lLU3N9AMdNpLz/0/IU0xxu17Vb1cPcuvnpzQLHgndHXI+2FIjKR
ChdMdjPbr7VBZoI5Cr/ckSwKOBs+e0C7AdGNpYzub8aFeeO5ueA76bUR/r/Lif2M
BfLCfUhQmqbxcvwzm26q5A63edHG/MvyhQbQL6X7I3F00++XOU6YMD4r2kaJKDN7
cKZKx/2f4kSNSdHsi2AxaqMhVPlFFQEPUnXk5YOAfOlvzGgmKuH/g/o7rdEsUrHc
UFYfZxvoPRwadvwqo2sHcKMG8ZhCIynTymyqn2wZIc/0zD7l7LxreJgSodQFqtIR
rTUmNUNq4WGo6QM/x5ipQKgTxF9EOlFqj0BsUpcmUuYjeUdhtrA84XC0+NEorW/o
74BE2LzvJCXkXTpBXgvDYhvn4LbITnraNtxNiksU2OgZA1o2OwgtuNSjEb024Tx1
A14yC309eFWF5VID+QH0egiDus26hAFJM9q6nFXbw/x77dxQUUvhWirhwIqPRA06
BHOv83iHh3XElPivUA8l1kMziIcaRN/5RUt+ymHQD9maPvguawlPD4P/CXti8ij9
fSvRKIjMNQ+0AVsb3XRvhrezB4y7kw1P/LGTRVgnDH8kgrB2cP74j3bH7ziAUHhB
yeESOsIJabZYIyc0472BbjL748odwlhWpqALgqvHkGBXCUbx33Qst7r4gZJL88cC
k/0UeN+oL2ajryI3fEzvg2z85Dbtb00mcqBk6yELnaRvx6aaW4JUYRrOEtOldbj3
I9kg6eqCfE3+8XX64fUYYLVVwmByx1i2qZoyxSfPs3jne6AWP3pTkzSVCArXLom6
a4QLtL8ykbrFKv3ItfGldv2O9b7rPhoMC6+SzfC8a6khXxdR3waY1NfahwONSsvr
ITBWBHgGiCb0z8MnSjnSiEel6MWwr+0g3ayawXq/4R/U76sjILgGmUZadZ4LTjBu
mb6BS8rrFNXthTgRUNurOoYa2Pv9Pi7QUsbp1gdrjuWNZMFmGv8qKc/t55Fcgl3q
EPzAOkaA+U+zC10AsltajoF6jCsMXVcdNOC3BHowfg8Nxrd9WDe6cv+kTTuiSBJ4
J5+4qi00LQ1+uowB2oyNOSlI8gK98X+ii4MmUgNyFKJVrpvY9Sce3zK1CpCXkaeA
FBo/K0HEwxvgFzC0zVEqXNNTCy2izST54VgfePVCBL9LZZfqdMRxVnYTrKho5nL9
E4iLCosOmRtHtba5ibuFHAVTLJdeoEcmGZpf16QY88TX96IrroYy0T6fI89gUH4F
6xT0hhGCkX3yAVVXHN7s0nZres+npx0jLe4Gw11w01RF63hyhNzzbjvuJbN0IEzw
pQI76OlxCLz5H/OrjrMukU+kIdPiovSO1+kvzElhXWDBoggkpnGRhlzVLGL8LjEa
/cZoYkKuLnDzO3tc2NWK49yf5zx/j/uie4MWvv4Omh7W5L+7csIVeUmEWhg3c4o8
aB24AzC4lY8j53dL3+A5Xo/GpTE+3+qVFxXpELzyJcdv+CfFY4Ge+dbGQUE2ysFF
kGh+3P7UM8WXKYISSuITZCsri/QMcfx5vNVl6k9svh0WQr68N8yKpPOmVjQpUyjk
tvMS5aKheVdj6Ct4T7+LvRrI7DlUxnqYP4cl65ZynUBPh9+ZY0nH39igjvgg4MVy
A6jndvCyW/hB+qCEZqWB/N512T+WC1N0lwwGbfeuNQoMppl1cewkIKhMzlQMxUJs
DRbLG6gXTBEEUSbJsc8laRokoOFaM4q3pJXuwYatccv/dnN973N6IYxplYC39XCf
LCqyAq70BWMrbGBM46DwO5Iq5k0v4BK1x4ZeAx2JJ4yVzRYA6qPaS8LjXZI1hzAL
QP1j4Tgw/7y+/ps1Tmrs5vV+vzozR2GVKJk20QYvShizcaQK1A9KYLQmpWvy+Zyt
7F9HiU6U9p2LXpbwwwVBouZRPkDXzsX6Gy1V8O1cuB7DM068NrkAJNOCfWiyAZ3c
75iaWJd+UbDb3iT6lfDBjzNWKewtCCXp5PS1TBbwbHdlrnwYX33ECPZAS2sR+hxd
7jJtSvJDiDpBMJ6t2jZJlb5YYYFJ/c2kxY1Scip0UuV8WgOo+xyEFVuwjo4z61WQ
/Gbndv27YvmqIAQmMBWiet/eEVjh41mIqjE0SmRqHyELJXIr1P4JFXwwDmAYyXH8
hcuAycP9x43jT8yCQ4EX6AHsBNSdQ4CPprZPHfyRkHKgEttWk81sXUXf9HHlGgMO
IkWoEuJK/egF2ZmkUBiwhacnWNh+oBRQcsHl9gH/gXLFMZVdM0Oh5GQUh69u67fG
O+wwwAbOSwFI3jzsSyJ4E5o6MTC6/+LoxWWJqbhh7cG2/AVykaacJNUDAefrDiZu
yD5MEgS/gBhr8Q5oL4oHPw+a/yFebvE2cQCbEldEgSPrGY4mQuQXYhPEnEdtr+h7
9nUdPGE1prfhItVJHChU7QF54JrXbdcL0wunGDmlEAzlcEmCNQgKXe4CovFdFCmo
TKSTjM2E3lUIspD2NecG6LGD4hFKXODoj9nphVjG4dhfUf7sEHQET3LYiEs+jSqM
CZPqJcs65BesU5x0/+IWXE6e6SKOazhYRslqN5GIUtdEhaxjTwTc1/rIcu3ZfxLE
t4xBJM9XLLkBag6EfeNHxacTwzLdkugt0Yh/0sn+6ZSAHS9Z7PDAmBzlg+YEHVgh
8fTnAQYY23M1DhjkoR/DDaMLz/oau5WKDjrFPVrF7cGEhnWtskVo77shsDyFCQsv
Cf2q060aF7b9wwomZ9Bq2O04neflqoYzlc4dVsc/yOiEPCxFa3GNoRYLZR5wadjm
pmULBlqANe0opFvB5oiKtQsAZDjFvdfayo9vT1bhY9hDrTbasM5r52sEHzxMWg9h
VFmZt8CPmsmqCqhAWJw/EJkR7za6Up6EBkf/hiVYRgw7FVzNkpTZgLGyJE/5SEnh
O5qhOYaJ8zTbiqjypK1nURZT9UTA9y0MV54k5YobSOdXPM57Xr3kWAbhd/T2W+N/
t7BZ/z3TduTCQ8dCSQSdEPyjbO+xjZRgNQnpnJ4zia5/G/kkCuNymsGSbKwjeNTt
B7WlTdpHUpXa7VLPGWjT1qszgUFWU3ke3KzUt0Jmu0saRUdjfAN4EVCp/XmvPssl
hveMMcrVat8wuqzaao9EfUiusfRS7sqdJs0ZYEZAZ0BloLof8u6QRt4bUfkt1sIV
OVZkb6fcfjIVPNiiY39JyJDJr4AQkslI3enXY1ei7qOVgu3xPH2UQYO6OKJXo25X
oC3An+3gviReKhK+R7I359xmeMvuH3nOCAxWMhLWg3qwbhXOzdcpL1zYVBzmsU/w
S0sZoNjXaxbTo6sG16PNbbQeVuzgGuC+s5qpo8aTpJkMYaR8rBroBNJOkV2q//Rh
00RWqx6GMx2eb7NoE3R1beMaEB7ZnoP+DiECo/C4V1OvINtrPrqEP+ltf/tXjDqV
kCizQMsmhEPPN5ZoO0H8SzEQTqIaiftj344vicUMNIy7QpWn28vGB5reuK/Rnwvw
E2PHzqX9bSsVN0H7iVNCLkZiB+1TM1o0l3haLEl9FTmzme3pl0PIhHNZb9WIlGqp
VMlo6ow95NuF4CotJBUYTWEiDfAVX454vqFdvRb2q+QBXDcVl+/ADJXcZKiMnZie
svoPrKOidVPBvQ1Os8xXSDUACqJAG+ZBJJvt7qDKiYG2d32Y4rrgZWmR3zvLBKYI
qpbII5vRe3+sTrekenkjkCrXGJrKXmOl1vDPLHNP4QqeeknKkkV9Jb+atP12jeZz
Z2uV+m32aMSOx9Ir/rpyAtF2WP43zCJnS1sygBSMsMNubT+88edRy6U1zMKkiwzy
kp7JIYzeTUM9cT9eIkCxAX4i/8AaRCHTxCtjDdtP+WkStmMvvNc8atITwn/d67Sa
9B4dgVt3aogowdYiWeU9WNaTK9WjTuVcPjg14+dzmf60EjZjoKgvbQuzXFjpsHS1
zkgZA+unRku3aaoABE107ximzad3SLN13e+kv2u6/e7MorBU+8uOpsDdqoppI7dz
3X/KXpChA1iV3+bK8T6ix+AOqRB3Xk9qJo/PbjRQRaYg3PqdztpYhJXcotNQDDvm
S42Ja7ehOmSbRa34ufbvIkxFVs0RvZNksp0DbHaacVKZiceA7008xPE999tfnW0A
1PCFJu32F+/ils1k3KEimZUfnUHx3BJAnp2PuWZpaxal27Y6+FV5FmXQFy+As82q
OLm9Wc9q6ymzgYkUs9AWHQdL+vW0aKVS3PEmCmmErMhko0D8uwPev6+Ptt3wZC5C
sjIvRd7U8b8brPkUPzTSpkU69P38YxtgYUiK+4Cc/Dhjd7SGlamMYqAut8TqEw2r
0fTV5P/UrgXMyhQQdgF//v0saqMk4IEctEQqIwaoAFwcICRUTlNOToofMqxKdwtI
gyKSPKH10V8e2EdJPsBqjOSToCPTHM1OhKRuQN98+cz7Ed7Lz6u7azIlPvsuyKJF
Z7mn+0WUm0w5YkuijkjIuRI89FyfKFEjfhrUuSvi9PoHOdVK3kZUTqs0cTv/EtPx
3XIj+j4Q66LOJ6NaraUpXPyyP2p3FoFAGz4Dm11wT70Z+1BOM69wT9nvoOz46dIJ
42pDqLQ5152exBk5A776ZAYFT3H9zPWClVEKppCblHDhj1NpM1/+z3yyNM7Lw/zR
e4xUwyAATVB+Zy/fAWyIdypBnCzNLoGiT49LTIPIYsmwORifQrMWp96qnVHtns4D
f+glWkK+aYs71izK+MSG+2iqSOzo307nXoRjoez1ZSo+xaWgNlD5R+wQVgA4Zws2
N2gurmjWzX23aCsc3CwgFkq7W/sN2FuYmBzdfX1HsY7hFHw+6DmvEzhOhAZYDmq3
F79LpuqWiBHvWQGALx1lFuaJdE8UL6ZLZ1K9QIUMrK9PTxyIMI6GnIfqydFFWkQK
9WZH9enNkP9xKcceJDF2d/b5dE8pDK3YjAWi78T0K2O4By4fyi3+I0BOorxJsi4A
H1XUu+KPoxLTWGROQyTBlfx3ui8JUjd+aqaP41k8HhZENOqxsCbmcmizYZb6TNnc
hSMOPBzKNtkAzUIxa7qO27dj7CnEDYy+QXb6iY2nv0iuGcH+a33hraWzUocVtKbz
1oun32/DP2U23f16ge5ZW4T2Zljtdqo1j/xw56dwQMPZS6MPnaencfPTDph41gcY
bhVeg2Q20qpiHuBjNlAxh0pmQG6hQIID+mdviLQTj/9R6qGaelt1y9z4BK+wZIs+
qZGrqJiVhvgQdb8Z86VnLYAmP0snZP9p2fn0Gol7hVmMcJ+I0Bx81PqRcUPLK+AC
5DAFGoFtFtGqAN0zHQsTMhKPWjFgOnEOSQO/xeKs0PhZLi5QiA42EFEGS+8CdofO
6RgOod639dx9Pj7nJmAitZRYFuUxcWhtgwkQvw61DpOJFoJ9EQmwD/nf972VN6jE
8kDpmPr/FQGhEJ/D4KJCxRdCCp8QlQ938r7YKKJqVtf64cAFcc2sl7yaNAjAhfhU
f1cVIWnGwR6/C7/BlaLlyMBLBKEYs8SPhQKvm9D2AZvcP5EwOh9yswOF7uU35FdC
qX72wy66MeVckCR0DuC6IosGGWunD3toQmYd9X224uQK0JJNcjKR8JNqp59Cf9RQ
TnVXczBGzRpCrKPKdyMu8jvPMxgO39WmtmIDFRoAYzAD3ikQVQosd+L8dmgyTwrV
1D73HiQr3t0qbUHasTGJlfwyUv36/7KXIM7cC9sr6VlEoCvazdMnIkCbLkOc/aIJ
sslR7PLu2liZ/L5zcTltb8XMe7cLhnbGmwoVKetNlvewQ4BVAURqDpHzDmmAeXwl
mlTwRT9I5eN1qaScBYh664xoqagqOxLV9GCSskdjr6yPxwFcUl78p5XBOUmTrdg4
sbcAtlwo59DDYW9Fv62OVxY2hUTOQ3p1aTaO1DIBY/6Bkp51eT/xMqxU95DiAYwn
HbOpO/Pi9vSmJC1uJatp89HyxkgkOtPwlJjrsaKADaRFx10IlbJSCN7qZUZzBUeo
T1jXuLmceP6YS016vQTsUId/enJvO4P+RxL9GjBWSUg6KbQ4mgac9oVBkI6pIquo
UrNWNvJEghE3k/qvJgrZwpug0CCPDPY3M12qoOPKBvM5zDeDzcbf1QUsRZDHbp6v
awkRr/SMWN8XXnD/W5fdKpARyYQrwo0TeAHsCxLm1pvVAfpjryA1SaQdlC6lZpXW
5fSbvJj1xGInrr+cHsVBEyp6FcZYS136Qp3ZlyBOt2QlsX739xLKhDCM4CWv5xCu
YCnjmL+JoqHC2/QjMks43BuWftLp7QkXcO+dsG93lHzaToLhj4RCiPC2sgEKWnKh
dKvKoWXuSijXXpDvX5FbUP++lPd9rKTKpKvjtw5rXwxAf31UoECT6xsV2a0G1NoF
1HVH5efI8sNYKsber3Mx3ExBWkPvKigMP3f606IqjTS4T0UtVKA7aS7JyP9iAxFt
oOhHRyYGqqDnJloXOK8iGoAZ+cWwuaaG0n6RTicZ3eqXHOGM0q87cDqPsOtKIzAC
WVn//kLFTRQisq190qvJEQSwADEH8+/1jzieSu4eY4ntWBKkDWyu5qoDut/DvLCX
ON1LkxP6jHAW2HC/w+B3pH50EzqrPf3e38LiUfk4ijaTWiJL5zVP9fdHpQM7g4yx
9qIMgMX4xe8sRR64Qz0Qvwb73pxXQs053eWNLixOo8pEte5D7DPBNrTj1vPiUjdd
vCPb7hXAbXwK31s7DLXCHB1EcrIPWiVtA28JBwOkHD7MCvHXP0LDebUjCruHdSu5
LRSvmqFb4oaI6WmxXoa+zp/mRYmUwOwVDZZ/X7hSzrlGTUcql1k7rvg2FX3Qv5oU
vJArnrkAQPo2hKAcFxDLKP2UErejCSjTM2K3X8M4MIi/PSKNIJTbhpGPwUDe5orf
DjqooCvCrqt55Fj9xTF9kCjbEO2ZiGXQq35jOu3Z2V2FYBaw+hL0VrbNwyldW3BB
tWxBYpbSPP8uIVu7P6gRWT/WlTOm50xkw7JLZOgjwO/d4GWQXvfdKHYboLgaTiVs
CQdWWsZ035jfUpNkBOdwOI5Wzsl2Uzo3CghO4CIxdDb8FlVHtc5poEa3J5t04DO+
/pPaqhQTijuhdrjaAMb15xXOf7SQnOtDdLZKUaYqlwNtIw7hpNXBDcbUK6Oxscli
CMjuwBkDWiomG+G8l6CTca4Tf7HikZFdrYtZEkmgqzY5fTLe0UNKO8n/TEO/nFmW
0T92fBUNge+znC8lq/VeHEjjSgYQbduGrn0PXfgDn2tMWpCZxnWlfirBNiYcXBAD
LtPAAMoLO4jtERwvgAwB3Hhfx7h+2zoTp3TeV/HlfhzgWzntKp4tu0J0H4WgnG7f
SGUiP3gtJhhWFFJcdq9X8BRq2sGPQQmTEyzFYerWGPW9L1SBiw8fcer2uVMOAVOI
bK54B/f9Y1vn3fL3TJR8NpxsQa3TDZ0XYQIwPxzH5tgsPifPJzRKMkGGpaz9CuwK
AJhw6spzWWHO2BaeoYHBIGL/UUNtYw5Kt8XjThYIJeE4R+ctE9uovqjkDhHQ0mdr
jcnJ0mQKbptGcRc0Bm3R7EzSYYjB5cchaUlr4kcY9GQ98RU9/niPsP6wL0zwSnmX
X6P+9vuEliN275F0yOr9mqzSjOp8KLc/iGN8gPDDazBe7Qy4Ddpr9eAKGI1k7yLW
UEfNqUEJL1kjp690I5QOL+25UbpOZgFzqzy7gl0Prb3DgiwPrJpVeoVzmlya1CjN
747DHfkNVpBmW7dt3jyPsfjQfwtRQLDOuZS5xn2rQJozZAkHVkoBBdmNn9JOBc7/
cL/zp4dcRlfj+Ldru4ZXx4j+8AW+d4PFhr6gCv2EAvFHbPTZ/0CmJRsQZlR8WfSS
lSAnthjTnW/rPLpKIQJnVXKY6PlSWvVk4m+SUX3HP5W4EbxNi3OfMx0jf5hofSxp
Wtg2i3HUfGIF3wh9uIMlETDhGAlGHViVeNXlcuDckDcQEzN3AtvJmDDj45gYEYzo
3C41qwcM0lovZoJSKe8iVUKOgBEE6zSFe0PEVjj6ZxFVG6fJjhlcJrNPP4bOer0k
Nxs8EWvdGOfP1UBVSGs5cJ9aizKCpEP1+NTqhAVDQZBL7hStKTceUNz8dF6/onhy
rFXzBlVDcsaIdj1QSwzjDPQPh9Qm5TMFwJCH0xiQ8tv2C9y0+UhKYWZmFvEf1gcs
9vuLBuhqs6zIkG7bqppBXxDjnY76E4Lw2J+0RgEIWt4G9r4aKyV7I3qRHdl8m8Yy
ZEMwx2oiPTsPQuaPvuvouD2H8WCwdaS4wyRNlWzS5xyc5Hjaxehm/Pl0STUovCIX
R+zOn2RwAZL+W1QF8o1xBmGoIC1NLfRb9G0jwpQQqxkyI4Y8md08XxalLn89vGJK
nXtef+1WWALNeRzUHNkMfTrvB7zi7QbLlTj4ZdSr1wgMnBx8b8XKPpLZTanyGAjp
wEDH7GTU9r6/Pa0A0hxcWu6pQdHBg+B8KRkwXZ5afQEQRFkICf8i2+bqlfGB0sbN
ienxTozE1JgRQvx5k5GiaWYweR2MN1cD7ojBOS+AaL+r/lcRFr8K+GiiLnNNyeAR
3vRXVXwZD5QDHil0uoylGxqDWp5V4R1qUAWL6wIi2QXMftJnzs1djgCSYQIFUL/b
We4aFzyZHqLumYrALtuvuBiWvrkaxkBL4z081GL3rVrnilWMJMVoIbAsHoSyRB0M
yPRt+Mkf09E9dCOwFGTi5P/bVvwVNP+MzPBaNeEAB2Q4sTXPgH47Or9YwEwcQ1TZ
+YiW1xAm8mtmKualgVgrhmDyKQcJbtt27laUzOrsryTkERZWYCxDimGW6EhmpRfh
RxZzfpwmSJo16C3M3bPE1efEhN0G+1wZtrlFUb2fOOAYbU5Api4j86yOVtAziYuU
jefzq07npTu5IpB0ylcNn1TYWG7WR2LaaRbHqtILZ3anietdkOENOuraUQJZqYd3
nOiJ5ndNop3vCLxqpEKULOXa2MRiEJUn2MzehhEncY4R9iCBW6A0cyX1qzbw/QwX
FQbTiOxN8PVlUg7wlIOIa94F6zgnxjadXqqb4uuWpE+Yy4POOpxyyWoxh0W70wXa
2LPv9UAhPFtXj/16bfI6tDeJBZTo+ius/7tTbGyFfP1nXASJIie4pWeRTkvaJ6j9
rBoZCM7GhjXijXprKdX1LMFKS6Ay16RqevabhoQA6yjXgFRXI5IGJDOBbXwCUZUs
nasZ9gPzyS4k6XRdjznynLYgGsGh4eHP5rLzEBPZwJNZwFGq9zT/hCzCp75xUMN4
6s4cpWJFw/8fqDNgYUmhxbC5qmNuF7xffdaEAKwT33htwamc+EsPY+HfmIS0u5AD
PyYoscfF1BEv7xFZBNXWSJJ/HlFPLsb0BsQJPy1Y+V4H7y14R1yX0VOInlDmRNrH
xD6reWul0Ms3EJaO9gjlVlS6BTMxlomdfo7zzyf5bXKYFomva8akFAS7dTUpFAwB
15jwFmclxz1wEBBGhE9iH9KEDu66tNy2jEnM8xfK+nFKURr+lA1m4niv3m+6h7NQ
FU0KK551EZryB//KIzkTJEAYN8Axm4WwUxK3Uzd5Cp1skoGVvFs3e3+msuST2c8U
LswNER79sR5wqvpFuyFmgT0z4ZxMMdWR+6VKBPhpohaqhlOBvEwOrF1PW1CW26HE
ugfMP8A7SNSqJsYaYh8LApQMFtzFaFak+opsfVQ04jeB94tV6R9qM6Le4kYC9Bfw
mzXgUfbxqwUcj9NTKSxmap7ZS/tKPFg0sT9+Wb09PiTOq0Ka0Cet+rDBOCAizbji
myEcDZ0vregEMrmmnukmpXmgUDBYYO5XnNZVkRg0q9mGxNDR/vrzEy0j/lghAqYA
9ZP52xMOGhcp4SOTEhdwb6g4KEZOprqpv0Zwtd6yfnppLbneL3kNTETxz1s1ZZ1Z
eMfqFVohxfAkk+3ejEt97+3fWyBLysPp7VKU5I178aUihGdN1oCFFIET/cJEdOKF
uEEGVx2VmlBpPvuoIFTeqdt0fIotIQ8l8XhrBweb06zcOj3HOsMww+wbwrEeWi0F
DBAlCFFtGK3Hv5RdoleD/JeNvmZpyYwyfXckf+cCaCgV2rL8ZIJTBjczcR0sHBX2
tXYB2JP5chQUJ2unbtmku3ZGluosekTrEtWkH9cBj0wDxkmtxYvysg8wtlk5iups
nO0ZBOLng47unHtBOwFjA1nbxhtrPKRyGiR4wJdml4zBoYeZ+zOULf8Y72XMnnzZ
Hce7ydTELT9zHvqVHjufPVrG2WFDCiLE+e4GIwK30VKK+7a5KatF5EpQSGCtNWJg
gl28CiLGSV6UIyOaH5IO7m5wrCY70cN6niTQ1Cvw0pY5pfdt3bwzoYvo7T/I+R8C
/1TGN6mo1U2oscDTvlhufUq465kuLr9j2N+78EKpRjX7kjLujUM+wbv5QCQW7eDr
czPa6NKKqEXYZ4iqs8/zg7UV9zH+NMG8aw7kS5ru+U7NrJd7j0lNf/jHZTU960AE
PrUODTl5WZwFYo8Y0c3KKAOVT4U/Cj72ubMtzftbm7Ll0LNIXYw05TuNvIHshwoC
ACfNXmifaFJ/qSizZTnytPEj5x+COGXcGlcPeYtDeEkQ9GNz4dlzM6aN0Pe5g9qy
5rYSczarxNNjfIzMUGL7Q54yMrr6OXZnmwv+Nd3g5UL+iJMPy9aCiqkMnIP1lucJ
FBz3kgiiCS+qsvUgsFKct46Rof4QF/8NNYOYtuKqm2HNzRIGY937EW99A3kyKw9N
HMSoVpy8xKVEb7kka9XpRQg44M/0RJLVpFB52dZgjfZXzM7hv8v2fecjg3p+/Fw3
p4vMGlG94UrE/4qkDAxl6hoKo9Zwl3qGKQsRgyd/UIcElR3vZ6sEKlWpH6zAu/Am
b5P71TMXZfjEC2W7br6yuwlSONhOPMh66KmHMKG2luxHYRwbsn0F/TR7V0F3XGjl
laIu0aIoJnKqh1TILhh0qEvUj/BbPaCGW+FT5ks6GDa341Xc8tYOiNf8Db1o3azT
+9y06SkPaxEVMwG+djlzaSLJ7MQgloX+nGnSNsulbVUPXiaYHp94VDa3t8z4bpbK
ksnAYQuGhSE7ikMb7YNo25A7lTibmvXLmgo4WksvrvUpClt89joeDS2odzE9vVVz
4dicrPv0E3zBuSIkPgIspRAyKJMICpuxpzPTbvWgay/sR67LSmPstNQOol57GuVs
LGiS9QzYk3g8upXWUr/gvkljCHNeu3CIi+44P5nDFiLysVpLBVJkx1DYc2ynL42W
cXS0TE7Rgv6yKSsOm21PfvMHt9kG6rcug7Uv6VqX30grfkfMWOFQQ0JqwGUbIPzk
u18JhjBJg8b+f0WEErrn0wE6X+AfeQv2Z2nJW90cqAv39Ken1HrVMyJ9Nf0U72XY
z0/y3RdbnyMAUTgn2DD/Kz+0aVmPL9F9k7PrZLJyZ7AxJ5fldEiBE7lYieRLhVbT
2ol6VQmuhHbGmsUQ/pHW5Gg13TmA6s4L02F7sbtLLxE/A0Ek19Sw/e6RH46ydah+
cewgQWmtwn/DiuOQ4qKzMZpQdAirxYE1hYxoS2K/wwm6sEvBC+0mAYKjq5WACEfr
Sbom9tNY/8Rq9xY/ffniLgnHsqkk6fm5h8pMv0VEuyg1hKoZaeSg4LB95ld7dYVb
TakvNxfPlyuvUmkpGH2tng3/zrQUDkyKIhPuAS2eo2/7HupQqXpPHajv2/LAUdtN
sFSuuTuAzGfvtrhTiRlCGV066zTb0TB/azPeFZs9fHCDRaLQjqb0ZwQIIvc0oU5l
M4HNuJEnRnPwF9smEi1aHdJQceuPZkBEbTLDW4eCh03YwGqdPOfPqp8d2Ey+hrlo
QAJ4XrBmyGowb2RQ0hbiqfLh8rFhlB+o1nuL4VQPsBwgZcxqnk4Wzv48yXQ2Njyu
caXU5NPxUVl419xS/I2xp7KbpnKI8GfFa6GhEOcUNDzAvPMounawqm+gfVmUHxmE
KAq6k1Z7NPYtyhdx4xDdUIzWEAbI08DW8NvnUMfGwvE69ctivu9a/hg5t6ZCvClj
IOoP9tXm5s9reNelF75vNzPHjeU5MFWmyXDwNNGJ6HB4a4xGoRpInvUpjur5fFgZ
VNbvB0WnylKBaKzNDE8Ehjf3lI2OYR5xASRJUZlakOxifpou0LmwmhdrLvl0M1Hi
uF21izbprFwQSljrNwTzOkTiXvY2nN2UPlr12f5dZSEEkI7D9mic0n7kIU0o+99Z
8pq/Ybr/gdI0y82lREzZ15K1FiliUjdN+BIRvbLunguvLwKSQ3BlO0G+G5HBG4fM
4yEvBAMWN2vAYYDhb/EdBr87qT00OA/pgX/+XXd6TC8RMJyfwQ522P0kO1r+qSAB
zR38+3OseQuZMQ2DLmoArh2PIfrf5BO98g2NUMjtUknGXL8V8Cbjl4+GljQmu5R6
+q88DECTm9ToDFgt6OnGKxY1kVWovmSib6r7mWjKk73TqBS+tbK/GQYL9p2uRy3z
PnJlzz0tZzMN1pf5jwvpjBpTyHRKc7Eu2cO4eUU46pkADapGwKtKGVdVbFa8TL/0
11gsnQS8l0trn6EyVHD9uM0FPrmzIO+U/9Llr1zv0GO0GmHfyBOEOz/vgsGL8cRP
HNanrvxR34CMOonJGZqlKvsEOiluVr+8cJrzvjIjkDW/G9Qw+PVCUXTEP68ON9vk
ofdbnq0/sle1JH9YXJkJjBw2Ew5zXDUG53YEgMj59N3xhgI050AhonXeBx1vbvtC
G6VPaQZx/YHhdKaqJnL+8FFtyzJWbFv4uREJ0V2Lj3wAKT2DCZnoOo7wWCFZYk45
/pnQx0dUASLBTOVeoQ2+1KQ0OozPFHJnTvMOaR/KZwDrCGhjHpnreNU+Ho6FKmdD
WqyPiCBLacetivK94KuaQJI1OL2TDCo9xxk/o38cZp99nkaP4CY01zz7ZoUCQOKU
NVnNJOfIImf7B43fK+IW5Wm5i3RKnQNvJN38jqBi47m0lPFaQf+kPJOutJyHifeM
5h/dXq6HcxWS8l1xiWV5bsdVp70bYqH5C+Rvf3zxSUl5H/+FhJM8zgMHEupI20R2
2SwjAhheyoI3ivTUwDghROTF0wPCieaByQu0UIsTBRwhXVWVbJxMKxHs+PqasH9M
j24T7g9828l2N/q75iUdzlsIsCvhJNTYwjlzeDEKqjcQP01DtA+WpIFCJHMxGQhk
VB0YRmOZYCOkmrndVZe03O0SHcUxUCb8XS02vkU7SwIx1hjk7Dnfa8CZ1czz8KDF
sWsQXaMbALjTJLXdSi5br62S6MjsOw6yn+/x7PSvIYoRfps+HvJP48sxaibTMJrG
Rk0SyWf9ylcBUUSSUoQehOVbU3QFADS1O62PSQEFoV7NdUkRSDKn8CBH17Fx9ydc
hK/vWx1d12o0tHl4lRfyn0VhSPtPu0dZXUCgS8nH7nacon/TUo86mPRjeQfNdz04
cl+FTwxsvbtrof0PkMYLpOnfnBJSzceygBkLJ03Otni9gfc8nKxqKleePrqNs7fK
MB+dRGaSu/m93JiRns+Oc8256X9dO6YV2gRH6MAdsqC64Jd1YFY21ozQwn+6zL93
CF/BOtft4LQ6Vfnsjwr356KAMJhFjI+Bly2Yx2OGWONSFiiNlKTRV9HLvScR2RLQ
DXR8tuYm5BAFUVYzyTHEjv0GNUXmy7iFafMXrCCpoV1i5ZXMlCh65QoCl0CJRW48
uDoXrBlXkae1A/Mvbe1aWjLt5cxeJ13dx8o0VgnwuzQ0cQjVObXto6XFU3EHZx3a
wKixEVFux5DCUjUxLRBhHd35CIRcElgWYAE+0XwGYd6Sg/b3Mq5JWt79u+ofsXV0
SjkjBzwXdzlyfpWoSg9WV2jqqUxTkVf4mjYyNh2FW5N1ADSGlORhhyPHvVS7n81r
gDWC3WLvsuDlz4PXemVGBUtCvjDHJgwoMh/l+OaYYERArWDEDmDPFXQxGADUfTZe
ipPTt2dFk8fetjEBCUypGVVOa9HDodOd+eYEBpC4JR7A0cA+2ZjjOx+hERh6Nlhb
lcxThZPLyOqExlwLdHU4179V3yNlfrnd4tetTSooCUEQEmjTv5zGb6ucXmC9c2L2
0yYN4rYKHmXELs17+ecinOYtnaIrUKr0Uqq8UTGJik1gkY9H3mFCd+lwyiEf6pwo
mDYZ5NgbzDnnX6VEf9quSM4VxHPvsAMF55HcAnJxY82a2sFrF91E87ln7H8+OE54
Iiax+BhJPXGH7Ggz88aOGOvCuh6/V9zsalnxaxL3ForDnfHhaMcXE6/EPRzZhPLb
q0dnSfG1Isiit4VWrXSEWTHHV26ZmkdT06tdF0lkryFmYFKYh5zf0N7YXpgyh0jE
ng+BK2XMzfz2Hsrwhn5GtXPtNV4CSqufhqQV2g+mjXJg9hlRwjczpfY8mq6OvDgN
TyWQE8qatdjmdiiy5b4v6QaDqsa7gwr8laC5cuMcs7kebdtuhtfzer3f1vyzaSw7
acGgJQF7f4Er09AABCi32Z759EqZg+fB2k58ZHZNJubfX3cWOs0a5IeQEsjjr3Pl
kwOFokYm57NuMD+Sgkiw4MqQOYQzAT7qXpPpW2Rbf8EIeiRnxKMfcR5MlVQu9XkZ
M+2vGSRQ09lSysEr9AGH76c5oE3R4MgpB0R7xdrtXQW0OSSGCbOEZtxSCP7TdswY
dgC5HbOyiVrmSvkzWAIviyebOx4rEACLhENAEl9/rY9L6DxyunnFCtwhVL2o8g+d
bW1yylrU9liLRlJdIxoWHwxIqYvabn0NYDtE64mJySo9hAs/FaI48Zzt2RilITZb
tUpE+HtJ+n3mQzO7wTrVckDVjmiDJj5OFRr+kWuA0QKZ6CQNhl2bRnbarsXMOEQO
rKq/z3SiNp/L/Mkri9gF155H+R51rJjZ6N9t5WbCpH8kyeIMeBQ7jE2TmD30lCkx
h8u+fOzvTHbQ0icb7Sl9nhW6UrEhLSbiRYpl3efKnH9vo93yI1vcSY0BLoMa/AEE
5ADplVDkOD6E2U98LtfJBFZ0pUg869ayldT8XR5cVULJj9txkeMKN6+arGu7y5OB
Ta44P4Gvh90j4r1gfDeZFAJsT1aoqE7aI9LjUtIXSs9mbOGun5vLENnR1Z7CSz8d
ARUDLLIpxVD1VyUV1uKgYIPxeIC4Gl/kuQbs5XkO39rBz1DrHQEKvsHgFTv9AVdz
MTJLye++u0Z18pSQUiNYupbbq823xCwxlGuPZ3/NKcpJQDXiys8ituDmUuRxnMMm
Y6KGd4w7GrDdNt8ghk5wUnIXUwJRw9yjYSiNJTAIgLihJFl74Ww6wY1je1OiWW+W
IRKtkFYIjhcRQNujTkkgVdLJyg3jmh5dUK9SclYwMNsM7ReZW6reS3ayPcVoVVmH
`pragma protect end_protected
