// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:22:14 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
luxXqZ9SfT2P5COsKeWszefcp3LGYiMRvpdK159kG/0onHpCFeLcmsEAnenXAxHh
+xECXis9qgcciJVt7BEz0xWbrPYO9gyiy0pytXC2PfrSg4U/V885L32aH6UcBBUT
BhRudqem03LgdmhvJEs5gAbZbTeCDn9/xiziUl3U7Ss=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8416)
dqVtjBoife6tX75y4QY//x2nf8lSAKMoi2OQFc0OAENqbUZwj7sssKaVzSyElPMh
S9KLVkx+CIkNK//vpH2VAR+7FdxN/TccVs4PVhTKP3Ptr4BRwyII6XYnb6e8tGXG
geANqsKsecFGkruc+dNBwE6Ma/2Re/z86bUzHW4ZZf8CXnxnQ9qz0VmqJA0A+odm
+RdUpd7A4tQ+RhJ8Y0IcvGvU3FzLobScHFioxg6yUi+UvDsYbanu3bxsnPHA1+O5
vCSNW/A+NEM8W7E5mBupQramdWiC5mDqxSVepu2w04mWTzV/5bnbu8ETT+6btdkt
OWwEdNXEngcnSrqQoAFhXVqzodglGjwWJ3hfJa371YeErXvgvW+MGFuzOKshdxzu
CGoGzrFl1lerOliPWbnik8d9MjQYth1qi15ww0qfCAWB3KekzWr9kGAScaz2d7yL
T36TXyrSo4h+HogIrMuD3BMpDcQpMO2W8EMHW+VUnawhYS+NkOhOk6WPFLc1LeO3
YVOmf6AtgP5qfLEdW+Cnjp9LwE7xBCDFnSyej2T9aTJKXhnYjWrmRGwz+CoO+cvO
GqbyjPEZK2MzNwoBZA3wdRDHFwpHZLVF851TPEc7m63+njNNpqXDlkS5qTFSjJY4
y2zPSaOFKaIQyUDJ6e+SbkPVMlRI6CJOlQ8/jzVnlNufJGJcb/EMxs90eMFcWoNV
RbPkxXA5kjrt35Nf8isQusYqA4DVYrZoFSv0soAhovQmuAOQXxI9LtADeJRgeZ8k
gn7QMfMpqWf0HQMJeNX0wfkpTc0Q2kQPlSNTZC/9IJvotYni3FOK9tJRrzs9lmXq
3kFi+97R1cwzZYCmyDMg3aZ+zhqDuXL5b/WIMYNO8XtW9ew03ZykTtYIvqHu70MV
jClA3ONsftqZCrX7tkvFXP73kyfrYIDUTiv3uKYyv135twn48pRh7Y/48xCZi+ZJ
4wDtrPBbRbQMZDrofjIftq4nniLTNtko14kWKRyFmemWhTJEvzevLoD4nh68A32Z
Cm5JbQMIEkc8I/n8i1AQbw4rEE01OsRb4KiFVxHOJRFdMoLozxYN4Dh0Bf0QUqL3
bExeSDAvVg3IZU199XC+oQiTxUdky1ti8uBo18pdby7DehHYjoW/3jdL6eyWAb+q
cDhMrt3i54du2M+TSwBD0YBjiZzkAJSNH5c6RM2ukvI4vC62mAYQwnv2dOyD3U/U
HZ+ABU9r1zWW0bgdhL/02pcfHalbyLHn7M3JAMCMlqf7K8hOaMzGEbVPYlrBs30k
nMJVUoDrecDCxCD1w6v1ZN9r3fBMcTSzL8uOteVLWvz7TBPkEU/YaNIUmP1WqjZ/
yOmZrI4A5pSJFF3WE8y2AKf20D5TPslKYgoISTvjQ+xOaDTVNu9F7dT5bv+GCKsh
14JVjUNEsds57i9fEfwD30HYVE1jCRjNO0JTHlqScImScMqWZVyxvEVw8z3RiBxS
YZEwgvuiwSDn12dHmdWfVUrLpma9qvnyoQndMU2uT/LesEyRBw41+ssNbyPd2AMx
YmgcnfO9gwnpzO09gqaabu3kTME2dmIY7/VdRVBzowBPxlxx9se4YWdxCtpW20yB
17ucYOY/gijXAvotkp9oIwvADTLNVOtl4EKEtOJJw06sTjYhyOZLcfWoBryK/kce
aniiEwC4/a4F0YzTJ3E/ZlizmkxiIgDqC5ASWTtamaOrgLKnilQkXO/qS4yUsb/E
m8rbkXC6ozSxau6H5MBObWI91n/MelHO3O2pQlPOHREixl84ssyg29GLdpZnKmmk
QAFw4HYJo632NI5yw5ulWZyedQSEXdEPWp99MHEybjnTAghBT17ZBTA3WtoC2eyr
gTuwF6QqvYHcVK1s12jALTUOxXiZ1+YWKeI2/8uYftkUKikjo9fDw3hFIsOOP/Jg
1qwsK/uGBygXut57DuC2TNkmMSqXZ2+U+5CyEIjYYGHDCVXi+l22oJ+xfDwOpQtJ
V3865SyZTr9ebjpZIk//lfcmjZbe03WU0ibjitFX1OI7e6DLmgvD+xNZ9OChxzGO
qgM7XuWhwCyP56deX+ThUo31OIzLKLVpwQCsvM1XlvKwIyPh09YdYY04ymAC5VEF
FTO1g9d/nh8dE8cw407sCWOyNGSPRZregl50dcLAX9tVbbLZOGKiV+t8+XT3hLxK
Qv2aTHM3qjAKsSpXM399Sz161HgizpxAutndgRc5qNVCjgLpjgPAxGgFBNgjfFhY
ZKdxpEsL+AgyqqXVtuD7wN+iCzAicg8CIMqN/etJmwT4y9IW8PT0Qiaos6FOS3nR
DKWMBgxWOllNwLmPoQHmz/dEFdli4B7hdpBaJnjg6zY0xEhGtlMpFQU/EwYIPMxV
JfR+LxfjJDNeXkzTZ0jb2LST4oQe451+FvNcsmr6l4VCLM47o5vJ2OI/dnj2K1K9
IC268UG/OQTGFYqyOPK+nLM6OBbMdLWHhmvCbL5Z60N8aBJarKKhWAL4GqmDmbBj
nO63PARgZrPWrnlICIg7eaKtm4NkwFADM2XZPbr6MmQEL8r/xdB7bq7Irh+ALJ//
LRvobEoRki2W2mQFBBvaShYAqG2oHZGyyhIMZl2wd/cVrcpJLO03w3POkwzPhilr
zlL834VefU4VeiqyGbNE8U6nntXD2P6Zr2LmUhQ+SG6feNr97x+XKXIN3fUY1PpT
XBR8eIIVLeHMlPADnHc4nPm5iqFB5N7zOUFxA1eY3qWxzERMPbQWg6FlA4hKIJFG
YuwKDehqrs+YpmHKjXiDbsJFfJ0NZJOpBJ3MtAZe/w2efVZ5OsBJGsP8KJ/Cg3Ca
YUy/1PsAjesWNFsNItmrGUJamk9BTgORgZ4uFVkoamAXAUe/yTzb1Y1HbJ2IOghC
IxiWpmcDiB4n69YqjQUDOrOVJDMXSgLrMdlEmRlb7B1w5Q/fb9kygdzcwAD4Sz/B
6qfYt25ou/zAJNaAsCSk1y+45UZeSJXx2Oncl2RGkFWFqQOZDL1s5OZwyFiVduKm
e77TVvdKCPOaHR+p8l6HRae3IWKjXRRj32wpRvl84vsyxTHyC+UnTOdTt/l6E4Dj
PyP+eSoqfRIXr4NDQP4ofB5WbM9TnKy+5fVfGvTFgIHb+kRTXctrE1la89QEAVh0
5oXSdKSiP9Emogm9BXqyqvwI1aZaV9TUO1m+X60kc5tsAxvUebGr3oNbJY5+ZkeS
IKN6uBL7fgO0wLzOjA7KEEtZpmX66+yuUzF5z9kuO7zXtw82icMZP/iD8tzLjHdX
3R4lhtAOrUOT22KYjws/faHtY+v082p2VobUYjJ/RxJiqDL/N8ApGboemp8QmHd+
V4ef4Iv7yvNE/40f5YAaGPrUk6sMjDwBWvxJqzV5P0Np5bsNAVFc51bdc6S5Syhe
vy6cEh1tQund6IY8L7pBgIw5bvvw3HUahArsyxOoFm9NTnbOmeM1b4eovDm11vhW
u1UYEzjFAxFLhezxmqDf7ctMG9xw8uf9VB84tDuPXw96Y6W7e+kV3A19ADG2O9yd
fphgmWPiwPCDH5N83Fu54do+8zyp5ZDMmiFyf8c/4DULbiDMGKWC7Rgxpn2ibvcx
eQ/WqR4aGl+sksXPY+sKu9gGfzvmiexium6p0a49AZkEkuv6Ls+Iicx4Yp/QHRko
FJ6yRn5Cl2lPK02zwJ0ZA9bho3UPb/UcXnuzotqIfQYRWLJrKstc1NTz7pPgbnsM
fPeP7tuCPs21sbjYHnmYeq6QGPRLYXVBqHDo5nJabGLGDbdBOdgVJzRPS/C5fZLV
E1B9qy7iYC9Dec0oKT87yTIe6a+gONF9rIiFf9cMSyHTcW3q7PLZkk8cYvzd2Uvg
eLV369zilqpbDrG7nguBvTISsuv/aCxpMl4L4NUq6OkMt/i/mpd31ec6JFP5qJrR
S+CaA1bQM3byzYdB/ZFKKiHlLr+yKPCWDRWjj/lejcNApS5UOr/hsUfS12FQeF3V
dtinJgxOyHY2+Cu+kHW1NBD8Nxp18170CCQRDVOn3YSnCSBDz9p161fXEMrWomzj
8VroeBmL9dLSOyMC0ujuLOTb41zY3WuDCg4OLR+6OVemrBPC+NZCkIigXUHRPIOW
KKxsjP89+Q4eEVyGEl6ZmxWRId1jdqbOdkLXKvCGfeK5TQZbaxkDE/r/MPaPIapo
KrFj6aCFs5fd0I5KQDsPxvaLcga72ElkdmrLJoTk+ApWACwIxKbXPdoBStmHzxnG
wKLNNZmgskvbVkcUFZoaEc9ss+Ry0udDQmbRDejU4NAmDHImWTFcyb7YjS14L7JP
yxOwJBk5DVXJhLaxo0vwTW+e4XIcWiKhGe4HC2syA9HBfmusssUxs0v2cIPLDt+M
EHqGm5xWneuoI6RmI+gj/eUFx/ulkJJInpkxJ3NrR5KsEb9gzkGI6s/h7t7hvYPb
4+rtlw2wLlmDUhAxNJuwaOH6jhzDnyvwoA+MP+ao7vsIwbuau/2rNyr8mJ4nv4no
R/i6Qw/mYJlwwyy0kJXAUpxFUNA6nsAhWIDz698FOaTcnIZ8/yiMhyV9hZIkEgNr
ec2dFRfBKkRm6L2EwANtho7fiHjFAhEttCTiw7tbbSTXpcktnvYmRicagSol0tBe
cQ9mClWjBZUJciIS5J6P5pUtrYm46REah1mKrT3g9Dj6JfGKWRNNjG5PegG9Mjl2
Paxkwsok1x3pRxmycwQecD5mSRFkfqQ/jxVFm7fAvjK+k48IN0nFHMVJav3928RO
+O6WwWkUAq6SHcJBDV8UDI+XgnAzS3tQ54WDGfxO6SOEnqPsD6PCsSQEvV6dlOl+
kz2MQPbS80T78O2Q6d/77Rk37KbG5m9hhZoJlZsUwpKCD8Q29reye804vr7WRRI2
7WBPVwuwEkRir98UA1UpMeEL6GcQdOccbMnwiuMOC5BrcVS/ek82jiwkffCxnPrc
DBg0TX56rIhvQtjN7TA2r6x5opj6vJc7VGVJReI39kIm3PWhxn81gE7yTSz2tBsu
ww/fnxBhV20C0eVjSEpxyHS/UHtDmI0DxraJrvwfGeLhn0xTHRv8+3YA1oguEG9n
4WnEmyzOo3/2ildnklSgwkGZIt04/vKqYAAkLJUUEWpGJfaKXKjW2enstM5+loe/
etnUuCYF1NWJVTnTQAa5JbCJpeGCyyOhSSMocljNqBcaNqV2yd8ePtDOMa2Gk/Gk
JS21Q3KN8NZfmkg32BncFGSmCwCef6a2MqREFW1PcigUzamD7JVZF/50u2ajD/Qd
IfdWIkKxXFnGaJ0H1zlkT5uUhJG0HULDp+hUcTY1FubqnMw9t80q5UKBK4VjMsIw
QYkSD4IjMyJwiNTw2/Sq5PDvdv3UpUE0IINkmuzeEbLLDkt1pSp4omoYWkWjjLLA
daO5Pc5RloWhO26h8aK6v3fVwz86tuOjHEGX5U35TS2pzTg0for8RXj6AIvPgI1N
WmhyWFUus6xeG7PaWIIqToyOy27a+f99K9Gkgjlyb9DASMQB2UjQvOWosCv7Tfy3
e70TcM+fcTtvuEbx03jmp9sXUKhWOcBbt8kUhU1ZBEG+tEBKRZpMRi2n65sUeHec
NREeT1gdJ7jJsJC5j4icDo4/b0RxhpqiqaQUyB8c7SDAxzMVbis5h5cIIwANYnTA
1exTA4SmKwAJPvL59g00HT3DQ4eQX/Yn1Y76pZ4/kID16Pd/VA2DMzXMFykVxnec
BrESniMZY8k7ecZPNNCPmAFjRC1ow8zyqV0eCKl3Ww2Od6BaAOSY1KPEBLEpgkFu
RMfU5lkd2PFjsEBhrLapylHIon/JMP6z3LfcgDWXws9XHi793/uD6PfxAFCzy7DA
ggWi27NY3YyidYtm6KkdXnnYGgBeAv9+OBUygTCMgh3mhdStsldYh0/aiiifNe28
A3QOYYCxzshA2HeG8IL64vjSNSY645RRVMRwMfg7RwUMz0QDX7GeUdG7Ury4pt0i
CxLeWn5oWzPDLbhcfAOVOGoo6eM+jYhSUjvZPsSoVcTZdW8lwuFQLQXdVe3KQ3fA
kfnrqCsG4Xdi8wSfKBOEr25clYCjNfw7nR/Ww+dJhipsy1hfTuu9XRLT8dhxjY3p
44XGkuZYnmeSCvaUKJERHHtCtlcq1kgtssppATikaSsCWZhECY95T33n1FpDvuU5
w7VVlEio6EVemxiIHTP/y1X37UjA9jlosOD9HdmIaFmNfco2zrm5C/u05ozatlzk
BBt5AxmXoVO8GsFafunuB+/7Reeb+t84Q9O+QgUq94an7X2fK941mditCb0cPajP
xsYPDQx6ecprN1gkvqibE1WwSZkenQB9zQNwP0MxZtfqwW9WadmnEbi09hQDcQ+E
dn9Qw31rxX69TJEVShJM8zwCzIpUnARvOfK94B01cGMQgYPSVyaQFXQEjvJOki5Y
eGh1qsl3hqu7EoRRndcHV0CUI1UGlQoQH9yskS59wrUGATaSOEZSqoudxZ4g40r1
Rc/rIpBzctBNHVETEMYiecgdCsJ2N3bzqJm9uDxLX1CSthL73nAqiSQ2fwzgMOaU
OfzpB5FQMXnULlXSDTD1APS19YkwO4V+VzPvkBDqdob/bQkb0iGgMTlHfMnv+GYy
cAmZLYT5OJdypYgJt5q/vpYY+P4bSbh1MmcZBDN/eS3VI6lpaNG9Bu9wf92p7ffM
rBT4jDlV1Iwvf0f+QOnrOx53ge/kbMV0vG7ndYB9Y+/QpVd+dRSRolzNUsUiADSe
XmWNCtkE2Luniay+ozONal4kx3WME2ZKkc/f52yN98CyiVdVDvQq9L8ZIGJH7aIA
93g4wH+n0v15FOqGjdqK3Ahvu2r4HXbrKSKm4w9v89lSHhEh01z+JDano2xSpuvs
aeBJZGJP9ID9Ov7169N7eqMIYoAd0fhxGt12+WvJyFyxID1wvdyBccsPMKrLp7jc
PhkK5RpQWydWDcFWhU16NfklKotGLdCt5swy1+lEKLu7j4c6CqODvqwgONwNMypG
AUKZsE3iM7Kx9tS0lFTvyBroqyKQO7QwVL1oq5yi2riBcSvjWiWUmNeo2q6akKvP
bbK8+uvfrRE1mpWGhy+q4+AUKMO8iL3BdnqHYEW/7i2fkCyliH1wlyzGYAoP1Uvg
F9QQ8Z6EWRoYsn0F86gYLTphG41ft/7zNDRGauACFaL/ojYHa2PY1Wby83yRO5f8
L0fswH8FTmAmspzIc1M8IzNy+8BhsyxqJDNmzUe5acVpnnhanRxQxOHm9Q6jICy5
ZTM2axqpJNQLvXdZ8a7ZlIwt4UrnDKR/xRCYLIormOkrBzeLEI/qoMYfMduVi/eu
D3RPPWnik2ZJvmtb5wKV0R5lHb+CwQ5rWKoYz8dfIb8V26ZvND1MAte2FtE4RZOR
8pzgfH1J1GjXWZoZQhoV7suMbUXVVx4apA4FRaa3L5ntsEUatrB6YVGW/tx25Sqp
PFJZ8SyvTwvokp6IdTk0oWdTGD+D0EjUs7tfJDlAUTTaYJLRh+usq4vgo4sUphB2
Phr2MVaqjOLaicrwS4uhPXv5MLxmjrD209OIe8oqZSye5klcCrfEdz+YgDwvhXUC
LVlabeQvGYNUReWwt5i4S+X9YN5DbRWlrONAOAZHbxVJiIFosL06cMfAhj1zRSvE
NjPlmngPq0DwQC3aypck1TcTGqgcFdFSbEi6DoP6+0nxydD1fE31afIAUWWpEMML
1PwQC9khUKIGVQFgEMBcp+w+VQnFXwNvgEoApqTnF1mqqlFERQ8P44LI4gLB2qQW
jrKNGNl7GNOZVy1Akw2hsjH1iyWvriRUyS3blx6UfmZ0vKs8mGLRStyiwAtuiM8I
3f2rfz1pnT7mnUZfHwWDzLoW0ATsmCyQRhDNyqAkt1oVlrKrmGsaeCmSUDSynSjR
L3B3YAL21LNeTy7IMJBBMmQ6UI8akbSlvraLblN/LRKJI9J4G8RFe5YZIdQjYYdx
v3XJgGOMPi2zAvxGlolzgz00acsSfkqLJm/Dsdx61VenNO3Q1d3W0IE0th2W+NtF
5apxBPFWW1w2qme4kcYuSFMkmhcwjcoiuGEu7xiW9U2RAFIaRyrj2jXBsWpetmH+
hMTbDAOzlFiLyFut6dn5UeN0V66MLY0xcTPrS4ywge6H5ru7Kj/aucPIhupE1IFI
NB44CdKy1wynYLeE5PpDwRMzsv4AhEOdesVF6UXy9Lv2wWTxQYZvCkk9clilOjGZ
9lZzFkJmmS7k9DHyzO3u6UtjCLAe6E3uh4TqgTFUaPOEGWnOV5PUjhUg59dqg7WG
1G06FqQh4cnwpvtNZYn34bju5FXDq8OL64uH7pu0SW9LzYMX6+fPjNw4zsybA8+Z
bmlW2cvPHZTgsu4hgMKlSKrFDY+oqrzMNO9/ibRvZ5W6E+r123GjHn1gnwlGMcv3
C4P5rNa52oUWnLO1vMiP8MEylApjcra7Kj1CqSfG7yNOe6Kqe1k/7+NAWw2tVq+f
8Z7lvnJ3Gd9bq4J+PlV+gIjecvopP8m6iB5Et6Si6FV0K8GzQmWvFe0mupfJqVsQ
OHMorTZwZJAxZb2cJm68JgfZWFmL8ntxqP6hpsKg5Z60+67hyuBOz5p6ZH7uOz8R
BTjDe9juSVJcoN44tAoFvNFN/IVZKW0PmGTVGL7G0JIiaHOH0JDde651Rk+1fiVw
XG+1f754fqXL3RTfjTkCFg+aKf7gDHH+Mgga31Wuz6OCOl3jRadZJrxF+Su7DNoR
8BXjgHRlezoyk5oliVNC1WVdlUUBWj1LhtOc6VWrgviFBo1l9kUGcZTAEvtbTjyl
7jKTtfoz8HD+t5S14AChEvBGOfJhiwgdGv83a/fBPbL4dGYEEWM0P/I07u87Ninb
lvJ5BevpnPpSomYLVrMfAPpLDTBYTDIUGiBq5EH+qONMl5gelDzC6+kZMW2/ngNB
AlL3Y529cog4476n5bE3UOEBchmMuVVA7W7+xrjcSH5GQjlo3aqjucMpzcCBlnYc
979lbW+1Vn9EJ4SpOIIrZDOcEOAYjet2KOKCOJBck9OxDppV/ddOzo10r7wHYYYw
JZBe8TVMpj9Lrs1tG2oe19/chuluKi2fIPYNDD2bIjFnVLcVMhnOgLPgE7GmtSUx
ag3S87HH4ul2BhG6ALx/iP1hXj4nbrdGdtcr3bV+0zDyn1OLzLkIjiGb6J87JBSD
XCO53VVwXCkeBSoJFjdRjb9mpbtOs6NG9OLg0/2D9VS2oEnpUpFJ6LmBMVcbvFHc
l9otJhGBaSxUlzqMtD2kt57bhCmZWNgnMViUP/nVAJXBsMDl3gyb42VJej06lWxG
LUINotKRm3mvtl77g2Zgr3kn/ICCtze7XfSa4Y9LXKAUwKtEpTa0r9/TxoC8A3PU
9njkXSt4wroanxXcdjkWMu1Fhgiqziz1NGw3k4q6hAKHeE1dEvkSvYX1AuXyrt6d
AjXXFavx9Wt9/4NfnlyA3uDjfD2kT8Bs9/0B5U5AF6K9wz62fqhwz1OuPVHzvuVh
XSBlWABiOgcOTX+YrnNRCiTnB/k8g2Toi1Z7vpQc931w0bWRgaYg9z28QSI670BA
Pb6qN92iFZy1TAKmE9Rs6nmO9jaTpuENHJJifvdcZ8946jmJPEwQfx4KhYq8g25F
vqAL0WzcqJ/kFpo+Tdz0uj8Lx1VA9u6ZPDBJtCwRL+6ip/Ud6iBmgP4fc1VsWr7w
NL7+yfVBA+ttDnKaM9Goz/uYF39/iphllO3eYqvJ568zoM/UTf3eag2QrdtjIc2P
xVcLaotF5LfHumuqOwIzLQ/rRvAWsLvrSWbKGAMlAIxip+HdHaKGoNmHbqlZY0R5
R6i77SRyr7edZqGWM96xH8WzJELwVT1fsuYZRwAquJV4oDN6m/2bvCB1Uk40iTWn
ddL5qZg+ROLnILC6NqEFGlWshEbH0hPdRUelXvfuhj3qikOV7kwjPSF65KygDI3J
xB5VQUUY0tZHIIFkN3dh12MK9lHoViDao88pck6SCq6CEo4PTh16g/og+xdr09q+
dE6jjVTlOCDRDUKYAFZ8fx3KfOWAHx7lKQihmLcUgKcK0ADmLpmP6kS3GS5q8YNU
lv2YT29QrNVR8AAsXIoi9ZM/6PX7fnnABKm6/0Adp0zOkBY3Nu+QGRMyt9EgW+Vx
tK8kD7xAVweVuwKrM5CDPr+oy0kAtgyziMI+/WTyZSLzqUwcvS/3LbBtQ2sfsHrG
1lkiay/1EYTSOy23rURyW8iZuPkLDIavqrMyzsA+G6LXi9snfUYn6gk9ZukrQ4wH
GX3neIPtmpLKbmChExhM7Gzm4gqnwkJy8AvmiwUiWAgNyfeEJAXA1JkvEm5cvG0W
5bHhqOnx5OsrkcwrMGKAUQaeaH3fFVr2gZe+WRQ127rs82CAnoGK5x0eDo5LIh0y
mUTYfCisWanqee8D8G35/frpfj3i6TCDkT4jwB3HtmUpyj/Qs68qiQRtJqGGSXDo
RlSuN30l4Z5tW5eFDClCKyt0knzvsfEI0pKMdvJVdJp3pSW8y1FYIpeKIKy6LX8j
VrHVBgdqVMONZCnhf32IIR0TJhPE2u+K1769xlAB2dUe346t+glcOaC6T/0QIEyl
+TJKaJlVK+D1Hiht1J4rpBve4nF7WtO3vZqWOCN9gDU+P6/U0bo9PjiVVUI4YecE
FFvG13N3uRlhfz955mMeUBp0UaR1bOW1XdLrY4sDqcGn8pVHXtSFT0GxbLWhBLLH
rKeTdbbHS17ctOIinu2PCK9xRGxpsGEbPDBbFfKsn1rwS2zMAAQ3jybeX9h2NcQ5
AKx9Xy247O+MYUq2uDczMY5zLokHFUigQn5K6xGJom9KyTwFyNYmA37fCT+/DgJA
Ae+4vHX3mq00IQrKOD50as6hUIz/lM5s6yhM8XIxDEFEqzXFeadfvJP/27Y1PUii
PjIxRAMJqul64IxvlpBCkcyn8HMpVUH2kGxYJorZgtPo5akcDAiFwHMD4PPpmKjN
LM8cdcYa/+7cj+SJDg6cV1OR3T8pXKKEYa8G9AnEvfZoI2fXpxM4QASe1azmc6KA
eiSiRrSBpgQMwji0ZJrMnZI8QNXRUFP6p3wAilAL3q3dExS7c4Coy3EbY97sxZ3F
XwfqQZqIC6aK/+AklCuaYhC++BfbMMOCC84zAnAGbXsqBJHQCxxzsXbQYDt0dMMQ
oeuhyppXdYbuJaLiYEhOC9Wl/G9vhH5qOfmuytP65S3lk2Od/hV1hNT/Ny+M7jdZ
KaI7gs6pI2W4/8fkbtYW7w==
`pragma protect end_protected
