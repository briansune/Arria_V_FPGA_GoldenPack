// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:53 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lFuUsviMkERUvxt5PV+G2TDLCc6V7kOf9cWBZRxL1AodCg30yohuTVvNsQDdWa3T
FK+sa9eU3wYYmOIPLQKZrf0gq5kEH4Rf7XW/JevN3LG6WuWKz9tkW8kjhCUE8xww
T9g/T3OMb6yZ3pGHemZ2v0aFig90pngPz0+jGnjmVUI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
SUrEEvK/4VTv6AQyu9eZOwS6ecLtSz9Bl8hVcf4LF3hzmQCOB74O7VltZ4EoJw2K
VFsxt4uWIgED2oSP0OiDcIYnC35jtmMj595NC3X2TYITTB6FBmMVBfpGJleGT6vg
f0hWJBKdu2Xi5qfmMzk2SB+BCvPEYBN8QaB022Ft3HYHXELsRj7ZE68Ij8Xqr2Hl
zDOkWBQmrXfiRlBGT2osisjusDsm1beo3iU+SHv2VyZ/9Gcqj8oMGKxi3EXI4Nyd
gY33oZxFfYDdJd9vpKYDJiLcWgFRw8hoOPa6LcJHE37NtB/QbEl0ZASa6RchP5WZ
zZu3yEHNXiwaGbSEy9hV9z33HB45f6ev4P94na9pgFLDUOquo0hUz1X24Ns7am3C
IeiaJBlWyFGNIDKYmFvXbbIWeEXMg1v9MdZi1FNmIycA5WiRdNaEH17UCv992bd5
0zx9EnOlWRjFTTcKyFaJXXvVN0Xir5IjPUHQmhBJqXR1zobTiHttAkar9m9k/qc1
hJqz3Cc4/quvhu4zY7fqASDOJ/fWMzHV8wndUSkWMqt80oLIJsfG7SnS0g9/Jewj
ZwRf0seUHD9nh5Wfjcs6WZFsvtFy8bi8tnvrsMMJp8kh/rDSeTewC/lrJTSRDFtM
Nyq5O5E+9dQqld8+8aJx+XEA3XXF9liXX+gzWZC5tMM54K+1UA1PS0ESe+nW6H0d
npcXuBnErVm0T3urb7unqkUsdK4t3EZ+H3FNCFGNTRLR1JZ6FIGgddutV5ezITdi
4RfFzJVKv+uc/padta6LEexFzFgKaa1BOuSA5VTk7f8kfs3zAmUueiLHGiyiazdP
NE0mYrl0nEUGLPfvyPL13KHOO5iDtirkoY13BpIARZclCS/mMNekvZgHoBtnYRxp
XD7BqWGg8MKPt+0WLcuMKsg3nyG8dSZK218ezQZ45CtQA66huDZLAayX3XubyyEa
gn/pTtmQYjBqaowFkBoQnMZNVFbEg4qzYTi6sQIRJj2WB9Ic5Hj1dHVT4uIj3oKC
ibgc2II7PXhThYal1wAmPixYvlYHM8n3nogwzihncVJC0Pj0b+S37Dv/ooYTqVgB
5a10N96CxinHKCBLMxS1UYvN6ZGLE3u97TmgWxxUCoYWkRD4yKHIthbbhmwojUdQ
Guzibk2xy00S5C/gcFXMgfF6sbRyQ2GluHLaPipJaHKUa50P87sMxTPq+KDnjMEh
97OvBIem/m/F++k2NZH9iYWIDkVy4pQ2//7FA4YyQFMSHbUgLGWCVKECjNdLrFbT
vLe4ht5b1+OXMBZI7FOtW/0nZ4fY4O3Xt/92r4t0M8CdjTbbakXJH9jvUjU9or5D
3T2JYiNh1LFeocP+tUxtQYL9mflxoqQiAqEgonknOlyLcmoAphgR8W5PDXhWv+Mg
UJtVBRKLX+rZ6ohBtjruceO8rohAccZA4erh6Tmvj7opzg4fsZRZfLPdTAEk6c64
0BbfXdB+jD4EqcMl+oRYsFkHymAfUWv99Bs6hZYpp1Cc5D0GniCv0W86xmOQbQS9
AjoH9CJpY2yrL0D+Xr+lT/9BNizL1gDrwlb/K9DLCK33H4seHvZQPvYOJuJqAaC9
D4ziQmlXgdHOSnzIK4EzXEyivkXGTGCcljejgkoiCqJtqwBO4D0Mzve/fdsklXSn
SShepi7EFmSrSFaVV7tzlN60cp4uLBOVPPEFtiWJvnvhRc7xjqnCN+VFwUW/qY0B
pVOsMNufO9+4gmbRdntsuaNjJxwFoS1bKl8Saza0yHobKCknVgNdglEjdYDju3Oh
kkABZdogIyJnOk+u+2jtBOnGH7JNJMgdVeKlXFrQbvMbyVj+J9JmGvFMts7NLyVc
cNESDIru0Bt8GQuWNF+6qgf9DAWqi5PAjj39UhfoImxFkhfQ8/DfLFola2adZR96
d0fPeOdQm6vSDfrocTy1dcmrecGykX8eLxfeiBhnK8Xqw8xJ93Dy/ZoVAem2aI3O
tgOkS5QcJhzGwdzTZ2RZEHMmFTW3U8VX0LZyMmBLFrTgeBKT/B2pU7tRU1wtzUMn
hpLaTL0DcQczJBdSn0GHrh7a6YMx4nIzzSieHQd7aBftVl8vaPAV7hYjjERAnpYw
2UxrVDmgAV5FtqVWL0rRybu2VSnuaEOxBi6EAUVxpVKJF5VOb8tnKjY+niQWzdY8
+eUNWqY0KPipRUMmWruQ2EoohADaZRAOZFVhTOydvyoiugPqmI+xeoCW3Q+GDLUQ
5S+ASnsDqqtUWVw9QgKE5y0KR0NAA5hNSbh9Gj8CcAEaXBaEThEO3t4nuaAkvslW
JQ1RZuaSXz/1KD05lj+Nt3DzsK+TCDt5w6lxoVwuL7cdieMsQrlUKjhH1ZK9gvCy
IrakomOul99IciSbvHoc9kj3lWTw9rvAdvKFhQnQzIySX0/uqultqElgPLzVlfWK
AUQrparsLm7NZ3CDJ2SmQPHqVMJkzyH3+A3ewPNUuD8/B+HJQiVohvkiWVx2nD1V
J+cBxgZsMbgcIW5ih98h8Dj0t/kZQ3JGuOAJT45LCMRrTMHd4sPFe3jtWE5FbfHU
pEesxkcB+hJKZqYPIQ2Eo2Oeb9s8WXnrGHIDtK7w4pO11y3tv81zLMZnUzsUdmBJ
2b/f7QJrb1l15zAQfdFnWhm+IVveyIJEba6H5dyJhUcqJeVwqO70NRNAOCT8QnGR
qCzb8DNUrbubijxbPKAS2l+pcWEaWpu47Oo1E7h4Homth/ytR4D3B7I7Ek+VINXo
nG0PA2Jzy/y8orHh33f3VtvkaN+mVTHOCG/dmMLjUHvJQ7m2AMMUyzvirAflkG33
J8zYvp0gl5trG0b8DdyQZGvxml9wkAJKWXAtGV8JgCMjA0e8jZBlmDotjFe1KJtL
wZ3xKvFnzJfNRtT9Y/WE52Umgo0o8/tMMsNwudxkmausFjf+OROreIDMOCWAOGWJ
hChdwmKbXHrMrFJ1d6wjni+hexusRHLd6t9oqJdW+tMY9iOPUJaHEnwvnvmi94yo
E7Np9hrBfALmgAsrpcSaFFLVx5eNaSHudZ7z15hl3w2ktRqXM3eE4/xYKenWyZrJ
xvBbRcZGgDnd3YTulVTFjgK1fDodWGBk6uLKepmq23gqrk2ATHOoQL/sRAOmiATm
yCUnHMIn9kNJIXfo0ieJrvltYb+MHmXXBE5Ou0KBAfiefrl5HCq1853sn26ullhO
9XCY/u1r6sT+EJ0wRyKT2J9AgdeIQWW1KWcdm/Otqh1WFjpDxVrpcYqafCDVnhkE
UCR3p4iHGtzQCiX1EGNX8onawLjoH/h6fmBF9qaUhqQOpADUQv52P5QEKzUitK4z
/N9a9ekFCfRNtyhZhGk2zPRFWgKBAE/zv3mZ817bIVuPXTTTOarxOqPkqbm0b6/C
26XPeHxCGNMJQEGeN7gXyXOuOu9zsd5C6LxhimJU2oA3fadSgbS62YvQEXUHkTtd
nH35x64veMfSRv6/69wssDNN+Q1R8dEr5ZCmw21jYyloRNSAtHWvDQ+F/oBrfVtK
Vt51KMBgOC5jqrXEZ3QNZzBtX4oQm4T94C/eisgee7OEHQ9v0ttXYYi4haS1bMNR
ASx9/ZSG4xdHDbqug7fOROTqyiisdYDVNrv24COupXeIloq+talWa+K4rzlmGjlx
3fSx+AvZR9ENaXE6Y3A10obGvArHi544iymNJyVuV9H41CjPTFJJtZC3QeFTcemj
dQD3RvftJnR3nxIuoYGQ0DzhuPTQqkffP4FTBsnKIqwO4WSVSfHKBugAySmvfNxH
EYlegG8bbS+oPZ7vUU/eUfrndp2QCgpE57thkqPTprdiXJ1hSXloWM5zViwTv6ed
ivURMNS5fnYc5P4prhKvNBPYaiVdnRDnbJnctfOMNYv261tuSPjAosWo+Noxg3tz
J3FvNaWuCxiI/9Gxow/iTPqE/ZSD0K8nPPCaCxnV2MOvYBrhD0kla7lhFLhvIVqg
5d5p+PsDhmBxOp/FtgJgn5X6bbrLAxVwBAJWGAgSgEswWY4BgUWfeH5IhAwjLv3v
ghEO+ZY0OZ3M3e8YtxrX5g==
`pragma protect end_protected
