// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:28:07 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jOfoDQXRLnonOExzT9ic5MsFvOEd+tcayGp0mCp5m4K7QVws60/P/n/Qh1gXCDag
TuLOIFBHTwT0t3g1bvuNblTn4uv3Xb3fjSNpypCrjzSOH6OG5Gp7IWO1jyrxKWOC
3RRj462T8fS00ZuHvXEk+1Mi2ZtLjNtItWGQ3W2FsrY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5856)
SGSh+ZqqpJ/9mKeWmK1R1edufl5hV7uh2/G6ERhJedZEiiiYfU6tlJzSGtGsErjl
PnOcPvpjjud4czrJOYAEgMjqT3IoChbpXOCsaYxyaYE+wnAcRNCJ0s9fq/ScMQjw
q/63U5eph0JLawvHMoYaUmTnKF0zmqSbHAnraxVllfPX/DrxmY5AiBBV0624Fjnt
9Fm4Yg9i08B2Je97kR5Q7cDSgONupzI2J/ofqo5g0FaO0GuTwg8jBhrwAtZngUNB
2VfnKeIgjk298Ocj+kvgIvoXjG1+xBL/aFpiV8Bl41G3YkSmhrtBaPgtEZHoMLKN
Te6WcJkD28c4SSL4+inKSKr3VWowNCZgAAPLac70dB3sS2Iy1qQNzOYPlCm7g9JG
paMXiSKp2NoK+7BZzyuMjc8fNqMFsRlPoYRz60rSLzb2g9XZKBYafpwiydut9eEK
bWsZqOm9fvnaDn0lP1ayksGyKGLz5PrxfOCmhq2+f9BucYStbjHQwy24RaIIYN3w
MZ4W82W7gJyPK95pKtU2Z5/jqynkPajZTFmhEfbYbX61AvnjmvlktjC41eq4UmfV
wphy4nh7PE6+HqPzacp86krY0ucyFNHeZmkH5e8J452OiTAVwEhc6NxNzxoRBDCH
72oOXtIZxsSuMH6kC/f4Gm8LnhgCvK6BDUTLlB/76pumT2bhLDRnELAaC6VY3Ajw
Ls+icBx4TSQNTtoAExZQHdXjFuZcZBfiw66Uwe2kVYl4yJ5Xq/7AqxtoFUCnRXiV
ALoldjVaLs42XuCNq7Q9TLYeKVeHfjWPHV0d1OtysHQtZVSQlgNXiO+svzgaJSZs
gvGsdoe6atYulZ9Flsz/irRnOCXV7dagQrOlcs/0Ce72KZJJak+xxIZjhOaj2IDe
TYXBU61RNCti1HXDY1/Eg5z+G9z/zB2EkZ1H7uiA7BjLSs6OA+lItYIQoQsOXXEg
W4mExXowgwhhdOp0tz1RMM9JZh4w0eyjV9rSUYQyIrJb3m2xqnmAwt0n3CerJgC6
Lcu5wZ1uWPBbeZI76dRn1xwKDI/pdwmJ+bhzye3jL5fvfYdIdq0QK/t5O7dEPMno
wRIZUD/zXYqndzJ+4lahcTGzloTnveHMcQW0HKjwjiD1myVur9umY3xsf2zl+MW/
yX9DEaxOrjn3ltHMOGUby5iNeZeiRmZTi1caYh+XR8G7M8Y/cNAQjQjJd8ko+hRX
R/iRzSIAX39Cw/34lmIdKqIhObAHho49CuQFVXOOSmVno/bmOzXgISX6xV2+3bug
ar74rVtlU0w8u4A2uSgIM0wyzbBhWZAMxgdqL160ZEoqoVBIl81ha6yx42h9U0wy
mlWqRyFcnfmZg35OUImIeNRSo7U9/XS3yPTMWT1V85z2TfZvSqmF61iA9U6+dX6i
9lLsMHOknQNAhVVRMzvGqcBwE/Nl7j+AFg5bWq14/JexEmn0a6vGLF3iPLRENUzs
3sE6V1Dws6GFUpmhO7H2JA14uxHhrPIJcu6euK6jwliStScv/oAYDbHE5nWhpYuX
bfKuPkSIiFDzzp5ajVYLuOYmd9JoJSbqCuNQE1vZJLJnM498UxVpCNyZN2dvGIsA
+xijaOddIEcbVR4/CFNxfjAhKcZECKgF4Z98r/Gyz5aG2sunIsGYTHRndxicqxle
j1llc2KO4/+dvpR1Pg9XNw3UfqFAU3s+ShfdUeOn0xtsVpawQtHSnoYa8uPnJ4Hk
QHFelmbrQkxZActCFYXsGe5YT6FnfkQJw22Ai6u5OmpzXWNaMfDnsCGG79g0bv1E
iU4ZgYjDDyJAWNsMdYvzp1V3zd7GiGumqggoqryaZirkFreId/6+VJte0lEeqpBu
zKRzCKZInfVbQ1ALZOojyTdP22D27mtVrUJJ9nT+4/OfYOtM/2Z62CaS2aIfgl0n
UFT75EGTTmEqkYFaEh28t2qgZ1ISXadqMWqldUuRgbJFd+mNbuzWCYUGzApS+/9/
w4VN1HuVEkVRKvi7JwmCrhXdP2eORjGRIJsoMc6hojkw/IgtA1e4oTvSiNKHMwFq
3/eiZ+3x4g3Y8TjWhjk8t2QeZney7zcPONzFzDI+JgOgtTohf7QNYXQdmp5+mCFn
JJ/yZxEoY9yLw4Yu+n8brzoNOkvFEKkP2wR4cWnH4qVeJi9UXdPWqhbz0gbXgFMe
Rnb0npbTRX+2mZcxnRFT8D7HxpVBCVwQ2uSrX0xcxVewOV/V1+HkLECPnj7yxAaO
V2sKzRgHtHp6G8SFX8M1I9gdrWPslHcWzfIKpEwfUOLjTJkrr2YYyjURn78oEqr6
eAe3WjZz/YjabuJOpqInVGOkA/vzbTtqBYY38pB0zh/Tbf/bTr4M6cZ2z46ZbqOg
BXBlACFETLi7uZXOC/Rqh8hWsoK4jXy1HNlf3mn21FdL9V8TRGe/m3w8wG7wCnXs
Yk40H0eNoK9O0Jaa9UaC+Fy08mvw2hNUMhF32aaehGZdlEKr1VJwZB+hO4Y5Zyrn
mKlPBKPoOLIlP/ODVyFMx7S5Yee0Ryp7IKSJ9oBaeqZzZzTOub/gt5gORvM2J57Z
zRayKvbF/wNnzaDkuSeOyvOzqOjva9L4SurYg5Z1gbr9Bv31jRdfyEKTCKecxgTU
xtpDvNdHH7pBHcS8ThYAiPi/Gm5UwcVcykOcqZKn/GSn8+s/+OzZdEhseNGViB/H
daBVeQZrRJne/7sO31bWCOOlXT23PtC+WQ43c34g+lFgiMVnfUCKzzB6gyiCDIhY
WEovDO3akNmz6WX3UMNBbv1BYUcYK8A+TMHkzMb5H9ZO8V2d1Hhiao9ny7ytyWcU
BF4ni8DCuQYtPkyBG1p2iOtv6QUYMI3jKN44kGoJDfiDePlXNe8ReZWXjRLMAlg3
iI659S1OfWqlsWT1s7flOxt5QFl7MmEOFHKiFZx422lkQC6svOvrGtU87mwypT4t
WIsP1lohUEnjf9/5o0tpE8vY/mHGTx6YOjHCDH4D6cgBPL09OJwmkXqmdS/ykuCX
Fq0s2o2xGfyg1mrQKH+6txI3sZq+R3RKjzmCtX6ofBbW74tGYCG6T3DohH7sggq0
M2sscLXQ76G1mI9QZpSjZ0fvurCU/9o+G/5P200Ehq1U6g7Ny6TfXnk5WLhAe8PL
fnr0GB/YC841gE+6KvB/nV3QOhAAZI+r0qyr4EQDmXNdYWBLgGsKeBykkSAmX9CX
Ido8Yc47Nak3zyNfaIb4ADEIFWs4WVFZwkt+QtqJDXdh2ZY0o2zWQjLHs6L6OcqC
EvNQ+eXT7ZswgV+jFaGW3NwEHkrHGGbjjTkUVWXUZ8BY27w4KqIMRL3tem1cW4o6
1qzvhfbFiQz+6BvvxxYLR0BtZy62lOxd6fO/gxWM2cFZsKWIXtZ2o7lp/FSzwvYJ
nOnxUzFTlnKfw5kNOyhWlfg3sizEuwyGAVRSO0sQDB+pRJ0y5tNnWfkIacbZaYcM
HX2rk9OHTyhDLRn/GbUqAreBbE1/mFSrAofE6Ko6VrVTJkwcWtn5V0sEyq2UwDG/
F4ClRT6R+pr1Z600Zr4R6J6PxthHfU2o9VGZrr7lIzEbPIDs2yAw7t1SEuWWYsUl
3rrhZGHLtRxNSlYXS6922QiJETUxCrjIOdLo9w6rFM0jTLmhUlqxrNQIgb2nPYJY
M8uL0DmrQI8pg1cdEChf6Hv+cAXIx3KQSG2EXrGDl2g7nUt/gCrBTyfG3ok57LEM
o36KMoLnWMWI38e/xbpOjxHDu9jGLHH/joJgn+J2jf1i+jTBeEtrh710cSJGAVTI
ay9SaAgrbju07nT+Qmhl0XyJjrQ9f7ixpRivmISRQzQhmAc/PEdy7fBFoeQ5A4Hp
fCYyxoy2DGX1Bn9RUzGjdgLbaNls5DO85JWDDkRZKzGqQK49ih6miG/GcC+NvxOS
EJfukYDsrgAerN4pU4+Px6TZNQr+TZW5Ip3SmIwo4Qra1K2YXroVbYyPd9YnlA6x
M7SrAd8m9lDGOolHftrFrYM5HgsjAtxm4rZ9mBlFQL/tN3H0R8r6CEEDOD/JaxHj
2B8N9byWEAQu28SEFEdqyaeXY11A797doFCNhWjw16+iIragHr0ypX/q0dQcvyhS
ZnZP3a8jlUp2RHFnH+sXO0YbcAgF4IZ82q1zOwY9im5Rh8GZ1D7tOvxVfKC0Yuiu
BM89UwyGESZy2b18dk2Q+Yk+qLylNY2vFMIgw925ghy8ZoXCy5R9Gq2K9lUXvzVb
3K3mCVRxiZriCqNe+gAv1BlVwTVWya+HHv0FrZxeL9S9jli7nEwKbiYccKHQG+wZ
ck0A95Rj/qmK2sDXGMx5ckhY2L0DmigVHqX3JrmF4mBrptP63HByeWAnJ56pSNqW
UoAhRyNxvKm6LXN+m1WsnV2B5uigBYsnT6fTzG0iPfcqFblLrt7SwBPUz3nA5ylK
LmYNNKJKX4umarrP/uiVXYLZZy93F1xa5vC7lNh9C8A/TI0zELgtaPrxwdzb8Uhz
zWtgjtoDRwsd5nmu0GtOsotTiWtICxp5VzItbVHVhs5c8zM5e+ubq7lMZEcBFD41
6PbypbCpJkLFt0Tw6lv1PUrVbE/lJfr23mwJXGDZm3tppqGpoCI5RDBx1aaqNtWL
8m/kgf5j8zhN7YmB8Xb1cfWznqlHP81Lqb8kGvU803kxO9ldjQWp6jMFLbToQ3Xv
9ysai4oEoBKuR2Xv8nrmekMfYNpcxmgjDLlAs2nMIEC8OZWKEt6+4Sp7F9yjYDMf
vd3cXwgT+Q7AF0E4dj6SKCkukIwXwsEFzPCUpeUK7jkhA+83FCgMqCrv0co1VoRl
E39740cB+R+GUQUCuoHp77+ppxI4Oe0ZhWpFHJIKFHTvGDFR3TKXYPvBsf/KkiEB
MqxxDC4jH0ESexmvEWE1WroYFOtZLqMyFSKtfAnQFIvBZBvzcN8SZptrTDx2sZyz
TGPydObiddnEBRfKYCw+0ZQ1Dbkv4w7lFhIRAYtSaWVH27npQxxbxyx4tDBnI1A6
7fIpOqU/zHVOdvqN28VJUMmSXoYRP8psEA2cn52VtDP5Uobijmk4s41iLFIQXcR0
WIZowxGz1xJoZLR1hTmlyOwfHgRZjydMDZsesC49ADYFJaCnh8uqE/ONRutvPBcq
72LWEzrI8exoiEraYw86fFaFr5Ggqt0NJmY5IfKwTKlbg7WV+uyaZYtbxTtZi66n
JxW+I/DV7s5BCgu1LFcysVZSBzc3YeY4rMV1eqHFnozb/uD92sJhusvkq4Mtqsl8
U3SjNGPdf0teAxcv8pCZKTZEH4NjvH/AlaSKOVWIM5VkDn11D7Q4+Jgc09FNmHye
fNQH3BzVrAX2yfqngLE+aXvIYBHrlh/OwvdxgJmQPHA8kidFXJS2/1Q5JVXK+R4S
BL/1IX1tokTyP1VLm2hz3pxRfy/7JqKIQ6U9Q/s6y18OCd1301mgu4dJMJBpe9wg
r/i2XYve9FEwn1waVGsCkWzfDSOjleDDlRiyFbJ45b2AXgBXD5WDpdXwT0YqrUH6
13QQN+Yx/MvwjNFKqdUi683sZY4yHJVSShjZ3xomUC22aGjrYFLkMzpS23xPUS8e
TIvzBB53vzy6eMpVMBXn7BwBXHzRRot8/KnOwKa0TqiFeFxDfWGEfOut1E1qKyfJ
0ZoXWh9fivFp8tzVLxskmgEeLpYYHIaPFkjncjzqT24WCoRgNQIItdwDou1hHhU+
BNiHcoDMyIuK4UpIXHPZbNsCa+3JnMW2hfYDXo0zYIInCejm958y18CLZ8N9tWb9
GgK7gylW0q7TJapL0d2r9Fq/Kyh1L286XRnXdxDaXXiG+MId7tvY3lWgUamDSjRW
fXUzWAyUIXIg0hrGvDTJh9NL0EFNehzcr0jRpD2omxLX3iJ253SfyyXyUueU7y7N
JcOTsDomhEs/k5p28Qe+c7UuYt6PPtKQ3VCX5NIg1mT8VPH6mIjWkmq5UiSshwN5
1osNWCe0BBis7Hbp2Cayt6JKyu1q7rd6Dy61AEwp9ObZyHOk675y3gAnwu18VBFY
d6Ul57XGoqGVq58DVufjeg5Mc6ctlmgYTOYuAC71CxQeG4+QO47IQHBpYbOrYIcb
GIvdbl+G9cLTBwzpfI6TzkcNqyUk4oGjXtBt+MKVSKnyr/aT5gVIyfvL4s25EapP
gqbFfFJwkRxzr50+kE2orM1vMzSnkjeWBRNE95Rwi4gMgKVGsIF1THzcplUvvZat
U0W/Hm4m9oZ3nrWrYePk94Aiq0BixsMyr5EC6zh/vJzXiLaCHg3KwfCsp6GkQqxE
WJ6cdochbHgOuu3hliQ8mtBwQh9l3Xj7ucyezKIXiIDRYir3T8tBFcWnNhjJ4hjY
CrmqA5+BFa/XQLF+VEcnI5Aedd0uDmMbjNNujS3PhYnLnraRY72WCy83YOk7r3JA
8I7qjGkLkMOI8+dqFYH+IMrNFT8sPlgN55pS09eHgv/DCE7GlsKTMUYKWtKFEHAn
sNxUPspN17h2/Ofvz1qLLPREXNxsCaXHohkmFM99F4/TFDMnvh/5HYZpoYgYtsvV
e8s3in0nC4tXhIVVV66otRbiqGnyNViwNKLGl8dyr2L8OH8FniSVw77MIeNfYPav
UXFw4ATia16jF5Ciw+o6/ERLhiFQQwH13UBAHq75/ATxfXbfQ3D/4xLjMkgYWukg
81aKIGPkwHQmW2Un4vezS+iRclOI7W2rtnHwmq0FC+euNwnAAj5jbcG+rFr5CqfU
2RR49nGmXKbvf6tloCDvU4ryCvcr+/2iN2cDouB2jnt/5wCSnYDW3xu0cVc48VVA
qBGI5mhy2lZTQiEFajJ8Cv2BhbgcEXuAH1kwBERRyFaonYf6yxKHhCWJiop7a/t0
om/0POumU3wWqgFhodzwggYwQYmB5uuptOJRYLi3poi7m9FaHe4GkDSUTUfga+DJ
FA9LWWN9G6bRGaNLk29huY7T0fv3uySY0H4LUqAW9pKEjniDI9G1jTqTva5swDvg
rFMaQqX/oHHEvcSX+O3VuYsp7MJX5jcl4liJLXV9JiVUUGBOF9Zd/iRbyX0h/xkV
i4tIWBv0HvUFNOcgFaho7ZSZBwzNnyeML669jWfx/QhU/3nAXQUoBuIcTzRl9jAu
L9/Mg9PqzUwLe9ngTLyJ2+LecCaR+/0Y9rnDn/yczlQCzKy89DntkNm9tfLmv15Q
qg7UfoE9tURiYvGQc3JUCAAYhCFFyPPn+e3WbktvUQYq228cLr6rrCnbJIxlM3uY
ZHrbyzYo+Lk0qQu5ggCyxDLgtgYJzaEF60euey9JtY4EzCrTUfqMJVaKXxsgZlCN
NVu73FBfB/v29SsVqzGzKnp/ZnEwrwd/Y3mw+Z87u6/EoC5yax3oEvwxjB8k7San
oI5HrWFZ/7sl1IH4rZXkDAkzBVFONZwKUkLXAr5p+r2O3Lo3ao7bUNoiN2pT+4CZ
SCQenfWyJKl5ppg4DqqjFGgUAADGV4WVD9lCCOyGjW8zIHy3MPJWM9Ti/qasZA2C
XJaRjQZBXk8fHn30CZYhvGFeA/UaurwV/R2bSUI8KLvkPpoyP8HUlQpDVeabKS5J
ihK16RzRZNZGp4FweCbV87gmpkMRaxCgWhx69RLD/CkEpyrXIpROMuD/BmqpIsTq
kqvnuJGEQgXygzPJUuYZtOqb9YcTHAwpwUIf8+fdGd4CrLdiw1tJbqqpXSvuQQYI
RXUxGLDgfr1qPF4U29FAnHiJGWEibNCgRiGcZPHyzszQENR/KxRYhB08CUnPCggZ
i3pjyreOgZlhRhZpAThytrx2wK4B1x7+3O6CJlJvTOr5f8Ycejnk9Xfz1PBGwGwz
`pragma protect end_protected
