// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:28 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HGDWH2fJQXpNppSBiq5qqEdA+C+IzbiDR2CE9ohjkOwuaLhTU6SXSL8SN7vwo58l
bhOzdgOb0NGYq2Q8yO92Na1ki9ulFXX4j2j4QRfox4EUk8o9RL+oFHhtA6ceRHYt
h58Ndyj5GGcjI+8HDe7hsOVWIOe42vJSTaPMKbxG0Ls=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
qgHoDkz0i4ugohIMLs4opWPgbZWmgI03Wwzu2O5o/QVhToDkh9Z3iiiuLzh5MLDV
G4lCgvxkb6tJY+u3m6MTYd2a2R1+aZKVyCm9CtODAMY/Q/PjUL5RFo4qZQkjW1l7
7tBr7kPAU0DhRK8XmxbI20uwAqBIKGaJfcqMzWu/2rbdO+AmHqr5FMjTwnHQihAd
H3ObDO0pumqXOSAtACGGfcXqm7OYaFEI6WIROpKYvmbpNlkrQJVK042NgCWZQ04S
ixYk78lmQZ5Lek+k7KwFGsf2J0DxEgLqN6qyhvAx8OljuCc+9VyrF4KWBbOPjYaU
pJDAVRfkHUvaSDqAE64R2qxdB4Sc6v19zXcUwgI5t3Uf2gKsJMZaCofAHz17okS9
D6rP3wk/9FjFV8yXMVFTHE9ndLWHn766p9xgo8loAv4WuDvhW0qx7oGvOI4ArQ9Z
1mF3VBz/Ae0YrJfFh0afppHgx6MdglJUZxDQx+0aSR/EM+ueEGos/ECu0lsh39bq
muodE71TQ3+vwF0TmUKvhgMub0RKe/IovxgKwGAbSxJ+GB1vTkzAvm59PCGw1Lbe
xVZFM+AjPSKS2bmWXg3i9ifdHbivEQLlqMo4FGh6laSXT8Q8u2UAkEh/kt1oZell
jDSOmCXedQ39W0JyoBAwezOTzqqVad8IQhd02p/eCYzU+n/+vMOR7wK3al4RLaDe
T7t2zoWpEIfefy9c/paSIROTK3DNd9rzei0d3o8WvpaALaks+JzU6D/2VY7VS8s1
Qdb0EozqHvrxjjdgtLeA5xz+XVsO53Chf689p8btQnLieDtctBQEAgpnfO2GAh07
ntFYTFcSnDN+cKB+h2nlowp73MFN6SnXB19ObL5X6q8XS4BdZUYvVtdyDL5QNdlo
AEU3BzX2TS21GBlvwdwErjnMTcRcen7J0gJp4jYXbLcrNCE9h7T07WnTui+D03Tv
J8n9Vft3sTfJg392fk0gX+or6OpDhJ6o2BDeAWI25AlYXoKZHFOmnlJ16ApSScd7
QjBjOcEKFzp2Wg2ZjcQ0Q6akABe/0+E4JhUjbKtj1pmLrUfvamTOq1SUz1Dqaiqz
U16Jix0hS/j9Xc3APmSPWJmVgwQfUVZ/Zl3iS1Vr2fnwjYyXvUDr5g56Vto8K6nU
eZQm+uEPjXum9Cq4vvrRX8PnD4LqT3aZrSyW/ODkh7YKUH3eiLTTEmHF8GnMUSAX
662KdJ2qokCWo4KpQNUisSOjifbk58UrW0FO26zPNjpKyZVm2PazGbTVgONrw0U3
yKSZWQKg3rhfbEP1bfjs+zeWOrXDcguQ5jVYz5HWJic/wbMXQJxra1wsqtcEFiDi
+7LDWK/njr3eDQLfFZBe1JU18FWAO5lqi+VJOYsDOzd5rW+CaEwgUfkRzmfBXA+j
cXQKFdxKOcgNg9GHxrSs2+1tVaDOa1sKs8BSErxFLaG5evuHUelMFo4o/jQcyI/O
apAS2DVCGC/bRQ7OUNDqE1OBLJHCawohAD8ar2azQG9eW83IlrmOkwjg/lF3bC4M
oKq51qR9J1zPrjuQ19Dkz7PXKnLZYVu9Ubo8I3P+aLrMk0qYXmtYSEt7ay95WXba
CnjNxYjEcswm3pilmNyGj1qtHvh8/LPIAlJXs3eeRsuLJP6B9RCpCn7ph6QS3PH5
6csqUxH7O7CZWgjYVM2SSZQrR5XCFEU6Nhox0By0ZcAxXIGgJf+2z7cCR6wRksxH
F9Mx/ZwE281ov15l30PAWDOKTszmuD7jS+k+XFA2OEnAP/AQwCfyhCmxtVQ2MH4g
9AA6VWt0h5e0zwbv7P5g4mqGQq2jz6pRR8t4xvUEYwcKYQ5lqlzm7zdSrvbEXr6d
/VTJcJ9yzjQWGGgaK9SncIVuDAbi6aqoeukmjocsxXMQD93nid9I3bZDEp7fZGXp
W/Nj60iGbR6qSI9n+FH987gIbEwoyT9rhJig9kHtwQtKO2/GQv5wNccLW4gQfIB2
oA85140BHXz4SQw9tKsnOJxhPMftTfADJ6iFQ9QU+lGhThThhcEVyElLJdcXObr6
+6D9wKj2EXECkTRaxvupoE0Lcvz5IDnkKGNw8CTG49EqlteKgzNoEygd9g+RcfLK
7Sh+hhCof7V9TaR8hB0qlsKPmgQFYIXkDifqfhzXMBdsd2qf1WOeqLL1rNn/ATUa
awIHkrXBWHAo9UD4afYEG2cLSGCNDqhtbkT6bOCoW57IBChEGOyycdbKcvoTqjD7
irjYtVrI977H041vlbhzEb/XbOOMnIcqslyR95Hydfc3Y5eZuZlGmYG2vqlwdGgR
gcmMjmY+/AEueGpw/LA1xhFVKF1Ci5d7Lmwh+cDfKwUMC4kBTlQ44AjYdLtMLke3
awqdwoUgz6Px6AvDY2e5Pi5a+uNkRRo6e5aXNNm0lWwXr4/CRmui8OAFod5v0IaX
8RsLbNSubwOd/TtznqoIvAU2Id/ThXxweGXoouSBAtlwwVgCbRpgsEMVxMQrzk0Q
++znTd8d9/acBErbIpQX9hSEMm3vPURZ7xwECPfA0Zkd2lzZTvsY0I9Xbt6d8g9w
tGfaieRt3dd2C8aHBQ9oSzqY+rq3ERMQVwSHvYMJs9uWmCjBs7Y5XyQYnA4DutiV
M9488WEm0t8a40nYz9IfmV2ujhRjeDZfWt7TGp7BrW27xjoavsoF1P40TxLjyTXj
AnRr5cZoZSU0EA+3HEt1A0+JaoynavaxwidRe0CYOToKRs0Wv0ZdAQUcnrepgUQ2
/Ln9tB+Vjb2DeASe1AZjzTFQ8bPoL4HgJ+RUM4lswyeQXX++uaGD4VX4SteT+B5S
iCF2+7h8I+ik0AS0yKb3pFBFqv9ueYNp/W98+TdNb3EVkCqS3R231fShnIQ0L/1V
V4mIXgMRw47OCmiio9Q8AqqTDzC2j2F1+7PhBqEJtE1cPNhHZLYxn5u61q5iHpi7
rRL/SNlJf0l6s6nbmsbJqOF10fQDa0rTxkv4sO2oUEaHi3Ak7VF2uCppF1KhZ8kt
rhpvBo9pFxZ2c3B7xmGxv1wGHFsA3jjji0UcJjEeCeJmw7l6kDuKbcKE0Nk7nIk0
rF4ES19AGMNHUtmj2mXRPAYILiMb44LUDRA7wIDfjHE/K8ddEVV/ZitI1j2E4edH
+snvtU1PRccMoR9eDFD+zAdrd103Jb5L/xkB0ZpeDghzlDjx/aKUUu+YAPOLUp3D
OtvfPsDyHXR23ubXgJY0BNmkdQPfq2q0bwTWDO1FuiexThzIBGBpzAux1CwnJbs0
jeGCGKQ24PoXVYBBLvU8L26mR2hPq/thCF71l/5F17dwS57CyMFLTuQgqw4bq96W
2qDfbdd5bXYFs2jDguylbfjySgqmx0iiW/0Gq+K68dy5h05BkbdSzrHxYvh4iufb
zue1LXkIoGbEaD7+EEHojol649D8OJzTqoVvGv/CejSAEOYDNptr0gtfX1N2fD2r
Pg5jiZperIDANk/Ih+ARY3NTFbKZO3HT1Elm/8zJQEFl3tMjXtccSxslfW6gyLZQ
4Cg9/yP2wuPg9ZGowNROoc0dRi1g/UcFrLir8oeRTeFiXBVDpv6TEjWItRIDsoga
bz22k+S3JDNTjfCM2Y0ahxArujGrZ5os1XtNy5aQspsG3jUbr6UNgq7RM5vdBk3A
a2UznaSzZQz8lmtqP0cbx4dd/vcKjjd/VnpIeeWLvrlB43tqLabPEHHnZIf8F7xk
9uXz9YpWB6Zok/nYtIc7/g+nJbkzon6sX7Q9qImdqh1ubAgEF4jJ2mR8Z1nhXWst
TFt1u9eoHosZeLBA/0CcezCWTJ9T9uRI+XwmJO8rgDXfDdrsm2ydtoVlNdxmD3Z+
Tn6GkzWZp3IsLYmqyns8UsvnjfKvVi7raLLbuxdIiZUDT9vU7779qeieBP/CgO+2
YOyD1P+YgwzGh0PksWxqOQpX3daJgRqtwaFlSdd9Bh1YahfB5tTBwCWboYlrH0Cd
9c7MGTGqT4ljDCdbvOGot3mXl/DhoFIDpv0xsIVaXtf9yPIyDDyM4mkHJE0emgL6
rmOlPKEOll+al48YxE+etZja514yB/8W32VTdrOdkIHICns+wI4AOGLctiwjIzVs
rwRAnmdv8hjzopqtqqYF2c4yzFcTmj6bkNVIlw6a7LkV3BIUXhslAO145mRBUyyl
Qe87SJsjQrs9B+5E/eIaIu+88cw9bqYn7YrExJv64/k9RMGCJ9H/vWMF367cC99W
mCPeMSjHZl/eW9/YJYYblLNBY50jl1U3BxrNf0g2jo7dovOUGFnoV4+NtDHpg2Dq
rQxBfYohJMuoLIMCEPtk3mJ/jf0x70gwQz17ia07o/S93l6b+HjgQrC5l1t2oMTg
YdflaHlv8rwuLRRk+bjMCHAB48IW22K/C5N8m+VjzijQrBRY2z6dEOtpYmlDuPP4
3srmI8LfN35QjWnIVru5+GZAw7b0/aRADQLhRFBCA0WlO4t3iZpQ6Fjj+ThxF2kf
j65MxgoAO+5avY31DQfaZ1UEM5EMZQHcw5oMUYU/ifTHw1TL+4NEBRiZ5RCt6+fy
XBVMbNHSqiiHGyQsxCUz55gd/Q0ugkxj/Wchx1G2Q7+BsNkm4eExxMRxTKs+ohbo
yFR1S+tbfwbmLkzKYs+onZEb/8cE1qi126Df3E4gYmHzcc6+yAPU302a1PQNV5b/
GXXoItZFCsZjjwEfBxUGfaFSYoi8gBb6RUsrk2k4lBzjmy2vujTC5y18NgGoYpSL
Zz2JAJ3xWQ0wxOeGuLfWK4wXbcw4gtkLIoyU4j7wVMgkAMUz5Wxd5+qJXGo4W3Mh
mLvoDiiKSu0OBiIX5/Bf7e2U3+61FrAWkgf1AscGqaiu6RQHxYnKVGxwE1Jvv6Be
Dc4IY0k8LmcljUXWRnADUXxdROc4HvH3WlAGNxai8UCB37jRemmGKRFWwtUQJg3J
CJ0z7KUd1uDW+TRTqqO4EWLgvbgDg2pDW3gSBgmyCL8xhbn8nVZTE3tyDIA6z6WI
rpFOE3yvSfjvvFmo+byyA9hjCun9aY6u5sL5GUb8e71bBLqjbDpo9Iq2hVONqcK7
UZiFMfH+0QEw0oveT0nlPclhejgfogHSpkatnAHJKcSlMjAGeGCTd81cUiHCpNK3
W4+oMe9ifiA/pLE/CXyyT8j0xpfvHjpaJux+IKnI6lra5HEvpkfyrP3m4ykgwXfy
Sr6DI7G+JBwSc05vRdbPfPJ4pn+LT6Lg8wp8UzmAPia3FoghIZIrFBWTc6wTkZDx
UnwI8Up16y5yEqyVUB/xP5HHEScEwFW6K1wKUd6LTKVFc03YulW88mFZYh6au47A
F/Ll1rIUGJBeQG8iLotBUhJh2k2wlX0pmpcsV2giLG0fHhRPNNLPwNAoZWeIBusx
hl3VSMIQJl7HCCuMPrc/4pF47jEo2pvBHFv7qCyCqSQVzB3qvOuyLg6OddE0Klqc
7HegfsSnGisk2yfiPIYNhAGl/fKiPLMHWg6ytSnlnHe4/u9FY3MP4EYct2rGMmCz
VCsp7wEy3D1JkVWZjIVKrql5DBrb3frTzm/LySc9QAM/IDXZ7sZowo0h8SghCDz+
uewfbPmyTbB9TUlg5ojl/koB4GB+qOEpb5YZtsdwfmLEqkvtmJrTFDv3GbWBn8dg
+BdOudGxkL+5eX4tzMJrqqdB6h97S7KqSy0x5kfZ58AoV6nnqaZyYUvfM5HiD9Xh
uVyftE998Ejcjn/lJOZXBHu4LvtYZqeC/wEkvdrWWP2swy7NqwfX4iljeXkmJXQU
4SQs5n1mPFwpKUwVtGbR4i64vdWhcktHRahVEXys8P/YRYEmdT9WyFQGe/ZrS7tG
Y0MqDh6CH7ITOIMsbFItgYpXXaJR7LEiePP/tjpOF5DSkd9kSgZKCrounVd3is18
lZQ+rWSYfJOujFCb/6oMnsGclxeo/7EzWys6HoH4lcfOkeOUt1oW1pPJpu9rycAA
6L4Hx14mB7ThqOAq2yre6o23lnGgV/5ncn7afwPGY3oWUQ6suHGtQrc8GOk5PGOq
KT/YEJjywkEcicyLq3eKORbNr11rflOTNpk0Vux6LMBlDJK7gHzydqMuddBQFWBp
M3h9AJwUBryS92uTVX7hhalXFd7LBH09goLDILC6+autuW+x2e18Y8bgWxPvZwJd
8J3oMNqfaQ6vt/37ix0LE1PjOok/vr3+TBmD+IOvHQZ8gdeeyK1jjHhvbFhMraEd
GFBeEPOo68XaoL9LphYGq8d0n8laVC61KL2hGBPtvoDgopDG7tPEtdwf4b6BZn3h
bNsGHxgdUbcZz3Eq9iBWuRX/s1z5Q9+/CmOjZv2mvrgiI7++TVXJzVPiEgmUxt6c
5D2c2iXSvVsJAdl2Vrl1ZwKsQWu5hU5NCN3iqrCa68mrHRJKj/dOMo4dLjZIx/ql
Ie7hfsH7OzoYrlThQwBlv/tGbHQ41Hx7k/wPYbaYbbv7Ykzjf6zEtM+m5FKhdKsC
pGuNQFGhcOia1RIGcE4o2eZ8+/1zqRWWUjZ+0pDRcwAghvH2jQS707P29NyGK4kx
XEUFDA/r1IvBdXZUlewdWYL/EGEZ3MbvfmK353vow37eFw8lp8+NETsgEhLyaRZZ
0/ADbUqIfs8uv5FC7KZLxPUi5KxqPTbsr9G1RhIniCm4f+qqQ5CBNXtBCX7dU+Z5
wkEPnRoLAynrKYIuYYO9yIbPmTZI/OfH8vxQ1LrHHMcvmVKq6N2dKLXgZtiasFnl
t2XuJqnszABLlHLjds0XiO7SR1OAWy0QKvBYKqj/iSL6zPVcvHlvRj9OLtbSkJxg
VisKwY0395z23rkITAsErjLQBuqI+imMV1YBOWugsDpMHLIae+1KWViI8EkReS8+
U5uPcJy6Xso0wUnoSrC0H+op44fFibofJZMImNbfBlz8PSW5LKL14f75nDEWIoLS
+0yW4Uajncc/smSzZe/AWmtyyCTaBabM/pIWY5s/ouqzI/VpZCU2cR1QVfk0Uq6L
DT0F79NTEc6kibS27ThynJDeD0rJbPUrRz5HOhmuif535JAP9x0uXvKMS+HzAkHd
eR6oT8RVXgKuuV4zeAg9QJCe8TgyH+/kzgM58V4PL+8YjiI4HDKDEgCa6xH9xjGJ
2Kd4EdCR1uv4jgaygQw6gEGxpYEa6NW7180xJC1j9326plkJaBZcCw1K/+RxHaUY
fOwElY17rxuNVJIAPSO94o+Zv/nVFZ0wbCszWAUdX47mDUTX4GYuRLEwefuYXvJ2
A0Uo1S6gEduz3zoDoqrDJ/hG//Pij2T3FnA0OTd1efvIhtHS3p0c8tGnSFM5/pzz
hwdp7akYfUgE9HmGxxkXlt1BvKIwv9EBYJGBMqfiLxTKHqveROoZt90etEsx6SQC
JtJaF1q4QcRtHSASxUu1VEEXraFVT4H95u/EKHAHkxN5wsCeQEoJpYxW0jyDzVaN
ZI8G3vQulJmNP9Av0aL28CqvFXbu47WJO25FmAIXZtYHi6RU+/ptpaT2GgpYUPSz
8LShSpalQEbL9uy8IH9u3EI6G6glMnKnMZ5IQyUdOv2J5hQaeK/cLvGyrl3Co5/f
aO6trgOL5SAN6Vv36qkOf63C5eNEjFbLgk77UxvmOmytYkvL8Xz69JftlIWJd/1H
VygAi/R5fYhOJHswyEf28y0LDDK/DVOwplPW7x/OmVfVaWJSU2M98zI9ilGPeaxW
AT3ePJbdjRA4Nf+g6db0r/gSgqFIrQczESylC3s+8I7cKVFC/NzMJarEBCv49HD5
Hm7qp7TPvivWESfqWIVoIDW7GaW/LnkPrvbdqZHVl+/4N5IP4VzWtxj+E0R2A2Dw
oJxgZnfbEz570pVV/k8qkPH6iPhfwQW+kZyWyYjM9mORThAuiUvWKdJQx60Kmu4U
FIcn9diOpPRgO3POTFirWXT62+vMpNAl6nLurOtaLzuvIUVU0dLhx0M/w9ueuY1b
oseYyzfQ977sGi+z7URKZeLrylB99PhgfEH2K5Ofp9FSNQ9unNMqK5SJhOFvSc5b
RW/GTz7Ak4pFO9e7epV0gV5oC8zAVdoRWrpc2GPiidWvPDdpb6K7V/fxWBdqeIp5
RocPlDrW6bBSjzfHDjY2glTBgHrA3J4km+MFdK7ez85PfMEL1dNtNyEJJf99/nBs
a/KCKuZUnO7o0cV2C0UkxM135ePG7y/Xl4lTWD2PP7M++ML6qiI9r983oy2trQHB
1KUlBOChz7qQDSQqZL8dg1ev3eJsc+U7HEJEt4RgWn9ZaHG3Dr48Buai5175qkd4
C9lxpGZ3ahz2t+K68ZiOPyd9Lm40k5IbICFhY7848Q15BIRIqs8/Gq9bEe5CZqh0
8J6iP9e/vQuHx5tUhTI1KhH5IswepGv6TRFdXDF64k7Lk3MA+ePNlMZ62I7qUxKM
GrOfVc+4ouDNGPiDc05XK3W2S7wpaUh+qozLZ+ZsA8hgskCoZQzp7qmOEDEZ8tMe
g10nJJoLqO54DNSpp2Aw7QpmQ+3B8Bpi3n/6+o5EBrSnhZT6euJF7dpUEL5jGw9S
ASzZEwwbHOQ99L0SiniS+5rdeCJDdpM6jML0ayX/EwWnm4Fj63JYKmfrRpIRV1Sj
6X7itRlS0nzO52GFn9YMrnU/AUlepoBQBEnmLxFNgLuzooqP5Da+IJbe/Ech/+lw
OX/4ajT4SUk3nvVGmFxk6Kw4J6X35TyhFXK6szbxlsDC0JbQjiad3GMYJO39PAL2
Qo8nB6cssIkjBthK7McBR0XJEZRLWAy+sHpA8v/iUuT/ZziS32JLp8SSbCmb070F
VzUoYWjJ2LpaheBWspu7bKniBM9QghTSZKmFSzf9bKjkqD0AFZOg5TPwxyHZuDs0
svEpaD7nTlvDJevke2ZD31pwxNz/wOAaaqjcMVBOvo8tKcJ5eDDIviUsPfrdZ5oP
HyYFOF7SPvrnkohilAGSS69yc2dRjBPVXMv567kvUuiYAoYCknp6FEZuv43xQWgl
hdszWKYh0hdWlrybGkl3xLH5qdxT7xu9Z5qFtHKqq0O7oOOCDjQda6rAZ2Z81FQP
nroj9zHT+1m46hXlIcEGdyt+m7AtXDtZx4BhS9idVlyPfPDKy/3P+UWEcfJnIJw/
vs3+Cq4SQwvnIz7oZZCkM6P1xuQsB+Hsjof9cNLGmTKZmx1ovtyqlbmtbezBGjRk
TmYvML+8tWZ1Akd80pjJpq2owcIUnSH7yjvCGWje9RZfXGrRz2Fv4zaZTKIAr169
/j1upvhMHKaViKaIwPldtXiE28+Bfzl1/B2St1M0kCNRUyoRs+01kz03HgHX1xWt
Ky2rkKrMUTbxQ+PKLOEY/Ki1KqdxoIUnSuWgMQjlbjcnKTpvbrTh0N4qO7geesxJ
Ohayt9eL9RKvnSn0Ni9faN+YipeBl7+cTncO3OH3HM8HtJyV/yl20wP88PC+n2Se
0bjI6/FWdXlBU5ZEVqQMuCkMYlE2NbBqAr/URYhdPvUnykKtNcC61GtZ6ZWN4mOE
dfbBwmsdojr3uwTeysjQF1vnGX+H0EAuvjjigMGYyzndlr0ULHl4EF364fhzVFni
MY1iYbGvOihTydYvGfHVQMlQH6T5uv5I+edhPWmo3PGdyS/yu7VcWDkLpo4KlssA
/sKhW41qXS5s8LrDxerqa/ahSHHkpeLgI1+CdlwTg5o2EKbKKu399YKmSPiniJGn
TJR6TH0f22asiPJatu2Ydxi6K3mGvOdYWVv1BuwKpCbePgM2nyeG38q8nE9egPbL
hH7ybKUlS4ivblTT14SJUHAtFf+ip8+auvxhJ3vzLxInn9QAYrJ+5i4Bfv7DoIO6
v3p9AmHmWbC0RXkTKwUr8pjMV6KFR3eJAwge7MfLVmLsO2sSDiLhPcQiBb3LpBC1
w4VO5dZ3Ag5wJK0iRJ3N+rlTxK90VudtKKTUKlPM9SYU4Mc7fROLLmipXp3gOn7J
N50bBckQnI9q1XSReE8HwXCDm0uUwWT9IFbCsUfPPY/rQRcZoMi0pCGmUXfHpaY7
4MCbVV1ZMrUJcPMWgQhF9M7pDsJ9Mc+xTLSB+N/ZLGubQnzZW5JUiBQHoyyZMnhW
yev3IIbo3ynrg4CXp9cfcOZFZeEmCKtkEvvi4dGC35vgnQREnUf/YFZJwrfYgnBw
4VDwPkxyyvSFN4GTzo9A2YlE5jHnpJetj1xjnFsQRTmjSmRJMKW3uQQJirU7Ggn/
CdjT3wr5yXNyH0bUeoKcCRlSuWp2u8tXIb5VI4VNKARxIePJJyQpinIwrzTKqv0s
sqe2HMSKYA8gEZaNGvvedLHVnnlspPJnw9Wgi3FkR3t5Dhw8evVnP1Y/noJydcX3
Kyg1rAbwydba9isX7GffMabpZQ5zhRiw4RrSZyQ4REzBh7PxU0eYRS38wbF7cWk5
lkJ3OcToaVXrGqatL8ZtWbMzvmn6mJSvhdz7/1ScAZ0rv6p2HeTOazUdu7/IUtAh
PfJwoDlyhlLazN5M1TI65TJ+h3U9LJLvp5c5KGpOBPSrY3RB/F3IPvyK1cvo2kMP
XLQpRjrYW8f7MM+n7sDKTg9Vi5QnYKovTAvEYZHfj7o5D/6z9i7dFG7l6+m4swv+
8NJYj1R/Ap+zXQB6hBRksIGWKVMR0zbFcm2bRAok2EIpna/QjHDNeRmcjnqKIVGm
Ctz5NT7hDlLccIYcCVSaxLdO3kWov0gBB+x09R/s8TbJ+yNaSVlXAdQvNOPDikOe
ymihNlnD9YGT2t0NCy7oF0IX7on48+mzilFUPYoA7xsDI1TprCBHOuqxiexkMwDL
dDTYaylbxOkYIX0778zu88ekmA/OO1nXDLI6a+JkFyOjQK81J5DQioHXrAp2Hr6F
n608k9X2j22pUYcC6mIaks4DZ5MCHETW9KciEs8ovZvI/5y7D/GgGHCOZGOsN8Xx
eVlXG5e8Jkq2Uw2FSeTrGAigeH6jVR2QbBw5XSRpRbhtCdMgeKG3kOUvbnq7xa6y
bKOXjcb9oDWoKsU7d4OaLh4yo1N80lcFKaiwRr58DXMTDC39HT3irw1REbmSxIOD
1+ziWUief9eSnMa7uCDoBSznW2e1UTNAt15K+62yqSTVvHtELkgFOWcNDBNo6wjs
NjZIyZr8CN3BR4HOBfLD4Q/dFTE+856VtTAOUzShhyABUf+gtCiTtU+28mu6eV/U
+/azq6sQKE9oDq6Q8wZMwli9mE8qXof/3J1Md50XMqszjShjpX4f7Pj3O9IeAtx/
0saKIw+55YBlucMPrgI+M2RDRJZ3vz93lIvhExSFRfcjK2mtqWVur5lVDFU2kLfh
xDr0RzbWu1o6KxEl9J3zhiWCVaAT44hf11/d7I98foq/lh637Opun5FEaG6UsGiU
2Y+mqp+6uTeMTs9k3on6be/vgdns8r0xdKowlgCU7IrKu+VVev/RKSpTyfPv0PYf
HnludziraCdL1GAgs+9/xP9cffSeHFHrEBIBDWgk/VB43/BKPErMSPfR0TdlhhqR
f6XrwH0SoeNMgSYXtQtuF0Hdezk7htSvB7FE5y+/EHuLVxlVS+ToXkSsfE2T9C4C
8JQsgc1Hvb8Cl6m8FIXo6V8PrjHB3HxQVYFfC6njBhMKuE2Clsv08mJLK7RXRMN4
qdZGWPkzcGJ6qA24BHwfGRjn9nshMBWfzIrvEoN1tdFWfyAI+0nbh4Rc92ibI9ub
l2mQjAUKP84L//7RL/i/zEEhcAL0wUGippLFbTehF7y49LC5FIlFeySEEGdLCNUf
G2CI4YMnuiIUXZ6u2dWfol0PKsHYNWm2XyyfEwl25QVjmRn9p/iC61zrxCmLbDAn
JnVKfNPVm4rjhkYGwxp/0kacTnhL/o+RCrYWow0PeYT9DxjLa+Om2DLjoqULvmtD
F7SCKsiy1frp8JuWjKojuOZYucx7/+5A/2EXGs/aBtOzlKkOS+x9rbsh4IbHB5o7
m/P23N6BhjxDKfBJjfi1FfvyWOwy+ZwVVxECAfXjyzZ++kG5WRqa+gTepJfBf/og
RGwk4BAWsLMtUbJvpahpRL+PFIls+wq9Z1dWQt3FrlMwC8pt18Att0nSkmltcCP4
5F3+faWBfyBdWu8r2Pcy67Aei6Un69sTyB3AUaEhr2liRWxm+DlafkJBg3wy8oKz
+1eT/EJoSBl+YzOXv7/T6N2paf+crKb+k8rexeXJGLRAffdFzmK2LCHDmYWNdgJm
e9vjrVLkf/y4mNHbWfXQBSpfuuPSx4P33dbJtCkvmJc82PbMI/IFYmre1iadBt5Q
XHIerie5PI/dWUC/wEvuJshr7Q4frVkUEPYmmbPOQsINUhtMYLRxhQGpEO/mWMtQ
hmJffIyFIi6FcAAg8Lvt9Fm6IOvEkbCQOUZbwvhLq4GTiChW66CUaa34YZDspVx0
aD4EXCn8USerwXKqXcuUO7+dlEpj+j2C+qEIDbFjBHoHRcfgPHuEmElsApPL2wJu
QPYXvZBSd3NDLa0/WgsGQ5iwcx5bM1JE3wXtqLM0cSW9wi2Y/Ofk5JVBpsssBf1E
4wzH5ZtH1utx+hqGMeo14ANJq2mwVVA1pCelqUAg62G/CB3gtt4vVPRgpmdY2gDF
3kA0HumJz/uNB33sJ0kxRG0RNMPDyduenayt373cyS0O73TQPm9tBnZpeV/albby
jQg5j0pAbXQo4OsCRhaG+LsHUoW3Ht3uJxJpAVzOzDE1wzU+EaiCYIG7Srt8EH3k
kcsJ7Wtq03YKC+877344i5V4SL247k8VxGO5Svj3JY9ctpdwcVzcNggP1144Q+P1
bX2vTxMW3IH/jpuiy4S7Lp9hLk6ZErfx99EgYo9BfOMWAHgN8xqO3EQTbBKffrjn
E+x2bHL+cKTYGAkJDpHkLUvlAMxc7Dnd6lVtaZ0wsprED+cCZO0rgq4wig1TtGPl
zCzUwPUtXhyJ+Xznv7NC2wVj7ZI4KzMhPPNXFzmlU5A0+39uM+5l5rUAOtYKf/Ca
z31GmC1Mhn2myElsKZotj++tACtqRnrmVpBEfdO6dczbsuA2EObsS95nMiD24QJT
O1Oyoq21Sk9k9tLXxD519um/hBSxnCeImeQF6hK10ac9DL+Rln7GgwLBcbb+9Ro2
EpQhbDY+amlKDb0b9HG8rQ9HR6il15Pv80GjATOp6J9dMtSwRG2VqvgDTqebMmFH
`pragma protect end_protected
