// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:22:06 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ov0UsfGT97Kpck2pST7qqLuRXwDARkt6TPqh7mPhXMi/a5UxCWNla+VXWUPnbbjQ
t+SNiZZJ2ug5xTLyTBoJ0yrjGtcR4lJgTEhHJfKuk4etfbaGR8aJBDpi733lQse4
JkyZH5gA7dhoi+O+2gm1mQh9PBHL/Q+9Y04qxpN6+7A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24288)
oUEVT2OjNpV6+nObuyfHHrsA5M4cLe9XTFgtfMpvilKnurA4oYDTOFUzPPxFhDbv
bHszGGaAp8+pphhxEz3nXLvDHFv+EZdGhXf0txdHUCZ3DYIkOv+MjGOjZnRsUobA
rLICiIesKwU/JevYYAwHVvF4X1ldu7Z/atuL6coUnVt58IOYMbWvythoiqaQeCAW
mOFLqq3ZFUuWLplpfczqV0DsTPlygIWvwwTt843m5+SS9VpnEz9eZcycjEoJUBx6
oK2TnIyYd3ofGYVGzUFLiV3H58tWbvxYE+5OL3/AxQOv50/uZzDhNYxDO96sg1oQ
J/KwTtXU3L2JJLkhLLSmndqkyPLiPRA+cKmDx/9GRHlhVVPXeRyjULJ6OVmF7/cN
9uKBh4Re+64qePlIc8qcfyAcGM+9AFaocYqvRKSHuFyh1RU5hMjovo3xZtfPAYsz
pp09Cn6OnAxVoeiUIm8fzc5M4jyWmyPDyBiL9c7eStNAXmkFx0tTHmAXxdusLJnO
7Twku403dbDcjnEUcIYQ2dE1tzjzjg0pmFM8kc3Z7JQYM3XBW1dnIuN6n/BqExA6
vor+Kf1HSzEUbwK6IdEtUOlxKEKcgMAuWlzVP3k0BeXkA6tB9ETloXVrqSBd8Yox
nwZQaqrJdN3HTMIOAXqg1NYDxrB9EwADsUEuyXv6FnmnVMfhAOKWDdSLXG7AUQfx
hWxR+1acLnqYMCq9fwLDqplNu4dDIwHr62ymBFvbfp7i1odt1YjxRvTaClofTVfK
vT5ofUYKeUkUgRxjbE9VhxDGmmnN5G1VeyVfJuiSha3i+FFHIiOqc9n0MPkK0xNH
9aRgJiYpomGGkxHJcc3JkSDWtnXErtcXWWYqV/fgMyCDEAlKUYe+xrb8oNdM4fmW
MMSAuIKiEWAdzrn6ls4KAwyJFk2H0vPDf/eFyk0uhEvjoacjryfJ3fr1mxw+amfB
gmx243pUscJ5QTcZkU+nHM3vfZhoFmqc8Ub1QUeWFhuE4mRPuisqK8+FbWfyloU6
8FgYQtaIUw4Rkkt83t6MeF9QNFVOQy7D8Bn2TNdMzN5fV0zCIz5hiiYZ/Z5vBDp4
vTRhNOD5WP5R65pn2rEMVO5U+gmrCdiwR9i6X+nnXmyCJZl8FK2Tk67O46K0AGKn
UT8UKRJsoibTPh4lwNmYSfZYG+PXzXPmG592phKqGL4ed3vXHGwDd7RQHO6UXWmK
zuuxG2kQDmjZponA1PFqoBCCYsJR7WHw3u6LJRByhtXZYbH1tW47zS5sljmuMvth
g00weTDnXTnw1M/CvKVSrm4X6JrR+ZlQ7cIfyrCT9Vsat5tP5EuRnonIyz1nGS3A
4CvrPeSfhbwilIlp1ECgE4FWzw1QJAr1Tu4tHT3eUSTG3AvzQgggxZa9rLlEnUax
lMb0/jI6vUXI17xpHWRY0NlmhYzxGBDr+uXfh3CcCf2wMBHJH16kMrLm0suCAHQL
K82ce+DZFFC3u7QtGjxZsqOvx74L8KblckG1DHIRiQdVsON4ClYhsGl76+ySIeZo
phxP/9FbEv9hPxMtdMv37PeA/2lyAxldljNcd2FjRsUUtma++MM9sP3NmPiFnsMn
NQkvtI+rsXes5DWi0gRSbtxPQ46z5PuUq0SCNruHoTncCxHc6AjHtD+81YwToGeM
A7uWrjfwUZ9cOiSSW0/Hrt16OpPyVZY/AnXIjVu8Z75gWxMlfyl6rbdotAxLSX4K
sOkHPRRjMjnpOZlsnTYGbCQlWGFkkCU3DLEuGXI8ZLPoY34SwW7nz4KOpxv/jgtg
YK68gjFNkRArrFAg/Qf5qeM5Y5H0mWIvZYKxg/d9V8sAbYEhhIe7gI4g8Frbnb2o
EhuZm7aceixFZg436mZR3Pgv7cmiNkpG6hP6JVpYgkCMmGn3EM0RyRJuHjbbOXph
AG1tok1lMH0hxHAd2pi3PHcZp2kC/maUXHv5FHdaxfdT0IZi820gAPqkjsQj0+gi
gvoC74WErviR/mjHVOaUtYHI7XpeOhZyQKFgaER6oJysGaiFImkbMulLoEPJckac
Yl/0KyGGue57WdWFpOJFhLrNNWjCn2M6mtVmTnzKPfFPuQZS3gtl1cXemxvR0gII
ZNv2/rl0DVa4wQx3+8KivC5A57Exwf9kqrDSB56IBAzk3povb+kysmLHdK663dM2
FxBwwTvMWzVDR77SBcwaeDN3cTvg+yF3jbsBp6jsgw0rfjivaTDaohDwsz6uvjU+
WW58yl+nq/4PoRnAXS/V4BfWyGuQfqo5V0seGVYJRi5SpT4P10Y5dhpxz/ayTc4J
9X8ZWYdcRpxAwOMW694ZWFMETRncBi7sn70UHqkhmIj7hnUQ2SNAKpsjRb96nWOj
kkbVGKS/kuXPcJKzW7XRJuId6zKa4+PiCGBzT6JjGT2x4deA/JOFiq6ehMU7GBde
rK9ekz98W89ZnJfgkV5+zyDrqLJ/ObNZy5FsKzYUJ88omNbear8f65FeOLqPUGNb
MVUf5qQCTWSgNISQ7HvhHYv2Os1iu8pNOTQyEieRJjl53Np6be0FStdrnpTl+9AZ
t/NfvwtcwoQ/fLwzeD+ix6ke3qY+7UdcQWBfaESo5kZox0N1aVRnQEgyO3SrLRTq
HJsE3oXEnumAZq2qR33AlATx9gszIStIuiYYLLNTcoJONoCN1pkBAya+N23H0dX9
Akc8znvlpogi5iajfw9oJZrveH7uqnt+qWuPDN03mwrfdyqykuOD7/2v5FZb2AVU
eXdWQkAGiuOmcchPwotkwvVN8ecIjeHNdRin99+ojPdD5LCqfnn9i063HDNNsFjR
7z/xE7ATe1ba3itgPWOjhud6g64zuCl9YiDruQZujLsAjW6PYQ+3/eXY+TLB9e8e
cUUtvPynV2Imm/Hdbjkr2jYYu0lB/u9JORWL/PGO5/9i6mY0zywijmu5WUq20cIn
guGs0ES/8NqWKm2xiGsNmKMb+3R9nXNzi9ohFpnSRi7YS4D7bL6QekLFsecv43w2
ZDXtwjxyolBYrvccB1PxVpx3c6RHXl8CGQRHEY9CRVEuEsWNbK3LHfwWGrr0d3hO
SBxCqCDV9zwuiogIqZzy7nN+c745w1sLbz8rBDEKxDhroGyZyqRUY/bX7a2Jr/76
XppuqNSVb79UIAZNwPuUXK0+p8JbTy7dCQDV9g5OzPk/rWzxBIneoCqNJqE+E9R2
VxmAAojVj275mXkk0K81XM7r/tDC5JdKSRUTwz3zSirX2yDFiar3ZJqnCjpy+/wj
rLb3FggrD5/wyt/+h0WpePQtXl4x6Rfsl0iFQnquze/UqDdhR7YCpJfj9Ps3DeVh
9ixcJ9JENmUa6K+4BABWftiAjV9K7tixkohQ5MnzWDoV7VyvfNEDQHDDHQJloVAE
AJxO6QyuIb9Cq0O76NaV/kojMXTpiVKQmUTdktvca5dgggV8VL2w/Qlu7uzLs2i2
+QvHlRcHW/w3/h2CwfrtXByX2sP30hLYRE/A/7dk3j+1lJrC+G2ZMSR67P5IRpmI
ADwan0hQ0oGwcJ2srLzBlQGzPKne6OOPtIvZLl51khdWsfG/D8kjKctRxeOq4M9E
cRnVVzIPb8zFOu7dmJmPhfWqCt61VNJNQciKbukStE1hENm0H0V2g4aHpG9R8zHK
5rgWqD8C25wC6y6IaI1FGjnoSAVSV7EAOJKnwHbTmjcWmvDGxeeGdlF0aCMQNIyO
etmv69xOenPoHuMHtPnmLTQHG/wF0aMH+hBKdtwIujp02hPahoMaGsyhrKljLL4G
mAMNVxTdowxt3ENhBg02lyRlDo1pE3v8HRyJ/7SwTQDUF25oL3ANSxGRlB28sXa8
SB7nlYTjYuK81lc/Z5YRckTMESKHLqzRo+HiKD9Qaa9kB+jaGZQV/AmyzmVw6W6Q
ZFUk8IL2QATaJkN4sSkYautSdnfMN+ldRFWx5yWnj0kZUeDFiCC4CBa1Bau7+i3m
dQwRZlL5VOZDXtQh2RXjsV29ObiNjUYbLQ0fnqSU2LappwdTZBeYSeq5ctrHbPFT
ejEnXhWxskaal65yuLC/8f2aCTjM/QnPE+xENavk+2ezVRfVFC0KKUQpWBeFx+Uf
jydg6YiPVJnYnQXmDlzbdfpCqUmc7EB4JJ2boK8YyMDIkT3xQOAqL0JHsJ0qA5fR
+rktqtsO6PiNKaELQO7SR8Sc8+7JTn3GbT1VgFq9Mgj4LuwXRHhrXPxLV7DPylIl
3ZGUiHeuXAPa/RjBcGKNQ4QktpCsXFlxOCBYg/NnOwVsffLdSxU3vgwgjB1O6Lis
dnmsEqVJTzFXwTWHfGMNxbL+eA7n7VhIG3eYD8cJ+3bHvUR3TeV5JLZJLMfLgWNz
sG//wXr0CjwCOiQvjmowdipDqfV9mAGGaEL0BjuEgtmR6vf0D/IQ4gW0ywgT79nH
je5v018vUr/Qx2zwoOhY6HWikdQTVTLOOvgNBmfs8ayGbN5BWkkRg9QCov+V45fA
Sfe8+58RdeHUTRS7+BJLuUjKXsMzAZcbpJ/bhrzbOdTOmG5jzj4o3zYBL7F3T1XM
t1RQGvINwZlMaqlZoXvKjws968ujBcNjXOu1gdqF7l7SJcV8rGMMgLm4KTTL9CB1
Nhta8i2v9eawtHapqJfseEJdRBG1MFNKUnL5tSAah1k9ho6MJCr3N6x6Shn1Mhd/
NwUzYVbZMml3HyvwTiiE3Tw3e7ezLfvTB2Z9ezlHgqsEChUbnijeByKSvP93M6lv
se+LSfqaQdWu6d2lkbX3cG1jSJRWHcRCXkN1gh5mffjZV3n5vbuebW0QFYhZ8PXI
ICq5/I79dZre1Sc64QY5/j+4YQSOeifVTRjS+H+PtaR5HyjmVege0QhMDZp/8v9p
kTT+Yskcy6PLr1fg/8qggDLFfm5Hi8rpsf7CnGAvgDZ4TyYUPWalnOM2HxhWRKLf
3b4OhXcoGqX6a1MXRgKdEGP6P9ooWT8HfVtq5Rk8NAQJklmm5ZxrWrIS+tT0e+3m
MOESpQ2YiwEAq5kJpdElRMtTsjsVZ39Dmx/NZ5WI6lyhC/yvgPyqd37G2TWzpuyW
7jdBEHD6CmKGrNxqZfOpfH3ruxK8+83hsaOfngyxj/8rPS9Q3BdKLT1lwKh5dHnm
b3vBi4iKY/4qzMFAE+W2FDYtirMFxo8u0SdWTdNPq6OYolHDQUmixkqmsEq7M9D1
1FWpDXwhRfUXYIuXEEma4kIN6a2XTIQAGLC1VXKNxR2QtCAMBkpp/KuIrHMxH7YP
/TRZ52hFV8YrnUfHY8/CFwJFwTxHlF3vnLA9v+gsbyvMr9HxrpvTKzJJ4oe2xDU3
TM1zw62Keo3qENVwc1zd2FZYDN3MgU0RE42l49HdRWccXEbZwJBeKR4s3EsLVSOi
Mm9UdxLBv/o3dNuWYKi6OcZa+gP1NPCnA+zEzD4rES/lk7G1k2aoxTHwZ1rzTCRF
hvYLFkWfvBtL8rXAmUN4hZKRHBAfOAwcS2+J8cgWHg1Nr2/ZW9dKxCTnPHQXLDCj
u8cFQ31VsOzaP6LoV4wDDT/AGJWU7xsjvQeGSk9NtlHBohiY7ev4uCHjkv7dRwTx
SkqenswVbGG+ownTyxWmG3HCdF1tV9ITmnHHP9CRtyuLaMEElXFhKsrp6JGzKMRf
kPMbmMI7bYTy0R28FUPu4TP6dWgGVoG+/ZtlW6B4shb4/yUqvV047f1YJ/7eJSzx
cN2BjbcWxsoaleiFVVA5QGA/9RPPGKSfMDZvuk5mvGAtNmBs1WV6hY1RorK8WWlt
9j9/7XgaUiNGUSDE1B8CsaTlTHu5tSNmbEDcUqhgT9NSK3myUj4/pUlWdjXN43tk
kWXRbq2tVb1AQtgS9AnbLylUbhMc1ZzeGoIhNAyUE5IFLj2++IK9VCZ8LlCA1+rE
nBhYqgJYo6nCqVONS2uFBEZrPjPwXhTWxugPk/0BQjypskcw17u0gnCMzHlrzKfR
tOfS6UMJSVDRCt1FB5MzGSZg5jZ6J+NdE2hrS8jDLZ7QlUH+XH+ruQZoBKA6hgw5
6GOhptWfSPF+qyDL9D/SD/LGiBAjKLvgQlv0u/loFIAfYI+X1aZlq6moEwzRc0OO
5QSG7IdAClBmV+QdMVF9NpCsl2T6l+/g5QbKe9SZoVTxnmmbR/Rh1aphVMk6O15h
jXSdG5GOxMVU8DJSSbOKl+BWHix4EvQ/7BEaNzpczL3JVLeC/IBxbYVHCbRvxidT
CN/8qC0dtEXbOZD0OtjiGC/Wv72Uzi1HPHhwmDZP1hoC8eFPN3ox6M0qaAI7fOak
MC0s1/X5kxFRHQcchi1H6MB0sTL7jupfe0EMSiJAJ5FpgKNM02ZwU8kX8pWLkW60
3wOhO/c7LU+HHDNM2x6Qofvbb5GUiKOsjqcWfmy3XqNN7aXDAw55mzBLlBKP9VbO
mvDUos5T9ySfUBHI+q5jDad8SRBvKV4HI62mWaUP9wc4NXPXlvvL1yxox1Kq56Yo
kLflpTmkblmNDlsJTIe3HzrSVcuLcdVdKkjpQ++t0zHeLn4+UjM9Xad9+tu3/lbp
MPmunb5I90Zzvk0ZaFYM/ID7qvfmmc/CB/nqj+yQdjfVcFGSelroq3fi/e4E6vdH
2njibbIyCva02oM9QKDDUBfdkR07+vP1CQXplUUaSCQaKZshOzlJzEOdi3aV/pRX
jijksYk/n1PZEoMSaSfxQJmHxZe3z511Z8xMmblu0SdtG+jtkHCmtE/XgS6oGBRa
ZPm9XjCptYRzmXFBOg53R4K+3VD5O77Gbq6x03SybtnfiWtjtEivA3so/SpHhNJY
TDCzMkEyaymPkIAUNKhuRrelFSQHt3YUvfKWBEiA/50QQuoUqrPLn7VmGGY+Dqvo
CbibvAOSt7Hu1vP/37wt6T7c0LuCnOtiarr7nRheQJmP+BMOka3EOBMPMNSNBPCn
si14dnOv99qgNewd5nTkl2AVQ8gCyr5WjdxZ6hVzpsH6Z5tpzxrXmh0RC40XSYJd
97sKoCi+dhbYoQXpO9PiREGuWqXfEnb+5fcNs0Io92FX0V6nPOYyoGQN+fIOdw2K
heyQ8NQFQtDLdxx8Lk8PBzw8eRq1QcIM5MTrL8AHRKxStwhfhEr7lmnFvpTm8on8
3b6oTtwbNW11KvXgU46DLj/R6/KXGItGxQcs9b/CCGbwHC+pPeo0SJ4dYbCioIFB
bL7TBr0OYfyDt/9vUsUGODH2TCA2SRGr9PFh3Jo65rsJvbktl2ZkjMPI1dv6EKvl
aIB46EVO8hi0if/f+dr2zlXzuZGPBm8VN0jwU+duHps9qr0Jt2v/PYJ+sx9pMBuz
28NxvhOv9LWmOmh1WbJdoicURW0ifkhjHsqDncB9qNi0nqOjUChymkYBc3AcSoVu
Jvtm2dPMQaFg+oTiMvErKGZ+fGOmcUzRszRu+NlSsOqpij4LAC+N23S+xNWp3NH2
f+QEY51xhhsnAAlp7Ov042V6Pmw9UnuX5syRu/vvLK86H9KZqvoZspl2ZZuS49wY
/g1wSLhp9ZrsE868hJqyRunvKHdAgWyPg7rEEWBiNYrPgAs57tmDSdDqWe7wK25b
PRDCRo4Loq3Q2FxdoUKtRTfbQ2iFLNRZYsnJ43eXU11lkhyNAXyBEtiWz5cmargo
ohQ84Fw5CIacFtCww0lXOwxjSdy7n1RGU2W6kh64FAUkYpAUXDLfKYbiFbD7IB2t
RXoMY8VaYDfgXRGZod9KeEjji8sTm1cmDPRPylKcNZu12m578uyYqUK5OQ8FLRb7
7AuYJyYeiWXvlHD7jlC9pi62acoh7WeWlZGwAaf1Ii1vQtIWrLOCwu5j+ejhd4/t
YT0xqaTARwx2rKl/gg2dNSofakTe4zhM4graJ1mpgwnmzPNLY/ZSUS/BnrXZDkv3
+bY8mlC0krioz/ZQhE3MkHfnIEbpR2zTMIixBWM65+bbCYtpxcAf0i8c75SEiO+6
F+lF7USB6Gd80qdrLXdhkaRt9KsK94IlpuCnm5rSL1x52WcAnshgdBfWbl0q0Rvf
r3MZBbCEiAEJlxRU+jtUp5Bcd8W/5bKcc4+s8a3axUOw6JrrzaWNHyuE/pWbdEKU
VI92LIPHoQUKu+gmS5zUnd24tn/yXRzmfnrD082oEEyrtbRP09zo6Xt5utvPtzO1
bsFxBZ0t8ElG9TxGUs88X3oNu+DoMpCIjt91BTjdquPH5yNGZGgS8zsQ75L3WnOj
ymq+mLsLAR1YTkN3syRsqVYaPb6TUG8GKZTneUfAmK3oH5wOMppNPjC0bbqHgFA9
Vb6rykVWvaLqXstCkFZRi4txvSxBo+5NiSZt9fDoqPAb9igFiuM0HJBD2RuMsfMB
vnjR/B68t9tbZww9yQHmRlJpSVzie3na+Oy47YwBv34/C7tiq8uSCrvMBcMDngq/
0wISMhkeX8/inT6khzF1mqj80rPJ3gf6uNUXDy9blokRYumfoOAXJi3teZc7UQe0
79zD78z5fzpBR+cCO/feRDtgOlvAs7R3suM+DfpNc2CaswKU+ovcmRTIlyaYgzX+
AGQ3DFH6TDy7D0xqrYbYOidH7PZmKm6/gZHha+nnjSxHDKBJvhmlgVim4NHnae71
jW8Vi9J6rTYmdabqd/6xr1qjsJVZfA7ed2HJaB5FkWhCRWx7In4WxbvY1vhmUQFQ
PAd9xf08vxZ5LAk3H/Lb6zUYNp/r70C1sZBxmE1D+NLig+Pv34/gN7G5KoYv+oWc
pkCDQLMXjZSgNuR/mzpSJW/4/F7cEoSLsekvF4cGi/CuPyRGEAX7LmFMm6AO3ClC
pvShuWW2MJR4Ri/5FNJsooY7wLg4APFIBtZ89bQnFH3JN6TI8sdfLNJl8jCC0ybo
3MCfR0tiCSwSRKXWkL+/mZvce6tVYpPkvob22InzKWNCMEBOF0cn7Zuv7+HK6zVJ
TFVLjtuO9Fw2S8GbcSpft8IX9tthMrSZ2xpWNL9fbO+r6sMhwYajylhwwLqfMHB+
ASzNwmdtc4OupZyHcQbNsBTMRqz3/VkAgzF67RxGrbigpcEk0vBILS4IZSn2Dil7
uBDQkWgeA/Dldh33+PW23gOpTr+fYSfqFjTDGFP+gg/g/p294jT1JgjbaZ8sYXNX
jis5g9eRV0Ub0O0CeUkOIcYS5ADSKlkkVmWGK5u28TOOp1zkz7hOdZsw25PfcDPS
G5ery6LK5QWHHO9c8PEr/V5q90i0TspGtfOwG9Z5xpnqVTfKLQ/m3/9TFGjiUjwi
dXquFjGOj2YHGKp50InVwX2W6gw7c/HwOf/s0dT3yjBRugHBBMhr/UiEKnR/RO8o
yTKqMf8TMPirWtX89qHf4Jn+bGbkDcpFjeKCXJ2yBwckFcik0a8A06gLFsRCWyyv
wDKoZOpqcvGkfu5ZihAD+SFqKEfYlM4KfkrIHYUytsMaJYTQ00iKqegtrDWHXlhq
y9YDfEaYAYERARebepEYP6jyrQAabRAw1cTsN+hC/0NXdgDh7OM1S1k8OjFG7xrP
fbQGgfWbcF8mePPwf0mAxXE5UJKxDghGo1WhegtYol7DzvFMvAPs9n7gTdl5bfOY
Ut2uoLEH7m/NL9oF3WNGAlsG7ubEJwES8XXHhiZfaevDBM8scfOI1hxgYM69WZ87
k38qUfmsr+6qzYvtMcN3rK8DD0m7DpGgM4oxwo7aadbHNPLJObEZ1aM6OJqvldSH
tj+WfpE3RwaqqJ7TlKgFiWcVwLji7fR1FwCDAQO+pipqXnVABkreZphyv1jpf6Yv
wvZLFyPgP70owjGyeAgghrzsIz5ifU6x6gwrfiRq/iSwqwBclRKHhHzGEtYzbaTR
GO4DsB9MQcnrE6ve7ZYN6S8zE7RgLeeO7xikd7NlVcrxBr1pDTKTeu71T2YD2ucR
zgwAKBvqTobBsVhJQV+NtJz8KW7BmDAAqRSzgXb+Rokh1P7SwOSsxWbSV1cQ5z5X
C5Pfo9MlYG1i4Jc84q82DjiwfJDITbjxNlygEhXVpwwl+s0X5F4SPTMIthbOmfXJ
Z68S+vhVX1hrC7g3BEg+LEwA8ZFtP6UKi0QiflDbIGqqNGj6g/yKhNeq8bAGgIvU
9rSPihDkB6fDqNyyTEsZW/oNPYv3XwiSv7qcAMGEeffMXYeH/Xqj4O2MrOL8DMtm
Nw6JER8P7tZVkg38syveiGf9TS9a6co0t3q2+Ne6aA9gEWQgkuN8SS1D5a3yQFOI
rRPC1MNJUbdVx0cQlxpy3yCLVtzuydnfPDHErKKlx/MQjJ5QRuu2WVHBzTob3El4
0ou0V7XmOHQ36AT+SGHRu6vxPMNIZ5+/jSPHLnhuQPC0TkgMM7GAKIyJpre8YKJH
gamYF0677Wt1I9jnuE0DNIjSS7opzWFf6ar7cGONOLmR+ikEopqxdNvojVKbJVsP
2jtpXeiZs3Iz653dt5bkxLqra2wWKByN0lqYAwIpQOUq6C9cJhZzY49kS65aPgzv
52MHQc4kZ4zc+AR6ouTgxSGg3sgWiNGoYxgMNR4N38p03QKquzBHhXRX0/kMc6oe
Nqr8Jje+y4TZ4yrxA8LEo0ub2QLlZ0OKVEi8VQmNqL2nmZPp8LRP1FioOlr/w0In
wmJ4jSpKmNJR/OYpQxHADOOiL6n35kwD5R8jBIE/uwXh3KfkK8YZ6b7pUuzudwLD
O1wY2Wv4+sWXD2tzePbdcpjSajsotn2JwySx4JBZiJtlH7dOeVDoXCU6Cp/AaeG6
f+bqQaGU5RlxHhOuYSNyuoBmkB9G3RzjEWd86S7RbV/2qonTt3iULihHG+IdNUTI
Zo6J7co1jlnBFV7EZnhROElW4ah1bp+OBnV394/9cunKXcZ+9DwU8Gnwzlvd3lbZ
ARVPQX7dE9NMWl1MLRj1QcL+4uAdz+jWEnBYGj+HvWt59dSpibJ6FfKU8V7P0dGQ
iNRO4ZPgTvS/QvKVQ7aNhbdWoR9syp5NxOuYWSw7IPEpsfWJqV+06jjccFOzl7wP
EquxjxTZpTXGRqx1F7WHPNd8GqBBZ+YMphw+n5rcs0nkfsMSXdgg0XviPfUVxuj9
lNYyYNtW6RZuQ40DY7E2jueZQdMibSTlmU4IV8G8UR8vU1MmZyID+1reSf6+zvvh
Wsmyqt6LHO6cdWccouy1s26GBrVCy3/4UU+HNet26iMmUZW6L5OGeOenED6hd3ww
pbzEql1GRyGWtyBTouchlaoQbaAWOdmGn1Gdh6P8FfjSnv5ldqllHFEwjhv/1Krk
cEmx0WyP1X0e7hBKWFUKN3R9Xf8uM9ETKLuFxQdmUqlbGM13BH0FlUWU79oOLD9b
YGZ2PRknQ0lZVTt3wh8FFWcq2kKixhusA+2xKKAXhPnf+y7wzwp4eheBGqg7pZ1I
s8BKZ5lVujg/Ehv7Fz/jpa2J4z7z3Bor8QTj9JsYiot3om6cU8SrQ3y/5RJpZAVz
towOY8fZ9k+NPDBbiUQqCOcDgOQH9m2sKxQFhrSm9Np7kEB8CEQP8YY5Egj8LroW
AyBDjj0u29PGvqfjs6/dvDuReAV2vDIAIJvXCmp9IT9c9RjNRiAUePSW3zhM+/13
0hGugb8D6DBXbYBThWIqeG5neNZuiitqdPCZv7U6BHWEZZoisB7bZFcWVuTDIe2M
nYLM1BXTTIbX6Rf/2ikB1rhktNeAcNf7zTHZlXXXebRnrOOa/0ZIqq4zpC5/d3gv
OTzvtW32kLtUl6hDZVq8JHbh9R0jhk1zUQwvv4k5BinSbwMjjr2ciJFiiUOG/QpX
0Sr7H6UgflcOP3AMcqSVUNyGgjygeHfHHzGg4w4YYdUzjmTvkzXtvJ29HR28qvNm
JlZ7SHkG53DOpK0GpwHFZFLt8xZaXMAsdf9KIn9Y57xVjYSd96sYILdWYpEiBFwl
7OQCfcTNoMKeRh895xv9mu3AgKZJ6rHCP3NCajyFEb/AtZrK3+xErjAk7xy909mK
PUNl4Y1vX3DP2aKQTk6up96jP4TKuBI/rE29mmc2Y0a+eahofb3DDP2fTmXWfpn7
BxKTOLM03fiWZeshk4sQc1ZvlLcLvDxW1lJyWT4euGWswfI9z9gqa1DxUZwWiD9x
/Sgsun1OJ8MsoRCq8tiXgUhgpA3u4yKBgMPJ8/cNUnzo+CDhjF0t9FNIbcB3q3ZS
lQXxpwsuoJNmvCZQ3xBqoQzS5Bb5+1wGTYxwCwVVxCIq6qHoO+q+0JwuzYP0VFK+
ecXYVweexom3hjEAjV7q1Z4hyfXil7YoVk3JdGjozqJt0ZQVj/5p/eZnFWqma84j
tCYZbtk7Ij9f7XThBbYVf6QZ0LpnR3RjVTdKa+SdmvM7EhyD6uWGTe4SmIcSpWJc
+D7wpqAU7DkWC5LZ1QbCxarP9oW6QcfDW1YkSk1Pe9bSrB1N3Vq3ZdrW5A+BFM0I
DGUmHTRP9X2kL2r85d3u/5J2dnsGRzpLRc6lSlT2SHF93oE6W5q1m4Lj9eOxw/Y7
qrBQp2ktQb+XY6sACzTTpviyHoRBQ6HvTTOXVzGZM6u1La5+hnUlh3VK6rsXV+7A
W+YvL1kdwVI/tXK/tPtCMFdvR+UqC+pZO+2phV0y06i8Obtw76Oxn2qsrdlu3aQj
oV70uSjMeMQK2qbQP27XvjVjBi/9Kd06iM8lZz/QTn3Zmr+hJSH48hih9sEsa9il
uFY0t+lVCJDE7lppdKRXYr766g8svdFrIF5wHpFrrmr2LLxqeMfJzhMmlSfLwgMW
Y6MYNoKoMW3KJ92Cwbmzebo7SWKIx7N/R14f2Ynv/w8aRcCo5y1djQsjcfrJkYCm
ZRNQtaixsTPVsPAVGe9b6ogjF68UwLNv+PrX9Xby/DfYIwPM7tw1NhoGpv/l8h0J
Ic9CUdHf7PEOWowiZFxxcabOBzOy36OVWbWXjLr/q7JPTibupk2zozqRs0C2lzov
vNVcqq2rN45D4OLPRFv+2ld06+qIj5oWUKp5E/5zMhn2WOOPNUYruXMDEz76e7Ee
68Y7berUxCAJTwWITmXxYfqMAw+T2lTFdN1/78IRXMILl2SXXgOLbV+p0G6Qg8JZ
by3eYscidnFJYRNWgBQhZkdvw1QCq5D9vhAwWNVOOUTH65+WXUJ7fsE+pzLaCfAM
anQVMgrRKfmlrzcHdNTuS0k99z+xvBR13dEVn+Kxmdd8Sr7MLmLOnQqWRMNwX4FS
68gP8d6KFOpURYHmL3P53jjZT/uObIHO1SRJ9o8jTgTubUNArOm26HrAttpz6Xkt
pm+/oLfjMwq+OLRC1rsit/Ak448z3WkMEmemLqZou9o5rYDztCOAXyDc9nxC7Ynl
xUGabu+5q9mzZemx9ySP0x5ZLas1+1pko+3A6xWdzsxgkYuUw7A0ZpYzIOOf5wnp
+b5M05YoTyECFvJxhOm/R+VCyqWASEMEssHseB+Kf1qQXWosdEdFGqRyldC+mtGM
/OryMwGDM3sWFcE+7i3NKhlSr01TSZbNc6cHZvheeytAjhjqGuKWQflc6jf20hrc
SzWDZYxcRigeaqp23B9BhO3Bd1BjllWiPUBytaaR5as9fBAsffBWOaijkesl/Muc
SXN1NLjRGnRDzHoeoMO0y8YC2QiRL89PBKv71mKyagdqc+hfT5h1oyy4swBS6k3m
enLtrOzyx568QV2Os4FOo7OvszlKrk/w37L1XIeZnYZ/l6PWXiAi/JRqUf1kZnl2
7HR9eM/42XcivPgye/7ouEuqxlf6q4AAGo+xUD5coj3U450LwDi7sdfi4QNpSbJr
JEoGkpFWbnR6wuDINY2loyb8Nx1erN9s9uXyLJDXdZcr0jyR9KxEfxpmWC5MuKQt
C7CcushPeGKRnwMOXgey3n4nwWJiL7fgZiu0Jr3oNKz6rc0mcYsW9tmzb3uAkSU/
jXjgD/fzyHfFNrw3Zdq3XwoWmefIJD85GWW+4DKlNMY+e59IJ0cUPniuIcE2av52
VI8U3YHGhEI1X/SvKWssjyIkpnZ5ApJXFj3kHhqqj/DIg+9wPSK4PCTNzd2vh2ZQ
yiLEIw1+r3Wbc9VJtiH/Sl2itgmZzQ2YelcX+dvcE2t0e1F9YVEImLa1A4uvTL2a
Buobls0jFNEMGY2JChVJ8z8e8SQewBPLEDSwLNdOqrhzC+oyMrsUAyu7hBF/0fix
JehnORO1UvUM3pKkt/V44E6qJM2HvGjXzokicAnkTgi+3ncCKXxh+f99pTPJgjDO
MZDNBzTMSNAmq8M9zWlUMW7u51DS5BQ8THT2cTk0/jDBRVumM3afb2ugJsb9H7FG
1n9rqRjtWE7x1ZcAms40UOTG+fCykN28eafeoi1+hCtFQdLTbQ623EP4qzLQi4xy
dHOpGukiG/NlfTjHm7AND9ygnj9nQ/+hGK2NPYUA/tvAsg2un+KLDPjnq6Egcce/
ocspD+wcx6w0vpvwxLyBbyiqkz7Q46LUuD2xdwwkQwRxmpHfg5OrEzoCjM7EGVkU
eByA3/UlzH48dNRCrdQvtObjCfpaAP4PXJMpsSM29GwboGk7cbpUEZ9t9nHGYqEN
xI3DxdSGILOCVoEtgUgdts0sAgV8G3yCxxmdeqn/jwURD++NaS9+HdO57JEOBPHS
EJecXxJZK3ZaCtDUxuAYXZPYBGBuz2DPUME25f1rkxgrL/T1TK9MLVHfr371lbZ0
Cn4feNSvhQX2oXVcCdJ+BEtz3xdJGXqQ1UU6XVIgwVlkNx2KfwqTul1GgUk+S/ag
3JFgOSPXJ5o0yAnRNNalVGpybji7O3KxcNG/IPPhQXobV2wLyRk0AniPKrNy4Qh5
60C3CarUQXZ/uaZwceshiVnKpQUzGxOAn0dTt/GfuqcVvncMzT0R8raHD7WCsmxS
Ok5y/Ck/5UuMEhyn4ePLOV+ntkmqhCwXh0nPaMsrPWYowLayBvMXfeEVH4XxPx8T
FTKzfj+/BoMVk88+64jiXRTOfy4WRGRH3dWmxy1/dbkz/6V5MjfJSKn8tyDqOp9w
PkvGBYvb8aTdu0P184DQgfiaMdlGzfi5ttPpw5IiiJtcbK/IReIIaUdSM3skTk9o
jXEH3F5LtW+7qXHYn/tQmHPVC79pnpgrXUEhI/RAm1DgwuiK7/3E+20BRjD1AbUq
ZCaAtozcZZ4YBzKKV+SeAc1BptBhah9VJm00soNsjHbgZtxb2i9D/1Jw+49TX4iv
K58Kgy9KNRC7FfJzo6BVPvBxsRh5MJw+g2TLrW+C9mpf/pN+S8JM+AjoQX4O4Vwt
04Vg4yxlOYe93GvQrCqthNtosOlldVbSJwRQErHvYCyflOA2eHqH4WAQ5i9VPmAm
kSyJRPRnveP4EunOfV0ns+LVPtoZ8BVgQGFg7N2q5PjKJWgIPK/R4X6um5HSHXJN
7wth+vQNQ0DHWlyzhhUR5Axb2lvSPzC3g2cJG0V3y1l+89sW0FCweWGDzwT5R0b+
mQU8A6x388DQsGIHNzgT6wBooAgpHFTkgEDMkVGwvGCk7EyPnDF0Im0OoT6BgHIq
BXzv3VwmbuK8/0DQTy9n1lhEQixOnxsILotb9VNrZgJkfeTeHkpCLGcuazDu3Wq/
0saUFLFniQPQCzi8fnqouM/neQxPI44VNZtCni9i3YHdLZ/JnjPRZPyjDPqH/4z+
V7ynAAG0Pk2i4Vd0UheE6u/67Ui68iP6mJj9H1kfsP3UR7aK4VNvfYFjPgL+YOQP
27H0BoM0yo/oieuqNQPP6gyS8y75U9LyXu/YYDd+0MDAehtnU/MnqSsJH5ei000U
He2FpCJUFGCs7aRwHpqREj3B6qkl6LkFUFm052nBQ6DMPrjhn+m3tIG9m4rCNm90
6amn5C2RIuQfiwJqmRLvXiDo06zZ8GFhbBM/FAT3URfmCOC+eOjWKX/zj5b9Ui5Z
MBSRCBsefdPozoX5qo2zPmWNyVDOtwfuu2yuS+khvzlqZ8mvUnLfYamFhzeNa0OM
mHd6HeoiN1LzUvyIKDcVTakyS392tLvY02VYONxQy/XlX/lGAU5e+DAkO9etLFmN
boOTFzSlHbcMvd4s4C+3tjQnCJ5sSNC4UVQ9DJToT9zf3Xqbvvbc5gxc4dmtnsS+
eMEqlIXffNFH19PU1YJiHHiPyAmg3NTj+eQIpXn9xELCn5GZY9RJllpjoZgGgz44
APsi5gcsOXrBJD0w60J0kfhhgsjKR+6YA+CekZGZai2PYbeJNRWdsfy0zRX9jGIJ
H9M6MIGCYl7chHX/23xKrVPDbXO1jYZ8dLbhvw8UFFPvsgSyw48JlBtA16+tq2Kt
gG6L5NAcSFVEQtjugtDH9Vjq1TQbPVTKwbdLJcYw47QPD8I+eJnA2s9c/8AM+xBY
ztMj1v5tA37qb6rdkQSq5ua0nSN14PJF88/fqT2G7Pwzyvbif1X7y6IVQn3l4qxH
VXmUj/SZQvUglwEO9p/kMvOeuI28aiNt6RdDTRKsgXTw9O1t/KnAWD3p6CpXqUXN
WW02ub0T5fuRiPGAAAAP0tBy85zQ1vT9ShMBZccm8axvjUgNyto+Cop/VSPgoXPP
6786dKrd9sffCYNovkZFxlxZuXJ9gxGRn9NuFOGQ7nVykBjB2RXjw+BiZOf7b6bs
rrRI+hRlMndemseHradSKyilyHld6LAxelBXlwKi4B3ANNLRM+RHh4BRDs0wJGE9
lQ8WMO1zV3wh7/II6cOPpOzQhwVX38rIoh4b6GVVE6fZUG8shhYdktWOaoHSia8P
kvrt7MRck5XgWK+VxRiiCMPrUAaBkqOlysXGT6Zh20I994HlA+wAG7HU7b7e1daH
U+XFR8gEk1x4k1URmvgVfdo2ZRJUvEmnlL7DcCcHzTkklTL4ltbCaV46jLk5BB0G
bSYXs8/HSpZjixuliaMTmcG6WCzgDJoP5jMrc6VA+99W3Yk1Dch6jhFdPN2QjKLU
f9Ru1n/VBvT7WwLkIXS4hVmmQaY/b+BV+U9kpc9kG3WUnCeFxBtka3UV/ZSTa9a/
b8QCxqDIhlhtxxE79MgiaT7FfB37kiGO9ZKYOHry9CcnMhmRQEzW+YxsX0s+TDQu
7eKXnjDu7tvltgwF1Oppx95HZefHqaEXziJId3zbWnGJ66dzj9jc3kANc1Y5inD2
uZLVItiTzgFSVBscyl0qH5KrKuO9F+txGz1li7WHpArIOktf4mK9m4TEYTk8nUac
1A2lWty/GjkdFT0Rc00/5//ID2g40dEjMcx2cz7p823fznhvW82zqMI06eWa+D2t
nmzLRs2kFWqbNyhIgpPA5FfOwcTqQo80OKhTnBS3/EmYSBoolvyNxsTjHgkQlLJm
Gkfyae3UXq9LeuqGdO0qoEcUFji3bHH9Jz6IyjE3ZOHPjZdBgdbJ/KVuprbfwhET
UGlqP5sjtqSxDA7UlOJoKhJgv6nujiGLCaaxAWwmgOrK7Q+I/0jWCbLZezoKDwLl
LpcvLa93/LvE8QWDApiWY9+yzKogc/w2jXl637RL/uN4zYt9iNP6vq1V4jHwKQ+R
8X7y2dP3BnWXd1/QhkFiEZjOH8SBxxjC5zLQRmeeTB6ZPll7GrSvHa7BJCauNgI0
5/mb1GldMbdYElC5qsYbbkWCibU33ofjMLXxiPH+OY6adBYY5xgSUjvh2zhrexg/
/51aqFj5Jqc/cDZr16rq20xZBqyBYNqDWkTgk8Zp2WqyQrU+2dOPwnQFUsmH7RWm
3Dd7NM9VESWYa/YaxbYcf2OAhnZbYyk1CZFKlfTQ+iuDOw+y0FFKP97HfwGaqanV
mxRwar9nBkpVs5Cin8oOiBl1b5Wo+vZzHKRI+I8Gvhs0bH5uLS0ZpUg+5XbaZNqP
hsK1MqGt1brQSUwF0FrNdMbYqpyKvwac9avKvn9RP/JcMh1LKzMaN1wXXKCj18+P
LUskODdoEKsyXOo/vw1hWYEHt0Hm5TLWueOmSob48rlRjkiwqigPfMaW7L2en0TR
6BGO02GPX6avHy+5lvv2seuJeZZZbrRzGc3UYX71j4hv/J3V0XvxCw2ulx8/gkEp
vGbW4Tgn6Z0Z0+mNbnf+VGeV6uPyh+dCTNDjyje/yQYe0euxdGypCXkN6dKGIxUZ
Kw7i8jK5TI+42ydxmizhfHFKAVjkpgBYuNZgIdB1XglB+h4NMP08/Q2yOaX6er43
xPk/zeYu+Drf5iuKo7TUcCJGndDGWzb7anzCRqnhs7F9CVHJ2hBKQE80w1QGl/5+
b/WeuNevfjRPsZUXpsJ9q+ENVM9lllvb0F9kQbFUBJvPAeXEX18j0eAS/OTcAOVo
FdWK+Gww1twd9/TOfDKhnzrIAMx3uNDcVnB8Qx/wMFaHtBsoVLbr0ADagyf7S+X4
ONOxdnoaE9xTsqH+lUAUJDD//87zOhWwgxrBJZanhODVN7nFllnOkLu4QCltNo1C
Jw4cOqD2NiltFU1AV7yTAATj3LWM2iaBLmlzBqmFyODBCkR3ANpVuct1CrLh578c
wNJh63SmLU1C3EtKvH9e8D9FBdoyOVspGxTLa7HqViXDSPsBGiHv15237hKq4KpP
dZ65noixGVTnh2Tm+ZyasBRCSVmPjsgWp4j28xiFj/fYUYk2HOQ2jqoKlMqQNFlR
8KYN7/48wMbZEx2JAATaeSJZGZI2riOArbiRqg5OEfKxPjMU5g8/2dNUyjVRJkD1
b5uS6UqkBOGQLetqzXhGKgZnTwLi/S8STyESSzjg6IAfeVllDXKrtmXxXcUw9EsS
b1rIm+SZIpYPqx2qAIoQAwSjMzUDbu+GWWFf1LvnN/TaQRDzXwvpFRTHfFW1B8BG
/NST8lxqC5GaKY2r2IxL2XlP4LybndBO1fXAZG3+yFr/5derDb+1wEMC+L4h8InC
qbiJA+xnU5myYQIEyWOFZWrnpZy244W+iKtaExCGDSmq/+u6zZpAuUmh2uy7ZbxD
dIPfElJ0FU1VBL9jt617T/jG0mI5tjLlLMVyKeKjL7CQLDmPeXUhmue+Ul4uMWoa
U9j9j154JDc5lIzifTAKkS3yXF0m1dlPBmpZMIpyqJIZkh3aBsPtupMwGOuXiceV
tHv+Urgbf2+jBsfuVDokmLoU8UCW3GB5RY+UA/SQD4pWk2W43goL+lfJ2hsbyRLO
WBip0RSSqeBayW1zdJaWevIeRVkWNqYlsypnjSHwaxu023A1E11zWyWXLD0DGGX2
fyt+kiZB05LHI7+WvTY/+B6pcq4dGi7arcds/ke+kv36ZFtc2mlmdTQ+Ghfe2ejD
MTIGYOwgU3PZThy8bAkaEK8qKpyJvPso+O8BRfEqDdddKzLg/7ptS8naKtEAS023
3q2aaAKqx4djz3bxxDAaKpJm+sG8yfqHiB/43pAC2yYLwVXsnq53LyLY9eC36fWx
jQuGnbLBg4XKBbcLmf57++7z12HBwuLOesxUze5PDOuZycxhuNBB129YHQiTd1z1
oLRdYBNwUzEVNnnr5UNWGIzcyqXiFgt9w6AR24/+AC43okc5NQTk2yaCTXZsnRSq
59Z3N9mbtUlEsiy8XWql6tAlmp+zuHCHWqXB5tD0JoFmoK3W6KVlAMcYTYX/ZOeg
Jh7vUJTuedyfwb5mrwXEJWAX+oxLEyBk2qQKRufzaYiB6SUXxeLq4RPCOpmysjCh
k0qFxwVD2t4i6MxJzIkT6n+qER5mhBhQSCoSImQTfRxDzL5l4vD+hzAqLa3iqsGx
il5FQ0uTb4Y+I1Zy1Y+J6KJm5RQk43a36O8HtsRPHVmpJjUoGyaM+90eHxY7xAZ/
vPv5PFTSdAHueFHDJ3lCLYoS8K/0bYLYlG7ouP+NHqYv38wQb+ZTJX/WDqJzRmQb
CEIagc2NF7GWqdjlM/tvk3OnR9WH2eeaGzpcNBPHWZvw3KVxK928Q8zhYu6oP45W
8OZ0y3+FCNhFfgX91zoRXSfgXgYiQFWQWPhkcXtODcpZGuXlQsEnNtNxlmBZjdSX
E1dV0R8AWuQBMvhqXoXaf4vvqCDCZZQUIklFL9oooYCllXBHRdM0H1FY1l1TnB4H
HmxOCFkQgVQbZHegLBL7nohZ9nBtNW0Ka4OQODGRFExlJCsPZV7abGkrukYma0Mh
Nfpm1pj3y523AcnxRFzl5TycXLwMdFmpOUmQba4OlixD+epmBpVqkZl4MOvGLf9c
sZikfvlB/f/qNZfTs9Vo6pHbEvgbwosz8THMn98dxFsLtZCI9KZ8ktgVF4GO7i4/
T93ZIIZLKDJ+I/yrbBFoZB8rpu8g8ZJT7x/fgkw2IZq+Vm2RTjshs/R8UbOwLQD/
CW9tQ6SekI6IGqAZjdZCw7w5n7tBLo+R/AbVkfGWt8Xq7xNgVLGDwhIQIEVx9LCZ
7V51NmGloq3SKTdLmvnXQtDT4SzgN2BrZkD7sIfGiYyt5//3S4kCJDjWXMp36CLD
fS9gN8ws7FbSKCjgbXa/0btJfLYFcPFgCnhRKiX5V3yyNpMDwkN/pLpN9kAxN54n
bcyqpzegzZn/Xjl2vrJDxDoPijFq4euLgkDertWGbEdqTdQKYG438oCER4DOLlcc
RggfjjAr50xJvlvDGh/et8+ZQMRsPtHvmFmSWdpQgyw+17Inrk5dbHfk2wQQXgb1
lChDPWHI87OF7g1xf5qTZTTlHtZC6nn2JK78z1hZteYrul8vwMLPvhDYgBNkuST4
Lg96f3nbjxM8eUwXxrwxVODRNOPnAoPJw6+UzRiMzxHlQmg6DbDMYSnmV1q1wgsF
c5eQF1md+EHfteeuMiuuHLVRbrJ4+267A+1AxIvW+tRvc9svO15sSlZQGW4je/YK
8H3jmHwoFa+7pG+zjgySgEOBJfryYRSC6Dm7TmqWwJV1Ng9G9a1p/yHLtm1tRBze
XmhBmwP0llqsE1EyTIBKpNaTzAy0YzpXtIj1eI5keVrIKzq5262oYiGk2tZsjQCE
6xnlktjnWF9to7ni2XP+/a7X/aDrmHOqLMPlNZ7OpNC7/pIpYE7FymkdCBG4oBAk
aVDTdppxQRZKbswo3UMJXz3QvEi5BAhl34xe5c+t2ICtWfijpKmi6NKcUbaMZHYI
sSriRDXU6iwZw3O66O4A9Jvr+NtabV9McmLCDIx0XHu7pMqA1a1v+7fis8rwu5yl
hn86UO9FBMZJh1eTIYtC2iIs6b8lUpJBTXnzRl2gpJJS9MyzmC9kiE2SQaPHDELn
c8aVLwm8ZjVSJMjeNSSx0/YE0yWSvRz8ZcvfNjgx34+pUO1/y26YQdi1F1QDh9ss
Muj6Vs4UKuCJTKBMN3dYaN1PF1GRq2Ta1QOPq+b+zVMq0AnqFskDwDv8Vv+0iZ4j
Khl9HpAG0yWllfJsGL9n+TJey7sbY9/h2pD4LimoapeNrT6DRIL7l16ZFzYmjMdj
FCMreldXmtyPUfqi60aBIborMuZADJoTutJXEzHzumcqRwzrzyfdeN0K+UKnuW3l
PYQC2qThT03Ht9wfOfCiB5xN4LiQ+MnfHTPR62gBERLASXzDAX1ATWwQNHgpAG65
na3lUBARWJiVdIcM7AvRixnRilwV/gMjOJmoZzNubqIbCI1UNEK3JVHcn7Fpn2eV
GGNqoQA1hjWZfkiNSvUuW1Gj58w9v03j1+mcdgWT3TEEchM420W59ef+NsQxi4fL
DI4I2WYfX6zgZW3zIxRetqtYF8xZK8Y78OsQU0EjpGGEMNAOw4128yVH/0uwp393
YFECTbOQ5I0pwhr6hXaOr+9WUxmdleHRw02bd5BgjHIwbMdmMS53inMPG8lpsaX5
FsxbMXJU1nQ8gVEjzbvI9qEr7jWMw0e9g1kfZ5ZiKFocqjN8FLsUmfa8fBrfN48T
YCQl2W8EnjFwtFegyo+XWoV9U/tMPvy8rPbQmR46HhMYLwwZBO29Vh0wQRg0USBk
F3fQJ4APQRxXdb78Wq3o9ef7MI/HtYBCtJU4wNzjlSTqnfbe71CJntHpumwDIiIW
BGnWZvbWQ3tqVWbBVbhfGeggfee0Tp9HtjGYFfr5hG4aMKLh7Ixe/3EAQNDESvFw
BjLxrxSbE0voz/6Y3aOLPDdVzd3yivQmNIA3zL9xoAkiAvft1L29H9l+5HaiCjgn
HBjtBPAMM/sRE9bMbzo9CZxmtzNq4RC6F2RHJZTQMeNFuyD7x17CKF6YoacPnpXO
5Y2QYT0ye9Cy2o0of0NHFGYdPS/uNEVqnIpnNES7ObfRUIsKdr2fb2TohfoA/I9u
GTFNSh3+zhZ9H/pjwzbEV9hPafeMudlSOSMDUhhxqTpkjXKAHzTEfThkqj4wg9lo
VQpDgxV+xHti1F24D96725yAJUdhxGb5jTN4FWWoI+pxVuq5aUcSQzdba1OaC1X5
acgF6kMp67Ulm3zsP3kx2j6208xZSvvk1p/SOj+52DUW+ZoLibB9EKEU2zZkXrum
V+YYjjmJaQGRWibm75v1NRfSZrPeg+a08vzXsPq53/OHRn8ce6gWN2WSfE2mb7PW
AGoC7hLflXMXV45P4DWzFNgnRiIMb6oGQeA3KN3azZWXS2lE9lPOcD9fsRHQjOFq
x4K+PMJZWU/0gmnPRQ5Un5BoGkpV4+2Db1X8jA3UU+a5hshyIhMdMI7C6aAt5Ig4
qt3h3rInGIaMcU+dcKMk/pxh8JnElrh8kdKykowPyPInZFJdneWo7K07Ol0uRXe6
2g6lZRHO55tJan1svA7NEXn1GWpaAYEKTHUfHaItjUtzCpWlPj1lWbWLXKjcbeUC
Bd5bVlOwA4/djDC/J+nTHYmEMLtS2iH9O0JqlbFhg29u5HdudgA9zl9yj6fth7zv
rNlmM+k59MeQjqC2V8u971s3aexsqUOdzV1gxzy6TwaczXh8VpjhGjYxuqTaj+1f
qPogMVlsrOxggfeUP5Iaw1bvOZu3a5Xx8wALFiTme0lMQ8T5CsnhftD27PVeMWtx
FqwYkl99EAXzR90G/r7RMNJmohth5bOtXQDAf8ajqqsB1MpI3gRbM/E7YS7rQbDh
rcDrwdF7oBHpLZ/HYvTFOG7P4/bhndYw40o4Dt0wVv9xWOigQ/5r9O6P661LM6zL
Gd5D3znjnR+cbb45Y5IJB8MobeasUArf7snn2je0nkzvy7Qm8QsxpIoKgNBmumFR
AH8ONsomNOSEQiwInqIEYqvPXZPOwS99bzkxwwbWnOzHK4OZsSb5FEyKuB2I2Rcm
/Q7EdovsQMFQHkz4ewWNajHwM2NmUv/WTXn8I0E59vbz4QLC258UOdpc6AA6UXLb
x4lxQmde711R5cgc3Bv+/PGY5lsIwyZcrWg8xyor/jBc30dnTqBNXfmuCCs6+/dX
LeprlAkHnWnrn0XK18fHqf9s2qnQ+7dPK2GChqUXxdiZYk0jezboO2BLp4APbS6O
lbyx092remjmQM76S+ZTsW1Xy1u4JkAAhDr8d1kM224Upogs7z5yiR9sqcDz2lPW
0XSQVDrosC9F7QeZBodVfEoKPf72AGOOX0gMpSXsGs80JRr08PX5Q5mn1ehUajs7
4NzF+s6SevCHXW5nxOcqjhjhnoC8vJjyzdPzLm3R6gC+1w4WJaXG33cQ7ddznnSg
rydr2HOIx2SQdkIP3g+ZxZmDIZUlelsHvkO3NYbLJKdwVD0m/86YuRERzwOacIgd
fasdA0oM14kdwQA9E/ovS1aUFTdHAjrTe09LRBABlkeLO00+b31+sMHU8v5CbNKl
TG3WkckNQGUmBM+QDNr3p8k60EOcr3oxHlfPK1PBYM70cw8TBtjalPDZ5RfU5rxF
4WtEIfxN16m2flYxb28KS/Kf0N67EAL3dUkOGJl+jgfHWHnHlbm51B6gyDlG1jVH
vFhWM4628QU19C5Y1pGcbLWvxaJN6GulKJnmMahRpRMymwororlKsJPPzr9J8T3H
uzEAY2QXUdY8mq92+TJp99PFNbJmPcz4cjAF79L7r1+MZNpCLanwE3ID0fyzlxK7
IN+ghz8jRSnguR8DumZlUXq8KaeYKF7iF7/k4umgruQoc+Chj8DKjec1DGAMmVo8
aO8Nu3jtFDrV/395pMyY7c9VdgI6n/RT3+ue4moGZEfWeRMha/0RCxcjgONIIwNK
RqxAp36eG+O1D1pHXuNyz+Ztaa/sip3WKAJEQQfxH6LoRnah7hW60FOSez4NVJ5n
d0kpSuUm57UiPRiBxDQqPvVUrV8YTbSm8coy36nmU0NE+6evdw2PvCH1zQe3Vlve
+Ykio4c31Y40f6Zc8ZL3Fh4OgXwDyNEUfLl9otVGFX9eq9eLCs/0Qz+WRIFakFUc
tNFTe6Z858Er7Izzeo7YIcbQUqWZM+N0GOSQiYnOkBDwVdL4HOeHdOF853M3WFL/
cbpqTMQIRSJsuk1FVim7NPAqRbTNwB+gOR5ia9siIbLY9+IzXfklhImfonVbWzTR
Fk9WX6CxG1mWpXcZ4wmRD285IU8uGku0qnJ6uonIpWjxomI2Bscj9jsS8dC776Ss
k/ksxnlf5fvfZgbajoWWMITioZYBDSsHHXEmxpsr+dk4vFdrKP/E1PwdGVLEVN5m
qWN/PifeYZcq4BD7VXC00LVbc656JLA2ir+5e1h7AXWuQIX37yUbeH7TeNO2GGhS
sxJiQk8SRVhHyvJY0jZgunJ3AkUpPkvFnwRa+ZwXx2bamtI8epfYrmIkf5sw7AzX
MFkBq+keYQncNV4sD7uSbXjSFatMGvCC69fQ3AzYAQUbshvpegMq+sL0zelYS65a
/EQTNZ/ImhTr+7gPC7ElkqxTueKrjOV1HXCdoU/lbJniUXgyg02RKZ3UBW5IiGNS
q/EqNuJyKkBMN2vD9/tAL2eHIDrpjWzjUPfhk5l5RXJID+4KXPAo0bAhf8cQ2kfa
l9MJ8IjtVvsvX/sKsbJIhSqdEX5m9gHrDe5AKFpeYqDXJ3GtMaXKDFMTwuMK4v4q
xyEVWl8QLUY/BrR0p+HmPFT/yfZZIAVgh7AURe5wYsbMtxOExUtPQHqPRppfdPEq
1WrSc3+B/s6s2XtLQ4thGMQCqgrK0LlO6x9GT/FGAk8GJHas/tUAEddCzUgzUWNG
RkOYPhPO8JBxp03uKN2w5t3ZhYSjXWLp3Xxxsj4zwLfxRAKuZxmXprJZtKIlim2P
Irr7Lr32qREgObj3NP+xxgrzcgp8kwowsiEWZy3TYxZ3FGpB5p9ambFuPWFIG2Ef
k1JshjtP19EULSuzmp6QYpD9XB/BVcA1ufrccFb6k2hkeDr/DdR49AToKvEKh4sd
uV2m7K01Y/zEk/WTS3+DjrFgMbitl8CvZp9sc9QY2vaYmsbqJqf+Q9oyGRsIjgZY
2IzGcJRitzhfqJ3qpI7J3lwg5/fEFDBeD+8Rh8ecn0rYx1ErIJCJ9arKehCw6Qn5
NvwU2w5Q2VRagw1SX5HGvqJ5vS7DEm7Ny+gp4MBtN1bJ3GK2HX1osN5YHXNq3d2t
M9A0sUWZiPpNkTUUK1mECLzfNNsWy726L3WoBNkKHEEESveANEn4k+vP9qNkV9zg
kZ6mLpHhcOsN6pLsB4GUQfrLSEYAkYQkq+UHXF9iRtOmrfFyWOjLxykF50NotoaX
xXDLNEPB3ogwYkzKDkaP4zGb87fqZePIOVhtMUSN6Rrymj5H2NYggQ17ZZtV+UON
tUszbnSbkOlKHsK7xxytB8iJ0+QvXBjkfrp1CtwsU+4YxsYJJ6BwQ4WHtnB0Iufo
41p/APNDri2GiNO3mmcFlP2fhkMwK5JomMhhPtCKHoX4cXvxzJIHQ7/pNNIbmtKn
MzSwAPxfJLPjGr5/1NZIUos0jBCNiMNByi9fwK3wcWu04f0fU9Eic/ZuwEAoaGhM
K+z9dG5TmzlogsA3CW8JPvhrJOEsY7yGaEU3fRBGla4KveSuKHa08Hi/5qTk7NGA
mrp15U0yXooe5etsc1Iz+uffK7gdLl3wYuxvCl90oFQFTkkTzHXZwyUxKAF7TYVr
p+UMJU5NHDeEJ3M6dyjYF4snncgx0G72hhY/m1O/7nPmWX5Lv0SRiZUHkk30kNgW
QBQJIjkgSxvIz7xQZf1TQRaMKd/rVDQAfnYoCQ1giBYp8s6M9jMi7Bi3+Bq6pgjb
5pewTXtr6dbaiO8+biE7Amgxfr6Z8oIk9nNtppgUyxOqJgTLKb6HO675N7bsyxFM
5hhl+trMZTJGVJgWaCS+1LY84AWdmaVHw/Fjqj8wNAfkeZjeJw0vD3SRum1hGn/V
l47e9lM5PLx5C9xcPW8iczGM3LbK2IfVlQwfkupDFZttKPtaT7trN/6riJTc1Ed0
Vro9lilOlHR5KXA8ig7Al/Iq4J2hX+BHgR2SrfNkkKE2lyRenCIgX4vQgBCNTfxd
d9gBRnt4/CJxIU9OibC7+90v1SYIadQwG9/FvbgAckaAbm/xEAdGh+DI/8km6qXX
ojwIbyNsKVOEuUfbJ6dCOG8Imz1ccRCc22vAFIV9OpCBhCGt4g+6rav3sbJ2Dybk
n2AwxfFGarpUI3w4HItniurjQfpOMvk0+SggfK6hbFUhzNt6xHIVLfbrFTfGqe6Z
aW6B6y68M9VGpTKhMgNiV036oXWxEwMGXhwA97Xl3BA3CRVk9Z/JKMB4Bs1QPEbt
h7+ryDb4Vf+/lrpR73qgS1+Ua20KisYEv419DjpyWK5BYDRrvtnU0EnOltaY+E2+
jeNPIahbJJIxoU6PXMoORUJ6E/TBjeb+NxLFCcHEZS5p3RItALs5tR+LzH3mmA7z
hZG5VFuZK27BBQLsHB55EtyZsr/xyl52NS+riq88agWfapQx4EqqcP48wxo1FKJY
9OwPoQUGtTzaTrhDIZMMQEtaWSG01dXh7h1MDyKLkPXTeh5xq7jCD2pw3m3mNRWC
IOgW+sjaaTeVZvxtSKTbggf5RL2Zx5Ak2DPGAv3MSOsS1FJ7fF0jMnEij8P//+l2
uJztLNkc2se+PH5XmHKQmon3UZlpGYB5gfx8vUtvSLL3IymkY/XWKaTccRZhJbMP
sZW1vng69NOAqTiVphH7R8qCguQi/osNpxpkinFekZ7yCkSXKHsylkS+MLBVwn4J
YO9SWOvPmYKGA+2D1wfAx3pHMFrnkMICmPucNUfSOlsy3ihEFIkoBTb+yhXbGEzO
KFwu0he7X0R+n3T/YqQLQZQDFAqU6nb713UoOfP9ZZaUuveSJWVEZD5ja2wQ8zb3
Yca5f3uvZ+bqy+KQwLuHZyHxnCPppL9uuqxeWOPzpYIBvq+Qsk0Hnd9qJ4ODIXSc
dih1TLOH34v//s19H7b7E1hyQcIZuDIqZG+lMmB2tz6rD9LoYMvlD0CknGbkZtNW
p9kMo+A3jm92q61eS1cmR+Oau1aQkzCvgd6M0l+VuwgMLlWlwLxdrqYc+bizkDCq
7fcj4f7mZwwS7Kx7PR5Uehv0TotP3DoSap+w32TdmEUwQn6OqkxG2M3Lkd+0IhmQ
7skRKm0u2TDMx2f2SGdTd2QquNV6oTTHJd2kWt1WmTzk2TbBte/5G9RInJ1I5xZl
oPOBaQDSbL4rn3VDut894zdVZqShDF8NZ11ersACCdzCf/W0dSqoF5Zsk+tLsZln
+9JYWuOju6XrIz9MF3vBK0uOCCXT117kXwbqIGxxU9vu97bXUnJY5DYfW6vxzd49
iMcqAbESq0DocDhkETwb9xpbvo+u3Jr62nSonIx4xIexa4XoJSQWzapjZP5zjZS+
ONrVK11e56VQn9/nUf6nbZQ+zS5QorTQ+ZdyhQ6AqR7wTZ2oRKlMhWW297ikHguq
cMwULn0PCagvJ+wMRyw84y36rWlT3yUv9JivgdDy6HpkEMnSeg668rioO1T6W1Hj
avxSKj9J1wHZNCaJBSH9YjJQ1KjTpjb/k6VRPpoftZ+kPRLuR0l6JgqC09EC4iAr
zEe6u3X/DrN3xkZeDS8ZPoJmafqXQ7DXZh/nE24upz2DnCQe6Sl9M7jlFjEi3UkY
Q1H1XvKk6++ms+/d3uJjyrp9eMana4+sSO0XOJ6uU8feoRnfw76xhWIc+2PmzRSh
38frTuMhFfkX/IuN0fGJoE3DEcXTk/9U+yj5OikItqysuV4G9E8hK+bSEySGklN1
hxmd2yCMyU84ddo7Uw4QSLWnZPoKtU0TXfd8JZi/FCUl6J1u9QW33X6VL4WgxG9A
Otw3OBBWacxeEEfFZS7O8U+/5s3uIb9rg/X08smRdttX97Mt1/h349pFJjfkBq1q
P5LB8pSVS8oknxD6avfi9wu34GNXz9FupC7P1PEcM9YLsjqXXGmgNtmSOB/iXPpQ
1uXwaiettQCAZL+oPdEJmLDLxERygTSFIiF0SjP5vJnIAX1aHGP+j2gDNe10tE3R
8a31j63175Pea6xtb+r8lINc9wJSGADVBbciOnvd+H7moxR7EcoXuubpDI5IpE11
k5EI2eZGg+DSrPKq1Jgp4jO5VnmB6tqGhIGmh2JzzDj453qFZ40GyDVJXUnuXeqW
d4H8xAkwnSdh5Pdb8a+dc8WCYQGna3rauJ9lmRs3aKCzMUKMJnVmZ1r1M6sJrfCN
Wf5c8iR00a+isgpCcjkArINIgle4KjKFIHedp2ZIPOnk4Ol0YPMgF2y0g8mpG46Z
kESzExczBfb7OdHP4wSx7xLe3QJgzHja57JMNo/nzJ/Y8zn88NGhhAmJGIJXEU5k
FEnWwg4aWS2VNRaiRHxqimivpiC6sTymiMvZ8U5QWiHpkCpki+T5l7gdsvE80G5t
DgzOVfUAYvAU8zYEt+ig34UKVKAxKJ/WxZzKLgkEIjQqhjXAzClPWGPtTn9lpV6C
MLljNS1Ki2eQBzIzLXdNLaiAgJmfPyzgaazQq5kPC/sYeQkVwE6xJM+y1cduXrSL
LYAP+AQvTtCuIpxnxtwfQnFAOIi/OdN2NYV+0H42DZc417LZSCzcmozzpIjOLIKH
78vsofiLLWs4K8PMurj7n8feRM5s90CQjnJY2n8X9FbOwk+U4r8yZg1Xm4JVSo9t
DYXXRebmlcnZJQeuc/l4i4TSKvShMIHz8qwijXWzaUQJfGwsQHHYIjlyi/HQHww5
x3x6zcuHUOSnc2PgfFKmSkv7J9a42lQDP5jFq0ADDlbE7kqo7thjzrZfwh2Q8gKi
SN8fwtrM4PNdpkXoNC9ijGHVC+7tozcIGENAa4er2D1hnLJvyaFdWxperkwUdDcZ
gLdwDCT+Owj49woSXfWuZBUe9KvDttzZis5Vv9/MdbKa34IPvsSTKTtRds1us0Yc
Ia0XsXBo7B9yoYtl2ls5CH4sD26zb8ho5j1qeFt9BCpl5Gc3VoZGLYiWqOiDfnM9
CPoWYEJuooFOo5w2xZ+CCwO5iJwZv3NyYwHyyO7iSO0YQ3gQXcZI6W3JeBuGG/uc
n56etyrzsn/SwMA7/wJ5RR/QrJ0GTzBkUYtDK8HB65pTIHAD9D2jB9kaTrIBgrqC
V87rTG4GtvGHdMegLho4wM8AspkA2yXQ4RNVNpyvCIOQF0Gjuk+EKrmCCVTAurFF
cQROi7Be85IUqDxXcP3WjygOm4qvMAek7fbsLuF7ScPdnaDg8HCGH1KiPbFkiBUv
BxetZnkQGr4M7E+cITKjwXGvQFRN7TpQZJ5fVaBzdw7XI/6K6+DYrQ7ytbcijLEE
hPjjdCdWnVV8LS8AXwuGTAFCdceaUnm8/6epNeZRzyOKstcND/NUiMqNz13pR+1f
xGSHc0VprZcDrXoNtMOLIH4Yv/28ekU4/dpzVmXlw2u1dyhvnXDUgm2NaUHnLlNE
92spNzj4XkovNKspQp01ws34+nlN1osu1gwu6mcDWG4Xgi8pD5JqVUPtu2fc0aU5
P6zrD3Yv5AgRfb71UByUIIU67B5Uvw/P6LX+li5ThXFnC/74dPWPoX5JzrEotNJz
E4/Ba26XycW3uuexkhjlZxrjR8RIpSPplGcgFqFj3g1o22xNk9ASf7HeRptSBMLv
mtzC8qJCeaFh5UmytnZjwLlp0R/M9Whz+KhLae2DxmZEedhR1RUjD7PDbmBqRrYm
GTy2sgWAGSLWTFS3xL6cm78gsSBzgs9IAXV/QC3Zvt2qI6lEpPX+Ns5ASIk7l2AS
1DCgXC+GMs1AyVTrSFLUa69E/G4C51LVuUBPcYATMzxkDQ4Rk4Bxi6W6gQX9D57A
XqI3j9cdeUsXM6b22RL/n4emmy1BNAt5+nk2RO0IP7PQAKsjM44JavWjpJ0eDPhs
lOg5x724efpSsuJCB50qFn8yaO60rhc/od1/QDCLL4J/0nRqCkgowZtveG3LB5SX
Q9ec8xQxvBEwjlbC9NLbSiioOcVhjP+A+Wb9MCsjS9yLVX1nJJz2VtyEMNyN284n
z1fwdUYq2APBlEXfPzUHGIrOxCuCqBbgs7CgoZLRjEgGoCy8joC3LoO+zf9vyzBX
botf4PuOFuBBAx8miJ/6kactzWwI8iKdYFc5Z4F44lR6CefUsGYgdXVL3YaYM06H
HSFcMawYsxNcMF3B5vKaCfO6W/PV54jqOzZJyc49PlkVGTvjfTtAMOamPcz0vr25
mDgtTnZqzP+twCR4jxQOikmeeY5B6eVEJmtq10xKR/vtykjwGaWvcs3z4tEeYWyF
4faj//05Dg7g8vQZIuRSKVtADuSk1klIYX5meuIGHZS9/7o4Zjtylvvw1IjgitNv
LvG+ymydlxNAgzipcLY3mwERZhhFe/RyVTcFJQJUljcSBTnh2SNVWAnEC1f9QdSE
lZIbZUXCOqC9DdHkN8MlXWzKeIHgtzqSO9Y0D4iok4DYv03Xg6Uh+j/LEw2ejjyV
ML6kd49Ethk3wzCXBBUsSiuOCDb/JrgQZza4d3cWuQNZJv+SZOlod7NLoj8RMNAw
QqiQMqGnWic+1jO5GrKBmm3rJBRKeYiJz0Q65oNbVKoWd3JFVMcvZY/TOcr/TXs0
27FVYGTGECcaZWBXf89ppEX/n5/EXmTmUqeUhOU98Bx7iUoZW6IHv1SdMpA5G3V1
r38WYakYNcK+ib+O6ALn3ea7DXN5JJVEGO89FyBUha6CZ36bDe3nApMGeAn3M4xC
M+r8I39Y3NUMGwtVHeTm/wGTjtgJcVPPy3RDgoNsSkaJn4koakc/FIjXiwh58sbq
u3bouCXzJzYDvyNUCnNm7sjCs3CMtCJaS10fUUL1LTZV1FQijji/Va31LTM7T4pL
tdi6kxkoVUKJ1JdO1YIIMQ27RY0u6pSkgqOyp5PLnAlIAPeCeaz5vucjeLea/q/i
AAKNTWHzFULmeZLozgcjkiD3AOXMiSdkOl0mskvWa9xu/pr/I+fSol61m/uA4TYK
NiM+vD5ypPDjpmAAdoLEIS7uLYIiVGwoCQMs0qNP3rzP1802JdIbHh5dHnHCXtO4
5PqplOrYUNi6O4W1R4dSnil+eymOCNTF6mAKNv59i/i7B4bmNKefGaUfpne+a1HE
Hs/anl/cTYJUZhDJXH5byHBZOeWFXbqmgLdSivg6TW3IivbUBjTSqMSdPT/QMoRb
pdr2HzfJmYf6x0BKccQnEhFnua3nHayaO06wIBTPUsh1g5jJnsUzpzCtX9tSUUAQ
fzlPdMhVQfx50n2uyNkg8PFyAazn2w9krcXRCiLPtaYjEON7UtYIQyT1thWYOssN
1fXKd9z0uS7Q9YBH7SFlWWmKpTpeK6+H99Ay3pUfJHZsd9nV3kKDxivJT8geUfr7
1VAHhl6LLS1hvnYS/O7Lx2Ln1fGR4Mr3R5kLYg+BU8vuI0+dWQV8xvXYKfY1HYh8
zSYz6uYPM06HYRPSfsxg+oAtmT7Dgx2u4IqYWxJBSlRl9pYH7cNPYYwNjpYI39tQ
cAcilaOZvRlzfNyVUhS2FJlI0zPz7WRx/bEE7deVFlrz8gC7vbHVthe8rnNiCQ+N
CO3YAN4AZZy93ecBiI8gN/a80j04AzGGpzQSxb797JFbhWlx1blCK6cPjUbEbQpN
2LeU29jwJxCXb5RMdiudEMmbSWg30g1OwMDc+miGNGDHvhTocfKPDl9S9OYTQnpj
267DxafQyNXhljMLrVez9BNAuKpzt/DWyEH8AsVa+mruv3FPCo+7pu3H17JoqYA4
MD6FETeUHT2ukM2S82MBaQnq9J/jNavdlrI3JthybLs0y5FWIAySTJi7I8y1RCjx
ppa3Gvn1r7R4HOQreGntejupeCAep7TMxh2mBtp1j6NuFuoIDF2f/EgM/OgAxlVV
Q/dXVU3oknoPCF+jVzi0rnMNoNNQxCWhJFieC9F49Kd0bqHH7yrbrhV+j6hNMjwL
sjBDVm1kVgPUK8WJjIFgI5IHx+Zgoq2zb4suMRtRuuVfu0G9b+IFZueox9Wt9QKh
3hbY880qnecD9QtqJZhm1i4BoOINAMDJ+rCagN4y9NZ0EtQdltSXvxAPr30nxR58
hvVCbxnZ9xhVIb3kQxeRw7sta7n+NfxWjxbVPTbytceTEk9D6g/wJX1yZNM7Mrmn
AGMDbKR1M07VHlR7OLehui6kpIREW0WNeFUVilYwfUruMEVYEQXancXFmnXdmZC1
kjPHse2Yq3d/97KGR4vTiArzZ3Tuw4+3BBh5ZCyfINSffZcYqpmaYFrvrhF7tWp5
`pragma protect end_protected
