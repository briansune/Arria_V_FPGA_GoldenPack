// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aJ7bf0r7T8WRZ882rZqTGo1DBF/SI9Ucz+lCl0G6T2sCYFdDLBPHuPCb9Dw6nOSX
NMVZpHXcc2Kj9GM5LHtb45ZPuoeWEE75/4U5t9a3rDvuHjp7NpNC9d1a9H4N7znN
120Vst1YjNw7iS6rk8bM8RW8XqoH9xUjTsYehyo9NDc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7216)
laCmVo4aNz5wmyEYD6ThYmIE9bmm6MXP8k/6AbhsgvGmSW2hpg0gJ058szP4bEIp
1bk+9l4hgz8CcMA3e1Hubek1NzGj7FNTLdtg87GqWRkGcgqadxEtWVFo7YhsD5Mx
sNdq3ZaZ3BF8v59Rh/dYCKi7BsDEG0JKghbnkPra6evDUa8a6pej6q0qKGdRGPEK
sQYyXxZbddlp+yDd5raBHSRD2vDjZX4YYJrXd8PrLA9+mGff+TgOoMIEX6ijrAEe
EWFxQd/5mjVsqcbXSWlVMDVHJXSYZLahgwrunym+UpacKdQLqkgIsDGan1zB3CYD
Qj8sy0L82plyACKn+/dXJvhPzCKLAF4vrIV3jyqRGp6tGAjX9L6wSBZy82AeWkVC
JcVPAs8g5BWBxKiEwjjjdGpw6phHSYMJ3csrbBQ3Sfbia88euEJ4cRjeoUbawxGW
u0BV2E43hVJaYD2DJUVv3Yja0jw7OTJNiK8SKYCt6vYc6oStFds906aTQuDg2aEl
lFGZr4vKt2PShJ/v+zltusRDkpQCIk4mr6odH0XlCdzKfqZBxd+UrFRaHgS3za6V
sE7wSm11NWSAIxfSlkeH21pupgQD1xDC4waZKYlPqSrMQgfeQWO/oSntOW+bb7ve
si4DMnKry0mWtbK5FztltGwhGN8k6uOsbwEq/2zWK63q0RcDHkoWukDMLCo5VTZI
tMCGoz/BRyNIt8nW3aw57QOVLRtFgLtt6vrMsBLMngdBFanx94JxVS0OJmG/mS0r
qda9KH9cTuS7UpGPK6n94cVDPGTop+Kdd9Z0th0k4UiEcJ7apw4M3jKwTJgOI6qu
jGMI+SWcKkH65LoiagQkY+FENvj1Ja7sL0eA35vd5phZhq9W47wkmR5xq/NVSN3B
pC4RSTnre+BtK1mkrUqzDIrMG4rLrGbWV2+9aS9KQ7+LNrjxhSafN6pdqNoDLPne
nZTUdhD9S3SQclEdy6TD7Udlu+UY0l16JDZ1FquwTDSSz7/K92TABfk5R5n+HpjE
vbXjk/7BtS8XfeTsN2q/aaVSAJpWMIOZteqaRUpV+OMHPHNE03zh1umXt5ChnCCP
zmkqR5IUTR650uFMONOKY5dJd00xnRm/FQesvW8qaRJIc9M1LPrxpFYdhY0AWn/T
SEDIBIzuoj3iyUiiN6lmME3tiTJZ7tq9fj94Ax0ayuwzZjcZNweKACGgsga0b641
xLpbebGI1LhCo53XspfXWcGPxniy/KnqPUKJS+idRoVwIk3xp/2+sQLBYgTXYeDv
XRQpoesUumA1uTR2UqonnoiiATL6hr+0C2sGrV2GOfOx3L+f3lOLRAv9OjD0Og9z
YsjOcyitFtcU0asGGqwxvWF4YsdW/G6bfCKqrdKVGFEa9aUSQ2Rhw+nsopiyaRZl
gBV0GGvoGIxL04AKRxn/0K8dycgvnyvP4EmZMe1Fzf6V+hYaY2Ch4aK3upUWmvcq
bb8Cxh27BuOsffqpEaowJof4BgFFpfB8kFxarhWekpceXYDO2jdVRsuChobz+6Dj
mGvXskj7+SheGCIuhwNsZN2zVqLrIlAHIaSbhDL0Q/Cbo+mObrv8Z4kw7M878JsV
v/U5kurAhWVZ1hguJZQgY1t38oy0um3CF8p35JJ1E69qc1wbsvGwNovr8wJMPvud
1e2T9ZUMOnGG4cz9MxqEv05fzjWOZ9E4ojYJ1ewYRzo051sc4aMHVJ2tIVZDnmQe
hAtU4+0Dxv4nDqyfbNYRI16TjEkpi8GVlkQRmNN293H/M5XdPAUM7S0gJbaI3sIm
rkhZUWVZFZ2Pc9svJXAUU96NCFPKfST64DpF6FdR+ogi+VmTFv3GtqMs1mCOZjLp
ueNnQ82cbIyLXFl/XWf6vBC/cghLLy7mRfMLRngnD+T8lYo4oztIpM1Aao1rmeIl
ZM0AwACambmHJjAkJAnlbd67t6/1HIcAu7ZU2LKLEQADKoaBNILVYIjW32FLCyPM
wy7ws/Aof2GRB+arC547aboAQJkWXPhxjeKvl6watcAaLTe03G6TeaZSSpdtenAW
tjrhpckDaNS3dApAhSxWVavUZcLkECdydG8LQlwGnVkjYWq76g0olo3/SHgcIVJQ
pg/PV9Tyi8M9eNPPqYDejbG4Zl8SZZ87N7NrPu7U8yLxYcXDF1/Xm8Pkvyv+/rzv
eZZYapVgsGwmxrqO+WUPu/VA5RpQe2depuBt/cwfhopPbvSz+lxqIGhV863DRQ3A
TEJPgxU8wDuiINHqAb6nLNn22g4CUIbKvYLSIzXDBaneQwyfweKqIJq/xc8VOg9w
sdSf+Ci35q0vtBPrHpOt09gxwGsOmxkfpzuqOFxtrWsYGUA9clwgWokdt28W5lXt
N8wG3ODhqOPnO7Gq2E7fgM2e/c9pyL98hocYSP/HMOTUptcupOIPEQ3vOWB/QNmU
+Sd3ngAWJfnC/53oEkDfY2DMq+slODlDQrgulnAmRDBoz4FCr4iXDWSaqTEAZKKX
3PqNtrtVd+n8VskPvSRKKNf07J8aKm9of316Fs85UWV3EjFKJCrb7BSN3Uz9r/EA
CNJh9RA0GJG3X+vFSRba9HT7RpfdbkixVePoWWbKaoXmNddi7hjrr2+7/DPXhVOW
eY7scpJa1jJL0W+27oInx0oDD4YKCUWtXtH6zGuSAYIjSQqfkWKjh1dkwYo4kvWO
eGrxoD72YVYZ5dpgiOuhVLt1KOD9VmZeJyGt0PmmNYPz90y/yXn4j9hsfwYlAp6G
/Ub0CvGX9qOipG6IWeHOi4QEbiE1NAec7ZlMvAV9WKaJAS+UeyFGg4EQZpqjQ2XO
XefcdvykdtqWSESP1W6xqorHRLSts8JGCoJ9NG1gSuPe+tMQQpnazUQ05JcZdBo2
mCQ2fcXv5r6LUKaf4h8scW7y9hmUW/kZW/1NfGSVXPPJZ3UAjI5szzY+FIm/Jc/j
ZSJ8K4VCOGzLaFdwiorZ/xGVkzdWJfnR2d7rKp0xpwA3qKi6I/XSMf4orgB1fRXW
2vmCu50GFN30b0WTzQKKFC5NsgYOFjdIjhpNyXMJjZ4zYvjyuxzbIthpPpWMDXGy
mjFrcDUbWyoQhe3HoMg71KWfKpaT4VfogW0kXB64fmpza2TCjxZWKNN5dOVbd714
wR4O7fOmaGpZYftDXQGSVpAgfuPt9PRV2IFNbYcGT8muHNFTNuufe9iUzaawlEnt
mEtS2WpOnT/uKj6z+vZfT0ze0s/jclA5IulzgAvuMBPPvvD9wdT4AEPkkXKgGb49
Tit2smo5NN4EAkM9qvLlObcXNxyi1ANklONGzWOi6TFgDgMKJt6eWJrVgRN3EJ/T
5qQIHXJjz+/ZiKLI3W3unVmvnijfnjQUEfRHhrYfiP5WfncqZyeREKJmbmfNY273
K+td1YuMC17cXa3gqt9g2Fl4uHaum5NdRGTzi9km98+ckm+elvhJKhDaC+J3ut8t
QMAXktAAHJRHUeFlIU/F4YcLcNy9Fiu2KSKGd7wCJdRFVXTlOz2uOtnmLFY01+3l
pnihXgwqxkZflRAPgmQvAPJbFv3eIl7d1wFBdTEHnwa2O4d+pe42JFyNZ/vfsJOU
kuJtFG+0nS0dNq2uExyuNeLtRGdmTpx0ffD7aYRhW8MIJm0MCQoHWEW+3bCWacWY
Ji9Gz8m8+9aIfJLGTX6dwjDmOGwP8Wdh7Zm8P7vJEzDfEBzMBo/JkReGIQYyAxCL
CqGL/4//oU0jQtTIaAlR2AuDrPRU+JMG2DosbyoDo8pseyx4bgyQqU7C4G8jIJnC
mEQmP7pd6Pv+B7q0vfYRdZlnp8YYWuR9STe+wWU/wXhqugLCq0w0f/cvGRBktCkH
e3EU39WUl5Hq09OPbccvuatz8QGM9vgAhMuj1R0mXGSJGr3+mQ5cj6Oicekvc2az
Ouknglj0sk9xwZAp7HNXTMlndmnWaEU7k5FY0IiO69YBr0gubG6OHZCQ5O489hYl
LC1GpyEka+NY/Hg38GigO4O/6P3hRlr1Sdn5u3uEGnfDTCdomIoRwk4Sy9D+7wue
dAd/Hgg4KfA58PH5hE63C268w/DbWoE7gtU7hbtTov9ERtH9fs8FGK60BFr0g3ky
r4oL/8nZz36wM6Qb8Em2Nt2+SW3gjPsbB2YfK+Ap8TwX5rcujKJQzpwS/2OiMUSZ
gTrKpjs3Kq2PBRubFtuw7UOOPPQoYmX1mR1vJMH1AV/MX/9gXWgN0BEfX6CCWolZ
0NOGXJHoNMjFPV22cwthDWVuwTwXxHuYM0KYA6TOXChwhfS276QaSmVcdSUy5vTp
Oo8J3+ub6REQovYMrsKPsun4mGtQNUyxQiMGZkLZFuEP0XE1Jm5rh3z8BiYDpctJ
CNqFG9y5iPwepHcqioPz/eVx3TAQVg7XZJcuUxaN7nRIVN3K+cGcEW7aIS8NzbiG
tthwunhYJh22KUPQEdVzGhU1MeVOI7dhbdqyGU68EEC0L2SeIHLkZVu7n7lGUTbw
z/a1rqJ92rXoYyXBRmhUKN1XRvt5yEzsOoYMeWKc6tw21O3XySGlvSkKIQhvo3tN
n7BgctpGDzHoBajVPXXy8Gns7rqSnLlFw7LvbFo+3h7XsuHcW0nO8Mz8reZAfK+J
JfBpLsD3o7elvWa85VO1qXrmLBVIs5uTCVtOrS/WbpqVcS4Vna0J37tnMnHagfHi
GX5bQ5o9ljOzduKoYWE1nc8QVq30Vs47FF0myiEun+yPJvzeCAzPZkPGDHYWNxjE
w7R43uI+aP3E4KCMKqxL1LDgdohQA0RViaETMdDBW4xkwoIpkI3rUyerKdd/ORhQ
rRTlK/rN59ZTlud7u9KrbZs+SSQzJW+5We6jQY7+jxDfVPdSu69l3cnBFLpIMJRr
BGO5b+ZfNfTA8MCaOuC2EOPAQJrb6NIH7tZDhmN+bC09wgeSS1H+QdwvMDR3Qx0Z
aUuQNuibQ74CayBDHNw/wDeLUnkXs45tDlv5vfmn5lfLmuGLjzKVGmPxd5Er9Yw3
MQslsbr28EeeKtkDCoxISmdb+bwyS5Td9Oex9dALDevjGqPmv0zKyy8+Dvfq0vGb
jDzNbH4Zl7hg/lsan6RmQrwqyGeYSvxlIzQoiVGV0byGQOVcfMqOQcWSY0QRWkP1
dtFHZF8o6tL+sRRfE29LvdWHd+FK8FBH9hLsd4OPoTXs8vNRFtk88DL9CRIb9ZVY
/di2JJXKYpTB4V1kF/BxSFhr85gS0sDWHaRww7QOahbUfYeVQlxmN4fU9CXnIbef
ovKvcRn8Q0TPHxRxewAMEPJY/V7dxqgJ7OT5G0o+ymLKH8o9wqLRW26zRdwmz4n2
lbuvAQYnXqAbKV+M+g7KeIPWoHk61TMZAroNPClK/76DvuydD+8vsiPIOE1alFmE
VmEjtx3HNHViPwmGVmfcgJLpwrlN0xxmGc9L2KcWVSDKNQj1LrBQQxumnlwtoTMr
G+OCfAtNUhIOt30XVqbXqt7qZMoasHaCiV/3UdlQT91a9AibRDsSNXE11uXu1ieT
eZSYE1Nq8AWSqb/WYPSjcCjSkxPKe05PO7IBA29mF5Tu9fDZn7WL9jR0nhKHZS7e
iE0kpg6doDXbk5nwyfFo5QbRezg0dscep4Pv2BlL0N75tTHlEi6iAvyv+fQKRADW
TRR38Ws3AJwcfMgtNLw+65ZrSpWCnMSU0rm2Do9LNI/EIIbAwauqsdLN2rkGdIBH
Gx91OebxaLilJ5svqyCaPoNR8RoyN7mVbnBXVBbBZbj3JzufTN66XVz+P8VNVLUb
zAnqWw/NFQZIyz3ngArIOXDkae52RJQn3MIB40qO/9UH5J41yZ2jm9itK3h0KrmW
5cK1GFs/ftHqnpIIqFfpUoCKkOarke3LvSbSwNpGbC1QkhBUcOFiBu12q59R40vL
Ac+EdOBfi2hdlHSJpAZmQJAYFrzVcM62W3caUGrPfI2v1vHoO4tBF1aLGDtyzhcz
zIlEUeJpfMgMUXXF8kvhOoXu8EHBFzsGye9bknf9G7Eaye426UjI9jyeplFxN0Gf
9CssgWo0Qj+TcKNy6GYhupA1AdWuHdfADX9c4Ic8AI2A80CKr1xUIlgFvauTS8MX
kZwajwE7Kq+qZQRWiLTMWRLhNMiqvoY5Rwmin+15j4XcOpNpw7Lyo2Q+nFfk2EZx
nB/cxC+qqI6/0LTtI5KcPSj57zhnh7mAwqSu1cc2VZL25eKoOv7J2KMZQ3yUdtb2
p22l49zo2bIJNhuh2pNzBV/SGqE+ZOIf1OjuHgBmRP62sfjBssm7LUX96PDhKlvr
ORxrS1aCtK/rXt4mBOtb8hzXC44UZZV/XdkzZ55oszZI9+Hvedjq60GQFiCFf672
tcHAeX5+D7M9cZ9h+PZP+hTQBtzdeUBDWhErSvxh1ybZPAYfvQ/voZ2yZojUWooP
4b6pruUzjDEM8sIzPTAqCQwH/cCajZ1x93XhrzpKWcQvjXZn/I/TiFCT2IFwfpza
TDzgJQ5YUwJNvb79ybqhqQWZna6I6BDYLsTU6+2ovZJ2nwWRoK3El3mYCih+tN9/
WuGlnuuYJBTeZ9bVgzNILYdNmzzvkTMkWaD9GmQxxIAU2KDKBwivcjrTxUOS2MjE
Y9pRauj+0ndbrWwC3cGaTI+43XD3DiviexeZ1QYC+yj81vAwyxLuhTO61wPbzGjG
CUP/2mwh85vkHXbS284iLcPOSBHfWV/GlCZ5HD545G8/lcxKc8Y7/lpPCE0pP/kr
GPPi9tSkDTj529sIp0iNB+ogUFkB7zqpAC37NSPeOOmtUPEPcA9vLN5m2clBbVaN
TAeNh3K9QCDOxa/PGGZqSYTtByoXMGltfH+iPxb4YIes4CSNgllushdELT/x1B5j
rgr/WISqAK6vKi/6pUoQJYRrwAfGR/FBd8+gQswEVQ6ZX5CvtcsRbKXiqfRqkZwH
uVeyTa+fovePQ3/zp92KfdmTpTrcd2Ju39Znj2IXEwaycT4ZhQk+BpIE+QXC9Chm
rgsXjsPfJXORN01qEn1jFqRSzENQLpEn5QFB7cU0FZ/Mi8bsk7jym+RpQPexpLQm
vE0ocFAfK656Baw0HLdef1j8L4Bbhmve1Yy5tRaVPqA9N8ax0uRf8iIGM0Ez7B+c
T7jujuy31NmIFk9pPrGtJ4ozbfQAOIu6+KIj8VdkT0MyLy6xmO76W87cybAYFU4n
aJPAOw/2kiFzUWA5tdrCWQC0yiO5bZYSazanWPmgadWnpto+o3MMacZzf9J6gRBu
WPa0Ju0mGxk+uvj90aneobC7ifmfVHmzXrXLX3SazilglWFnUa9rnl2cSf6CjdME
PGJPyh8pEXfgkwcjhHnhNV2y4YSlBD83DBb5Owga0KNweFUU+JqcTwfbq3ZrQ66f
ifV7eXyKHkwCHu5kH+9qJkbLWDVxLJhLSUd5FJfdv6lRatJuxmTlkVRZUZPVx+Cw
zyTOusrFSV6utDw8CmRcwMff+rQr7qPh7JY13QpULWrTz9rhZHyYMU2cUtLU3hTj
YJHgjOzqqHceyEN/0aPodTTX9/wRgphJ8/iHVHX5wKn7rMBHZVUG3fQCDCNAOZfg
UG2FjBzWOwTJy4eNQgVZmB0SSSfyJdUV80Oq/wO+Zr4J9LFthR1s9aa3on5UvgcL
9opIc78DdUkImcjK2Gb7MBoBk/WPXpokMn5DKZDsQ4d5mtGQbm2hF4FvfHC0wPxY
WV0lFbJwf3rX7EUhTEkiccBZWoG6jDd34pGLeMmIhg8lSVuO0uwaeZB7wcZiJm01
6DhMKYkwZe0p9AojaLLWqlLTbNAmLVYtrKSCH3dotdmAJYcGNQOOQZMugRUcWpzo
sEZgY6lyG6gnEgCV3xCA5LSyN0aSYpx+Gi00USrNLmeZteDxtUPZ44y1Jfb41WJn
q1JycZayvrnDhwX6Go+Ad6zmELN8FpGwx0vofHzVQPsBm806GvhYKDEm7bYM9guN
3BlTarYylMr4MrSJXiS9qlWSu2d2pD6TegGP9+lFEtGHJzcGOznaxlOMeWmnEE/1
Y0UmLJKf71hjMC5Xcp8khxz1piJvRh8AIsFVTR0d1hZthCY0kt2OecrfJeYIBWf7
krBe5HnZfxYhr6ztJq5LTBsXTp4cqYoV/c3OUDYWbI7zaaM1/mmgUL/sM1sjZRzP
KCPIxr7HvlgIytCfa24ptRXLoap2Ft7QnBC7SZmLo5kOSKq/LF74oqnCYXRQtyny
C4Pp26ukrUQGz+7U1d76EbAr8uEOFkY00CX+hGyYCpifD1rxuzckZ3R64WxrcxdY
CZQDFoyn+rYc9vR3QftYndTzPSVAudVb1Hj++Uh1coPtS5N0aeF2x9GEuyamr1V1
h1XN51rll5+HpZWSgbZoSSXy3IkksJhy+XPnJZmeeEU7cuDpROjMiXHjjeVsQvj9
TmHB/Hhl+o/YNRAfzLp4Iq1KVZtkpkNtY8N1sogK485ACWcSfZzlp+VeazGsMXNG
WlNhza7FJ4I6Gj/t62rZxqUwsqXr46lnekNRX5XkYAiR6lk4CvnoKgKUzCjvwC+1
k7LatrQdNckpVWfGFBs7tOsKahAv4q6X5lmS55+BlT1dJk1+Fvi9KzP2Fs5HsNf1
XeYTzrtPOZxcKWJK183XEVQGNtVsVISCdKmrHYx1gaLKl/N7WyxPFzQ6FNTSQiCp
CyR0PKeJMTuYgmWv+ECvLAlHlwI5XCiCFHOV+qT7UjWEsbCUyyj9ZyuB9vRoxrwb
W/goX7imsEXXCS07iZ+CKDJcFpJnePtDUBQfvH91jkYHIG3hFfiQPqTdkRtgc15I
mkWsEEZ9iM5ycDwXLPHCswF/hxeJ75i+MskihUWoDFHVgyTY7nuHW6ofGYCRhtoC
aI8If64iNPOc4MjSJyFeUHGZw6fl+A9rFTxZm8OAx9YUvOMA3M2ONTpBiAFdAszp
EFktXceazph2Odg7iKAwKpD0GCmnCrEc1krRk5wW3x9CM9QQGaXsz+xHv7g0iBZZ
q4AONcdXF+MoLxBuSly2Jovp9/6DZ9jMBjyXPbDkiZVNkp1EKwSeJvLNIXN1QUAc
Yvj+A9Zsp/dvVz+ZIwfJ9VKBLbkRVcRj8YXASVh2LSCna9jwiVX7J5N44Kx9Fcim
WC/EE66kEtDilJYuCaMlyW1htZcRQ8Wycyg2U3RHGLNTgkkh9Zky4/a7NbeUBxHZ
QjjnffMkHqH2OORW5VENOqVXgTfTljUafuEQWb4+sC+K8UGKsr2VwIboDDO+ZBwb
UZqpLpYr3Yc0/M79XZ3rjvj6fUZg88muDhbE8uhsUOvRX83DG37ILtVbE/ZRymnf
K6MbAqiA1jIxbq8qCG08DqA9p5Nyn0rrbqWe+fntloN7B56MMLaj4Pk8YsMaWDMs
FRdNT7idpmgiMz5N/yNPRPVQ6txJPlf65dT2L+dyFMYiHt31Ud3q3JV/C1aH2foj
UB+d8EgLPo/FfvnMgTh0LRbvA3sa+ClKDCejCEUeAJk6mrEuIgbLiPetKRXzEqcf
mEOLqJ2w95V5d/2h/pPYfYyhWMGGneUTqgUboYRnsC4qCXq7+puLngKQlIcvbTJs
pqdhethhg1/SiUGJHDnZ8+o9l4/QQ01Fj9diLdMs7oALt1bYYmbB3wGJ51KW/6H4
HU8q3CdD70s9fQd5SHTV/w==
`pragma protect end_protected
