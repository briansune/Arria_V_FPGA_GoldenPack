// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:36 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IfTvMinH3XAiLC4xHD+0qWO8VUeqAlwfMlX2FxOfZIQbN+4LTx3VdP1YAkJGd3Ng
A/HuhlOo1ZECeCidjlmjVMDAEdkI/JBpPY4GgvTSv+Iusv2FStZ3DYZnyCkKTKfk
vxXrWlaaik3PSsESJivw0g5tbFLOezsjAj2knej4zXo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8256)
lkP/burm6EdZ7HiTCQUbVzxE+SWJ+KM+xCpC36mYDBBT/TC34IK5qP3J8vCDqj6R
bJZ5M33k4UaYTNs1l475o1NYatQsmAEu8lvBlOIZ0WX8G6AFxgtfFJxWeWD9CzCA
oV+s58317fWPdR/mb+fYn2MyVsFxDdQ4qPugJQZI9kmmaM0MgShlfIcyItwY18iZ
xMzJpp4UO/2udp62uPvBNnn+GSs2kGJbEZvYK66E6SYL4Cv5Tno1v5kJ5/C9qsX/
v+X+Wsx1hd27y66wi8GPQ6AiozGQr8C/upjsjft1dwgZAZiQV6Ax6S+SWxJFA3i7
a4fns2jCvLF4q7lFCSJrLWoWM7J/iiY5Vmus5uNXRMhh1QS9q9935YOP+3JzVYTz
RQUIzYAj3x1SbxjufanVxz7gcAjnxIz14sp+8fQcXSOZ3s/w08VYaCMJ27Rh8IGE
kK5I0maJozh3AzaRF0wUR79IrVeGpefkhl5O5gxNXIifhdlEbk4joK4FU9l7pyLN
fxb88QT/x9J4f2bs5/nrDKSweCi268fvkZp9DJOUe1wETvXqL1E99yMy1tc5xg9f
s4dFLy3t5gqKxS5EyOIP7R2ojjy0M9O+10p/pzDPMLy+gE4UvKLXMAmbU91Wl2SS
l9yMjh5IzdaSZSic6lVvkUFzFEahvNCxOdymIBy441TVfTd24znnoglXDgRRe4KR
WbYkYB9s4yrnN5zy+DJFpk+/ScRnvbXeiBCq6lUQL12/n13kQyQqNzu/Hh7pmr3C
xhskiHjRbfBUv53ZtD6nmHnlGsBxBTPmJLSz8CmLeqaLlUU8N2N1dM8/ei8MbazX
AilRc0Fg1WIW0E1f2KevH+3MNUIvC4xJIPmpReDNepMgdkI9oqgVzgjEHI1YuEok
d9UU5AF6oi+5aUY6+/7KBQwUngwmRSDVmUd5tu20N0s6epVBRDoWkCTPO5uWL19H
EQGoX8RuAjVGjOlcJQKQ/4ytLglaPuDQni4kKCgpp/P4qW8lQNxYL986XG/LazxD
Ny8MH1L0J7yiH6wxdEOTCYv1YYLrNPwHo5e1G5g1bfyKIkfyohRsM3/QeF6BAGYu
QqsOIhY0pdwwzrQYmRTERlnjRnp+246FPvUWys1AmXgBSz1FuBPTl3em63A2FhzT
j73cS+xWnRaGd4isn7oG2na99n393LeMhoxLM6egRIuCP+zhs5r/0AgbFTWdVqZN
AGfDBoHRXjTD6tRj0elohsd4hcDq/5/By2DWmsziBomV8vfQV0BPJIeGR2JlDaHI
U2iGAX/qWJnV3WFP/KWJy616ZCaIo7yvLxUIkywt3bKP5y7KH722nz9V0SokNI5i
sQputJkXV044K/MznfZW6VRidvEQQ9tnp2p8kt/z+jnaLxTee968+En17fkoCGpO
X7cOt0GhSHFBU8Rq0GveNXC73/otb3HMad2LzaibAluLbUS8teFJnddJnoaVpY8x
iD7CyaWkHJIFsACXJ0XhP5CixrO9BWZ5Gam+bc1YzMWQvATylT/AXFpNzvkmw/BD
08bZd/rZ/0Vf435eOTkYXlj1CE0yd7opmhW7qIrug9ysdEnXApEx4KHqHLGXw4cm
BWOn/NdK402eHS9y6s0+piJpMTY83UhZPhr8IV6zilR6Eu/J+HfdCKi09l/jWOEg
36f9oUyt+BtgYjVC6pMmXOWgrvjs2d8Zy+2sccyUL+5ayNoE+duv96PuL28ppgT0
ZrBs55bq2WA2bToAxmykRqQaS5RRKNAT0BZEmXEXAhJsErmC5YOx45U0ew/jRNb0
5oi2cXrwXA5OwEPrVj8ODwm4z4H7JFp19/42fAn5IamC4/cjcGCOMr1DARWDPxoR
CS/kJum7SUYy4h+20sNpHjW22KiFrLNO16zz+P5/aDMS0ulM48CL+4SNEU6krMK8
DuSzpU0Z6n7/3UNzKdKmvHr9iYA/FWUeJod68kHG5YlKQDL81Y7XWtZqQvkPhv29
9SRcPFyOiCvB1pxsYjGFmXSVw8bAAOJvOetBQ13g72cpUNNCVerrutng1kx0ieZP
UYQjEa9KbZs19CYysfZE/tkq6yp7pTbneIP0kw3ogbomzLbci40H/5w6wAUb3QB4
Bv6qb0OEtPDYXup+rnXuwDHhpQv0SQ1zLowKOvDfoXnD4RqpfltDkFfz28E/tU7+
yzl2oVMi5Dws43hBDLuMJIh8TM9Xi9upIdZ4jNJIg9iaKzke14Q5lXGxpBwmm4QD
+e9Y5hkaZk4b9apPtpZ1vWOKUk4GU6yViNymRIhfRJ3Pd/tchjreZCKjWBn/Qkwp
oF7x+/C9SX7kuilZWVH8sqNHxF7m8QkdTHIog/TY1qenDU133+MmhG0CCq7f9SSQ
ZOydWjClx+qFuCH9022zM87MervbYVWVET7lfyPf6wi7jbyGUQwlFsSVP1bUbM+L
2FxX4apfPnQ9nxJQIozQa2ceRzU7gejmYiYw5vRQfFZrVVhF2hP5XopcyaTuOyAT
pKiBDT3MOndGzx853yTBUkHh91/V88qpgqfVy34k1e93O0Wl50D/zz/TCOcIJhan
6ZSbDs0//wuRgKcXlIZnwcc8nGWZPLwelP8gboFhHb3k5+ygr60odGK6JpOi5TXm
tEPgo/BAGWRy7EHDDncI87WyVcb3O3skteq8MP5AyBeTvAgPwk0bNibBVuhfhLvu
Gk4uaCTQTd/FDs+uhyJVycGPs5evK4Eoh9HyrsMoOJmMDknKkgbVu3wIBovRKzCe
JuRd6qK7l7S1mJ/H8sP2KZl/0oD1Q9NumXebXcCYhVLO9Kr2p4dhZkkvll6yc8ol
Hem1zykla0BqrZKQx927xjQLqlKxRhSqtlJMeiKNLo43svLhOqEtRML171w0VA91
kG+JFH4WEyUPZK5j/nBUV2n/guLe3QdeU1jkr5zZN3LlsnlVWDPAwb7zEVOlKvRo
FfvOjJ3ZZs6HWtl+ZsUXI3PbUpD+TQo9twQLBmg+LJgT+FUP0NPR9iJKLYkbB8Lp
xh26WWdnJ0DHqSwod03SoG+lZQXPdkU8lEECl/ISbxlD1Qmki9ctzqcrbBX9rO5S
Sjagtv7dyLamWydJB2UEoGgQTm40LYXIWEmTx+1+V1d9wlXPBmUGcSefoBewgTmg
EHAfYobpqyTr8LqLvVEGn/5h+/vOj2r2Xzv8706dFRPi2HTDYtU/cREy4xBTwOJq
6SL+K6x0bwuq/Lu9w/cOaCRPA20ZnDY3IaKeDstY1qO0Mjrht5ToOnYwh48lEeIe
YgkhcqNWrL5SN/owZJcN2dsZ9gJxC8HRJ5glAJPqF9JWss84YVxlnlCTI7oZyipT
t1hxCZnERRPFBB7Ih6/EsreGQJ4AsJCwY1DDJphrOC+mZHZtLA/vxxEE6olnXucI
MBHJGSNn87j4aRyuDhp14VYR012AwPy2AKTM3BZ4TTXPEJLXA/J9E7Put91oTsvo
+4XP202YUhCAlPMinIG+E97Rlz6Sy5bn+oVJo9Mvu3dxAvMszu9qgCqc3QUx7HHO
ZAmxxTY1XTyvFKP2X6h2/9Ar9RgIQyDdI8vPL3QvyzH9R+PGbo5RnUXjHq3+1kOS
DCy4/jdkzNxPaUQjBnCNoSJm/dREKbDojygzOadFq8kGitFviZoKSGg7tOQJXEkp
DIyz8MeANa4Bgrs7+hzYTpuusYEKlUHzoKyCflxDmSufMSoIbPdzlYKjXLUTubkM
QhvV6856YHzXSaBIna2S6uocV0Qql6Katb+70GZRW6kJjoECeiXIjdU3UoReTFxD
eHkMhXMk0GeBOwZGIpAa0KazlKq+QJMWwgWP/4zZ3r1GyB0JQt814SDqKCq0h0x/
hYDKHkCt05BTy4m3stuWs6f58rPtRO2c0yl8PZQAiJsOCxxpC0N2TN3dbmYl5PCM
1ZxdXmg3IPD1cJo/dWpYnknMjiPPLAV92zzqFxrCbumdFU1HDMQYq8g95IcJQXe/
vKRg2ZBqV5XNK68uBG1LqJhlDptBrDljqvJtfHxTXJlxtMPPtL6tQvzh36WRac3V
Z+QBFjm0SImxrQpQyk+alDMtQQtgUjnoIFeBI6mQ8sTI1eOHGrpBQJ7u0YmwDzwD
RSGcpIaNsZpnebodI8IcxPCxdI5fUNp4U6W0V5tORKOMeq0xm5/VRzYSRrQyRMFb
j01Ec5GxeHuduR9Wk84e9PK0hTkeZ3s0fzqtHnWR8LudiWosBEkzr+ANeXPB66v0
UxdeC3JedjGlXiNidQ9xxr6dsALdzxPa705tJri5d/NNXou4GfsNZSbf6LuBKid5
vMSNRgi61c9/xzVwjcRPMGpLrkEVim8M//0O4ZQm+wDG8JBl4zVUDAgINLFWqugZ
NnTZixCGI7s9Qzn0ramJeuE623fyGKS3sEB05IRBexeHVAz5w9sCU5awBryvAmZD
pDg76/VLj4cS44CQ4XwZtWyRZcJXPWDMBJWabowJivVFkkblOwYKBOX5KtzodQz7
zrq8ig7omYmFQneDF2fJeB2u/nd5m8Ue/821uR0KlJaKvhNPVZwyTsJWzTXsdEFs
oAdPrrYqfMrUH3Cq5iupUKRj0G1wpH4ujJsjco9HXMKVoUwZCjSPu8KpXNXcTfgG
URyT8BInaZ2Ei8BQk4GN6Du2MOZ7iEOHubSNf0wFeM0XJpS3bUyYj73TInWFQUl3
ERTGFnpfYGiRIk65TUvjlqIFO8KjfTPB/fcr0l9oLXBDZpX3hctl4NinFiLkoQrO
aAWiykcFsCr7+IUEShRPpEo1iBqxcmJrTtSflGRRnbm8o0nzzpDx/T6FHwQh3NZG
Y4Vieldtiyd33vIuqGeWQGFsqYm/DccJCLFGSCdKtKU6e6dSzQEz3iCaZkfVRIkS
hUrD5j+7Q5NK+z5dEQ3lW5/sWyQq61w8lFxE8za3EsLZxJZKVtVCLQC5Da92Zfah
s8UVQaQkt+lWK2cLI5BXuTDBiJNVEp8Scu4NsGlXmQP42P/Vr4glykO/0HUoXEbY
EHsh4TPuPWq8UmjVk/ngTVMkE+V2/R5/GWGDLFDMnB7dEhSHoN+r4yxS6JJiReRT
uKQNMRUlRH+m2BTImKU0Lnw0b0jVmFYafOyRJeGicjDwx/dwq0FXR4mnDsumhEfK
GEvUc2bgCKgE4pvQB9MOz0QAEA7cPfCtJ2yMGK2Ta7iAh7jRMvBHVMmHNPMp18n9
G7x1XLEjIOAhL9TXH4ozsLZPNOFzQkK0xYG9ksGmLsyFgiRseG5W9ZspEF/hJLgl
iOCpbdUy+pOXIP4ao55j7GzaG4qy/lGidJHad8p/lDX/a3mtATLqOeRpD7v+NBJl
6QD+bc5xFXk7ZPGTSU5DKbjxtGqqUPnL+jezhblkB4Hzz1dtoOFFbnk4QEEOqs5P
+cV2f1wzgc04toNQGO1NrXb9KLvnSCBokavQb99viGVhwf0pxCGMLKlwzGZWmzs1
Ya4VAlw85uiIrjr1rcu4GndI2RSvHl6qsQQybYYz//7xj8bVA2kbPz49ifyLN9/U
eBFpT4MBXVWXvk0O1fU4k3yUATuEh8uVXPlJ2aMmR9/JxXnZaqom2bZb0N2Y67xQ
tlHISzpZ3lMZ0oV7hePAXP6FInML2B5h+3TjsFMgufzLdxGWd2pP7gRj/Vzqr69y
XdD/iHpBTAT4mnUDM51Xze8prkEem5CZVrkIgWgsTH0lQ6IdkFGVt7+pMcKi6ROo
yLjPQFhEe02C0NFgIZfg+AbjYoKovSrNMlit5dCzON+R1/diJAGpTq4URJaY4Ww1
zlQD8J8JbMYZ63mjYtslrDuM9nrhuuX8sSbt++CStxHc/l6CORJnsZjEz4tANXQE
8yxa7wL2clcYGVjCDzHOSX0feCgbv2tf6RVGNgBgm/lXALAISUAiV9J7oxfV7Tvi
6hWEVR4SHRlYVqPm6bOJmv6zTqkkvovs+DiODCtk7eN7y1ZIdcZvBYWIO+cXw/Vg
BH1bjY5bC7iAfo4c2sYb6R+zfx9y2s54KOKDyM2urnzP7ebf/q0uv2FhruSzA5c0
+BVL67U25v8UUFtsdbpLaQ5fgE02/NcnYjYsEj7+xn5yyB0+9jeXMuOP1TELSVyp
wpDout0ih4wwEe8sQ2rDlsf4BNLHRbpNu1sQXXd/bFrZksleNq8lad8cnqYAQhnL
uw/SKTEJLlFraWQaTHbaGlUjeUxtyqkUZHf5DtpgmD2e3PWKm7LcB2PpKd8rCfGN
W1x6KqS/R4zYpKFjKApaU0zKvyEKs3FVwzQuT1yhrCG+N0G86flc28dlKxKvDPAB
28Ur/22rkDRPZELTjFvEGXc0cNMEyI+0FtKtrsnUtxCaEXaUxhkQBd8bY/Ypiw0f
0iS9h9ypuorwuuhaQUA+Qo4vtG/9knB4gWfqNdo70m63dHKnqZw7CGE3Gek4Z+Yv
l1IJLCefNW5/eez4V8BCTV7hDB/yZjAnA7qx65KU9BzVjk3nxl3rlMSdTC4NGVNU
6K9Q5oxyjEk6hW5qYpdz3orp34wA8jKrNRRkMMZzXR3cDLLLFtrNaczGgk6V/+LU
dDjCxaRZPZkHeH/wsiRs80amvkjHduP3INTYijvvzJpgAEvvbXR2qZ7e/MrTcZLX
s70sFSLvDgPpmd20m/tQx5qMQoVoX6HOwsFRXdjr3SNxyY8k/Tj+KZgvRP7bcfnD
dgOqNNxWobvKRxXKzZsaAjYcHNunR/cMRfVWeu7YAG6uTTmfe9IVFrbh/VTVaXaG
yYLqEF6Nu1Q+uEl9Nu5PmZ5ImEXmNKo+BMnWeCp+6eUhZ9tFmERyZDVeHh4/6hao
Gsmid3toAVlUbvAfJwJpLa28LJKjorGD64OGucyK+iSlLI/hq/Da5WN4Dg67qZVt
BZLyaLIv15OW2ms6GHF4tCVeTcD94mkkxlzYwYqytlEljiOXDGKTMShY1/gtEioU
nuQtcB6Que1BDbzNSbjZVuiCDplWjc0Yr/bCdyPMWtiUyFA0fFIsFrorq1Y8mVKo
zBxPPCHvmyNuMYWRo2QczZDTbbNXbtzCyCncSYX3h4x2qiQ3muvXy0ttsqwoanpf
czbpeckqZnx6+aBKSvQcQrtqJRoCCh+FNujm2MtVzyVAwYl8f+DoIEbzTKKzBbo+
UWDJl9fQBjm3LRO/PxkxPQdsXkfTrH/NYbdvfttxvteRwIRspkzKl6uoBC8JGqVA
c0oGMgEEOww2Qc2pkH+STsEQTlfJRE+v0tLG5wLNEpfQ8JKSFxh5U08C/2ArDKLS
huV6yPdC8ZUZMVj3mN9pbLv7Jg961EH+Zu/r73M3MbxIoJS4FFW24YMCQyM4SEnX
LgfTciTS+puwnhZhkVjYXv6H2ayc73AbQd2NU9mMDR5y+Kh9rtvqgr8vl3FvLjYP
f6qzUbprmUUUDtyxFKkRIa3eR7cpYZP8wT3AzIBncQiZ6MgY2pdjnlztTkwPbguU
QKHOct/UZlcA0MJ+tY6c4vj/pCJv1V8ZHZL+fLh2r9PYbnne1IXg0JSuwUbX6pm9
rcn4a5M/JCeR34GBTQgRb7emGRTTEQfrDfiL2bVb9MExClcrFAcD3B52bFFVOib2
U0p+PqBuS+0y0OUTMA2E8dl4tMEBMp2076icNdYkDbwvnIT9i/oR9sh5Z0MFBdSR
y+kUw7s1bE4eMvAwwqweRjk3JG3TPLC7HJE7N9pxFXek01v9hCq16NF0lUuMMueG
vViORfPRz+Un/CgHd4gv/ZVnXQjluCtJhkP4vxTJXE3OkdIWOUDDthe96R9L6AD3
3SXmcsqiLWzlz4U5ZYI4IJbZX2HmIbodezqrP0gjYfVoOXl8qc4QpjVmnScfP2jt
Svu6uFiJ0sLGgUaNGVESK9qeuuK49659tiyijynvMXdcLZDqkankmTMhPs7acvs1
hkBRiQbUFKNubrGoPkMJvJxA8hWsHaYtJabj5PdlfjWw1p0KLNkKgpBxgOlTX6pQ
H5wBeHOE9u/M0mbLmcuWN0Pf/33YkKQcxXGTNG9l5UBnmox1rhsaQ/LCe1sGt6so
EoZyCwafqxiPam+rN9KnKjZpUCv46baLnEDnBuXf1enmguFt9/4yo7ai8eKDYwM6
zZsadEjTy/NwI36HlyjwmOubLJ+BLKz4GvtmeNBBYGeFtS4oLT82KjvSSMzo/zqo
TBFIVvueIwkxWTBh/l7e437Mlaqa6RTFhWkNyzJ6DCJaq1ODwtte3jcwRhb3yGvA
Z/Z+RkMcDIEJ0g4KcNuFTVpGsyVfCVpNvTKz4GOeOuD+/eD59LhtHmaJMD7GGeBE
DqLZi9pwr5OLqbPbLAWJ1GZ17XnQBE2Sz2wXEk15GUbFxkno/9wR1RqOO5xtUON1
7kfVmuqPvypE0tCR6iV4PWAry10pJWWm24pbigseXxEROXp4MBCwvB6PjGcoxKhp
tIs4PH7NB8hCYk3IgTz75iszahNeDe3Gtv4h848qfFGRVzKhG57XyFCoT0q3Gy4u
0jw/LZYLQhLq0HciLbnLPae90MtZKx9KRRerz0C341F6PcAEtxYlx42I5EITmw+c
2fXgVTuuuPrZ62aer7e9DjMFQl1CoUKarA2rGUlWAoPRo64z5iYgyh5bxj2XEMYf
SWGMMFWIrUf+2WEcV4QhjQjNzI3nld5QV73csZp3gn1Fn3mDKOvHfMA9FZCKZx2q
6qwYxnBVeXH+wmTnG/KFBc9CSsRchaxlOkB0yLdeLJ3bpntoCZ6t/hRwUrvGt1yx
m/nI5j3iVEcpFw9lLhtjRiW/RJ1JBy5WxUYCYWkq8me9aXxO0dFgOI/3qGOp+3Pd
nbAcM9AyEA9iA/+j44xo40yARwLEbCSQ97Q9grukLovnRook5ToFdjbcJMaUF9zX
6icBNY+AW++qxHFKnbNYDOZ+xtU75GL35krVS3kSKp1A7M6spOwaHGx+u/fN4Bk0
xRz72bmZVuwhEVk1eRJlCilHjMQYfFwPFkT/Xevs83mOOos4h4C+i6s8S6k8Xcum
/3HfBAGeS12hMS6jDd9Gt/2E+DFYxAsx7l7YMKj6Qh0zVfnnwX6htgPtgiC9O1jD
U1z05Y1LTBCy3WS1LZ9Q3v0Q44Bu0s+ruhadn7yYuFjroqoTwtBM3u2G8Z7xWgZd
CuDEwra/yf75oOB7lyVCPBVvsfOsUX30tgFJ1763+tftoIHWHZBHouaESVb/Jv5F
ut1R8meKRPYs/LhFYDXI+eQYfWhZ7pzTyV2UY25mQ8o8gbcRfvpylaaaxIRTRmcJ
ZjCIpT9mEsAJOHdpJGVYBkj+Z/zS4PNbBpmz+RPz1HgxNe8E/1i9HSBuKWgRtxJ+
fn04LxVvM2tQFANf2iaI7i+2MzgzjWUtj96ZGbb/rUm2Majjbi79udGa/goU8fcz
DaEGgK+i7A1kiJkxKpYF0FC8I7PMJn3HPnd3n5NEzMElnjpqKuodsTNUM4esKp5V
jrPmzTDOlbF7ZZPPpkZOILfWVOSZx34Q1Hrl0IYbuXWXPOKYC5dPaEt91rclDc5m
S5ucRqQ0JJZlC1ss644jVT1T0yyKRNklZwoDmI3D3PzmuyOn5pjB/PibPO0K/Ios
j599n3iwx9D5fYW8B0X8U0gabdMcIeTrOqBH70+LeE6RM5NhlrfzEj8zTdTvSbNA
SQHnjPz4UVpcKPhUg1TWmRPTc9eiZqKyqjl6eWcY3YZpC3//MDJiWOpty2oewjkK
VS6FbR/QgW7cA2jhoR19wQFKaD2PRniCNhXCSBG5DqiBxDgyr5YQb1gwE01UBSGT
LXTkMVmTvXNotgZtzZBKackMuklcgvX9e0olQZJYFK7EhWDawvYgGrQnta0P2ZeU
vDjsXCW98vlrVNdGZHRTyB1FhbjtgdXBthJxivDOXUk9KARmrubxEh7ocPvix+Ow
kB6tsIycFPenIXwGhLUDNWYW2VkSaeZt4jGlGdz4t8NrjSzfmRoDJXD+ZQ4hDt79
DExpUmiPnatRcnUtecTMZtTv4xQ4QbrDusGfjA37l+22JqDm6G3lDlFS53q3/qFw
olFSG7VmIVj1ULJhQhc7jBDLpLQKf6oaye8c+d+r7G81x5u6tWPfMSLwqtVsfCcy
B5CDJtc34VPvBCjaHV2+0xLwWx5VanD1AQy+3ANOzpY3JLaTxdhysekgxTmMrJ9u
4ZuoGYeEdl3zrDMBVdn/j6yDbV8rQ+z0mKZmMNQv7DJPvIP2kH0vK/xgsNjOKhtU
K6uz7BoDl7AvdleOraEKkjY2ddrdgs+Xij4S4XCXf2gDwpFZG2cXx42fhf5RnpkI
4yn024rcrYWPiOaha8F7mTpqUzhFlWhv2JJKChLtZsavsfgFico9VQoL6VdT65sn
RUNzrMTgK351AR0JrNibo0QOOoffelHXDxU0yi9fZdIR9facKqUuTb1tIloKyOxL
QW6HFvAUk831OhHN+kk7kZJmdFaUPixSKdv5MeBokAbvtPOHpw3x6he6CifQo+2U
qDXuarp4mm7QQqpvUDPwnTG21ebcXISUJEO/MkDtQQQzWqjyneWB/LYdWJf4D+3F
A+mz7Cwzxxs7a16clbPyGAqY+pwKJ6UtUvGQvd8QXJbJWJt+528ENqhSPNjsI2W8
6DwwZUPNQbNSSdEnnTVps+3+xFuL7vtOCUQ1R5tI5SLoXFA1i9C2GbiIB4WPoH6N
GQsaZC8jFxMxMsuZDA2NiKQM3HbMsB0NeyTTno7dWXoVi/5HkKryFiH9egPqum1j
rQ7TvWSNsf69obaYShEo64wY2w/0S5ENcMzRiVqT2K0ZvDM8OoYdSA5flC3AWtMc
cAXAWgxXPHFy7GbN4q/TjJ5cKlljerNqSJHr/xE+r6gHjBOIW4kmetkGlus8xtwV
xgsuIVyoP3TR4LqPurjnnAxlpSE1LNfN3pbdFsyASlSuVHMc/cVjHr/OTiNP/m3Q
VFRWakXOrmo1R42oiZ7IHMSatWgOroOTI/Gz/LQpWXvt9a9WAI6cWRlyVo9IISIb
FjKhbYVRkKaWBmxBdYVv9jwgKP9ErWqGiJd/qaESM83LZtEBlFA5eKmLLgZ2YDtS
`pragma protect end_protected
