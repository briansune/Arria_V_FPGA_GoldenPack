// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:23:35 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jRJBqpOE1cC4CAdEP55dcJ44hgG937D58Or8tfb+v9vyE3E2iMKszaNc0U1Gbe1V
hMLeuhiA6u2ORTuztTIr6KX+wn8uIlfzLi7kBkaN2E+E6u42NIUf8zHLoUrT+rff
ZW9TuiTgM+fokqFU8ZUOWSJIZO7p2vGAvmNYnCIZ9KA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1488)
M+aE4gl3i+GJIpXTRuu46Tbxzb3DGrh/QAhGLZP3b2712polptsKKAFKzLloSZaa
Np2Y+EZfUecvFAt4APv2UrAlqx68ZcfFGNFLtEDqwjkDHw3NMcrKXywEbhTE+dYA
gLQ0E8stdmd9bf320z+3+qTLX5sTSE2zSkRWp1avqv5RzlMoWzcENZMKB70P9rSn
lgum9G3GqnP+k5qfI6+HnuVO1sKGDZUxkqbFami0VAgpNlxmLTZftA37TFGIyW79
tPbkoFUjlqNJnVRYJ9ksD/P9u6Ghb9knsZC4pGgv7A5chdmvIm/b/hDGImLWtOXm
9y/aCuhMgll+kQkmWRM7k9cpsYpBoFFBlWDjbV2lq2gWoksuZO0yvdnxi12/4pPn
tyiwbgO+Z8EABhwQ99eppnUrc890vQGa2irt8V0/iS0/K/UAZkRIds15fTOxTadW
ImyGBtSRmmaRBOvZ1NLiUkDo+e0wnhWys0Wz8Tfz2iyQxqdby9Sihwr8/EzJk2DT
txiBrVXx/qOgHPmb1dNB0IYOt+DxPT6Xy3lzyxWRuDHcTKiQyO7Xyq5K3jkgiqGu
lLrMILyfgnd7l/r6dwa+aihKXZrnSbT8BsdPrTA5WfiMHROeFJ9giY238sWJKjnW
QwDft+C8uyZt0016nFtCkHJPeIuvgmee21j94RfCUkYbi3qQjcjWXQO1gwOnRAam
N7fwAZWIpBqyACkNK6kq5jaGFGoueI9k7QkuNMVemM3YDJ4r/lpLqoOBmNx6RnET
BudxOLgofJC19flkAEF5hjPfkyw9/TdwNEz2geUHjRfKlP7mlciQvcIBn1RPKePU
CtXc1q+EeaBA6ZOIS7FfGxm/nrHeb+62q2CI2ue//w8hWHGjwGLkUMjjGli9N8d2
LB4lMzfPd/A60nJF8pZQyX9mWLs5EhVxLLnlHbWHOjEZTuhYXiZSYYw0fg4Q25El
9VH/STnyXlcmnIhjmiLcY3Um9LdkcL0G2vPE1XZcj6VVJQr65MSDli2b+YC8wJw5
rSM0IOL7nvnnULdZsX6BHXgxwIAM5HURfVLFyISuJBpZ+Xc8xdKudDz+GTpbNPBk
UdPTKYeyVMUZArhPABAbTazJ42l5tUYtUm627EY+qmZMJVAlFGvG7UTQ8O+otcVE
p2a6GQa4KMIbzDLdjt8a+rajg4rU76sRdONhyR4Za6y+r1imoPqfMyDgAXTC10ua
DFoMieybQ99vrQabqRlK/XsNiifimqg9cUH0fAMr3hOE90IbbKYDf8qenPI/HBKb
JItuwvXuLkplEvZV8NgDP0neLGCuR67iJeFZuahP5Q6Bk4+mqWNldMBCWldll1ij
eTB6aGK9w+6Oa01/zCCp0p5zVA2F3jlQS3a/TPi1MUI7sjhj+jdXa63kYZKxvd8p
rxtAa5TqoyyuoJLmN6eq7rnrNbhKGkhMmtJ35qi9Xxp/g+yTBEngHuyzHoQs0CsH
1DTBus36cH4FrKGtv5XmbQazFUMgVJ5VOI9WOrzhevAeCli1obiBzjV0kdnE1mld
7qY3zZgBVpD/kO2gPz1/swzKq8NcNx+72DvG/UourHiPB3KIi19cUXLUTJ7OSlD6
diD/n+zyAvCOoLU7gsu45VsnEzLF4RHDvDc8VJwKfuvcmbHTB21ADz9d67iPw9ST
csSYyiHgfyh5B00yvnKHDHYqNOLdDF2nZTeaGq9amk+XG88XVwAoH0da29SRz5z1
lADlU2UoVhfKSgVukIDIGGdLpJ+ZHFTjivyxrP+92kScASeGB+gvTdSv/Ze+ki3S
8NGMhCqboMMHxSjUOttYwzasoo+eBgxL1/ND47BB6R0J2fOA+mS2IClqYPwTgb5y
6+atN1WD58Jk1EeBQWpsm7I6MUSVtvUnnLJ1tjAcJulkCTTd5lVdOiTqg7CGsqW3
m6ancw1UJJA+AB/dKnqSdyjZH+75nnxT87jlxAn3P17PpsOayOdst5R+8RkQFSEN
`pragma protect end_protected
