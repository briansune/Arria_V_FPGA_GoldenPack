// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:26:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fuYPLV70hNGWx1IbWiK2vcJypefzfzn19YvWNo+JC5tCDltS2zo20C12W0PXSVtq
SIekMCsx0POckBFApo2SK0liif0IVWCHsTOD9gQAYHkQbr8DGUioh5H6LobUN41V
x2JEwEsoOQ8rq6RDCXw82vYxRl4V4Rca0ptwj3br2lQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5552)
LFpSNmAALnDhBlvxzXu5Zm0TlZ8w+2ZZwxLssBhnBZiY8v89ilggJoIevIm7zXZH
8fycP+hva62Ulb3X9WEyvadUlYHYhhFicffb8NE+Y5pPDEmh/x3wvB7dT0+ZD/nm
kj2cxD4UJwE5H7Xo2swAUCkIhpGBDLoiJOHpbQjVPwAbL2BI8fBTgFZ9T4VbMswb
xHK7zucSTTgmZj7H8D6KiLBU3PWAVqt9ARAzG5e4CWGo2qpgZig/9y6QA+61VM0d
ex9rm1mZlPioMjAGiM1rHnFCT9K6H0vRKMbpWOW3zKATI56yXXDLNCqG2Htp77Rk
iXEDyfPtbKoR2VooAjjRUDcDPshu7VNMlHA7M2CgOCBO0OWLMNmIeJqwXbo36KaB
8/Z1E0OuDkut7q12wq5dd5GaIbmJ5xdXjnoccp77QW6eCKHeRsZpQaA/8zSpJp8L
tV4f3OT0tm78hyu1OQGfF/0SAVTRfRWaBHR/EERhI6CWOPPEywwh9rIUOV07VVXi
xztGYxwi4q05xOD371aKDMNSWhPfiBCvm6bnKqe/p0qtpmSU5FetHbPqIIFEr2rH
dcM69X1y6boi/H2j+ut8JCLU18fdx1BbLqynRMzJzqfM9xWwgJFR7Dr0L5UvD357
uaRnLpU5IzQzRM1pFekmir3YVRb0xkJ+OfFypzRgduKMwsarwQ7JYpuxHZFyTgnX
iMf7g2wiSnExJWvrOoLjmyJxQUmWUQ2YTXyGhSCr3OeEZyR6Umu0dDfVV9ZiBOcj
CFOOzTjgtzvuYSym6/zKE8ed0nhOx3iJwhRiN5iUVvLnFLLDsA+puunjsQkWp1Jt
G2y8VW4LfzSB03EvK5YCNan1VJ2uxG8eHxl9/4sO+8JiZsNGQJoMs7+z+e8HsLPm
kvWXVHNJY3Qa6OX/DjexxKPhRBKsKSrGhUchywJr/3zTd7KH9ZwFvOQWpmfYM5vm
cfJdsGooPBod9MZgWOpFfRhzZd32zGqQfjzlKFfxpZv8Ylj5Yba2cyoCFElbjfwy
v/ZUzMTy1tXtc9ppA0byxwy+ZdWpjoC65zY8iI8eCLTVki6xogQKQIP+vEqB5XFb
q23WKu0dkr01c+hDqYoRnKqsQ5PZcHqxTqfyCp4XnmfPovlIYhgcJAYkx328uyPJ
vGR1CD2AbreBOP1MC4w+3BhaG870Bf4KSh15TM3RLsidWAFAmy7MAEVaCe8BObGa
yjA4dSur54uGPq3Lryl2dcq3WCejR/i9ztfC/THIfOFxnK/EfX9zwPUDOH/Qmq9A
Mxp2dBtoLeJb6jMS/Ie6sXXt2lLNeDvClh94HDEh85JiXId59WNj/O/X1HG3yH/D
XMahuWtaVwijDsrUh5jJyqO0N1k4xuiQAw64e1sS6mYKj2ygFPXAm5ueKcGqeZux
Omkr7AtAyuDnDRwXg2uUNlymrzQz5Sxg7qUNG4neIovM8o98E9TJVOyPo0zGRzE/
43vRocjbAan8SwFO5pPQQNZCUhi/A8rDV7sE9x225YIZthu/T50963b1lbF6A2bm
awgr3AtqMLtNEssYd56YSiv7fl50aBVLKANY3nc4jZMxoFBQM6lDiZ2YOCLa+qM2
V7gU5Hq1ovRTwUbL+MTORFq1GQQYw4ikS1YSod9lvaKv9wdo85E0b/8uLIVQOeWx
AljaHHox0/yx4CTjvCqQvu7Ad1ocUNgOltgUf7gCyC/l4aK/gP28rTydZ/7JlY4n
fik7cQACjYfgYRZnyDBCqCm7NLJW/E8GuctbWzH4TW8fh3DXa3AEY4lysA57tiUt
7M5Ekb2LBNDXhpUiu3OdXvTekJa3nLS9+cpopA8Nvoe8G8wzX88kzkiwN/PcA1SS
xwSRWfIkr5usc5Sp4LHoft3rwBtOmT3xaU/qO1h1ycFWw76qSbU6rii611ZWIjwE
ZnhZDBvP2ms64MXmamoeKotiT/ETEGvB7f09vYfoD99WykA6rw9t2xgdvBB+lbv/
T/BQtTB0cY44gq8qv8jFCew3OlfZmIoSQxBDUq7CHkBkEv3n/j3U0HjpzaxrMi6n
G/8PegI0QBKp6HHVeCQLcU0pMVlmpzXnRZhI4GyHS1aIlXh/wF0FT+A2uuMOIgsO
/qo0pRstjKYF9tFpmhieEIQeTBp+N6oZe61OUyWzP/AS8S5mN6f2Tk/IBLKjxg6c
bP5dQEieMWzTB0ba3kK8GEVB84ZRlpG3SqX1fPsV7SZNVK6Z2l6EO6pciYR3H6Re
UxrnFTxpNdk+1S26wA9H0oip+hLDxsoaN49S5AmIeeKgPq+KPuEUGc7T7hB71M68
S/WGg9qbBQbFR1Ffz+zpEZSgwDMp6lT0UIPrUUOQhuhN88Q6J9BPPBzMOuBBGLYX
mhMo6fQBydrsRFy1mKLibE/g1ch/s6s4ALCQ9FMSJ7mD6Lsoh88e2fyUR0N+F/Ig
LXkLzyzyJEkHLrxeLlptO0eCAzb6irSmQVmo4jsBbgLLpFmpC0MJ30ItbgJY6S/q
HIZB0f2IlZqoDejXTht/IDFBurJjLfnGbcnH1PBmoYkMu218p5l0kpbknwqsJ7vV
zxPlvdKkUUs8+4dmTFYiAJ9lNKlv4VGq+vvpIm/WcorlVpWcX/dX3i+EnIaCp3/B
GjDKoVUVVRI9PNqQdwPR34CVURhXMqg0VAdLwzyXsLPsaFNYfqKI5uCVcEi4VBM9
LZceN6DNlNE5w34Vu7dVkNyqHs4tLqnfvQcFPpXN70k9GBtzlORU7hincSizgeeD
7MD1oxqSo2EBVc8m4NLOMpkJkR/pUkiMbc8qfiaULSaWGl54BS+789zxFcxONfoL
uEGPWE0pvOMCB/ZmYQKyD8gskSLVFZ3iE3U3odYbU+A0j/4M4wnCJM5jGYNpqP+6
GYMWL1N7AoMh91802vjNnB5+IywCvdqSnDtp1+5hwdMXzpbSaGLEB6y1sg/5Gmbn
0gIhiAQ7H1s0ibsxFk4r+4xUOAqdlAKSEAnnzn9hzywZ+KrpMbKos4wNdX0KLsJ6
u5voCacWjNjf6pU5yueH3PkhJ0KpD6xzMh9RCjnDsH3WzUf/wuhXoD0/iPyCmU2P
bvhYJgmdzuYKPWJ9AT0ABVvftXvMR0Rv/iBC/w45UMup/312abTigpoeoeSTXhOG
EOgZwqikIcuIytdFLVLnnbyQ7fglr/Yf0KI/eVkM/k8pvMxEuWNdubDjZuoHSDJx
Im2l9pIrV3LwnLxIUqrovl7uxYfxXmUudvV177EJgJaxeMJWhSqEXb7NpcliPdNa
Bgl4nOlYdmYJm5eLbKYzeJPsXQHy2e0dWesWNYDp78SxnmEp4y3h8VrtNHafmPla
TRyKSDo7MGE6PoD6gXX8I8TUOj1uxJTwOZr7FREPs4fCqeeMhj18v3oPgU82imM2
VuRlf6WZzd+lmW/abWXs1jnFwAg+CGEQ6KUzy4sh6xDM5E83XHqB+STwfdwy8KV5
IQI+Ur8I0kdRMLaVK5mD0McqYsWDcS1sb/4aWemr5k3vCKCF2FyLymKEqtcNd5Qt
18/GEK068TauEpT33DqUUDLmrZQrHRPOF3Dt2BzO6GNbYyErb5rqg9zbtJ1D51fb
8Xctq803c4AHNgh60Brx9uHEhso9+oOBsmtf6SKEaNi1198kdRA+uCktELgWJmAY
zPN7YHYGNPP/pCj36T5iftxO0XGZ4OxyTsKjJmorv/NRUIe9NtGk8E+FU8R3D3pF
Q5zzi+uGokNRH1Z/jKhVVht+BXotykeusNFQO4u/fcx4XmlLw+8oZisCT8VRu/uV
C+t4YTG89+mW3PfWbVPDd5/EiPNgOHWqPZbnibm2KialNjqX9+Z7bRiiV2sI+t8w
dGiD1MKuGnvR4k4jxz3C1wFHbzBAQ7ytz98MZRogqjtlYcJd7RimtwJA5DfzCwFH
dUKsoftbUB+Thlnq9cAhqCJ1/46TcfxXIk7zzvJkCl0iaISvxgtX3IHNueo/XDGW
WnoVNLFjN0bU0HMSnKQ5n8YpUqUGmd3iPHqcnL62YQVDBrrZ5UFx8DN7RpO0Ac2t
+KLJbkQpPxTT+CEtu9/W84BNFclQIpAqbipNnSYlRaGCZ8ygm0RzPIsCBBgohHX+
w+FuM5+2rkGyhujkq7WloXj/ruKyIb6VpMV0ML1PkBQ9meISioPwCimRRWQ1tDZo
+FZWG2nT8WKoIPdvJUgk9KMVr76YgH2ZpnWkubTaWxRrdnX0gbTXzoGcxx2UU22+
cKYqpzymcqV+cuiLIdxNG/FrtcGlg44jV7pjPYSp7oBdGvIz9mEPmT0IWXa+eDUX
pQsvqV+Yz/ZU6TQDHzH9yQmJGV4Unao8Yq8H97MXMj58M0C2f9ft+p8ZWUtprMjI
2s0jHNhJDRMUBZulupceaXIKMpRr0fOnlRoRREofhiJozg0VsvWO73faQ5063Rzi
dpo2Udl1leJ3R5UmcagfIL+175ymi0ad0PvqdMOk9yuJYZe9/o2TpoXMKVrRT+Y3
yeYRQ095DFpLuoEczrPAImYnABd+S/BfMvuxld+TY3m93/H/xAaaciWcYWnee6Id
AjuX8oYViWYQQlO6BtCGRBaAMwvgEl3ONU4gdBQt15ZhNj8gVIE8TcTKvyMcTMJW
ihPHIwMQNp1GPtMkiOY/pKO2MDrmYBRsKAlQdOkasN//av2P1cst/VVHqlQdc7cq
x1leS50y+M7O2NLRXgpyfmgwJPS+C5Tk4hYAYV8ivNCTjsg1+a2QSp2VYTZo90UW
JYcNNkwmB3EQcAzbDossYDJn3u4SoVw3lRj5nZo6xNnAgQwodXtnrb/YA0pteVo6
U9dQSQMaPI9KnhWdWonLvspQhKVCJ0kjwf/sMybIgw0obwJvToWZksjAz659d9Qq
I6cfx8hofnm+9YJ8BHqURtUqunf0+wBR5AL9L8dkAfFdOHLduJU+nnmnnT9ihmRG
AisTtInOmpH8wdupRt12R19AWFD25FJF7F06SC7k85cBBSrwiO8t3FEISGXaxWMU
Kbj07ckeue16uB7avPrXlYlSBnSGepkxJAHLejG0/NZjpnEetsNc5KaIbGdwTnox
mGw7mpwSbAxwMGHDS9S+BMLRYFxz56t6/wyBd1Rs7KkDknvMbWkcOK8KFKNVaPdC
q8jz8WA6CZHrOc007Ek7pqDUcdMgHQx2YRAzdn1UfdBpNszwqqTfdXg5pSrvVDPv
CJyjoMqK9m079vhz3rgpY4BfjjmzI+baOcfFTsrO7EQME8GcPYWvsJ47VBH4hjN+
UG2g+9ymvJ+ihkitsVZui3MkI3tM1DUwl+bYEStPGBWsWrD7w+FLSGSEfNJzxU5b
Grxc7J4o/ZcqVdxzANVidbsUGP8YfShLdDJ45TEGSdDTd8IzXgYVlyeLto1NAoCc
l3H8fN4XNJt0uwby7AgeRWdeMUb9Z3ljUzZKSWEiDfMml/Z88dypY8mJQLqEEKRW
XQZtChOcHOyZ+mPimLGcpGcfT7Ww4oftilmd2lmsVSiJL4hLGPkvquDSuzeTHjyR
iAZ3nwd8BxxaFcuvOfKycUA/BU9hcl2X3/rwAfCfrlBQ1PqsmGZ0Ul/kZUPaH/VH
GKALiQzDdwI8D3FM3fiRDq7ISvYbWavKl+zfkJmG7RrMfUXzMzmGzkl5t9ArP18c
+0KMmMSBUpq/+/UM96FtDeL+o2JVd3yzS1V/OyhNE62NOy2xYT2m5Uo9nHJsKc8E
oLt6QKxRn2yfrEGt7UeD+Aa/XRN1clYzrEB/+DN2/kyq170sLh0QsrLsNrjD46CJ
ulhzMa5RoWJxkAEsHEu6G9qvDwDS+cV1BQGn9cAy6GVLD6Mww8cE1XAANpjW4bI0
pD/CjU3ZSMGAMbQwhb9fmQW+oh5wnsm68sA4DJFRWtz36M7Uvg+Nkh++3CZmWuxL
U1LnXTXyaK4KOsasVGYJu9krFDmAWPwZHAPaz2yTprlO0pLJ0aOHwFJa7HcIIUWq
dfVCXwk6V/3PiKIwgfZkVjctm2xYWNzmygYHnOA1w7LUdK4UDtM0V4GdtqRmtS3N
M2NDLmuPxsmVqkRXoNLGvS7I4557tEzaUNwhxQa/B0TTlqjL4Kfas4pJJk42bgYr
Z9a33XbE1Cwkvp1zQ9P7Qy3W/cAfAwT6WPuGI3ylCs8uAERhE48JTpU9sVvr9TvF
s9Ap00YsTxo2JCarzuVpjn+7tmk+1r0M6oPAs8BoVsHzQ3d1xdpukrouFrvTVkOZ
4e+9WS97jkZpU4ueqb3XrFWt7Cd7HSw902S0kh2YizaNsoF7BIgOCzg/P/+DKUmh
zELIZzc93kdVyr8Bfj9BAM3nuJkssbjMPFeFdsTIOt2FmBwNy0/fXoKmZv7vGm/O
URdh15hnjrJynRb8g19XE+HvhiF8Z0keKb0nw5Es2GzZOhJdt9kg/IN8pse37Ngt
eEKw5U+5mDCNDKtv9s71S08OiC5BZxXaODSYHHZ1evW8s+0c/aaT0bGSkmgkltTN
kH2PjqqxWh/hZSxBXmzCqRoxh2+7YuXcrmdA94ILXlTtMS/n8b1Kqrp7M1RHq/BP
D9z+I2wDFEhv4ReNkfNF/3H4TzjSUvGEzm0fEaljSa9xyejKNG6JUEDAgVd4Y2V4
7mCC0SHxpBVTTvLSSr92jhlEBoxZKyx+LQv0jjJZCtVvUWkVBJt0QPW3J84f9U2O
b6eHlzMWzfm5qgskaFjEdxN+3790mErWBJZp3Kj0dCQ1ju2g/8bAuKWI/jwqbL2i
VmhkrVZs2OXjX0fksXKuv1sAqNhb7jTLUUcVdiJvs1MyEqvHg+dO0m0DTgcpX/mr
geUV9jKxNQPoLDlp348wV36e1Yn0BtK0NKNIvUPEA0rnKW+czNxcTjgWSo1MDZp8
PQxQiksb587odKfyXz2eTbrCx5sxTe8QNXAGeRD4LTrrgWJNpArEJMH6seSdsQD7
q41RqSQoelTfpZxH/78mPuq29QldvAe0FwxHWce8WRvuGvO+UhCnqRnGcxkby9Z4
EIInIwNi937yaPHZ0qysoJ5PufDY9wPL5ss8ouUSGknqDlpGK5Za+SZbQA9oiCN4
5Kzisiqt26D4gNKG1gXMaExH8ulOaIa5MtBLhoJ9tCUVZ00+HP4mTem357TItPh9
sT/UqTqQB8mXT40xo03CH8d4cqkBx7IJhX/3YYpWKpE2TUgenag1rdYv4fQjayZo
a/s4DggR+Ok5o7tCzSsnwanirCmtDbOPIO7ZAT/mfDrIGGrqFDIX8xwY1FJPTiqc
BzTarPB/bpYmUDU6MqvaJWhUmP9FhJL5WV7PDkNhGpwo37WtKGPfEwqWKVaP20VP
y8zKBt0FvyW+XGWiCZRV+fwhlflsZi5AcNy6o81Oirv4F598aQ/KjmTgVGs9sfGA
T5vv/Ba2vlRvIRYVU4PBLtL1BVlLpl1FHNmoQWvXyv8=
`pragma protect end_protected
