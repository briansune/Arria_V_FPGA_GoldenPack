// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:27 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fPz8+NOk4q6nm0EMpNwJeGiGIAy/DcROHs0ku0bK7h6qBhurQt2TcTVUpBAk6spj
BMwloSCqFJqJVFpTm1Y8h4o2eLMgckSaOr/muVXU/hNNAIBpu4+yerISarEs8Ix0
r87+gNw7jUsoIyK0VmNSsbdK1isXI+TszfnY+bVXFU8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11632)
j6FcUk5ZPSnxcx2JkLxFZgvI5LfQm4+UAjHeDlor2/N6dDNfxsZzU9GQu1QMfTAQ
JVNiQ6Ls/gcwTMoiHn4lr5oY4z9GjOIH2eooPqvuo3GNx389UO1Erb+wo/4xbmai
TFmffLZpUXcgKetJPqa410fdSwun9GQ37gtj33ibtrCR35U1xUln4AY0YQ5fXleP
pl/f30WFt+R3UrDaA6/iN5gDzTxvqtsP23ZAA3iIM3xxNigDFdqrk6cj+a99s6zM
8I/oxHrYVmeXRIlxLUU5u1bOJbNAPoiEq/pAtC2C7QCaY6AIKHtw2UGDV060qcbM
M0rPgw4+gG0ITlDzP06YMIb30W+q3PLeW+AiW48AKg58P7e7fIqSVRFs+drDcnfq
LrVGMLWwH2Ty4zsZ92UQdtYWuL+46WF+3iMtDCO0r1vn231sOix4Zd/aRJxEDEj8
rgQfZr93SDyaCjuYueLaKkAv6ml/N9fE7t7Bs0XNpgRzbWDksIE/Nlv/lDoAnOkE
LNkOwV1Gg1NUbGyyTCc/3jC4/F38eKMFdD/LTLK50XThIHwEXMJFPhZIpDY77GxN
zFNNvH1fTEB9HbwnluKw6o/2xEoBZDzJ3B2iil/yXZz8vrOn5uP1FfU5n/eCSmk8
mvVUNS0jErp/P7+I+QrJW8QeDcW0SOsRuasFBc7u5ryVnmiI8PQJTfSZFeOSy0MT
/8jkp3SqamJ+us0U4RUOqrXSKW5gCE6tv46PSSjkSBdEwBeQO46NR4/ltM5yNwAu
lv/C2O9uFyC1cj/zejbo+DBj8YFcCAe2C2+wsGKSEEHq6HyrtaSpHmEeifDQTIhr
BaGMgf6TAsVGheFvdotYOCJ4KD24YJ4wBczqLQGNVCYeRcLkgzE9FqiG4TIan3oF
ZXg66tXZmnWqT3FGOj++aKiPDnBL4UoqYhOcWaqhfSiN6xHeNuNT8R4ksgmwiDOs
1F0pEYdT13xV6A2ErkuauWws8eVYSxyqZzyRngazTbbRaHNNSClEFY7uLCi+rJ0R
/dGzaWwzv50uUucdEHnEN+RvQLpQe6JDEmWnrac9+4Die4OpvEfyWFbYXvVC9r+D
KQlUN3Df3w1zNO3bJLmWoFIDperisNhNBVPMmV6JTaoXclrDIykR7EnJKr0IHeuQ
6tNqljS10qIbsCg9krhsv5nRj+zQ/yiI+lsPTzY6N4Z9rNbbaG6JcbzkYiv7aqI/
jwTZZGaBbK7zCiZwoFufWQ2V1ZGaXdceCejERG/v5iEH7Nae3/0BceXugYwXJ7um
Vc+1kjwXKLEFRF8G05OpvNb5Q+nPlgTATGjWmC5Z17fWvMLTNJfmiZCwKVzQ2+QF
lD87shPPNcNAePTAlqbFJ/Geml5lmGFHrshdz5C3u2ROuy1BP3SsR4SL45CvSv8a
meqIdXtM3oOxz7R3E42SO+Vm6GbN5I3uTIUXw9YNl1QASwAKDzh41olokP6LnuIF
iAE9TFH6x5fdU0E5m8anHvXiorwPmsdqXMKVIHdBlFvr4vAihhMa9rjVFil9J89U
qmcpn8U/r5XC+pwvhn8KZ1sVCuOqlk9jhaKDvu3c1u80wBs0lV3haXipnN5azkh4
HQ3IuSaeeachnnYrhtaSp0r66rj9VfORVYhWFXC4ozpSXy+HieM6CqK9zDDd8Omk
bKyUpHrO3AZTKmKG5PKaHqojJl7sAPTTpBZX0h6CweMbxc0lE6VaP6M8kmkUOoI7
CPWSKEhIoOp+Q9F5efGBn4FWFCHIQOvqSEK1ywOEHVFSdh7aJlFnzA9F+mY/+66y
Q3S1kMp8Nb2fRn/E3wwazBJ/RUoqNrvdHfeePHSsR1I/+bGSpQrRx8IwVmqV6n+E
57a2nSoW78LxHzuj0wVaMtb4AD5z6Fm1ACuUldgliP0m/Avf7kpetcg9xlqBHKan
pbXGWIbEzWjYXSJRHYiJ9v4IQpWsgglR4WkDL7+941dfXTRbN/nkXjI3ES+eVSGP
Goq4e3Fq23rdDgYiKLBUKITyaJFFAkhI69JIedRYaVAa5aphFySE7rYegmcC6t6O
7Eal5CrwYnKErwsSqYnqpbn1Pz+N5DAa91+Bg6hDaJCyNX846ck2DwYkdeQnUvWZ
wI/aHOaKDkQ6nzw2ze0vV6awI5glO2NOwVc1f7gRMBZjnCTE8i34dhyvgrGElp9f
fEL/45Rhxn2f/ojeg5nnyFf/g1gI6l7capClDr+Qe+ksJlgOIm/X/0QPILg4YcBC
hD1UgtKYrlUa6QpVfA+7b+yIE6QN4ARt5C5pfqm/qQRxl56gvD4PPMgdYkKAOfzF
FJOEPi1GxxtRiQOO5fLk/0XxbdwHDSFVSjjA24YGS0uigi71qprmLj6gd7/lUj5+
uH7P42+kIvvtRpeGnSOZFrb4PtYKA5gpsjU3AYPJlZNNIHXAs5NDaCMZmgoygOVf
qzEdOzp7cFSoKz5EDfwVi477V/GznLuT8m1RKuXSEP3GGnKn63ub5+RBlu7dTwqN
YD+HcyzqMHtyz36FWyCd8DfQb03Vi6gFXHer673UkTWFXmVoFHki3nSiT0codf6j
aKY3PKbXIgp6n0TpHxqMx2fpUaRKRKBjGtrwf7Nq2MNEf7eVyIvqJOdcVCxCMd7v
NiwVmPsjdVWmCUb02m3Yp+4TP4+14qJijTGhoSE8sAbNxSHvmBktHLpp0xPHr+h5
dad6mdfG1CT4fluoCbbS9TwoHbqApPFp77K0RqfwBQIZPWTdhoc3Vx9e4t7dQEHT
/RadpTTKAEOERfV4iCRr/ZXRtA6n/xWqht72yxPeGG2lvIVb1BxPLntfD71odFSc
jTLmtqhuCohguqFdALOYHIlFNBKZWda4D0g0h3lDgDejzq7YZTvsR91mMK3/EyOW
JaNEnexArmRZBuZWTHoYfTL0qBtC7h1qIAoU9No6KWr5/wLCtbo8vvNExHiMqkZ3
J3/YGygTLzMijmqqJ1TsoLIY/5JAPjQb7UlAO6OA3t9byRxWtECZlwdpDMoR2I30
YD9DbK2wT2UUyu7rp4DWoxAVo04DxouzHQEQF8pRXS92r93RE3hIQd2z5e1kdVCG
5WVGLn7aIWDNHysM4ruWLgYzabYve5ntCZxZfxUcJyVQFIOXuzfUG0XWNKL4YDij
LjCj7uZRLltn0jr04g8vBymfHt+XaEHoPiAsBir+ViG8CAji+9faVjhI0mhyCUWB
g+3QIVZSVxGVhaOxfSjlWWQHup1uT9n68gCNC7DsTmw/L0WzHY7QXMcEdoHyhtsG
/ZJDPUN1sjUI3TtSLDE5wq7yUrTohfd8WBtHBCm1FtZJ6pMHkPxtDB7Lnro8YQ4m
MpW7GuqUd2pT1y7B6gFYvquPuiBvJeq9h1EdpXRpquItxJzCr4Nn+3J8bZ57yaDu
gy7dt/YN1w/e+TBiaPXK0OI1SJgXIObNayOBsNatSlntXKAlKYs3FTaEX2mcB6aE
ho32MtGndALC1cQhdGGUewqczwJWTnHiTSd7FVIleoels0FXXJojn0G33YeQiw8P
oKxSsjzkdvVGs24zc6c3x/AOmuzxOihcLkKbcDtRjEhJR8LNxD3I4P/uX6sXzEf3
t9dd4/KBuEC3wKWKgpNvQjhHzRf0LS8bczob8diyQPdu4rAWLBKnU0gN5lwqId1P
1lhvOjRXU9rizrv1BLbKtTG88csIGbdyjOpnnvoZGYERxzEIvA/APRPPBuOcCcMG
eYaDhLvdtF2wnE6UXj1WWkADDy9H649pgCk4tNmhVxqmg8b6HCwi61px6PkXRuzn
V7kd0Rx9RVqyDK8D2P7TM8z+4TAd3hXy3xeXWJZwhHV+Qzfe1Mf3fY4b5lKjbEBr
ldWo0cRc+k1wlXI2PxO1cfokGcXOVsWAIGtDQsxQmXUlSVQcZ6tTO4nvjWVYT8eu
TN9ZddtvZDTsbwOIA/6QApfThKDfLzOEp9Vk5qlPSP7ZqXLF/vZu+Ms8Fux3WeUv
MpkzdobYtz/wVmPL4XcSAiRX54lRRIYbJhVkQxMliw+gOv7XF4nVU+b9iOzjNvKo
w30o6KAVYINSjcVpWEoq6oatsExjL0CCh3GUCdYpWsfNvUBzy1L7ddJw7jnIcBtr
WPuK8fcm7syuUnVjkv19NFguHo5LUTTdsu+cgLnfqDrDp3xik0LwqjO4cZ21bOkJ
NvUcDvtHI1mi6Q+nDLH5itgah6if0Wuau0siGQVzAA51fUpWm+312d9f9RRZ8Dhw
BcSYcsZ6d2ZIujJCjHXir05kYSmTwsRTEJQmXZr+pAnC8v8S+SY5miCRl84ixW5B
uXSnvuJtToAat33UbGKkvDQa04cdYH8H7e1i20KdmpGo+X5Sm1IXhUZhEDPeApwV
wcfjJ1WV6Yl8Vt7Kq0hxHjy+guKDIO+hprSX3ascHi4XWvU3CtvIuA9QOP3zK1uR
Zi/JdJdJmAIskrbJ80Xu3ikkevO74cUpQtH1AoDOQC3zXPsvrkUFHo7fPlOZVJHX
SFCm+ndhB+pYci22YaOKoLY2LwBS+obah+/jbcgT6R+PMfUNR/O4a5tfDFY6nvqx
Imxj62bIKdJiZzuL2k8HFJ8aQcqWTHpoy2h1n3d60odv2LHjKRSl1jmN5j4QDDPv
JLmQRjaET2S5BYXGq6EFrPfUEjXadO5BkDgvcQJmfIj7hNp2jI/i/1jeaps1aO4D
mmek/v/nLR0uWtkUqwUbLt1nDGgLcIJTcLCQofWg2ra/HzHFLNGeYCSI6GnOXXmp
aPuAk0hVOdex7PbCZQQc9EhupPStCZtAAsvhWRerb4+kaSzlK45BY5TFrgPTnK4H
8DScTWMqcNhNKNnZK+bVXaE4tFbW3mbE84qSU4tAl6pdwOp+XGu7QfTme8X1Zlvh
+X8XvtVUgu/Tu6+M3pVuosSLxUIi3wK8wZo0W0bPAc/ns31mPjKqkf8UKb34v8Ht
2dH2sDPHcC89gyzbLSxf7ZALBRjdljDECN8MPkcNQ7E7Ix6pNN587krhygOREPks
3IU6SaSHkD/NcF4R9/l5FvUl5v9efmznF1q7qEt5+ZDImWhv0fhmCEl7bsr+IrFA
VqCO6+Jc8lhq6qiZ/1Calg64FUs4Ra58AUJKMC7LuJm3YWHrZPoyhJkaQ/osBR5N
6s4H2+77qk5H4Kw06ygrhTBwdV17Ph1b+nLc1m+wT1jSoOqxR2rdlG9b9VLB8QIK
5ih4pdUI7rGkChXL82uRmKalmQTW305Jc0QWF1v4G9cw4ehBYCss9HiDp09CuffU
sVYhSYxErL8Gpt2IHwZK9b3j0izeMXRRMnsXdXq8lqG0L0GO7c2gx6AzfkZPDWrJ
WTIWEAg/q+9pRqpdX0jpxwOipFWFe2aAgF8UDmQLL+td79eH3ZB7Dtp+XkeUGo0V
fUE6iYTulvlA3bzih2DmDnW3TU6OypkeKj6vs2ToE5J0yu+RM4ZCt7MLtVAGTwpf
aIdSVGL+EjQEUMw9gJGappTdd47/tkrJWlqyGspSWL8Xk7JhjUDRIbZpazsMHuN0
VnIOR10+rQBIrffULHwpuVAIwGJHgA61U58U7mWgLMeYEEOwzentz1uAbxmks6WB
O7lTQDbaOVrkA/6GBuvsEcJohOdfox+VjUkU93ZtjcMAm6+dKLYTRJLGCuFN2rp/
H47ylj7YHGHEK2Mc3UgbeCqH6R38xL0k8gf0TiHtzy9fwclFs94qmPSlnisLN20H
Yu6KUeP+kq/M7OlS2yTbMfzb+3pkKQ4qJgjSrY5x1Uoj/ATCfTMpD1MOfzZiyRqO
9WynRTa0mCNQzNogImM0YK5aQzH730i6IxV4WDutNpIUgW39Q8mWm/Bz3quaFIwE
Njw5SHgLTz+BEwVfp+xbS9xiKPIHIgaeeKIAKwz9cqFfmLDQ2oVShjdbGpcwJDCs
utUakguE/fMIgIbpTY0XY+vYaP+H1GilnkCSBJCVYdgaw/NBkuTtYvrWYM8os703
t6WQLe9CNiB2DRAQAqltO3ErK0r07Jz2uD/wa5fGfXvcda4eWztBWf6ACBhqMa2D
65R5hiX1RIDdBKQlNmFtSnlWCyUvV7JPCm3jUbCy2jiCcvNPfRcmYcTJdow73Doe
UIXzXTRKX8d9rM0w6PB705tnKTxWlrQ0vSX7n9fCGike6JEUCkTZHiyqQULQtbbs
X7+TmQJmkBUkZph/iSz08apZBkEalz4fsfH6a0W2dVIhjHq5vge4zox4XP7hIOQN
MgtpaXaSVmJSmHSDq4yaulmZCxaHYyqB0OCU7M0qE2rQKiE1SQfA/R1shSLoUk4b
8ZSzdfY5OD5bc0Z7vIW0HKGwMFKNQYr6ZL1CuTBOhHUc1bk4YzdJr51gGHsuNKpN
p3JqPYdcNr/zaK662jtnO4J8wg9IMrmFwRqz9oxq3H0aaYEE3ZshoY6YIkWLKc7a
CXyhsmOmJm2gDjTVTU22fJcvd4Vgym7qhHXyHwLYU3rR5E3rc8MGxHeZDsLSGZQp
HRVf4JEOnWvuXhd5yAP3iMjqjnoCPdJ8+nrVTBkkzOkuoxFwiEFOBPHjwlZ60vSc
pwKB+P5FWorrjBoSWM7iQ+auDGAzuz/fNR/oW4Z6W4vMv5ofi0Du9MpR9IK5VB5v
UDHO5gvCeNlJVkKHWnH6Q3qhOojdJ862JK6Pzr7KjAUcyXrEwagLs6urBQBSf8AW
0NV/0Xs0ezSFv4y4M5eUdB0xvCsCRKvoKjwb4msdlEuiaO969Fh+NVk5ahBMYpEH
pnTZGDHeeGnJwzKQxTccC+L1oHiig8zDhZ3OOy7yMFu9shbYtOL+k18iay7cWnIj
1i8vBTXo95znrLJTRZfQtcnZY3PlDv3JfbOQ0r/rWW65QV07VLGdMHIbTB4Eel+C
sP3P+exvSEaIIwdnxo5pmgV2OsuRyuyU4Uh6tSnj7EoXE1akLnhDcIB6zrHqbdzm
bbkSuCC+lWcymnTXPIzBYM5nRqH26Vx6o7DBFlKXp5hjDzwRjjDxw/pVHhR0oNVn
vPddjAgIRS3G95Zbk60+DSspiFmGb7MUa+2TFMxLeME1wgyadYqEK1UFZ7gzP4v3
RZGT6N5IzyTIdPdvm8+Q2D6JvZVWhChwrqNxlT4PXo7pflxEyuPNKIfTT7FMDqoo
KCL8HMLSl99ZrhZp0mfZKsG1tqKFsSjlfJPk7iFZtcx7ugUtAoLcLTtaOg3uDQh5
43L81szk3mCLktIPUN9UfOTLGylbSv36k/PQj202y+XxHdFhuG/d+CDB7c+Uv+SS
CVvt86529EsfSwP6fGlnWMtep/hwgqcEGiWboS3AIPsbXtqSTstaS9pD/YSv3W8a
3H+aZAFZxoK966RPFGPcUOiNd9mruu38Rp4/44p+TIR5oyEDWsIRLxb1EX4oTghW
Cx6HiICXmdv2Q5aXn19aK1riFSOsAuALVkNlyn0jnQ5UF7D9TnI/AAA+UfsTpAtV
JEM1aBD9yq/4oVcsNSQeUuDPAPaP+HIBrAqrwki5gqXGkml5Xri9ycZ9MNACIym4
mEdgQIbIJCGJzg8MoRJi1VkFCex9brducS8RH+MxqS6vGLHUl1PP3bqU/mVf2Zoq
fwDAuUpaizuhliZzmOElDVZOkF0uZSKbleh4hOt1UKmoDL3+jioL9ms34ypVNhkz
oBcN7wdvDAvBFiE0d9QC0AapNujjtsfc3gHQlD7hxoTXj0MCojbeKiMc9WBFE9Uv
OHS/UCr5nevEqlk7vCVuVS+u+DYTaDPR9ukmdnZyOoRADKZRZeHyKNROFKFn9zNY
/pxeAVPkLrKX/ebJxI6EX6lh6NHPlG/8j6W5e/CmSznLCo9EWfURwLOvhSiZBSMT
a6zo5zG9qsj1MQGaqtozxhApxC7mNmusRUsOTLeeK3QpBfu96IEZAX5FGZvA6Y98
UT3susANHWYMEXs+vpcMGPqEr52OArPcnXMxIYdzb/CkMCq43AdVRAY2c6HgBKRb
/WS0QKYW4ajt0Br2VSs7tG2MixOqJN9F9UKY72REclgnH6PJr3WVZZm6r0Wpr3EH
1H4Qyitv76gDrfGgx/4K0bn0NMiNZLIeqGS5v4plv4IGq1FOZhmEU1Y7MRjDVjYv
l3lglOIPc/tAYnoM8Aq6Tjwzf8xxtyY0wFLRMFRXDeI2uBde/MqUkqPvks0m+3ie
1aH4Iwp/pW2ftH7N70XPQkGZ4BYIh8HUuO3+g3J6MwN/8Ghqfutwcb7LLncyTJt4
YAAzh4ODwPLMTaQSFkXpSqPzQMl8E/hehvkQ9gAhzL75lntUrQBrBXhcM9P4XBdK
wcPhduvMVOm8mzdLUXnJCI+tqlIPr3kKANqB9hfbspAS2AtQ4Ucn7mHOSeUM3Rs3
a6WeAdda1767gmHCzbyokgMq1ZasFQhsab+ZhifcfpadY9jbNiMnfdZTp/hflu6P
KTiqJvnLgZQxPWrNauZ6pr3rw+Oe++BNUlE334Yk8K3rdeXAujbSv0+i4DvciztU
aaC4nIL/6xoecM9kQezXOt91NeOp2ft9LVNkBqTEAi0gqvJOxArn5JLG3adVEaJM
58IWbhOIfHAqYFH/KtMFK7DUN4smhpGGfQ6LlElvhtsDW303VRxBCi/i4Ry06l4B
JSz9FoilldkNKH5RvXNr4LQQgWwBfS4g8zZ6369KK3NhBoHFaz3pUhMoOPud0WKZ
srMlgzkcSVak/PrendCCUd7Tjxs4aQ1mTLG7Eb9UsGLlx33mJhu/RuGjYV3k9e8M
A2jWnBktxbh8kuFuffiaL5TKJdar2Y4kJRclrF5v1x2P1ocriEdMzQDe297eDoy/
0Ub0IK7vhGyYo98MwiXWAXkygg2JtAX7qAk7DW/jeYG5BSddL1difpMcec0HOBbl
4vaoNcyERHIVoB5iLYegEyFgO1p5UeK+8R/rWchRL+/xTVM0g06LvP4sQ8mP15dr
7N55TZflQhn1u+R5nVO7nr42obDJQBhamdTnftxrdiOdP1u850NtCaoE1EHl9GH6
GBEvgHyVnKEY3I4hJbtH+zNDaIV/uXPXq3Tu1QhS71u0uRRwMdtzey2oBzTQfso5
L/Vdiv7KujYJuM4SpYdxnDkdDXyJRJOURUXcZIpVoFqV5JlMsqkA0BhlOe86YEx9
KmPlxox1luSEQxLQbfOTJp3cfOjTXqPijzS6cuvyVHnahg38z+9P7t1H9xxHQLFw
mx/a3etsASPpHdb9OoyHEhtDQzfBP6iX57cvytL7tfoJz30dXbqjdVmGsl4B0xDM
pi6BfBGmqf/gmDsiG7D629gSenfH9NoZnqFkHK9FISf58TMpzP7bdBiyi+qCDmlq
/g8RudHtwXqwpJo97ilLuoy2a2lPEoAjz2vEhTE1Va/+qkhQ06ZmdltXB6PPvRh9
zYZet7Bj/PQlyriA6y1kc7iykPya1TIUzMSGo5n43OHp5ky/giRSdfmw2cIzduXW
buG6QEI+9AMsRAfIFyqq8bmKtKzUcTazJ6d6+AR2wKyJQStSEP62iAEh/kP6kF0q
XIchp6Py82+q4auN4GT3i0yHn/uD7sEqZnt5WkdvUeKu6sYBLwhMgNvrW1r8E9G6
a2T1eFdB6xe4maXo/+qEGduy5Z1mqYS10uslr7+1wjHnBfIIXOiuFq23eD0pgHkS
EjfFYSGzoQ2ygMDkUOiciZn5Pn7As0UA2DEqa5MtpXajK66WTsIWoP15nC5o2fFI
cATphRR0D5fkQ8lKZ6MEo5rClizGltPcByBVRd84/MSHBtchXexxT+265vJIj7oS
dfILWq/L1yi54Xoi6LXlW+U+85EXRTX44JV++H1FXrDpaRvNK37VqK+aEyvpQzI/
TWkgdENwdH5DdTuBD2aoaASnruSzeIlz5ZIlwAfsGGA5taeXT3E+Ad3HL6sbx4N8
b5VAJwsLL9hMDjciLh66GTCoag6Nx2VMUiGSzl0tm8atAzgfaES5y17OuzDcDjTT
+aB1Eq2JXLd0QkcpNGewx+Vtez5ye9A7qdrtkQ62SBFwRUhH5NTgf+SObyInjjNU
ukmcOFM745DMAkLKNgG9SPDFEHQ5aev2gP6aDgtCUSVqZk7L94Ym0oxoUJ/58b2U
HNd4XplFW3mu78y4RCsCfYlvNm8GkfxZfiOtcNJvH83cICsDd9ML0uBxL1tmBdSe
Rmr1Gbp5rfjD2Ft0UJTk+4jzAPwuZHzhgtTavXbgodYcrl2DGk4cSZyTs6gJvLGf
vZmYGL9mghp563vxsIq2oALkRW2GNKirIbebUhzToLnDZhQ6fww97djWwQPqTEqX
NPC5FAEoC77rNZpvFUKNYyJ+Ihp/Kh3CqNw+8pPtou2dID/KuEy7XALntS7Sv+hS
4r0eQpeMBV8DRNKciy0lQ2/qY6iNIcvqnct3Edddd/X7GMzCgb3rVpby5DvNcovc
fsE/NILYrpPTD046S53pHoBXiG4Be3O0TbvMkW+0rrlPIZlB3znVVbjAI/83vBeo
DGcgYz6obZnUygeKH3iDMIyIMeMidjwQhSIX9s4/Ag6LswPxKzjYk46MXDIglOgY
cUBAywM6zhZTjFCfGYc1663E8t1i8JgXPNDbngpnMGru5FqdtFK3eGpp1OTSehIY
tPyISUMcWGa8yRItqvt6ftVh2SxFkDCkrZerh5zpcVJNNYcbnWm1SdgDNwa+jL35
+AQ6JF4P0Ql+HKWuELMunBylEOPXxsgUo7wzImjVk+/R3vAsJkkpqjSI+R0zBuTp
fdJqTkoK27ksuswPcslPq6CWkV7aRo7w0JT5kaNzuvhSXazNqd9RsHgldmq+vaC7
LmIKGwxlnrwaHSUrsfcFCI/oCyT6vx/JWdGsCTReaGi/sjc3polChR7FifJhTk2k
lhLD8YhvjRXJI1Hl5WeHvC7y8kgzEsYBv+zvt9twuQl5BjFBMdsmRNLwPQjD3U9I
SKsRV4C09kZBCD0I1k26ypNQITg3qRQQ1tjjavfRz26U8SNhTP/TOIoO6yXSX+/G
uF8S/yPiZA1BMBG0u2qyS+HxXVkWcrx+wKJWD19GjKQ7Zbw3U90q1G/Z9AlSxXpo
QLVZTSC5ARfkLOwmYNnpbkMzCroimVEwYMUx5AaaAPBbKr2iE55cpqmA0oHGjjYx
aR5crNzrF4fZRM7c1E5xoffXg5nr3u76W3ajfbcFa1mjqLhXi3CFfuHmryL74sU/
odJeBwFJvsZy0OVMlZBWIduwZRgU9k0bz/whGkc1WKMWapYATq9r6ivnK9rLD5NL
tEx54TzJ8KQU2wg/pHIbwusH/p+MiXK4ziT6SUEL8brYKvXvrV7F5ke1AS7ZStZD
cvWSbVKNQ21hgRP1PzdZhUCjFSxnCxBJJwBwQsIaXHrLUAFw6Hn+49P6YPonnFZi
pBIPWgLG1mpzChHr7d6+NohsoXXyfRZvqVAhbeSTpkzGUu/obQbc/Bx4kBu/HgZx
r4JM64Hs9Zs3rdMA/6d5y8kBPOIvlK4Ia9WI3DFFBTH3YV62vCtqgFLb4lhNMfXh
v2A2tQyhtBLvst5NYUvYLqljYDf319sER52WN9NbkP4ppYxB2bvlxEv3ftlQUb4u
MJiC5eGeDg9bqx9be3jFd5RjUnb9nEPACM3syzqGuoEoPl39NxFGT8XJ/VWUBWqE
7bnj+B/qE9pO4pk+QqGxyvBp+PgRRJ554bUUnV/BelIm7PXemt2irGt9Wd1102pi
+F7jlcs9ZQ0RAcFmNCfHqmERaYGsPUwjO8KVNchlOeu3XEpR9gKeFwyqEE7J7fyR
r2WBArgu8GtUR1jktv+kfdxasQE9FfUkEi/VOztnfWtxjLNfgEaF2HPMztzZBoH6
hT5waBZ3behdn8U9NkxxMP1aWVRcYo+NAZQ3D725sSIE1UazcdjBFgtbCsXWkJhV
GR0U6tUXJi9iKnpadwwFViQnVo7TWgPVplt6OhZBBQW6fcU+CArp7BEPs29nOvtQ
b33GY74a+q35p4EsYAxZ+HoGQoLtL0C7BBgi6IQVCiAFn1h3rTgw+DOTq9z0v9/9
UnWIp/WNceQzgIkJMChpUIQ5Wkez18H/0ed6lxPef/8H/9GHsZREQ6lcUZpZJUNr
CEt8ikCM1TpX6oCMq7yFYVt1vcoaoUrakfBzyu1KvLGLmG/RwZwGU6+X6wn/pApE
VLeGxueNZif6rl+EUmEPK9yRWOMTGYowCZbOsgSfRO02Rx0YZ0pc0iS45h9Vjhrw
VkZ8WgCueAL1A0Ypolqg1kfv3l5Re2bzaZ0DraSg+04DIjRE+DeIpnAbFqEZTiW7
SJ/7M9nih8bKhI4gZ5tYD+HyKgt3pa3ig7xO17ZNPObo5xJOUNGFtVz79zBaguuW
8oVxj/IW0v9VLSQMjiOIVrX3WNiWBJpeL9/5A7MErWBclAbMONJINasUm9dvJw7t
CxgXHRKhgXNJCHiX9PDTJ/AiMqILNY6ZUq6Wvx2amtqDsr/gAMhazphPAvuzzgbv
MXmS/Rip4CA2al5sUaATuXe5H2YB+iDA+k3KabtHmqk/K0xXzEVzgx95RqYssrTW
cZE3x1boVoPdQftRu9+S6OOcap5uqTrywfP9Si3xPVdKrEXyXKmmeGkvMuYfo8Ur
MhruW8r5zIxSVLxCn8+iZ5nffZQYp1ZQbBcuv2M4Kt9vFEzjLoJ89YC9pnpZz4dX
X4cz2rJuPLggCyzEr7pxdSQeeV4YINSoNLd/yihooLUtMMkecG/YuCRkY8FSKOAj
qnMBuaYuLkG5DIY4babN0mEGV2HkNlf9rX//HVCNFesOOps4tfMbWZdN1iPTgq8U
U3LwqwOuKo/liuIM+Kq2MPQ9bj6hH6bKZRCMJo9MRVcaeriy26O6y6qfDfH/B6QW
TwqYE36hJN9M+yNIBPJR+RwkajbSNFTQR4+pOBAuP69tww++SP5GwbnYKgTfl8ul
/cWZXvfeXzuF2QI/bI1z6wVi+8YFR3y92eJU0Mwl3+2oPMa0GOp2Ip4bdBVogfzG
pARVKNbCDxLvD2ZAZkyDp7l4L6U7esImRVxERMtkqVzJiOWhmoUEK87FA664OQpP
M66UvTCcD8aTs0Rv+/PqpeInsB+tmtFSjxR0qQTduAE+sU3EPHFR2rqJ7PZwQ6F4
gNKyI79ZxAiTmkykCCp6bd270MW14Vn3zDioiUHFOcJ2Mxdl1VwXARhLti1gQmMw
WzqFJwjZa6tIA8Q6NjIpBGm5JBnle8r5EKNau+HkCX+vvE6Woo8GhHeYrvsiXNPW
F/REdeEwo7/8mGZl75Mplhid6yuIGOexi14Ae00UQwb0mgqe5QSgHRAoIJP3air5
E+UdkIS1U4X5DbTj3VKLXdutGe1Sre0Rpka8TsENV4EpYW3kzaoH9orGsavoUOa2
GCalyKTT1NocrCE9TkIo0dbQmm/LmAfcCAzTzoyAlTKwUTd3z7yCmeopaFd1Bz06
Cc2Lq416cX7Fg4NyxuZbPPwVDoOkaaK/E991/eSfQMZfMhVHxEXPQfGmnATePR7R
hv5MB9aeXvGBiqRjthPoQwfRciEKXxsD3kLT5KqjwX/MwyUS7UQFcwPbH5RADtma
LnEfkoD3jlhuxtwbTFLoKsC9i2R2ENO8ikQlcErrvIXrB2z36XsDQl0cCx9iWIFp
+V4uUXiTA3xnD+Sb0moEvXgSe72WL8zKk/2zHdekFElB6d+8BV6jyyfUWB51YMX6
FpVpiqk0kogAkAYXWIZ5mqtekHUXZ6XSTPMgPHRg+o0DcGD03AX5G8c2Ji1DM/s7
XlKc7wEKvlDeAsLpiv6dvsVy8rX9+Y4bJBVNK6mgbU8Z6JujE4dQdTqhoGVW73yM
cWUOd9N0Bnxk8LrUt4JNwC4BWRo/WarXNZeqRABxkfvp5LRC6sVGMb3Tq7GdQjqw
dfvZwDkaBYMui+zr7YtvrHXOcsDylr27HSTCjGHI1UOU0cT5w9OqSvR9OV7hCcfm
E5N0c82eYMwcvw2TUZf84ynK1qOkd3ewO1wrzv7n1yFJKXfFt/0FY12Lvo7o07ym
WwTxQA3NEn4AlTiHVoy+6VnqL+TA+vYSV91W5W32xHpyuSKe9+xuG+ZpCIxD2mlW
eofqqOxfLGuTjKpu1N8EXLU1qbig4DQtzQnMyYKvPoDN3k+sbf4NHnQQEc7wIGZD
/nPf5cxDZuQRybciY2HfIkuuPsDAK5b375nrHn5Ea9GyHnOiniDObvRaHOJRrz5S
XDwsaofYTwm1nrvAfKVg0aaV/gm/bsfZfwdCloOzi26raMev36j8CALBchKTSpeU
f3l4hHbJQ2vtqnO+wGFFGh9qiHVnlsWgaqi8j0H67FoSQiI7QytXftcg0Zkg/Pep
Zr9C3Tn2zubOkGkZ1rvS7r0mE0gsQB8IIw+CC/3VR9DR2c+3b0X7Mr/tvMPAxp7g
jDmOlltvLjtf9m0yzeV0PGBxGsoCKrOVrL1j/XTHHtzuL4Ro3dAEupK5Yl8Wn1P9
WwiVvJzSEB52NK5sI30S5poE8MoHNGndqGCcq96qbBeidVujI/uB+njgJ8rnmkIL
Zesf3SIM9oal6LjA2JgpHGzHogRdYnVX4IFqKWD4XanrhOC3a5Av91giuHrt8EwB
XDISGWtm9c1uI8gz0F4q6vhrVGNLYYwGc8J2iFXr4VxTM4uF9TGGj4a/DfLOkCvO
invyLYPvit2kRB4RXk+5ny3TqL+pHpb2iYnMxNBtkB0oZDZ1ARVYWu0JnJNdAoje
JEL4S2TMMDJEEySWBLxE0mJSJl0Mx7wp8WlMstvJhbD1mQVQO9vwBEFC/ls2s1j2
7fVOBYgyUz2yp4GnL37GMTlFKm0aQJRpOkQyBAISt6FtUL12qUI0b+faW5L/siNh
xfC75Cm6aXSvGRy73g4fiffP7bwPc0O+BmcgqAg8kAfNlue62jYh8Abg1dZyMDI3
KBDB8b2F8/5xdNFsCwOM2JX6ii/D+GF4bcpQKaJlhAArOXviARw21bUZGoVc4WDP
D5egyxzkdeXnIKbKPuLD0Ts2z6geKeSr08qwf5gYxgu/HNpVVO/vmRPlQPAEl7p5
AmWx1qPUCMKJIXcDAkVagOraT1knwnyiCb9FTaet4UXOEsQSsObrbpudFRKpa6YM
mH2kaCO/IF7m7+yrsKcAmFTKZr0WtI4+8TmpUUQoqNL14P9YvVjTulQKmTjJoA4W
jBvXvyoS+YbuxX7CIbOYns6moGEEiS8mThy5m0hGiTRjvCVPOQY28ygfzANm/lKi
YSGCgrCTxK/rWnFSJD9A/1y0GEXJ7Wz6OeD76D9AoRUFN75ykBNvFe5bx4lxlS+1
DJMD3I1WIO+tfweNI88hs9pfF72pOuDqi/KoJEMZFIF1JFh8orWGPgOUGyjdnTp1
uXCe5z/D3SyDSmMZ+U41Y7OyAmHCnnlq/ChdspLBSil6ZH+a+m90qhTMCTwETcq3
sYyErn7ZagQ68+ZQimVgyGMKXv2/a+yRjuFSnU21vi3uwEY38VviEmBxcQ9N1miA
w+P5EW/u0iyTqaF2rJ4j92HjKPj2CtMsECS3Ng4naKy1LRUlWpMlhQJGv8Ejc35h
fY01GtGgkg1jE1IGa24phw==
`pragma protect end_protected
