// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:21:16 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LRuPSVX3OZhzgMZcUhSNapyK38a6CtxLqu7kR28iN1sIQdQvy4k0o4N2AYKIkTVa
apQx/ztMiYTs6v01YuB2VjpmjWFEi02jyD8j5MrCuY6+gQDYAEhfLWBUPUi+KpvR
Hlp/8QEaRjhWNgHrX5SxhspxgiQo1M2+MT6kIS+C4nE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9472)
VoHkhClfm8qj0Zic3t4/huVuNJtccynKq+FroCN4Pfwy48/ZShEDzH+zZ65DtdqO
OMeEHfRDXMwkx6hDWbzNDNlT4aia5zf1OtZScaSYHMRLZugNj408i3G0AAddcWGB
L13X8tmCoqySW0pEsg29hdBbuihh2Sgy+GVKokW1e0JldVAVJ+Khoj+WC0DzQQFq
VEgnuCiJW/jWThXYj2x5jKJSPAllv2uiOk4jlyJ7p1DNb5xZou4NgFyej0S84YHh
gbztrHrClcHplHohHw7qqK2GmyDYTxsU/TfBCESghTp53PFLkXXFuU+i5135eL5R
J1dGR+THbiufagF7aFML/pbQc16DY2qLbfR6VjYgie/k6KgG+I2tau+qCpxTpDkf
QRxsGT3Q/1ZFDz42nw31L9GLFl3Vb/vc1b8VwbP0+HV9F/0mkWIMgbArOQoELL1m
4FrD/t3IylYWjz+uJMJ3Lf82LdD7vnrJVyygfIW/L+QYB5ZjjIXbqUir74jntNvH
Jgjwa31llgK3fkJvofQVrEh7X373muWIxKSp+5p1evnymTob693ZsZWevFGgkXZI
8SpYeZTieZlvOj12HxOrIgtkFTYcJHr1mdbS8l5YyFsgI7O/6GUN/8q5Px6iBzP4
Z9O/goqSN95MesVVeltTWkzBukigwxcU1eX/MMHZBt+wvYABcruH7mUcQKKISLSD
0whvK9ENl4JlneT+R/Zo80ExO1yqP+yO8K6okRUs9Dkdt80U6/OxgkeGHEXPjQIx
gKWoMQmaBI9Y2ILhF2fw5s/lekq9LOjuKzwpnShvHDhms7968CTjk1/+ulSZEBi2
+RM7R4vC/PSp4FetiLCrs6gO1Oo4P8wYc9G9zIW6F41PMjQkoeCbRc2Ipj22FDdh
6RzLaZerQOsL8oGLHX89IL+q2XVuCISX159neIZxUWJ7VLhWhpBJWDsEqCHLTsDo
chxIt6t2P4rePrzC1HOBySZqdFae7kxJUBcY6o0RhTw4KZJYZX2tF3aDttO50HTz
UtiaHqm2QiQZ0Qc5Jixx/PL0OGbk59bWENqWyBgxAUSK0YztpcNJFrAof3+zKHvZ
Ph40bW2mQ7b9K9HcwXnf5WfnjUTz0VN4uOeFWKwg9Q4AUrjN+VXNPh0grO0OJndS
T8DU+eEsWeQG5zA2/fyJDRqlcCJn8YCTFP/HTKdFkel+WXFTpahe5u3LOgFlbgg9
vlxR97UC/ob2nE3TGF17xFc+bgTnj2vJ1Pmw0Wc8SNbSOrIXwPhbpm+waU4AQPtW
YvogLZHyGmPOC9vGBDgXANx6vmvQvqmi2bkb4rmt8JNjWtZ1EJGPB1CkwMNY/Wvc
JLQNUgu76PhdLzdCcD5rTP6QZNz8IlxTfKUnOYI1lcqMEoD2AXpxah1LpfKz+fDf
RIs3O/jp5OfIqTqnsYzK63yeH+Mdj/W7wJEpU9ZkVxcrkzR1jDg/kp6HpdpXoNWr
5XxMSyQFuhVNDxgLP/E7kFet5F6aOOGjC8Or+cwz2+YOQU87An9PezK/TSFlmeAL
V1t62BgMHNDtU74GUXanVXdXIBuN0D6gzR3TH3jIp9zfjswZp27igpwyAYOgJQvZ
xz/tQWSUPuG3RQo3ECukUQzKZlSiX/IE43MkP8n7+oVPXgPPIBrawvL7auiuA16p
NFm3Q8iSf8w0Ekom7qEvK0WeLILZT3QtihATBiq6x0EnRh1vNVB5rHuAL6I1WnAX
ipiEVMfdhLRh6POI2cDNOIW9TfGA1opsUDYSj74WTJHLli8/iJ0XI2BWjA4xmE8m
J5IWY+fj8+JgjAsp7B6BkkKlW31HAcK846YItH+a9ElktSb9rqWqo8cq8niXNKdq
nF3K1WEBKaTYo9FMvyTFf6Rbj4o8HXXunwXsM1WSGrakL8fMPJcHilMdBWoW/FTH
aTuXfC8NOzMEpHQp2lnxRTozLFBpxjpfn7zF09DLG73XIhsLx0TLeSxcRz6Nr+T0
G8STe70DqBCyU11X0rQWj3+lCRZ5sULVfexeWVtEa5DXjb34TM1LjjqWadBOwJbU
5B+JrwIJq1pg4AlKoKhx0TkTxfI6gFEsnJg7/U0gjOTAbEp2Lu+tOWiKSxhY4Aky
4TXHGyWbniq7/Z7mRuG2aMDSSc0Ar/UpDiHRQxkIo4T1Q5R2hbbQ4K0cb0Q4F4HI
1sXdRXLmdtjB70dpJDOLknEMhyGVRjGF8ZRklxZJ70Auib+Fu4aQu7ZQzcZwbQJz
q6lCSBqAMpng0lvCH9Vh1tqVt3zdGi5ktKAPSOpQi13oxI/sU57y0kkWMLtMZTXx
1Rcqyv5xDpFdlLneV3bHxwjX/8iRVUpCxiTbpvWB2ZKXqaV6ops3+vb5sqcD4dGU
tX1+kRB6m0dfSQy+yfmNxgKp2ZMqHmK5MpSKkVj6hEkLXKiBhYo8jSOJhmnNWi30
kenm0smVRZCnr4zN/yq55hqpi4kebbI3zxhZdM6y1v2bsHLBUzvgPp1cGcLy6dX8
XUH0gj1rxbjJOPYLbG0sBTZ3iVYyy5YfvsX7U5xb4GSuFWmzhVC9i6aj9ZyIr+0t
f2bgy5YnXUxsTdBbYFZHuzwxy+0IpqtS3XAItYIIXxo9q3ilOHEB96uOJbGQRaUy
vjeNJ81KMIp2WBYW9sahlRqvsaKKK8v8IkNEtHWBbxNvHyXTjD6onJHajDt0ehbn
U7i/5FDsKx28UaFe6bJp39hd9w2j4qOxPyJ+7LtAvIW4hwn59Dc0uNzVUzkoJjyj
LpFMU4kWqWItceYLGpybhyJClQM3qT4ihClTmehXLb7srLF+Q8ewO5+0DkCERDx2
oLOuGjRrbKAeWUvJmYa22n/jBF/QHnQZsHg4qJ6UCYESMLppawSimDyko+k0BurL
YfKxnoavjiupUd72zGj32qX9wn5PkEBP0i71d9rJA0gsBvT3AGBHySbSiJM0XKzj
TB1EttFXmr66UoWmoLDmOkTX7wgueCDqfOb6lZC1t+mbeXu+mp6PcnH6luy/V12q
AcHhPMXgf/vMqOg/JG8Uyzx49I6Dmq8nCHlXGWdC93/NRkQiICXCTUnxmnmyLz2z
hkvpJxhO72F7PesJbmlpdeVGXEB4nwCdGRkdHKdrCP2iVkQ1QL0uufSFUKlSAPc/
68xBLd22ofVqjKm4DONupEK1acMA/EYLACkvdHfuxvJ30WSHCFV94Rs0jlRi9CTl
gbEhNInR2pDlG0XCPhjdO3jbW8M4sr8XLg6PLt3gZrvqgy6M4eoa5yJJ0EuoF7M/
jvmIXiDRMAHoZEtXxGDepg0untOfr+fjONJlsmLCG4hmBLzPrdWmIUobx6LGpSs5
vfzrnkd2UsmQVYMa0lTnZ6/2GtpljNIW/wHc8ND0cEImB7SSg0hATBZH/rk+btFz
a17XKa1H5c3smbxASu2pab+a4UNCo2l3HFCfzcN7wNQJPp1K54thfED55tWo4rjH
Icvq1eBliop7yvirjnXwtrcZAH/NPMD6N8epEAOVuHp3IAOdz8XuOXQPHpdLYLhd
Inb7lYJRpxHNKhqD4Vw3RzOfeRki/kp5iMC/+AFjLNYv2a+6mFyJbwBZetp5IrX3
bibPIqbUEJdTUW2LmPHDxh3rj8zT3hS8chtut1lBfsz1DZQgXM0410eh65PLAwPl
/5AttJ7HTXTGuwiTQNcqv8/TYrVltH/VoJX1rNn/XyO/XDm5g8w6CPM8VIfh+fDb
nqc+VavSXYx9eBaCYdQuE/uJT0jYlJUHbqyt1e1+C+AXx5rvWYWz5MeS7/w/LhpM
WLfauK7V6WJnROuFnwPCMTvShap5s9vtNdsmITEmzlMEtu+vz++oYnxvhd44pPux
LtG2dYDxRQzNcOwIqSwyhLWeNJd7FE8nJ5FiDxygvHUCOTasQMsKBt224gtlV1b9
7wJCkLzmGBFmjt3R4phRKrgP7DOGGoQQkjFZtgqKCLAz3T8WY66OsjJAJwxT5h5P
WlXxm3cuMqZDrwfCwS+aiClNHeFuMnLrvet+V1zIbIyqMsGh7JKsbcsmRwlJoMkh
ma0wGuzmPk/lhNCuR+q55LMz70xAmr93G8qvUS/dDH+QTOr+FSS523bO1ZifFF8a
I5vjwT0NpiJ/IKnxWHRdT5wAzN/oEhwSOApkKUMY78FNnwE+bYg/p3QejUBpTeBy
nmpPkKCPMIq/rjfARAB6oFlF+beLbI4ip6a6ska14zHfVWNzuB/wOxxGkOlYf84L
3eCoqHAl6h4CfmLBQLbx2y3keqK+8vH3+7BmuabrGyoCLa4jHH6ZxVApDxZlSBmF
bu3FpE+VPtHm/L+T3vWPE+2/lP3nJuTMKE6+C9KdmYOBRKaQBzRJqS+ZK2kzjdof
d7vfNglTsNa8UUwUXTmanOjzHd05KYX/XgaKtWkk/bkypOlb+GoYEmqnMRLByXYI
qU51JHgLgF1WxY7I/3f0PW7Y+jBF4kZqCsC4uksZsczPJ/hGnWyInPsxvxhLu28D
i/BgzbIDvCMyO345wFzXsg2Bnw0HrDOyo0W0kQDSQQGHzJ8pJa+zlpTMuusIdGH4
c+OHw7sg5BeyS4sr+ipB8CUZettkyKk6of2d6mf+S9HPuCJ/dtr6r8Bs9Gla5nwv
Wmq9OOnNT19J24Cr7eZOimsnN9UXEyOAOTG+pkt/JQovloRx3+uWMhCjffBrfXoS
hFGIio8ixHglIzcECXTMAVwqHRcImCvlpPHqYV7p/WguliCTxHUlGj4vftQHn8BG
bSt4ubStV9dbfTZscNFfFN1M+h+s15pdNGUJy3ecxLbGqw5+b5ahfyK/VijCGuTY
e1ER2s0MYZeYyL6Vr9wHlBS7ULXSol//uYQwblnmy9+NOCIAia2CGoHj58p9aQkv
FoTYCMepM/Wr/cfAj2lo7ThKsJOwX0LAxoqB1BwUTOnBZFr14V6PlnIr1EI6Q/BC
914hqst7G6zrv5JY4G3jb2DGbRh/8+kJK0ANuzX9KOtQKZzzDorqbujwIls4W64W
Hn7494+1IoYY0B7xTBfdfzUKwA3m/uxIJN8a3MAcHdCwINiAyooF5Ze/04DR/FUb
hvXMkHE8A15NR2J5AEftEXxa9Qp5Gtkarez3Z/74Wv5rYWFc+QijdWKNLfYTLJII
XfQenzknx7/O8lumHYkkKI1gkDJBbIMTirhaXwwTpaZS5j1XUXMANuB9JXBkDqod
6b9i5wPUZgNp/5Bili0UafbW69R/7e7Wa1r5tUNGdTUJQm4qFe3hOl/SEI7dDg8p
ntoecLub4biKG2sv/czWt32TzluXrZvokbFW7Q1LLNXgNQJU8uUsOQWGZ24dz1W9
k/VyrP4ztvzbFnsZJY2aBilX7tOSIIp8o83hVeLuWMx1qi6wBXg4L8B8xap6AToL
VJ//kEepSL+ao7TwNMiEgWMWpCNIZ17qhnlPGsg9EWLeu+qT97jT7VARJBVbHRwU
BKWT2pND92nC7c3Re1hYynrK7Mksxz1HM3rvwQTMNoiLB8/oIIlVMj/PqRVXyO/k
JlcBNkl+HKtu92OdB8I2ah38ufzemFjve6ArMIytzdnjAnZ+d39uPFnon4AbmLR+
d42P5svrjCSLHt/R98dw8xWSMoFT3w/Eymk1eSwg0dKvASS6shgH1826M371FeP5
5gq4AS0c6TuXq9jx1kWXzJvgaG/jV1+Yh/WLXSIYH11RjnNtJCHzPvWEC7ykHi5Z
ay1AYXZMQM/N34gUxVg8r9wWJuZfZ2h7TBo+JJ/Z5eCXciwgsxl0yMvSobQ/oGoK
zT2ZiVypT6Ln4rRXrUl6gRoEtELXt7kLHzuWlvDoHDJ9mxkws85MxWhQU8+LfdWe
ZDzUgfSTa9E+jXD1ssTApoDrkPSPI5Tk3SwcSzNLD/TGftZTfhr5mU6z2M4+thse
MuNS92CNOU9vYj/9Qci8YgrdzQziXRA8/KyZgBVjHHl18o2KGraY0Mn2Qw7+BZn+
FZgLXe9UWIwXcfwKWywFNtz0WkvLgwQcI+vscy3UqXjlt2U+ThrAJRu7jzgHV7Yb
O8HND54oWQp8EM/43BCvmpHdmnTjmQfEP7qRRhstorugKRBq1N463RLiu7NHIWCP
NzQfHZqAe2dfc6UMYRNpv9sb3PawFrpYxqq5Df2VAEwbTGdIqa6IH72CmUqHtuP/
1nx2E9EYdLOYptv3TNebxTTLXdwTm4vQ/ZXF5qNF4iEkCzeu1iRgX2XbmVyHvaE2
u1JBRGiUKa5/lZVsDNTscl+0uOfL8Ldg9a2Ag3tnORmjfBimuylAsrvZSjvzVZhk
834v0f2GpQdEOYcJtLOZVhW2rAGpSRQQt7naHqeDE1DJTRcWuNPRJ4A3bUomu1a/
uMn/0Ai3tYciN93I1L7diYNRU8u71nAa0UbmkN/4baBBE+uCqAMPmb3xolRvauiR
PtkjSIS1Z1DCQhybnJAyiuxaZbrteye3OiD7WfhnAImgTtyL0LlvnBrefAanj9HO
hgLGMs94T8lx3KHafkQm2BKglhQrOguOfdaQHUpTVLnM/6IzOvw9Kb5z2I+J44YB
mfY1JHtUo0Kq9UsaC5RxEikIv5z01S3AHHdFouIExywB6dZLJo3yt6Hj7FyZskvp
txFQ8EnBeYY1p03L6soFoFz+HePh7hALibkuIzM/utN4P5HcBq3O2R5+mXqyFNqk
yMFdgU9ISGOXorndrEzMV1O+lZfzYKve8tWG1LI3Q6KEQABouCAxUcyBUWiTIRF7
n7JqqLb4agjT2v75c1//A1MHFinmUopLKdD4WLr09BJYQyXDJoAvIfkX8ecbpmH8
cGgpxIgnYGPSKaH2Mu+mvTM7RF7eKwsNZ6KUOFuh1Na2hDIY7C60ih4EoF9I8kuA
ofqMLEq6dDBtzW1TmSlHSCrmjk+zJagLQg13DOnyi8xMkV6XakI0xeNzZA86jguE
qhM4/Ruv4VJnBinDjr94gIyw4Ql8u3i5tz259G4Z1ZIvI26WPNL7kQJ6qcC6csw7
HmkszBDzy9UTX4X4aVIhHlpT7po/HZrwUK1cS3crpd7pQukplczIinJZCy0CRjsG
aBuZJiiQs1YpDA6a4wgZQQP1ad0yNKY4mPzmeKljFmgu0c6ipCvnC+kdr/7ZX0oB
F5ZUBCLykvYSRQ0tm250AF4KbO7grib2DFl4I4QSpNWyvXbY3V6MIj29Lsm1vHOy
nizt3MW+TiezPg9d9E6rb1ZiIROsPUZ60X/IKl89dYeGF9lGlB0VBHqY/xbdg6GM
RBxFdjUjc9LYKJUSOa/jPWSSzO1Ufi19cSjSttCX1dJp3CQ3b6uH20u5KauZeA3o
4Ez77JVxZ7J7aq+c1r7gGsT3teZN02nceETbPJk0iV44mJ9iUIkY9msBfTsZv00+
DKFUaVYGVFzFhAyT89AhIUvUVk8wQ9rwvInBZmRdzwJdDhv4vts60jjpeP96RVv+
DWbpFGlt0eN9Y7MfuXFHpyjT3btJ15vgZ1OO7DDBX4Gx7J7RxjT7wNIudDNp5V0H
lIwX1QHOjFcGHM0TXdRD/ARyUUOKYOv8Cphs9sRhUGZf+lOb4ELUCWa8BO3ev1oo
OL2vvWoy4r/9aG1ILc47C3x6kosFJyiVipU2dvSTpFR6itIvpLplsXOhK68pvzEZ
sbjWMD2qjsleQrRr1uC1mSBJ4NjI7EF7IVvk3tNfqYljAfTIhzELy2QkNAyQTwN4
u6N/EuwwCnnW9dk/CNk0UvK67q58/kKsfC5e2kBf32XiTpNCDdz8tKaXVy/247gL
BfwoytzPbzDOaOMkv5+CxZL7MHrT/pab0UOMoP8NdYxGB86rmzToqj3V6pBFLkXn
VimZC0CZzq487Ne5n3QLajugoML6t/nchQ7IOdKSToncdzhzu+hBsCjb5z1cPigE
qXyQILb6eOyluktN5dy7hW/mtVXchdBTP3C4/EwtO36S8gr4XKmXOvXXUWP5ZWIS
kk/LItD822SI6Vn68vm7LnF7SCO3lg+nnngRiJQekI1r7drKGVntq03FJaUJfJUw
1E79grLt/Vaq+Y0yN9XRXBB5spXUqBZVmCjHxIVC8ZjuKkWJXNtYN8Po+sKE8BND
9n3yNG2U6rtDy3ILY0j/ezs82MxMNaNGgYKbr920O2xfEG90DLVU7Kh9ihU+JTzd
Wkw9r/lRLsy/9YGht9ur8lmxU1KKPvdDHnllAN842JfxzX1YPD3sTMkQG9BvkFKA
KePhfIspLU2N1ZDzmwVLOseiIHLnhM9431Q1DkuQqrrNLZk+yk8ILdnKXJDC3gAj
tkmVUXrjwJ08d7BjcuvgnY8Vkegls4SaV1OS6CM1ZejgKlTWvCwG3FwYfThxl31G
YPWMU3HZRZ3mWdJszXsuGeHCge6AG5Sf72saI7oWIoLl39ouTbOZxMMYahoUyJ9s
kuymeFTP/RwdsDU3HZy4j9G4vEyXeRHmFMbYN7xFqK75TSJr6dtvtvB7JEWt9wlI
zPSCoZh3YpsJecLH2Q4QqKOK6wmkOkC+geskEN50aUGLOOD5N9Xz4CgQrmcqQN6P
x6IgJDmeoHPOEotf03bJj0pUnmEqBE/24ic1giEpVib/cAXui1m4pnIuSYxgYPZi
Nog7NLGROy69L/3Z3GGXEG3at6lGC0zkG9hFP+fvzgqChWt1GuOWro5MvCxzYLmd
BBRaTXPotJiwTiTuB+qveR8Vstp3zzSuWmle/It6gWKnI3SkZvrVtWCZZPPZgDiX
2nbPgFvi/MnM+KWiciF7rQoGcOtu/7MJkYh4UPeiNsiy3bfxt8clCE1qMfdRrkek
bp54kef0izSx9ccnaIyoQCYcPkjn548nEyAC3uA/12G1Baytf8jlrINX3B0RUSj+
8etqOgvmr/0CD1UV8uOV8b7hWWYdjNuKwLgRjYfZwO1CMr3vK6cirMRkT2/zTVxB
qPXknOCJncftADBsHfplWrXuFGX+zJbI5e7zXMs9Oof/00ph+AmSL3jfehRxIOi6
9Ovlcl9ItG32bAREpheEuabXv1pCFVWc5bN9VQQ88i6ggbImJR0+4S0cn2wNuVzn
DQvR3O2cMxzFW8dgvupwU+64yTDa5STJfltiSCZ6Mwj+MXDJ6Ovz2Xr1A5wjhq5a
FeaciARdSUEgHs8B50gLOyhBO+cXknhEJab0udj+3u+ScT4uZUCJzLpvbhtcksG4
GMYyOqGhhgsZuxP9w7mxzEQnrJwWNNrFtqcU2Ug4n6yq7TnyfdovtHLk5ktyh50M
CITTNS+TO0Q7H28WoGTDMmarGnrmZidJFBYZI8+Wz23PTJGDrO86BK3gqNGioHdf
+9vIK4UcYVnY7dkLKHWHOXcWvlWJflGWjQx0oDuS8iPH+T/1KF8aDugicTvZW5MH
iMxK/0PnLkRcmn+zP3qJax/DbggHThG+AIfTzmFeI0ETQNHKtLNvrcfLFsQuCYuZ
mrcCNqGfiCtvMPcpUrX6SZcOkWm6seQVzS3Ut1zsY5RLq0kkcyQfZ3ZtjowMoCVB
UtE5GOd83hwlaBP3n+0G6q5Zgy/EVHhWH1elK9p+SDsKxnUHeqZsNpvM2eRVPML0
k6AvM81neIu/4/vh5S3y319T6HbziDr/vZHwZV9bgxISqq9vbAcVjJxmmCBEr4Jh
lUlOH3T/ALPGUchnrrHp3GKEizRI2+RJtUXLCpV802VwT7rQeNo7bqSajeh/LWJk
3SSD0LvX9Jp2RYtd0oFENjJ9A6N1iXniAvRg6kKhjIf21W5YSs2gCw1man8NL+PF
xPNUrdbjM5sNV/DKfB2CAqy4ngcHvmr6ZwekVP0ZoFkxP+eWtDTRnxuXLjO+sbDs
hEWL0+I7UORBYlMXqahFBda5Qhe3Z72IiTaSGDCEvYDRDt4RT/HDW8I7icL6ynaK
VsDGLlFuYoMtMzYYQmrtiKeK4074yWs7JuLXpQ3S1LCCyG2Fzp49B/03giMG+/sr
mQ3YXWmolyFU6NNM9NfP4SFIV2UA0AQQl1lBMpwvSf5RDzrVP2BWR25rYuXx6EDP
S4YyyZ+1MJCgSNfUUMUlp2kDIRQa7q9zMeLCak4hVI/JOaGywYCx3NdIQjCqftmM
avFkgmFaEJ24Ox9Wrd9m6onqErOAnnHRoBRPJU8LlhmO9nznJyUEQm3IzVCsfCei
rVUDLgOl1oEZFgBPdi1tf42saY2iZ/2Bk/ojm1rFgsbhHA6lgjTt8Hlywz0K9XDW
khZTE+niyoWSGq/ib/rzxgDcduCuiSvZTo2Njlw7SU7bL4PCOLgJerIRwaldW4YV
azlN8KbzJ+R4et05XzNX3mwp8L1NHtlI9t1Y+hpFb7TtyVztz8KHEwPXuMcyqJMK
oFw2wg/tBrZWOZ2XjrWsoNi+gXBnUe7CRwskLOOhtmHsii0uPF7ZbCCIf6/ZNMSV
0429xSuoOgWF0w7vcKFheKAEvM2Y9rWKojWvo/LN+tO7qv6zCbrtk2YiPQb7+Klx
OUtybu8J6njSpVDahF5Jyv9d7fL8GBXxRitMlqPV+L+1myvTwqDa8JeIH5LxM1Qm
21uDp0Q93rsz8rNAByyjG8Ytany5Wx+8aFQ4qMuv0GHotLCs9hKSImZRhPbGS32U
kCkc1W+6hKYQCwzSeex6U5YBq/E4WJeyIt9joMjjHygo2eeaOMzyUAt8IlqPwaPj
NfKFF3izTs8ulxiQAOgXHAFxqm8+wIOSgl2QGZzK1t77s4mn03PKm8Hlz+7jBUEw
0yKCGtfPtgUBjaA/IuXtXHxxF5Vq/pUSPf49ksDdeQSK/N7VIU4T5EyKObFnG3Yu
Q6oQbk+x4piHJNBsjKFVAKrFgXEjemY038tm5YzNOjs9jb1XurOM1jgNjkES1j53
RbCPzUefZcgPDp9XbVqpJe2Bd0NgR8xAOfW0jNv7X9Uz1pgQDHNtqAGHW7yngTx3
oBOt8bHxUb9mQk+q1XyWuinNuFFN3SowO/Q5oqjKRujyZYJKR/5OWm3E5fmQrjUh
S0aH/DYnuyZWr9qL7d1rT/+ZlWysvEuDmuY/R9vysnavPyEp5AQypvYL2+QdQJrr
kdI4WjDtIHApCoHrSyCVPo7dQMK+Jlt27CaEgELYTKXb+3UtjyNUp56W1yBlE2qu
jOXgKKEQlKz8r3azm4W9FsdqoX2iNs95fWkKfV29fOU1afxh+Lka8aN1qeZQxCyz
R6D+YlnjhH6PtH4AUehJTT4EZHwowZWZiNgHUmZGS4eIdPjuykrIaeTMFTKZp/58
z6h2yBouKLhkyKa2FVH+4CvOdtWRVGcj96ciYAuHVjE7kcUPDae+xJ4da71phKR5
ni99sdUXSV8O8mjFIS2vISCtjjnl+06h/g1A8kutCHzDqMJHwr3tVblOR7RXj9fv
BP/WRqsOYnsrekhS06LceQD8sQmTb5gX+WeGDVhhdBNKwJ3badBu8XE5N8S19bmi
J/QMD3TAZfIJTVemDpoSEa38ogvn6oIKoMUhuzX9Hr+FBAZ8qxaALhv6jx+VQxQJ
IRxKCnGZ6CmjoKOyilpyhA7IfoxHqbtL64gy+PHzzJMlUxTkjPTJ8U03RTXl9Kua
rrrKRoKwF2mBQhWgBxva6fMzYmZ3LEXVvS8I9W31BnqqntblSs2vY98zJPZFb7Wu
mrlHsrcQymog2O8Nzl5hFDc0APGacUiPhCBtmCC4J9bPugK/iTFcZWslqeokjPWF
leb9/3eNq0P0BS6Lbrabe01z4i9JChkdGzkZPwHn871duI7qplmCstPk1Ej2Lr6N
+Vj9P95NbN4wft3zZqerTmJfuteNIgGfRkwnd4HLyEOyy6T7PuH0VroNViDHSUw9
xvQt9Za9SISEOP9QMd6nfbQdnVPxHOb4NkcM8nBUbjWPzMpf116hV3C9M1QrHdMi
/b/3rfWYjrCupdachibB1Ce6umBvAyZVvL6zK/cbfPIh3N4RmmxvhVpvvcLtvhP9
vBshFe8b0xQ2Ih47pqvuMyt6AvBl1OSyPXnprRhaRjZ1U2zTCvMJXUIM4GDqkrIG
Dulou2LK1P9kZo4Ie25tX/85+23JspmgAHdn44ciwwvBYH+tX7MbigZasHSVZkCk
Bg59JwS1zZ7Wiu5Ob0iqPy84N3XIDN4Fcb6g4z6m8MizBRQewfknAZJ3nlcoMoLj
pe23S15fWo1Qg+zWErk978U2450kLkh9htjd3Gtw+QzDVZ6+BIgrHEs5rSf1WiOq
v8NSRIL1ZZwHaTPTBUu7V2dyWXbjO2qf2U7vc4eHXizQRQFfDalCoAC9vDEAOdyJ
4j7arRJ/Dud9riQskq79QywZiMTooDpt1IpH229OYGN3y0/SdZRWwukEUZPsSFsN
Iey5aVOpXqLj9HxqWxrgScGI8d4UPozAX/PjTEIOVUfmAup8lAQvZaMZCMVFbBmA
0WJpqT15irAEPvjY8nWdcQo+eSXF4WGqC3RPw8RbVEpMRCUaamf93vgEyVoo++T3
7YOS8D8kP+PWq14QkDy1T9/2/7ZR8cRey58wSFhCLCzd5xScacTC4Xds1Ildshgc
0J+JuVkSM7W+H+PqhhugxvMxriNIrVcvIixfwgLmwU1gT089CjC8EN1ygPUeGJ30
BAP7RC7m1VDY/i7Jr4hIue74iLD7ZkCaz3zDqCEv6PF7U/Zb288Ybtx6Rc/vUSap
X9FZ4sCL7+pgwgzK8u6suw==
`pragma protect end_protected
