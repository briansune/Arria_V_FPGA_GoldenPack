// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:24 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KPw4ipc0jjGfTRA5OBgIZG/T1XR2VZfj8BBM71zUgCojfmwXfDJAXQobPBdwY5yZ
r0plIvjcl3sQRJ1v2z8DfygE33qHoLd93cZVuQEmqPK+1zg8ZCaKAaiU1qlz3FTU
UEaymSCNu3hQEkXtCKC1OSHB9rvLqDYT+bFgnFnTBz0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3264)
FXoDEXLecj5XCTFoqCbY3AGI/kKQDoB9tkE+xPKfH8aSjGiLJPS/BoZ7kSiLXKW4
t/nT0z0AIn3cVNElRJBppSzHFprzD6Inq2UpH7zDd6mfVlaE13CmFZ8fEcq/Z0yb
ZFOnfSyAkYs5sDj41W6RO2FvTYqmtOyRjBcvoQQsPnsZyLcwCe+GNLEQ492AIyI+
G7K79gJAHg/j41UhCt/bukksnkYQFr1yM/YEynlmojKf5boxk4ybOQChwIREwt/f
haauORJpgJGo/BXW4NbeunMaMnaUFZC1b7NhhI+WKD9XPoyWCroh0k85qaOXwgLn
ngE+m4tZmUHxBys5mTPiL0UC1z1KlUdMRseXvVoBK2vqrWcXG5hL5zwvc85joOra
edK752BQa2aZ9fzt3Xf1Xchgq/TU0LdDX0odd4FX+pXbvnIcSUR695JY4ouM8IDh
5BQ/QI7HTK5ru7WCTjj42RQERKfjRQ2Pzl63OzkN15ViZAj6AvuEmTIOj3RXb4zB
uyj9Kk1fa1kBySS2hFn5UMrcJQZq6nDXSiCQxTlaLP1iCKkRJKUxiy8x8h6iqEJy
gyzUbwee+wryeX7Shy7+hmu6wSARzb6V2ymNg9h6ybE86MbEnlkyctTx4ytIAtdW
C0abHawmxGxhso9BwKu475Beh0Dh0N7I0nDqCrDDftectPis/wT9TQAW5ncttEz+
LZ3Mi8J6TqKz6UebNZpeQkyYm0ylF3SfxMp82MSSVQvJCZP83RM5VIOVIzvar95z
N+ps+Eyps27rCULmP6NDC9vf0x12dscF1i3j2sufiQi1WJdOkH1Q4VdEoQMic50K
tRcYlNbSkYJ1Lc81NivrXf83OJ3udcluzdyBISR0qSGv8MTkn4XVSDxlQfwP2nm4
ZS/i2kUjnCyOJIytzIGjdXGCyjeMuUc6ov8aZf3Z1KBS2l7s8GPuR8f/JqLK1d+N
TgG16CKjQgtG8UofUsiNPKJ6aBu6m65CuiG3WGjf4NuyISeipGz2DIW+K8MD76v2
ZOg7qP8PkESGKgbPPRxvXrkCb0dqHQ2iZ/CMHAAoSoHy9xBeg6hgL7W414K4lcg+
vWQgoQXAELNfyujYSMuDXzPMrWoI2HP3PHkc3raPySMAKyUnAkleCHXVhvpUQ1Q4
bFrhVuQVdiXr/E/D7fPn6f2ECyVdryg6sgiK2GQ14kWM3LZE/HlZiD5bPxvx4S3X
5kd8v8udae+ut6Ds2RHRDRCWtqtEPi/DjznT9wy/BFpRyd7LI4WisZbWLrMCaovC
4ZX8b5lSlpFr7NfTCyV6bJIKQKT9MKVenC//hIahb6DIhdzbnLag8/biAx0E0RGl
t5j6oLtW+ambvbhKHlBqZt7l4C7wQ5CCrFvpVfZrzqJb5rEvvWu7HC0oebefkwWn
VFmM58JlFYLiqG3E5Tej6Xyu1VaMhs7974xGMosGgEWjy/z9IJr77Cov456UJDIf
U5NpNq2PlN206gNjHVUs7NhjNgs9dQvrKCwCjo1xjfrG1mOgFywso0mK0AWYZSGq
k94AsTlLJ1RcIUkGlQlwFMio68mBNRIzatGOV0jaNmsN3wHr//4nLZDldoXxDutN
JCj/2kOF+40qykvfETkPF3gsgue/81Wq2W27k4Gi40BRX+WKFgzhtGjxcnqVtRAS
KDk30qbgG4kCWHsS2i5NFahKgKoYvqFv3ymuxJrt7LTe0bSMAnUVzC9CNNWo2iqn
+kwK3knlCJnv4CymG9/HaCVRVT3r5iBX0ZJE6ghCDRa/f1RT1NnkSC8IgwMbpP+F
QZeKvbVYTIe9Ae3PbOyIUqrzG3zb7R8xXv64Ehq5VGNGUL5O7ufdVC2rCqrD3dmq
kI7p6oQns2UVTOjG4kcRbpTl4DYPUz+HfjZWQ/j6pO8YDEpJvICR5BIvxsxb+Ir2
IgxP4J2QnN+EfZeMThGMYdDvX9/pmYAwh+AfDeCjyQh1wB8qXYdZIveMOO82Eqak
QTax7FybMc5gtXjTj7MyO/eObXom3miAeoQztiSA/cX0EPgbC/OwN8SyEi2MP2pt
9gWuY+qW6zQGWzyjoZXQklUUpos7fDgwQUWx+WmOumj85Bi9n8Hnd9RTnk1ka6VW
tPZ4FEtAsAVFMCPuxCjBhdduQly6wZhl9NJUMXu5RYdqY/kvFV5PwbHlfylTRQ7v
9+B/z6Qf+o/76zbySHlMxE0Uc1n7xE+bsM8NMSk4CQ/6f5QYwgT1dDIozAI4e8e3
YBAENz6AtjijPAXG0kBKMPO0pD0MQ9bFWXD4i0bX5Fdj2FFmXZFWRSN1FkvIgCN8
1AaXK5nJ8/3PbZ0YL2tWBpCRkQLKToBhM8SQZpLJ+C7iBGhTx9LTgcWUdfDzM0kl
vFgaZCPtVoEqMD6ojlAmuHDREZrP/YZRNixXQliYw3gPYmFOq+hzV66d+t18dU1y
3f1qkuLXCNv7A7653xW/f86ygOiZh7Vv3IJ4RpbudC+g8zj6sDVC6uAbyqXCQhaE
y8W8EhjDR9D3iBd6bBGWcqbYZpxOkc+SDgWbOqX7EntxF2RjYXGdSYwQW+kx6LlT
OHHngUFWNpHDd8TToZLmVGhxeQJJd4pB+W4R77RhB/tkGgs0Wvdp1mdickGMYfDr
lCxEN9eEEuMY5z0uaQl6PGgki6y7niZpxL43tJULiUNfi3TfXomizoUFSk2cAyps
2NXgcQ3ofUeqtGshvvLjuspoWZtMYlkL2imaMSHJpTWqSmIe57l8DJivej0ux2y/
drZMOdqWWFhzyr8sok87LXIYkGs8AJtb2cpVzGh+/CtukZNhfV3vOLxF77JIaKv5
4/1bzZx6tcdFHrwkCBBUQJHXu909/EsKytu24S/5GUTmpyvZfOm3yHjIpeykHOxp
33kDyZxdzYvEqGftYSdhUyddVGkkZEjlrjwK64nVRWd7C1dnAlg83sOGP4jpn9xF
6m6qJ5MgIsfv2fPHQFpQ9erTzZO1vTLExQxgMGsQFfLiz1Z53nIbFOGgFSmuGDrw
4GruuS0aoc83fP/+LAiAhd5VnCQjR5ZjvmGYl+7WtS2WBxbNnH8X6gGEB5YJpMrk
APKTwXknv7UHCY1pOPN32VOoPPx4E5vBPf9ZVwNjn35Rs//J5rx34KuV690SYMPx
v/lSWgPwVMvsgVF5bu089ZDbqM0FfaihoZMZ9j5ntqPKNxWzaNzf3z8BQP+/UHsr
YFbPwIKOjDzspf2YYYot+23mTJ5zwZpzSm86qN5YQCrdDu8Xa/kfGJleWEPfVgxp
ts36vsMPUh2hlZohyLh03+unIBK3I/upU6Ovuad7Fjt/P3xr/IBbyNtewTJFm6Xm
VNhQIDz29UbubtMeV/WBQulpnYGz3lJ0Dss8sMEETYNOFebPZGd/4F/umgUSCuIg
EnEjBunLi+nLlcgsfnoOhON5QeeJyXEHfSI4pj78OyISRfWlW0UJ8NENf54yfSPP
rhU0Zmq7QbXbjsyLJ2mIn8GXCpn095wBsFPGItfMC5nqNnt80Dn+4BatdydiuIRh
dZK2N3yGYIjbYiaNr9UQjdc5KGpy962T97xFeXkLa9yYMGoyKI3coA7ZkyTd/eqN
yw195h9P3Oy07pERqAi4MGe/FwkgmhG3+lQatSiW9Z2aWtQVjkAlxj0G4uTZJxKh
5B+2UDs04j/xtQYvZvbZgUzApcKSt+EwD41CnQdYcJK33Y+fQe0t3AzmwR9vZ5oh
0k1MSvZ1zcobZCXPxFdaFhYPkdIRVCBT7IbMhGJEAg+lJKrPcWnanLJVkfkOIZHa
C4mrzKUNn3+l1nMjmliVHKf1ldi6DrU3igIY8ZKkfabfciXZQ1+qeGcGcnN+5sW5
EVBqYR0i3MsUBFtpwGE9hBp6K4CGTxj40cP6GQS7d5l4vzS9QZTFpxyBMjXtxEjj
f1XH3D7QVlSgfVLPyHz58NEw9dRPNQtCd6YFlGZ4wwzu9YW05G9zMVQXbhRE+qds
k/GwDkuLq8rTmkfIc/Y/tpcp/iNS9ST4XGTR7DaSTf1IMphLLHnIARVVCqnTqj+6
GpPW5+FeHgMWlYml/0oUKs/MOMVVKEMF0I/YSAc5dGI4lONDL0xm3CpGy6DiLQFV
l2OSG8bmJRLhYcRzLeypTuUaQu2u1TaDizV+4ecVA23IdC5RRpPFqeKgnEME0BSv
jjYzzM56C4Q7FPZory/m1l6xGSh9+euJyRpzgYXo++LtPAZtXLJMKoQWeUHYlp/Q
+DliFqqukMh9gjG9dqtWB6RHMYsQooS0WXgYMppVYTv38+Llaj6+BAcGyM40/7BG
1Lh3jhX57xkO0aZ/Ev6bGF2Qw1AKJfy4rZ6ExDbyx/1ECrV+m8EajdLCN4jnwhB4
`pragma protect end_protected
