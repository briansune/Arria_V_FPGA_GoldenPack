// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
E1GQ7h6t7RPx+woGqDeLPo3jC8m7IjTDIQ0OAszvcY+cALTSY+x+5NMhjEsNfV3M
vIPfluVS7+eHb77TQL3s6HwBNNideMZLZ0SVQxflKr9ogkt6088HhIzvKkbdxD72
igc9L6dh+GGZ72Z2rTf9YTQlMP1FlOFnRGinM+Zidnc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8304)
fqndsv5FxgxYu+14LZfG8j79FglvHkbW+Pa0wWBDB3lt6V1YJRKdyA7qct4V80Bp
xPRmBri3Y1gP7DvqDg6i8kBXo51RQViOhNxdzsy51ph76HE9Xl1jW2QTAF7JkhLY
cBL4HiGOhsDEUtMjAroyOfzhZDR2QGHHn8fngFmjCUJVKv3wBC/iEbX1YvhAXLJl
61tOmH8jvAmoWSHv/ggd6VtHcqNAkxhvfE4W5k8QDUS7rgTR1tIFjwQswIAYqGrU
WjPhvwOz+MbDzt79oSICuIdEip+1nAxt5Sj+fIXElAaBj3zHh2egNIuI38RYQtIK
OJ1LOJ+io0bPnpHzHzvX3ZF1ZuO6ZDxSFZrLEF8WwoNBBryVdVQVj2vB8RT4d+QP
hTrq57CSohrgnPUOOirttj1iMbzPHvIKV71w+k8lGHRu/Pv+hXVS4ZXW4PTNlq+6
9TWw16C8hpz1jBcensEXbsLxVwYjrxD1i6wM7GC6wGRyaY/jXAW6A+xfkihFarlf
UtyFU6hLA555I6olYh+qXygnwPF8XlS5zLwEwm5KzDLHH5ZhEUMiV032Ni+R74Oy
JLUeJWeNpb7kSFEoc22ZSV5Yv9IlsjaSDWOACBQfL8Shpb5cghtl+eqPA4ATFvn8
g/R7hTQL7dX+l8fu4cYPeNAP2CFguBaNYAErVhFnd9oAfNUF7jIh/VfT8xBQN6cM
7ope0Fe6dpuCDQcjWvRl/AtMNPwBn5YK3/4rLWDl2hadTBY+VtT5eldoWYJeRVg9
2A30C82PMP/gLWjnQbi4OY2THbAYqDYrdgJamNcKm+JmqzJ9PqyGNRAji49v5x1g
xMrMLi4vBzN9bLPTj+3CxyEatoZYEY+cyHBmmR2fSbM1FGVB4aaOHRBTwe64mClM
KaDEUg6ZfVmkKvC96tKgYbgLVM9RC7mOt0eZ79cMyd4xdvjYKcPOT/qC3HDksmTo
HnWr/2g65N+DaZGUWMAGDu9cpNhZFwvz3d+iY355cFpGlahn/QzPcYb5viLLqUkc
XiGXphmy4txMFjX5Wgb5gELYOYDZwLWWrX2JcRbBlb+qH8xzlDTPpaFn4GlUuvj3
VB8sMzO7NcDipZu+0zVPIxw/EiscwKE9fGMEZeg/MWKCgBycyC5l2VrkN+QvuKLd
zeKvYLTEczCHlGCzK8RIz1+BvuHvNXW8VaKdORrL+9yTwHRY3K42UHMysA9OwnyO
JbnxNzicBThRmj8leuWuvHl6T4nmC7ZC7HkrKTCunkLA3FJuaK9F1TzCjGGKWaNm
L3Q3jN3sAWnKeWO/YepdAXGIyQc0vl2p7Yzmgpo3Bxpqlo92CjPslOq+5nRB/Ht2
nMfWrKUkztTpKdOAbf5k3ZCqJKxNBEP53taP94SGHAQG5F9dewo0s875LcmHOsGW
3QWNjyzDWBJ3BAmVxJGd9fop8oRRaMsz3Fgyo2IuYDlt1hiW6q5ntEMFvnVG2m8z
kQ79inyAe/2mhW87hG56kgyAZIXGBzEuNHNndKLzTRsft6Reox/WsJ4eSJJ0SKrH
waqTdtdSFlzwsOXvFWJV1ZOlI4YwBeMdTqhBx/hMBHZ1oEOlXuS7z2ZeUN12PH/L
mKwGtY5XAyNr6blfJZQk7dbhGQsLDNpi8uzrewGnNvfn+Zahg0taLG77XhcHggmL
st3azK6q5U+OCwKu9DjCEKFIlrkHg8yPPEyXmLHtuBtnO70/+UVBveTLj49X1ndY
IdJf+4wMBb9hKn+63FfZJsU2eFQS7pIiJKqkispVEZt7sjbQ1LRaqbRZ22fTXtEO
8mWX6eIpcu+uuzmjnQiyTZouLpdWgeco13zNZXKHu97vVY7CnbWD0pMZVTTuQ0qE
Q1qMxKssAXyLw2tIueOFSWteNgPUXimIznZ6f5EIFMqmqLg6Ddrg8Aj2dkwzzeaK
2vRKrMEvLi+dLuEJ5JcPNPwJHybjkoVjWzgvVmOunGhJL0p2L4tji931d7IZUxPE
TXIj/HSowEiC0+E89ZQpfMiAbkAd0sZAcVwmXhSmW05Ha3ZK3fAUzxjKwfuYfzgZ
tPz0rCx8k0hCLDqCnc+LjVAhx8bW0O8chYwi4HiKeuckfwmmlRokc2mVR5Vgi1pU
FBZxEK46S5aT8sJEXANLvmcEY/flib1jQuK3sVPYRUJ1kmKVSiG9gSbij1IIDYsj
ntJEx2WwbC33wdpf40zP2B349fjx+CzM0qYL2RCZN7F1kU7G3nvaFWJNi4Vz06S0
7/HSFgokjTaYO0Xwan0i75V+k1e35JkAWtTy2Wm9MtmBBb0QggGqKioZ6+RyyJKW
lW7P9dn9dQdrSAo4CFrjycFudwLD3kvFnzMMpPBIahcOzIWkuVPGb/vsD93J1Y+l
fZYaaJ8A3i6WvGVA4Hj0Nr8BR9p0ulbrsaDx172asCRgvTxVdWiPKVIabhV1yQYD
AZazvjlPC9gp12JFOGplXIov9ofV4JXiFopOyQH6bHbGGysffbDl409oJleYKhes
MNVC/g0RJ3h83R45IfpfyMBMcDvrkaBz41n7sHCMTIaPS/TPLcXNr0q0nPeGEVbe
rn0nKrFpR29kmVDnz5+5vBPowtni5U/IjJlnn//MYVVkOd2J2/NTXowFXmtFH/xE
wLEqj6+McF9xU2BN/XIx88uFz3T+qeBsjcTCMDOPuYnXtnoo3jnJwsYiY460Iz/L
5DSGtQ5X34fxF0X7RUaOfHcSicN3nXRhmxrPfWTfLCwGtXaznzPANf4kPcB4JSz6
Zw7tKCdsI6VsXUL6VT23chTBcAyMTDcZ7Z3DdgiHjuadocmn+Dz+mrXF/0MpefmB
U1txugHE2deNhkV0dQGY99MFP2nYb7gP7Befz9wtuTzPCe2WL+fCwk11bk0B/ty5
7CQitzCuGsEfnG8zI9B+trCDv5/LpttqZyT2z2Tv3jFEjjIy/bnytoc0RHJJz7FU
dlMdcz3mLng0QywLL/3vfRV8Kb8PPsp0QzfdBThUttdRpCRV2bPGzrmD+jPDQtGN
ok/E1HcX9s/PXiBC+wtf6hbWMnHWn+SF240TJl7PH0nuMR8Edu6cw2jRRwc7Sllo
3CngacdIESQXeBy8OAtWvS3fraherDCIi3eiv8r6xhsb6+fRsLbqCGSGpICmo2nN
wv7aM4iw00Jplrxg4HLO5EQVOmwp3DnZXOU69yPyoloPwXOvk9QyK9HwFE/9c621
KnQG8stU1KIwlmbEZZR6AIAdlGbvEkqRwwzWhCsbAkR7sV721j3olq1ns9qa7esy
G/yYc4Wv6MJnW7Y7Q6oo2v35pW8cPu6Uc7ZShmEVv6KPyv8bkVnruPo8xjiwBv4P
gF11ysDGAuVIq1fclks1xOZSl8nvo/4iz6aB1qIEBTaqKl/7W/RmO9w7l+uJpzrm
zGUrWflMeMPXx2jLfpAe+GiQFyENWGJnFa7zVQhGOzLSYSKyi7YrqsQdhxO078qh
mrzUTXZNYqmpTpC12yD4604vDgQV8g3ZS0v/N5q9uPglbErdEZKMT9hNMU2EKFFp
5YvED2KMFCJAWc04BkXvzrvZSDnMELorvam7wcgAQGxuTyaDEdkM9Jq3/vsJ1pw5
Mnsr2fm2KZGIikz7O0Or2Gj4rlBJHlOu9ckAHjff5SjhTJ1SaK+utIpS38ewSGEp
ycBNOOF4fP3DQbuloyfVLezu1S5bDg8SrHe9k3kKlStnfPWosui6aWkORts14BhY
0cDxqfp8L6C1fhDBTe8y5XS/LHUr5vMv2Sl1UaiyyC441CJO2eFoy54juyEGBaKX
1pEPOz+mpxYvy6KlHvC8tj3of7lKY8l5jHCXfk/x8Tx6PGPKlUhLDCckYgHmdDkI
TE7tZovhDlu3yV1jFyuP9PulBkNiWo6bL49vS8ctrobaMyrAlGrLRL1jg499eAXn
ls/cqcW/SgfneSXsT8vU/U6oajeb1CU7+KWgedG1f5RcNLU+Vpetlot5IG7PQZQn
BS7OKwUxUWxUMpM2d76v+6a6/v1Wxt89iItWOf5a322J4XXJ9R9MyCOdT4MYkpvI
Q/mZvy1IuECUBGW1YyY5y+/qVleV5zn7q5AfswD/6skcIgRF0xIgft5RqqSPydXy
b+5DRX32nSPsG5ZnYraV5HYnF+cwVUjM/OE2CL1aOR0HfetkBkAK7i0k9l+CpjVs
JKYb2xqbgLhmxamImfbReqHDCcLY8jr1FwFsPnLBsF1wtQ7XQtIW8mHSbasYzTXO
n6GiBN/a55+MvWL8YWKXAFVdK/oSzop9EoFG9FANXKEQZBcMSlapcQGk++00mNSK
Awu0VeWP+NFHZHmCuPaEXbonjpQLxaJbr6yIcTFY23siLEgBiO8FKaMFDaeYP02L
MQg211pSUAz0PoCB1WQh1nQObvpjdlIENRoLmsAq0Nyz60OTX3wBM0gZ1IkK9dqz
dbBsX/GKapf85U+zi0UY3qy/5k6ph+8GtBqHs8F9g9H6KQliLjZVtff+ZjHFqkNG
aGj6ZImQOcF2W/okCqRXXnoGL8XOx1kz4Cx+AQ0BDuwMqyjlwhjYPrPBDoI+YttO
inPsXbep80BJddAPtRJmmgAxHkpCS8RQ+i18oXSCquRANANpy5O9zni9ytsFlUR4
pNJhkHwfyxCRRz9wWGNr8hbvGwr6T/9wyhOdE/KjbdXDmUxExtkYAeaUCSujy0i8
MxX0DNenruplIJadePDkU7/kTN3KPLPlxMZPGxWR7BWOJNeKiKaDC1Zba03qjHDE
n6GQAsaB2rd8ayQwWfzgugHYif3Qwe8GFglm3L9uY/+mqsmc/dTvwtyyYLrZSt8r
++gDY2J2arYvjLL5lr8D64B7Dzk8YX58DcdoP2nLb7DF6VeuV7twb57qDFs4GOu3
fPpZLXV87FgO0nV78XVs510tiEsnkak8AjAu2NTVHJAaLlrQPbnzFhMKQk0USSUH
uen/5+M85n/U5PzK7ti7BzJIVd+R+/2rm9CMerXIfhiQhpUGdFzgbHCbJeg1YI36
H+SKFg65uzQqSDf3GcIlSnKZ9cxZBOhjdUaoA1J7YLgS63hMDQjeuwhiQgpzbE2A
av/58lYgca9YqBIcfxkFDLII1Sp9mDZ6RF7hfKF+CNr1wj5DX6Ras4hCYaut29fy
PhdlrZwIdtB/ZpPbsScKiJSWmO5dMYAw0M9eji3+70JNjEqSWDFb0nzkNk1ELyKS
xvhSzDtWf0x/k4d2qbCXOLOE4YzneAXqY7HzeZDqjwn2kygksThVzeyE+6XnpPG3
NUfzxJ2QKl4KyofW55Ph2CVWabpr7IO9t0FJsGfkDZxTQUfLKPBTEGSauMNA3lli
tSFq4GI9qHSCsDnx/iGpZYlCbLs9c/SdGtJ2/hKvybWyYw7PdwDzEjuUx2hcb6y3
SJB6M9Jijyn+3J+0AjQ2Cqjslupi1LZQk1TO43irY6Avke955ckM0VDTYq7f7JbE
fPMqGNIppQSGRZUbOlIfg5lMR3hXulapI7rAlA4y5PZCe23c2afuRopqPc1NVw6n
ToqdQPivAf961ywFCbizEnLCcE25eV/nsF3fH8oS6U2LTZeDzTqkH6UlbKfcBE9G
hUnXAka4TrYGOVamYT9G3ZMDD+BsSqzga6QP1eai1IP0fPvDy5Lzl0pNyT314Ut4
9wBPYoE+TJC/+3m4h4eWx6vAnaf44onJk8Rm+97h0IAen6CE8ze59x0913H9kHAs
E9Nkn3XOMfl5+KzAtVPY9bhn5hliTFl9mrcZNtDA7l9z0IBaPinPCC1GZrZwfbfs
Kej86e65/tlZ+uoMJwCzZ0NTx9FmCFFFr4ah+Kp7nuKLkM2KgfbqxsG25ZpfKOYd
Wv1o/Llig1eO/9kUmDKKgz/3ii+MZTXYmD9vwr5JNmwkKpf42I6BA5lovCyeFhYp
zYO+t/8OahJJx/Nstk7yPBri2Iz+FHrC03ZQmtmahrmRnU7AW3v4vG5wdFLNc7MP
tAvCvJKB/nfQVWhfoS0cqaxHW6NfEQZXuednHoUyrR7IUTjQd4H1wwqG5mmWX0i/
eBSDwRia2InBIePMuiMZXZFM/HGimMUMb4jA4d455KW990OWonm0Oyxe2VPJeAZP
KzLVUVtLN/n+0cpwI7ZtFtTenMpXpItGQg+gpt3AxOdL7iWbjwGYhwi2o7LedMni
ZmLUIrrwjUW/ju0NZkYYB6Fk5/6JkKLjvr1dznOmvjYZvbJ+u/k5BdRla0qhl58U
8ykkLEoC3R8MYijWWN+KGDOPcc81LeGWLOyHoURiikRgMFS+9scWG4//H3tQtFbJ
kSWtxcZLl13+aD/U/slUSrhen8AoOPjv9dM5DMtx0rnHy8giSxd0G0fD3BsCM8sU
GZH+d/27bx5qgzNWpMSSpbbVeT5aNU9GY8cVSKwzmwdP4VI/nSfW9dZNAE93RluR
IOsRcQQQJIKpx6JTfrCvIOTre+IQYKxvk6HMVxJx/FcgZywI+cK36kHPS//QiIxC
UQHEcaoLzry/VPMwO2//nL4FAStAbBFo7joVAjYdjaMrjaYDv6c8ngDFjNmdMMzs
SQcU0qGjc05r0MNNENdpS15XFB/DgohOSjTAJc9EyBQ6ju5b1a8iNCD6U9r16Cai
sSAIZHaL4LU13CBaWYuRusjYff43SlCOfczV5xtM2yAca+GHPbi9eDb2DLGBd+rF
VZwK3/LXCFecjFOu8xJP7BXT18mQ2V5QElWqjiirzTH5BpyyCboXcIYE3UFaaEEP
8QUv+PCo9/iBR3Gra3oiA9uu1/6NbDWVd4hnTYl1A24e0CnrGJ50T3Q4eSmt9pTV
pmlr7RRs3HgxeJGHo00Xm2MfMYDIEeunP+g+CBxep6DP+oDP/OYLmQ90GZjCXIGu
n4+vqCZI4H52nMijUvM3x1Q9HCnarPSROtaT/Ap7BQxmDhR6wfxBB72jXK/2PlRP
5MZGQWtEgO/GlslGu9Uoye8luh60gbI5KRuYb0Mm+qdDU7+LjdE7xQfvWU0xHKAz
J2y/cykvafIlHXOdCcRndd8EdQu0tj17WyH7JSKk3tCU2siYCjgFczLL8ik9qbGi
SymPbRUZURbaVFePJ06TgeOQi/AMMsU9PVH12tc2fKwJBqQqrqJYKqnuRXSK9wIr
A8J8WXU2DChJSazPe/pgI6t5WqbNwDpJgYDOS6sFJd7wXHxf47bKNsXBx2PdDgOb
lUYvzaAQUYb0O2RcKMGDTutnl+JK3qh9phAep40h/kYHrM96vjklh2o9N6K9pAWs
8B8BRdy5gIB/yC7tRMMVhmSSxnme3xoyJ3Qs1fRg/FEeI6V9JEHGJd7kyyz0LAb+
ELNI3A6ZilarRd8xiqzzw1aHZfqfdZP9nfkRTyrOsOThukuL7QO0KQolmYkALKAr
XLq97+rfd8PmGrj0Nmxg6w/q0fB8mLkhmZxHll18Efp4StTUP6Qj/5zy/xHJzNPl
u3ZQUACFXwnsTIfLb7Es9NxRaiGe1DkjosqLi/9CoGIN7kxqBsXkPoYFkLKner5f
l0PX3ckR8/zvhumfXQrIiXTG5/xRcjFOigVYAIaBbGGX8um1/INRhICZU4wi70fW
PCgaG3FSkwJEDR43Dc3Ngi3OxA41pZIYQ6I0EWW8hVHe7Rg3zWXvehX7n1Rd0sMX
nZtfzcpz1ixg0bHpxfLaI2jThtU5EEpaz9ZWVJM9M7frf/vppixk3FXhQ3sOk0Tg
jlkMah+EI6mYg9UISbikessHr0AYvPwIejvue0qIAwRQyzKqi5RAay28RI8oJ6bx
bt8lMqj8hBB1DoOCaPEf5WYNZ5FLlUUB/qKnWJEdUxTWuBwrZuU7SvidWVBhjgI0
dinWKPePJI+pyW/wU9V6z6P7iEM8s+7+wJPexmFiZ0iOex56/Ahz5Mrlr3tYkV6q
LLCnNelLGcWQrCx6/VfY0CwS0yGH/D+4DHk3R8Kj8C8ruqSHNB/nS7RsU08VsBD5
a3PU/RZ9ySrIO5I8vNFdwJ9w9tfHcuzVr5pDhzXwuZDpTa8NTK8TYjw6YK2VFsMB
jP7UZ05MiyNxT5DnmWGwzwdd0wRpHHeI2dvfxDB0+Ha2O1Hm118G5LHr6QLQjdX8
tIzDmYYkXIwdHCUVt4hEeTQX0XS+ZTAbrkngrf7H4quot//6OWTj933nautlRji+
MoE2IDxWqMxcvLPfGVSkixhnCxYbHnH7WL0Xz3Gc56G2DBJJqgQchChFHM8qesAr
8WKB1at+SmP3aQKrPbIh3iN1/59HmROUkNLDto8gLT1AfFQn7wrd2pNOePQD9wZN
QBMvq2aq819c2BIw33YYrixdA/gKhA/fUjRlO5vMnjpJar2oouXeFg+j6CseY5WH
NvFO+0ZNRu4aRki0XOfkqwPk4LOPp1C9/Ubm/KGaKNYzybJ88J/zpNVx7WAi+nl5
L9nAsXBjlZJM71ImRNqr2Qf5+F+OyUmeN7R3+jTcNgqmWnn/CmL3EPQ7sPRicAV0
XTPLSuBVYC3VCSEHwkoq9/A7kqdBBCYH1UKqVZ/vRUK4Jnopt8M8Q9QVH6zwREtb
//RvxjcRj2mDLn2XOIGQaKYw9fGMREEctUxFqZ1ImEk6Sc064FD3YWQ81PXUkqtJ
rZm5SIGsMyHp9Biik/yDTk+OjbNXfgzbhX4GsNOyYIyP9wwpBIAayqFYMp3q+WPQ
Gn1bYDHAcclKPqPwqA+yIXQq2RXsawEuxkDfTtopjpOcu1pirS7qb9ir1LCwdFJE
GzFeYa87TBOOdt6amMO8pQzqQwvTdZovioTRRTt87F+yk5kb3vNaYd3CvUK0IB70
EdVyk18goyC8Ky+okguPS7tw0ARuBqD/t5boR3UPdrkqvzU4wuitqWJG2/QJIqzI
u+IczJ4i9fLB2jvD9If3GFHHeSGGymaCKH5iaHJfqT5T8iaaLldkMFca80ZBj81B
UiCfqNZkj0bxNhBCMwirVtfsPEiq8vpxbugyVv/4giukAiaIFtEtoC2GvCSQ2vcm
W71ec3r2QrGxiL7TTXl7oC8FQfQqJ4tbSVmdfPd3yL4x8B0D3DuVihX6KpO+HekS
gi+dsnW6u1q+GDfDrRvJxj3ORCNV384IfjClBw56j1NBHElCBjO36OcOk0wL1fU7
HHC2hmDmo500bPR3la7VeoHVVYV2KEhmlnuim80dWC92HQMn284smSYD6sISaOo4
XXqEIjuheCRYv/1hrlxC9TWhPJe3iWD0KyVOeZAEyflq7HYRiiMaUoZGQDmKTKI5
Xnbh/94Fjnjgnz5z0MmeVumFT2FmHivwRGVkigUyRDjB0CrqiGN1ZMrBhkmwVFPT
KX9PG/RYi4HjuF6ves6/HfIRfQebyVjCOzyTE1C0TFFD0PMa2CxJ/URxPRUIyHZB
RXokER2MOLZqVIko+X9X8cTK5B56UgaWIwE2srwVUKcT4U12atVW+yDR/NNJWm7G
A7e/YBhzA5arKBv7dGDEdrzBGQi2JfAPIbVZLZQwscSPcNcqJsFotZ4bXHhySHI6
eHMRrmphNRBygUu4IzVcrqCBxKB9nijwLQ2USC5ndVODsJdq+d0y+60IV1mIzDdB
I6GURwBKmlYZOtKFgH8Fd8VdWiW285N5VPdpBSaGJsk6oo4f/bTT4a7Bwuq1aC67
WkbeocMUP3QeVCnGg9a3O0WE6g3nVzcIzRLS4avRUsYPMOzVphfm2ZpYluLntOCf
rZJAIIMArVX1DBFWv94yiv0+Du9d/vVMkw5fePcNKyqy39oiG/E6jAPa25A/XkFX
mupaaJX31hA6WiH65g5EM9x8AcseCMMJVRDLvCsvJWbQkQHzspnlt4YX8MftLM2z
fLEJExnvkWi9HCYF4KN/v4PTrOYtGHPfEYSX9N+FbG3wRJKUSGE9ds7fb7aLcEMi
nEqjqUn9BjutZEd5fxqqBuiITWmmSnH97EQCtvTU+qyl2gbuH/3Ev96MQs5eT9nz
OMro5LWEiKp2+X4oguzh7qzzr0A4JI2ce812+LC07QGpeTxAHW3sqStdg7Mh7cuc
cq5aTuOw4LexhQsAz8VFEd498l5sAY3jSKmgqqBoe9yDinQVp27uiHBEHA3S0fMe
i8zIBWVUZDLnLzOkhySey6TMInAIQXHy6Bw1T0cHBz9TsM76oxWzfx3xgX+7CZle
lASMXk5fLrbhmcTToV2hYvbd9BTEtjH/Uw4MTWQ2pL4gxskwLldMHY3ruIoQQhUJ
ktWdk3gATzGaaSWNMHN9d8Ji4i4f0RyCuRo78ui/qtJccZB3t8ZhzBghG3KKqJO3
6GQCMygdOgg60LP47qGY1wfGhvVWyK7dJ01lq8zGa6y6sVyIFg3wmsgyzk+Q75ux
zXvkWY1WJj3ZfNlW7ucZa3vEe+ozvSz0ymxoG81wIFE8xRRqp1UbamkTnCotqBgb
lc+EUf6l3f2uWrhJsmLTqafVjzDSTGhk7vjWQpt3iJ45N6rZmOZytm1XTbMdt9kX
PmrWvlU0wjOcA/lzgqrwCSONvStpNr+CxWadxhOG93QSappY0Gy6xeVdgkq2t1az
a1CBrMjxokWnXLxqrSU//0lPlgrMQzcpMmYO3QKGAVwFSJ7L9LStMxwvnTyOBGpW
OAP9uw4eDCHlGAIQY8M5jyNmarN+a0oYpCyd5m+azib5XBcRlQ17piFZJCnRWKT9
8MUBX60jIi5kBX965Gi/jYvZmPaIWe/k8WMsZhy0oX+yzEdemKpigoSJ1uKZt0A+
fm1r59yDDvYfbr3z7dEEbg6dNtXqOoo8k9m283CKYeOCt90slF20qePIVAySUheB
dRIPChEptWYc1wyPwIuBLnDtuSDCRVK0ay/gUk4wf9lqux7G+hUnv8j1+voo8FMh
5+ieo/FRlUkRkc+RoOx12ijH7WF6VplEq8UmRufB+l2QZ5Nt90CTczuHhnvS08rr
kWlS/27skLY64TKb/84NeMGNUR8nI8VqQKkHq6WAYk+9qvWX4d3eQgdLlTAHyHuE
fjgy6Z6bi/+fvlaW1lJOiWsD2BmxA9fI1e25t2pTewL285EE9Uc3I8FJ9knG6GWA
NETbnDTDyTISNnzsCiHTVE2rJVLSKo+n0WCRQaGH3lbQOGgx+/uDtmk6zBZgoP/G
`pragma protect end_protected
