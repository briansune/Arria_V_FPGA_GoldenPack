// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:21 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TVgB2Xd+tMPejcNkQXeo+YN6kQqJZPUj79HVlYKK5p+q+rk4/gSbuH0szk2xH+r1
24tlVGiomdPwuA7p18RqvMGRUJE53B7JCeM5K5MW0MTdSXMhav1D5W9qxsQW+weQ
l2jMBzsdHvfrauCObEtfqy/Eqo2X1PwC4TsRlrhs0tU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15680)
HigBz+7zbbTnWpw51m0eIbMJEGt9Fzw3N5wEElffhJCdTiFLCiYzmGEMMI0LvuY1
5Go7gpDD59ZJ1Joh1tUdG6J4WaTj/KUKBeYZNmwOx3Emh5itkzY2g03VzlbLRY4+
dqPulxcfatvF/576AMj4DdHwV0BL5woxe72Dtax99CarelLdAjW9qIwWZPQ1sZ9l
5gyulaRHYxLiVdcuGp/LFLqBnn+OksZ1MHZZ+9QqqQIlqkanW0Waw6bxNj4bTzXn
zDzKMrSlEvlxLuOPTY8Qx69UG9juDcE9ieru5aEGQL8Yi8oWlXaEU2YTO6e7gFG2
/wvO4wla46er7dKEj1G2Xx9NhU4+PYfZM2oTYOdil6W7Erx7P/9eivg8sZFsaMjH
kxgRlwnCVAI8O4+umKP9keCJaHV0CedqCvH2KiyzmT440mTH0GclDpvfcU9uL9UO
wYZ8GyVdS0281zuazg4zaNE+1X32H6Eq4jln3H9uX2SP6ZDlVYM5DIBAn3qwl9rJ
EyZf6BVqNlLiUHBQRl8lDQVYL/W2skN/qjhmzYZMjf6Bggm323k5ejpyDtnpOCVl
kEhBfh1urYEcMLlmMd5IM4P670gpgTuQDJfGXdIN+qQuhj28LET9eYp+lhbcAKdq
41r7S4X+ksDJRliXV3z5BdJSp/q9YReETpw+7EqLf+c5+svpGAw59e0tOSWxnANt
4FL4BnvKyoTkiIMsDA09+V3WAifuVzSTE1n14RuwF455R1gQxsRU00HZtXhj4W8C
zkaVqZX0KJ0tlHLHMFqxoFQBEoXC6fi7Q2z0CqX3QK2wD7WLlA3vUI2B4dYtMx98
G/uIb/GCiQw3pSIy/uquosZXAYex7irU55ZDfIgNRvI9MLvLU+FVUcXg2gCRAAnA
13zrtVql7N7gvpCxYFeoMT4e8SMz0GEyIp8g6FJJzqpPJoccdDytncgKC3UjmrwQ
sR0YwAs/6Ld9Sa4EwJnYnZbSLKSs4jRiGXsslR5RgxE/T7WzLDNB98Bqc3Tp3wop
57kktkDKpYDfl7LVUCJVPObpVwUHBkFg1VVaCqUZxaekffoCSg1GtKH9SPWDsKnj
XcNmkc7M8haNcDnFGNMDqzcyN2UiWPDWbHx3nJGVw1AWFcfHpaSHKtD9b/WfGf7H
3CmXOMvkJkfAJIbx9kbd5u03eBp26y56ZtfwFX6Ee6jUFfhpKpH6JO3osoCqVuxs
oAjDIJzlY88bK/1EYqT3otjKn9SvT6B0UL40C2zMhJ66UnKM55ByJ/gN6xKqwWRL
TgqBU/nREL8DN2pHmH701KasaFKrfSH4P/wimqrDbvC3cBb2wuEfqIBPm4axseCT
jm4bJOmoYqpbOX22hbL71Xrg69mMlDs86WHwJrQU7JJasagZXMYqp65E5s83ANvC
9LzSEjj7dR3W4XwWL9Yy1pvmQ/XEV9ZTZRUja43SkbYlSC8/InrPfHT2tIfA/QYU
0ZwtAavKUz7z35ruPDpf1+U1eRblnNzFzPcy4ixyknHlwAjUaHPdpWqfagr67JyQ
Ta1K4o9b6ATfZSchCrGAauw3I4AvcAR7MD4hIE8jUp5H1ZW2bzFc+0+CeOH0PpWU
wHHaFTQ9plAmJJ/s5w7rrT4BfWT+rE6fFyqm3uy+qc5G9l1iQrAtsAQqppzxcf9u
Ix6TkTGFYAcgQ2cMUaoh2J722d/CMa4VWwawP9c3Mv+VSfEQ9zsSp5hg3pMHr3Ny
o5pW1DXishSDNECpUBNV9Nm+V3Okdss9tAS0GGLviMBa/HfiwkkeBEvLqvw6vEq+
EcHMsqnvt3viMS/3pR4vdXQvWXxA9qq7kFhu0bxrM4gKIILqKhdpXEaEAaEFmnqd
xFxEi2DF6AaV6qYlIMDRWjF+dawygE7DLymoPlF7Jb0pwtcGMejLufMOhNoB4YZ1
W8efIYkn0Bo5MAolNdcZFI04oiP1LRBidqRhdCDvIBbVNUugn0lwpoTo4UiP516n
MKWVgVVVLshNA82VOmj1gz5FlJn3c5FnjISw+MnnbxvCwRlSuZTuvM09EteaojDp
366jKwkauYHO6xQP91m0n0/AmuXQsPd7KBdmel84kUbyzyUj6qefqYFyzH+2xKsu
vsjYmux8cJz0DyCwQKFyE+v+IosIrQr0Vu9ISMYb7cYxJ+6h61MEOfiYPN9JoqlB
3wWdQWryZC/jTTYHUOfxBWtHwgYrduXbjrnd7hPNQv8p3yv8ELD335p1vNOgN0GE
SGcw9ZejvYOdOJ6wgYWJgVi+ZsoznyCK298T7FJ0tvlmeAr09pXSqC9vwbL0AkjW
eYhmRVqrnSMdDbj9lm2SKpUSNfhIJkJcPhrW57SsFblT1wCKaqMo/FnKVYjM6sFe
Z0n25d+bk02nwJpIyMyi50T8uV+Z8VuXvlnrKBP71zrpPTBfi50yLoh1hXgDDPX5
8kX8cSC1RI/GPseuOEhkhhgpt2l38JHvGIZbvDOFr5J+n7LdRu1QufL9ZBbgezx7
cXJp9goYQ3SnJt6VEDtfE1qaNtQMNQFmHDRgVsQyilTp/jxPIF25CqvgnxFM+Mbi
MkQbDfUFlvwl7GIwY7ymhPFvjzzKRYWSHUrfqqhS9kX9kuEvd3uNk2lNEGpW2gQt
CBXBQXul+E/NxWQEYoASlN2/QzPpQBeuxC8UIwn2eGTNubMXnGtFiyTtRngXJuV+
wCs1JQ0vLlWYii3QVUHZMhThZQfqry0Y+7rOp+tZ/Hu+5oAHHqOL9cZLSDs8A5u9
EsUmElV0i054QfjdpGhLoE1D2rLvu5oTbSQmLm3Vt0dFSqiriAPsv3xHXFOlIJ2X
2R5PHENJKe7tYb+W0v8tAbwEpB5N3Z6mljMeUZSXPOZH5O7YRalfFRgFFVXVv5P9
LsCNl8bJEwGYSyqM2WHEQrkEt4raKlkBsB23cPTMuU3kujxcfbJVlmpbxvc5dO9L
u8osjccIKw8+E1kV3JE5dg3D6U1uztTLa0JMC9rlDhAxi60zIK/mOHPy6o2yS8SY
D5mZcU0Wmb6xyvqXS3cxJu/H52ssEywAFO/lDBAmJVWmt07QqnT4fWj7PSDgvb+d
Xaz5rElhU9qgyIwVcL5AuekNxozt+o+6aTigURmKbrK5ONeyBGytuQF1cqqjjZ2I
+OHwEgK8ZEQziCQ2KJu2AmdqE2v7AycIcnH4b1VCFMfjF7EdKnCw0DG4uO7hw+pu
DFnJO3eVg7EU16gMWDoUsrAXgPMjBW49Ls3/nCVSzgpYzjsfzEhkhUHchcIhMd0l
oZWz8SjSt4mCs++WJ7vIYoHy7IaS2m6aZ5i9ba/+57Vwo/qvhnKvt3FPiG/B/NSF
lGdZbBpELNdWCJiXrYWSPtKwmA3GkQ1Fua+XW5dD28Emrj1S8q1nj7ORfjQjMvWp
CGyneqidHwqICJMjBkxO0uGuOS+g+F3R7G/qk+m+TF4fLirnrikElvohE4Gslao5
whw0Ro97ct5wSUJquc2QZ6lEVqxn8PC9YBbLm1j1ZFcp1mXPbTZo+2xYw09vu8uc
bRvC71XjWkEFhJcydVAeV+xePEbkGJzjxTvu+K7SlV04+3DoSoV4zppeXUVR9Jqy
gg0DFcxCwEAeyYKHeRn9BizjrW25ea64CE0WA1dl9dZ/24R2R6V69SMJjccPPHhc
wOsw/4ffVcO/zg1vZHRuHi2mnDL7KQZvS3EaSUTS+J594NBCW6Ct7Jxu7z1fe2+9
tOYcz8T7wnaF34KWLDF+MRrbNiNHW0wGx+POT2xD/PbYAApcYbU1bp39WdmG/7Vj
xtM+RCcAHJkGw5YvtY7FoM/cMVjJi8cJ/Kt4HmKnYGP5TSnvAc+TkYDaTNPBzuA4
jSA3M5n5CO+pbo3f2zRXk2ev7FZww1s5KKYKJ6DIWA9fIBC6zQMn31AWsVvxpB8X
yMCl3BUBaQ8U2z693DOwa0Dihor7gb+P+8jX7Tc9OZc1a91JCeq7/fizBxfIWxcn
zadyoJhn0qjS75JdPGkpCr+Bm3aDv/nT50iVc47L8/s8tPCRNHd2zKWJva/CdPON
5Il8w1OdfJUiGtXot76On9IQcxXyatZ0jGXufxwLIK5YTGIgLJOxnSXo/J8CQjKf
bQdqde7xqo/5W86voggAQ53QgCORK02gFkLXHRboQRjAOH68kZrGgXzrTVk7mtdc
hSVLJm0rBgqxAM/5t0cBA9gefVx6FKcKdxxCmJ27Ddv1ABVTaJtPK4akzvXbMCoj
EDJnxOW/civJkIHRdPdRH01nBN8yCl62zeI5k/AE7Myid6zjydviZ5sOfHh4cdVO
A/VM0eP5FU9jMcRpvHknJd1HBC6htGsyqs2iUqCpZwuvRXYvzKbg/UQiT6vg1L3i
D3swSQPPTH0kF3Q8InFwilQCEH77AiraZWHkA7FJrLxwnNzIsAyvZtF6teWH2Jdx
hdWZgALxCsPgGzCUW32r6QMMPQOy1Hc9xbpflkTCGe9anFM3G0H6fm2pM9G9vOy6
lFazVP4OTI5fv956K2pJSayBv/GGukunZDzfCJuATF6Cps2f12tc66hra/rbqSKS
/4tvl0rjXU7LGdQUCWIIRk7xZqaR8bVSIqKoHQByTox+gMC+pGMUCjaqAGzEmW0w
F5RIWL31i6Q8rtc7zENWNlwRmAUzq4LL9jO4oxzwv4NHMZpJsZmP1cClDpq5eJIa
r2rb1aNfk2CYIPIuJuEqkcSocS8Jr822A/IiCWMJiBzZdYWg+LWhgXtY2GSSgRff
Ol+RgJFjyXzndjFW/HtZF0uM9V9OGFAM82G/Dl6oxM4gA3KiNFV6an+Tg2M+27VR
h1hIDoqfItm+47tTspf4i/BdOg5rus4kjPXcj5g65omDcWZUkvltpepSbNmNiJAb
m6yfM2KOKnCEoh+pNgWFAggwrcGdcwt2wq2W5GMGmHFqGKrvicvVaOMcO+C79SSz
MeK8Tk9QOfsnQi4fkni/LnKPTSKQEtgy06IvLzVGay7Pb1Z2BIwaVCPE8VjOdAoU
GZX7QHYru4D5jNS6iEMoNOgQ2NN2NTA1lWuVtPFP1NwOCEbeNXkIOs69EuaujRrt
offQEZHcmG7fOxirOrD1ls1S5tUlegWSeiJV9QpRy4C8Coz+RMHWPMes0ppqkgRM
Pwb2tfiHOGJRDJAjfCBzd8DKlEAQfe/x9Pn1E4gR+jtyNgntv0ycElFsGjjQJcsK
uZIWBR9GSu55ZnQroxw1ickbO6pTsZdKORJTz+y/z4mSIM4NPQ/pWMQAsHLiV5Nk
CrLKu7oQJSZz72lOMlIplN8pKCjndfNDB2T8hwDRRK/Z3zUuJSou0qZHGzbVPniR
VtSKO9QFWlgPxO1RTiqbAamDTIgUoRJ9wLlQ107W/aiFtH6BrRTevf0sXWVmkkA5
GmYvbQVUtAhenfd9L/J/RDETr7IlRxH58myqIXIVWg5t6jOtX5imjuXayfbxU5eB
ZHzKQsNeNp9anKGbiWLrG5jL8jhnRKZyLPoclZrbh9GiQRYcIB50VNEVKwoznFap
hqcQCSMiQApXuXYfPaT6PJKevra6Mt9iDrmC5q2jXewEOWWJ/FNpz7dmoBeoWK8X
UmaULBe41/QKVFPDkppGfsVXVu9jESAAOrBLGN3VDS5/y0qtFWnfjx8p36U5bh1c
TrvWQ7C/+em3lH7LlG2IZcLX9L3i3i4/1FRyxDG+iMWKSaQe21nbBOCqZ8OoI/9x
vvzX0awtqJbqTND1H2jypnoOVkuvgP+KHNjEQ5w2UaHeFDL1qWf/cVoow6t6N/5o
anCPtuy2EKzpjNms529eM69aAa2aODG7IdDgxnMO6ECiIrrokQZ9zV+xV59dGgNQ
QbCgszOJVMvCSp7GgEoFIKizIEddZxRfqvmR6Q+0u/Ce8b4Qc+vc1FtWP8+jakQL
lAfRsepnPhlNkz1Fb+kgTgAMBqd+1dxaUfprzZsiEq829DK7W2s451UKRZfqhImu
0hD6wHPlXijwfUa8uV7Q+4F9Qb2kQBxbXFgNyLagBIItQ/ohHID3xHSQtpDXQ3eT
5D4hAhDy4Vd5YCdrkNpKRfMk5WJnTVT6o/XfawOKlQt9xzDV4F2GkHRju2B4EJam
RRxFx5PVN3uQ2gBndAddg/tHTK+hjD3smd1BZRqhSnUUIiutvPeTMKVx4ImanSav
dsfdvy0vXTkmB2FnXWI+PIQl1rDMIp3Qz2Lh58H1KQMAMKQa2t2xP9ZLBwKL1Hjz
Pkm8DRliL89e2B1mnbEX5tESVIftqwG7bDMxh4P0dq6ncNMDIzUzdMxEqx83vXYa
0BB7kjUpRTL+Vmb9tKiKPqBP835CGWiN52wCpk6v10vkzXmxUBPKWxd4cR/TvKGF
1mtFFmNNKedgfaeVhdibIMcKPfGiswZ9lisAK7uvqNJwRgsAK13xoYrnNniodbKc
pLbkOytsTmPVZASXkLVmCM/+eIcM1emxqCeb/S5vHbwtvDDA50RzI6A/cNj0qj1h
opm/vCnyOMVWMFz5YC7+jREJntbs8sa3BGhCnTxb/ZUcZAElt06SS89Hgrgduu0G
JmJT3eAtK9xZrPqVGQOINquHBooCHy6jxiYal8trQ4XD0OttFGSc0W8EYZfDDS+0
Z3KJ1SIUfXkG6X1hrWXNYprnKXchSHgnz5ptk27OpP7NFwkpr3UkHaqIy4H5sfzj
A001npuI1GeW1FNkJIMX+xzzBCJG1bdZ3si6S+5NduKj3I2blZmycPayqKOWthXG
VdUnO+gKqbX6NbBu4KwwImSQPXpCI4fPAKd8EeVyhQgu40uQ0cUm0UdobEIpe0RA
JAtpQN1/94t9j8KGKmmSo8nREMMPaLNoLg0dso63e7T2ZLREowLb/07mYX2Zgwc1
2f2SCQFPIOe240H7baXm+0SJONJVzNJ7s9EWrJcOKUVKyHtdzJ6Y4vWtHI6mzsnC
NFhz4pw+3b1r8V9TSNvSxYUwe9lQNSCYmqLdqMTUPstt02gtk4qRPZW8LIKASpGq
KUCOOB7Rdf6E4QlSWf8xT4f5SQKelokEHX/o5LnStMM9D7xCTwZ54k9nc750my24
phD0ik1cFi2vWTCHNZQGwuWA2IKmbPaI9L5aJJerUfkLPg6Lr+8nGcFAMtab6IZa
mF/u7WwfxvfOBvUUubsjX1ZCnILFkoA2vd+b13I9w3o/kh4BCxFUfxCbHEmUclF2
Q2u1zHh5LLHkHGhOk8HvTpemLf+SWwp6eqTpry0w+8YH+5wjH8ZHaYwZVZ0L+kAq
7l406ld6YMrxgydldCeAbMZX3mulEk13d+K+8aPidiMaR3Qkh5jd2ERPKWVMv0xo
+B0fc0GkYSbkrXCkyvmpPaKMi9oF4l7ENouzWB2w4ZQYwj4Mn7wqDVWVn8uIclkL
bspbM0X4OKYJMFaZo6FEAsS2Vjg6tjidQ1HlrBPtRI9+lTir74YOI0Mojl05fDsh
QXiMGfNicoHfd64nJYeF8l8hMTvAh9OPwvYxCuiecVOKF1aLx5IeJcR/oK2pLRh4
dHPaw2XYNiqVtctrMVCwkj8WS0otpFFM+AAkFzsHdr9V40sj+An8g2cSDVdmFWeM
n72kZJ7uRVFtNAst+AnURKCmQgGuiMn990Ua+fX3wA14BatT1J1vftCv4BgKT/oe
zP2Zh+POiKgWooVUPsr5YHZa+BLUTOmExM/XTws50Nc1JT215SvAymX/liES11ZJ
h0P9KB+eQOY9gKiGCnzKZFeOX+yMwqg5CQfqVFx5b+W3wa5iwqpth4BxjW0yT+ft
sGiooJUESk8cDYm7uksj9QqJxCovU3kZIgaTWAlE2URCghObMDUpZrGPTqFF3Lex
vZgC/M4Y7yDpJXHxrsFzrH36mfolEYmPET43V4xFzW2jayLvpZefNPw8j4vYv9WD
994fQzl3ylyPIIBTYdVtN5wIixRPdrkFAoMor0uapAR2iYN5TYrEIbnIy6RpnDbm
2FR8BiBj1cxxwX1qTrxU1CvKr39573QsjH7n+tDPU40cXW0tr6g2xrOgp6rxd0g3
xVz8vZPsqtGGkkYDPknUnGcqQj/yXb2+SCGxCtZMQAVGq+inge3fi1QfGXSd9B1m
yI4lWniLwPY7Odx2JcgnK5sLPcQQFjPUg8ylrNpUsV2ha96tc4zmEWxIvWnld4aE
NgrYxJzA3DFL4DHBMCL0Z2AG9BPHT9nMsXx+tdAI4NRhr7i3WJJAZoGbNNRH4gWV
W+TrzXTMs9sD37q9xD/kWTIFAlidzVgi5wLzEyquXIBWydvIgPPP0SuqQTnys3lD
3BhEiK+MMUv32q1Gd2zP5eflbkOub8kaDP5a9404zb30XF74NdnbkGDbSA+f2+As
lbUYfGGeRInMs86WgDhkc1y4N8M88ecTy0mfp+7rDWqDD0wdsha5zNKrmR9uZ5iX
0GkY1TaAiZ4oXKYc3Eq+xKROdrHZipJf0Yvmc3scSHg7Mu8xruB3vAs+edFMDDa6
fL1OGy4ETBAEQjQTamv+s1PkNBhQ3pxdXf6EO6/BuyI8SyBBJOXuxSYqirSi1/a2
DUsf/6cTnJaGqyqk7WdrpoonYP5jfl5bFN7S+Y1FcJP8I+JrOPSoQxZ/9lkiI4mE
Cj0wP/fvEtmcZhMlCKyy1yIqoMjE9VpgT/FreVyB78vV6N3jorG5LEr5ug3kJlB5
uPOW/kPkYK5VDVv4MTDJsUSNzDzkPFLXeqlBiqhGknOgjrKg1laTDXtN7F6ZzYUk
J/wLgv06DDRvw0PSUGkw4AKvRu7Pdjqti47RYYBOS870bxNuv3Aaw2yvC2F5V3BF
qZljPS9INHriVzqwY19BxgFV5UkgYfGZ+yj6/KtesLfogp19allWlsEOfmnctEtY
ULErn0yvDAHZxq+3bkoHiV0/beyywZGfwPtwNgNDByw6MGJ2iJlA0DsqozOiBsa6
sG6tyw5xFxvKABhWln1xDQdWjZDYOaANlxROjPJ44ZcC2qp2LeitBuHQKXuuU5CS
HON9BzB07JTOqhdXjmt7hK6i3q3l66aTkZEK4dBWNN8u16U7NDYOrCnkBhqeCtWq
1Mo1vSnEy6Bqj/2AgrR4puSoaiGYQJVW2wW7dyAXRlTqnj4XxBxwofBAOICBFx2c
p3vDx1vLbsb3ZvzGRh+3psM911R9E1RY/GCVXPBkYlbC/O1ivr3YKfePliPmu1ZF
XR9QTmmAAD0DYRLa320O0EXShQzlJvCX6TevRWSGlmcUrnOYs1Fz45ZCUrsmy5+Y
k3Mr3vomx1CGcacZsuJSShIRkcYxdA58oSbH8i6qYSBeToPXy4mRbUQ8mspPrqaO
guwKCjhEZb2fPn6d3CGf3yVrw5LMymZ3t0S/C1dqPtrDuS8CsK/h5t7EhJGskudz
cwIjZc2u719q376gMt6useZ0J6vtXL7gbnQm/NqMdwyRjiB8O496UHNHkcr4iURj
TRCXY0WFlxCLqDzZC2VzYCgrNbyoAKtr2ByvApnEyevAv3NUqgEVrTPZsDEe53Nq
WU7GCSYSzdBViVB7BlpZzOdAroIBxgxVq9V+ba0QAh3LzG0WQ1vswfJ12AnmhW1O
iNi0mqBdvvdfLKnYgErIpXYBvHYCgYyK4fwe2gX4TFUy3MbxZX/VGsgenk/h81Nm
udkIbe4usfyhZPlHFkbRz1qIOnxCxP+lcfaSHZuepnfjWsQP6opd7YpllVanDoTE
qBTMLI8CYnR8mlvQuj3P/g+MKYlGfJH7G/kgSidAHgAnSLmzaqSNxMCQ64nmCmMZ
na72oZIuumsjpgmBWsNcCn12O1yKl4qkNFPjQwrIuv3hOl0BgSpnZaTAva1FArl5
Kii8ihhjh/d97O6OkzIqsN/1GteFbmE/ktT4ZqXSwA5M6hmyCXtAjgX1wGuWGUGk
8hUhovA8YIX65T6L67VKcApcPE84k3we5ULjuFaL+Vw1fSj1Q1W+7t3VvrBpmUtn
IKyW0oZKWlaZ3V31LqDfSg/CE114bpCk02veiy++WKvCAGfYoAfnITcLLYM29ZQt
wLsJrLNR8YjI3W3sjXa7j/pN3/FXvSWcqmgKnHKhnW7eOLv+fDpMTV6gsZOiQmR1
cXE2eOYLiI0HiGhbcINp1oxd1qoW2zFYoE/T4G7IRXLNocO7o6vqItaUS9Kh8I2D
qTWTMmJycWuEYAnqxfcONXIhpuQWor6511feMcSDi3h6d0xkKOH4BtDI5dC9CT3G
yJt0y6HW73sbCu4tiRXAoWOwcT2A06vn44+0xOzIOki91BAenmP18U5UAQvBlF2J
V64u0w6thLhKVyNKhkPVfqOXwAysmaXqYTRwPG/xbH3MGqZqB8vHwCiRieqKGw5h
Enj1b0Sv0jdFcLBJowFoEz1v9GibqUj+z6IEqQGVxnyo132+7mc/3ETsVDWxLQM8
yrB9rwM604wJBtEFj5JIbzFOdvYQlS7juaXzvRO532KwPel1EVAVAZHxD87Zg5oQ
iZ8utSaBL5HykistdJFHNfsrujF03S4odQWKP5rpbznosFVhwfl5oYMfS24qrKCj
1e8zxu3elZW7O0oyVbOi3aYpigl7aLKDAhcI1Tz5beXZQk+Z7a4L2uZm6pD885EL
v2r1Qo8+p/K+YX61UbBUJGbaDrjmKnWNbjJwd+QUETrKrP9AOlExwrr98771HWzC
wJHjvMrdmtafbjkPzBY2YV2PfIMzX+inDNENnk3+ugbU327DpZqWkroExR4mhqHa
X1A0o8gYgUZIl1NV/pgrwDBvg7pWdxtvR2I9AwuRIWDXeyb+1pRUmxbkoEF4MJd/
5hdgxm2BwZ4BrCiPOt10n5UwS5Rdi/qID3Y0falasizgJPUGDKOfOHQk/IzpxoV6
9COFAHCC/Z5/vNCooD02+rh9PHF2BKLPCSxPYA575tGcOzXESjVszrdpeHzsUwkL
wcGhGLiv0190lL6W/3PE5CWIaB4HFSOmxbRuGOMAVUhR1PQzOnq0A9+0yVVY/3YX
HrcBk2yLuIn9Mnes9tu7PtN19LHWNnyZUcKlCAJENAnO23im2+oe8QDV/fqt9Ztz
nsLb1/QcMs5RqCEs/yB0JEsCin3tAfXZhTwCu3q+HlMC9IQuiSN63ktPPGQFMO6u
k0Mx6LV32/npjSEUM94ruHqfXn7xm5YpjrHwGZuvXwYqoF4iJ7kE+H75PdGO4G6G
HZgmQyoQBKITLw6S0pa84ctm5tALgc1EPPovo1XV6oUz4k0y5e5spAocOhLXLCu6
DJWW/1JlJ9/hvb6aQEEIcnRhj57nBd91DxWUexHF55PDb9VxJbrupyHXqwfpRUGx
pvyr1x8ORo1A9mPrDyub4OLMwnjXXQbfaTTVJXStxZ21qPlw7wtw4BoF+ip8WYE7
PWMvNGahpt1nz7b5b5pBwCMC+UjIX8C+jLyc34cayeZA0FHD1UlLJYc5bVh9tFPD
jS3spb3cU1HC7ul7HfSEAflVC++pbymPHpLHdpkI6nzR5IpVtils3uJ4Rgv7P9ma
Ayry+wu7JYzojwMdu17qBUakkL0EqF2A0yyODH1FygkH0bntk3k16SToA+dCp1/s
yMnyj82ekU9Xt6m6Tp+VmGVYVUvH+7W38Os1s0FBwtiysE0PXSF38Et1Txt8b/lC
fpaw9Daz8CbvPwJ182QxhJQ9LGw+1E5PgqWmwBDjlh4FcA65f/w6KQBaLI0zFB42
FIwYel492t+kSWgP8UzTd9OEnGU/ePwEchXBJxdxdKOJUq8ujP5ifMt54yEtH22t
3visz7ml4CxFzp4OIa3tBn5eYFclHk9acDa0S2+zMQtYjo2PiN6ZNUDAvNbMy8is
o2SSw1ILfKJ5iNYD0s4DYKIFoBai2EjUP+3kP6mLKOVHDJTXqJ/87pORHgVZLQSS
pVZZ42tXTf1+BJ4nVS2fcpnGCcfr1DS6HT7dNOgjvW+aGYYHTxZegvQXcaskifwx
PaOc1VuJnMeb5+alNanixsLK4dNOSYWtgRUfb3clQJ3vrUWJJHCGtUyFTb/UdOl+
EsC/mvZVu8KCncyBGq5ncyiaKaEOu6VxcJCEqXOpAxBs0RWRaKlG0n83zV4O8VIn
sDojFz6aNZw1dmODcRRBEbF1CHnAHC141mE7F5VCqeqtMHWJF6Pmht2Rzroqeyp0
+DNN2tVg0WwK7gXMRt3WBqvB2qvoaBLVP4mZWBw22XxR/NA1zi/SBbY4g91zdbn+
C+nO+ndKywu6/fjV2dzacUgdOpk4c+bZZbCFoqI58j0VMWgOZpEtgWBwWMNr3fpW
q7R56rw6+qvolad+mtoZMDrdoWXspE6BHCpa7zYemABwPmJuUQ53AnRULAMP99Wq
TRj364z4MFSBX/U5wPmZfjvsDlxDJaBx91ZX3woMtBemdi9WfYzoQxk5iXvH5F3L
n+53YM/+qXL2BXgo6DkLjYuVhB/EbwV07LptQh7jLe0xksqtNkt/YGWCyzWd4n+B
w7Js+Joh7AHtayjuY4uIcJvZC7VcX9ffPFFOv+prrt3gHkwHMdZjEOhNtiFxfs2j
IXS3lNs4UDPmu8T+YeW8Oz31n0vn86gUoBFz8Wg6jdYoEbfR+AKGxNCHjkxivL7P
eAR7+Zu8Jd79M7AgTC1Am8VsQoBGUaMK8dGexG6ksH4vIQdVVqJqn4EmbEJxThj8
4I9od9ApmLHyifQmNTi/CcmgFmzijItANxgQQ8smLojMgDPCn3eCvm1990DadQsh
HMfn66X37aYy0/jk8kHcV+CKUXYSErE9IOzCYI1NeaRsPMBIleSkAv0FZCS0myb7
1lG2LMyp6QD4QlixI7FjOTsIaXKcpMt0esLCbOk58U4i23bgW16ivc3+PPyeCf5A
2q2kWBX704rg3xACwPj3M9k8+r9M6pQ0tXz2bbcJ7vIPa/uPZxjVZ9rdLzo68z2y
k3cXr9okFpmIPLRp2jKTNFRrn/pUUnlM+uy24UCzyMeNcugkjid+GAk80lul4eUY
xqcbPPOR2KhHoiYjyxqk8WhFtjZ3KS3CVaNNSz5OBeVSm8P05bRQSMU1uZ27QmIN
SP3LFfxc3FkKOq7vTAgqatkXIz8G4N7TjxUab9MPm3t5zLubnSKtjFoMUvwPPTDP
vH79vYhiHmVINtS/EkI2qMhf3bC3VlXn4EFx/TNUBjO4kh3Ac99+zQLkMEUB55oU
iPIuQ7yF9zz9baMBbOpY+BRdLZkTDxge3Hq4E6IW7wESSzjIVRTVoRF+De8c8AXR
yJK9QXGLzwelinecS48bZHppC8e6As5NwdCrvayUsTiFDFV2entcF9O47AOEy+2a
emEk3rixcPJOTC0DkGWZ1FbJuydLDC1ya4ABdkYJWHUXX9m9lxSuQ/xMuP+abgG/
pt5SnFEijBGalrdapLZJudLpcG0ebJi277OHl1NjSZ+tuVnNgljDMIJn3G+F97r+
3OQDY1DhWKhE7Ws1F6ppKUjBIPeaapTsWyjLHYqUIXzikX8dQ4IEQil46W32Ed1U
3j8CjFknExrBuHn/3cieAuMMJoZuDnbBu6OF9Odtahk7BjONb+P5GkordZlVxDPS
8hqi5056hqK7RVYmUMJuFHbQEDYTYcwDUHiGpozjDxVFFzol5j42yh+QuxPxP3Bn
kyMGe6m3eVDg7zSbVJT6Rnl2eJ8N6MlODtsz1r6AERxre/7Oi0aDeGZBS8/Kqe1Z
uihr17oVdu0oPcKAmUEdwa18REdP7Vlqq9+LYaQ6S2dIKw+eJF+6o4YFSsvN9PMB
9TeExPqpOM0iWXdljd5BAgoS4s33JDi66HpZEtifFlpdM/XdwSiYS/02WnHs+1D9
+QxoS41/DKivC/ONO2ebmec7LYJsawqHXPhkmLz+t6XRfTsYZKKfwzoYup46o02Y
/qQS7VyQ8fwYfOmlBOEQY13t3RjG1lO4ngIOAGa36ZQYdD7/8y2NL+t1804UxsWw
cu7mNx8f1r05DfzgxUqsouoasEa77eRISf+hbPqn3kzO/jQE203hyIaODXJbYx48
PDR+DE9CoQfUuBYdAkb1Nc7X3imtCj6nqdeDGesqXkr6S0TmLjHQHZNLoFgmQ4gn
NjH1fM2aVmg6PHsGTWk0B1BjAQf6KJINn+EC3R83PCKvnJq2LATfyEbUAqf/hf1c
oilfYhZGxP2RklNI/vaaRTr8YCPrGkUK+zE4xRRunQhpNFzunvABGHnhK5dBZRna
e9SJVh19kCr2FAdNUAre1vwc6WfjfLvUVuHbQSF8UxKDQgFzXNywp303vB8kKypH
OMyPNCO7qI/+WCSv86x3KHGk4h4mYtXg4F7NY35JN7LE5QHbTL+vDSO5RkumP8xG
90ekYv6/UnviuuNNOWgpiOoesQ3FQ/8P8f9T+SMbClnxqGyPPVRwngszuev+eECB
2ZpAkjs8zUzcNMQe/TNuRzvpDmK+UOhXBgLqk34uEl4st+rr3kiJeJMmYISEoq5S
l5G138wlX+7ID/aUABxls8oGXY065s6stNd+0PUBX/GvcfUvpYWADSEJ+YrqAy19
zNIMiruq4oFOufMIaGROlLKLeojOYRpDr3ZfFsJdU8PIil3338Rv1Z/DVh+SI+Y1
MOBMXU4iLXjjzWsyudcaJq5MkzrxHKOeemAd1DgasieTRhYweEmZbAtVmIqGY2oG
gwZVR12mw1i+LTwIlVvc2Zldm7yB5LVSugx5vZBN8j04mQTmZAhAOYoJXGUFjKys
nanNyMljYxtweHuaEBQvvcVCepZvlO0YnJFjYVr24L4Gn3QB6XVgx+b9tuEfO5/J
SIFVFIjDzg0k2hmoJxANeCklVzFdB6c5W6pBL69pqK5/m/yZ/mgcVCugPB3zVKFF
/DvAsLsqMJkSYL4mi20rPDMZqEdr4XLYtekNUjvF5jsE/+1Kowue2DCJS/y1Qz9L
ANUQHFzO9qLTRIa7tywAHKwoZoJM0Oe+/eze9xhyMYLkqrb4Vmy7T1tkbNgzkHSp
IDKVjsYess4w5weYIBszer3UvbfZ8cz+sGBaAS9yShZqfzqxDDO4MjWACcGPbsh4
NUOmfr/x9InJRezbPQ9R1XSSqKLVwKhVWEIVPW0QV8zSW5Sqw+WwzBZatHkxaLTo
5ambzO+N/cZcQ6WLw4AJJtDG1wHxBLouiD2XL5JyXfDkH/odo5eumSR7fgbt7nQg
PCXvPETfpBGzPEsFaxIzO+I6shNi8f8WcCa8m4ZXFR3r/gLQKAp1doFq7/9d/LBw
O5ZnmT95VCSmU+MVHqQH7hNkHTxPZZ2PjjTOLG57l8ORE9GdzyNd5bsQI6bGfimD
6SA5uWwx70KVoBRJLKEpg8sk2gGXzbH/lLBaAuf8L/aryZOT0kSR9LwXNffZ9mWy
9Q+PPuSla7D3o8CziIcUmzPTbQR0FINpxrFjI7bAdG5m41EHyrLp41mhYdlJ9n29
Vcv5Ki6YQf2XQU30SuzaPNvWhxgwsrxYs+w5hz0a5INbyBZZYdblLyYbR4y2Qe8G
mu6jzYqnw1I+vzgd5+2K2Iu0GPOPIWVNZfNYKlh3Skg0Q3XWKig5bH3QAkCC5iB+
89zzUU1dD0Dr4Q89+dDNQTN/PVIyf/u199Z5O57sll6Iaepk55FYCi+hFiG181gj
SFuBRAytjEjAa+HSr9MfVCBOqeVrwtHCUSu9isSMF7REUvfJNt9aI/UJqWY+rO8A
elOBt4HNLRCllLeuguhFPG0OkDTjoZWRncf1OAVc7gTOvNL0KMnzX1AYOoNc32CM
SXAKgGAiZuJL3EmBFNfxDG4TurTB0dsm4Bw/k0KsoKe9yJ7uua9fJilOdTdq8avO
4GJ7V6u5zHGqFusetOOq/lg8B+E50X5pnlV9cNGDIGeqwJ9WMveWYbTsCwCAHQ7k
OBNS/YPrfElfC4PQj5kDy5pyKgjXLTaQ+K9feH6jJnVSfOa5/S9NFt//IHWkE32O
M4LCeJ8cCLxWedhnAjpyfX3h8G/SbNBt3WAfPJmmEXOWQPCfkVQS++u2tL+3n7d0
iGOzCiNYH8qQota6zjOfcWl03q1lUaLoDofhFCjXP1cwFVxcvGgDX0JqqOdc7Mb2
htqipYVOGZ9+doe8bTYfi9H3LmGm7Y7A5gROp3PkBpCyA4QdwcM6/l/qZecvNggX
hHkv5+Sz6nT9YatE88zK26JAkGR4Z5+bnTpXoBloBDTLbwN0V5j9i7NYp7XCnz8+
vYkCsL3kYsEp0zUqjUo4IDVIpgjPFfERRnd+Zi7uOXbfu9RZgEDZVgWYTKRMJ1tT
oGXk37XufYLa9WOLYrI7jcD3Dwhcsako+VZWCT9zA9zPdEiezeEvTrCzDq9bBov3
M3nN3QqluBmJeiwTEsBDw8jlQ/P8lBN5kjxaxihGg8G1z43a9scZpvvH2xGzJIHg
G0h8Wv4H7nHQD01ZZZVSic4jFndfNCFUTFYSWpueUnRZ2A5qQkDrpGB46xxY4ZVo
haceU7QI1kIx70rFxs5cytU/F8Ovd8ECkDETsgRhQ82Z88+MNKQD5Dbw9jUV+G0o
kjrOBbGb+jSsCzOEsHtBKLQC5Bjc37s3ql1/MkmSMcfQqntrwH4Lnbk7E8hlvnT6
764Mw9DgrVgZ2xnNYdEE/UTii2GJXY70uZbSa5qstIQ/brapbYzjKwg3T633ojhv
g6KxAsVwyXHxrbx2YJ/mG0ZoCB0l+7dd/M8FBuIl2qP8o0dxBf6GLv40m17u1Ymd
0XCIrNC6MVuBs6Jjhgxe+2UM5KrpVcr67GJ3bcl0T/IWPW21FTZa6IrQCtKhOgU5
FYvjhAoTePnNxACyz+MeL3LX7GHEcpAtaxK98k697NuSYGl4G7b4K25aMA7o3VTu
jP4tYDOtQo6EX3wXqyh4oZmXlW0ezTGmN2blJazGKM3ELu0bPQqqwzVCtVoEvPGq
be8bmBu6VgNGabkVk+ABQ4A7Yeb8hsUmakC4imX1npHUQI+2MvjdQs9GhuWVp6ql
i/KYKq3g5Ea0dr7VozI++SEGNkdnOwLtvwDvbk0b6Ck/IIkZBMvU4YB2LKXvH33v
JYH3tOMgA38K0o5RhDmaNTFNTSCRHk2YwjJiS2Iuco5+GbQEIayKSzDxvy/IheLy
D/zfMeQvvx4aXgDG77AUVW1LwpqEdP7j6+e8OiHCO+yApot3YSzfwEWqR/fWCQ/i
w64XPWJt7pwM6ye8vxrhHMRhcOyfxHmRoXG6oPdT72R7woRJwuOg9KTUpXyJ0bpk
sqhX9CYXGvAny0c2+CnsEQs7JZ4FhRcZX2AHpbe921MuO2WuZVyffv2yFHM2rvJQ
MwXRfOQLLCzoxKIQDAhlibZaiRF/GH7K9Ou4lfyd1uv8fV82YW45pfX+fZy8ST1S
lZFPMwVO2hlWIRqRMvTFcgVSNbYnZt0LpBDTjrrgGMVuq1rctsMECR09nwrVNdim
rXHTqFmifAl05zJaeG94c6r27Epv7F3sdwBldlaQxvBlhwza+m4H4nCAGNPRZsbC
LFOledZ1mGvUw0MgrcQw4d/9gT5xTHQUxFo6R5VArWvkFvi95W8zaSRBFGi3bjuZ
FKH0KFjWsSXOkMNJLrj2XBPDyTkijwIPa1q4nfYaxKJH8HLVJ4u08W4iusGClNCH
NyPIJEegIw6XmlPHQLI21mRg3mcwRjMOcKZf+iVZ88B6yG35PL7TK1NUZPptBuDr
QAcsky2jlGnrtg1+WjVFQLMPD+6e0PaC+dH+oKSdKMekKVhvTCUTLtA/OpKsH3Pd
I0pMehgXFEz0K+t0VhqiEnc+tynXrs7W4DhZEMw3fV3snnY9UuFQoXaW4qy/5uxG
YmGcQYxbExe5X/PefsWciPGGhG7AhG/lv1TINu+6UJ+n4EOU5yPs8RZ896IxizLj
Y42w3stHGl0rHXTdc5o8yvCS/ocVGFlmozQzDxqE2Ied+tCm0EpsYnWAq+eWvujD
h7EI1K8J4LPBbtmtLVrqqaA9V9bcFJrtPvxjr1UlwJxVGaCCE4+SqCgZAGz68HkE
R93avJC3AFHoGEc+syMvEBG+mJ6PdkwOxipO0j1F6j2hrcMILnsdL70c8W6wdxT2
MP6IhbG/AfuDW/6DczIMLJAcQta9ErH/lMoCwRZ/+Aez9ww/zjlu/cW8dJdMqCZ1
PnkaaY9FntMxDbQnocFKoUwaJ7baT6iMI3Qm38Rgcas2LbRx0eWRnrZpcBW4CKQf
rI1aJ3fLvTPscxPkEqbA5QQV1xqesMFLy1zKmPjsfisgiX0ndjVzZfLbxdn+gxBI
DxowsWGaS1vRN6TtQLU7X/owBmCtVCObMZfG2/8rmOSbSQv8q0vsHhM+RqV52pya
TYh3xAF+XIV+A8A9KFndAB6R1/uFh7Y/QWbFbPXHRWdvKMYo5B3iZlZzp+R9Afmu
JUw/cjHH4gExVNuX/yuXhAqxyF9h/FwfY+9cafFvJUl8Frsevzq/pzYRZ0XyK1yW
G4MNN5XpgNY9ayLBCLgDo7O3JsbRhlYyo9pJyBn9QtYxRAHHLQe5E1X9E3UFaexO
GmOCbrkGaOTplXbF2lZMGC4BhnF5dShd5dmEm6RCsaoapJqEdTs0kJCM0un9wVF9
bhoZqF8YVKohT+Pzu/Ia3IHsAcJmIAuQs17yBABBNWOkPJOVOlc9BD+YoFEVc7A2
BJfjnpVLCieMAmR8SoHnXtR6eADbMVyqJScE0uNQFRzfLPkQqj2ExQTEZeo3mNuS
veokp1Q83/JquwfKlE8k2bvnkmNu30ZXcK4741ua9buejGpxlmdJLY1gGFc0pefw
CSaDA7vqUlqhIMEZwvqQsL7Mq2M7Jf6wQVek6U4HYJdsmou5VTdvNpumXx31auQh
LeGII6qoOuSERVHkX5P91S5PqZ5MyI35ghw30B0GUVg8yaLA7UJhMPHuZuDmPqS9
D34An7k7Lb/sOLvJI+7TKK+kWxpgmU/9C4TdvwEeO+Pqn3AopFBqrEKpjt/BLHz0
WipRIaFNH6rwtfOuX/Y8a1Ukr/uwHyGe7OXGWsfKBJOFiYhH6Z5D/pLcfhYR/uDK
vRkywgNhjFNckgnCCsyzbApfFgjabGJws/N/hYQXA8juuXam/dfzTP2ucPcOnnaq
wx3PddB59Pth0E2b67DvD9PvM4JpOElRZWl+KaR+x+7aPxZeKkr1LhyudisnlQA1
NSTftSnfgcZfa1Iut8xwLd3hKJFkUP6MQudWmjT0Gz07zBX8OFqDbk46Bm6o0sYB
r9jODFfZ+5zqL7R7IMpWM/8ptr86IOz95jUZ/TVXTrB+SewvmwbAqEXoohDvrfpU
4k+mH+7E/mRGOMtPesXvUSAy3TAYMCuUqtbmGT3825iNrBlLU+FnttBoWB1t5dss
szFo9SK9CIMdqvDBX9f+JEpEKm+4QfwmHBGR4MADyrOy6fWX/qZhahCgseWnDcjY
qBwoTdro3+QO6cOHGLaOoaY3KNmTrABiPop5TiytvOs5eT5XPeohKrfcvjEG8o00
ZfDYOVoITqCGrN4Zan7sidJPkrKpPMlejCJKIqop4MoBvj84zNZi1TMnDsP9oiDf
+jdcTdSZOFpaHKuIYLKizTLZBxSUuZFOeczDmC/YL6uzSv0Z7vLJ7c4oBhSyHHhf
OT7mAYAEaDUrhY9Lhn7HbU7IdZm9VpCgMWYOdjbeMnhn34RjgsTlDBZ8LH1wvhcG
fOZTvFT75K/qlFllCFz3ljOGjrxDgZGnxTcuiJLJIaDeE8AWJwUZKcAEarLpDhDw
bN2rmIDRGvaaqhBj1IGwiIK855KZceY5/KhSVeUtTrmiEGo2WkZkXIkyyOw1o4e7
ftGB73NA2nnlQBTkkecfD8s8qZmoQ8eOwGHBYmLKVQcNQnUzz+c0hD/ehlr0XhL1
CzANv/mI6esrpM8/qWxLmr4ldfx+2WWbg52G0rbvHQsOTbK/FSaLh2AQ/gc+gl+F
rYipL0PJwUTpng/YqeUcYZaI0hAaBunJhrTIGJx/fI0vbiRH+VO28V2OLpyIuOQN
cnj1XwW+qPj3UyzLonmud85j2a5zeczklLnRqnCLdzLINKCZ7pFyJMqK7F0PUrXA
sa5wdKbtFYCufITkgb26r2iAF02/XBIp40oNuytQp+StsYMeS3/0z2shjPtjiE3j
o+ii6tkgMtPYyT5eGyj0u1uITdTxhFflpz8mpclLvFDEK+pGqRyRpRL38uhnFk1f
geA/4gXUtvwvPhKac5qZ8or/yHGwrx4iFot8wifiSqMgmULfp7YY7RQG3Go427h1
g5Bdqe0kVfkFy2pgpVwgpXnfXSVtPPNLlEjgtgERwbMDsJ0Ohte9YUQFWzqJP1sZ
oAml1v8/tkGaA7E08EjBvTrTxC6GWJy1VQVcvJxY3lPnQ70vnpGpptT+vXSbEH2+
UEAxvrRPifGUNTOj1/AzdjAtuLDlXcdVlh01AdtbwLEk07XRQkcDa8uK3nqghIuc
uZn3H7+L0EWr94DVGre78Kv3s/ndTbTrh8f5s6KqcaOhCDy0EvaKCdmshnjMTfFi
ao1zr3/ahGh+PD5lKNAAO5RQz8alS11OMsY5vwuFC0kuQUvFjBbEiyZhaHX7c6Ns
3qEZDBq+4NKSFsFy4TdPqAwoj7OSYVWh13JfeZPQNgpPvjviWAjwd17ZZ/VpYeR/
imM4S+hlusXIsnhfv4FfPBo83B5B//j1VPuxATPhTr5EImqyjFHTUn4upDq/G8Bf
t53SfrrnSVgAgJzFPXWH+zd6+995d9dRUoXUJ6Xw/6koW2WOpRwCDcPT2pMDIo1R
xQ10a07dRLVxgl4WQU9XMiGbgpZfBuWYDPoYX2YksA+JkwRah/uU9P2tUywA1YDn
qT2kpF/+iP7SLMaz0D1GwgtjZdbAQuGJdZMfJJi4RGZ2wgdzn5h985FscY5IM1Ld
7kG8S/PX7Drz1foS+PSE0yBlESmVkYjEm7H/X8RQj6GEgcEKzqsQFwiVbtLUE9WG
9Z+Umxwt9gq3Ng+33Vu193CG645qx28LhD7oSPc8YBQ=
`pragma protect end_protected
