// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
dNdz9JXBIT/lB7Kphm4DKhu1/vyWNitED2+4/5yvAzQrAQ6JUag5dQtDLTmZAmUSdOJbUMeAh27i
s2+u62iROYpW9rTY4v9xnXRecNPG78YcMqUckJipx45YAZEaOuFEGxRNFLSYPKRRHvQdW6bfb52Q
fPLwRqM8ioUEebmLVMegDf6EXzqUSP4o+9zztKPjAC5qjLFxNqAboAkrHV5bBvKuRbECPGPZzX2Z
6y8AvJKYtijRfSOd+C8m46vPcLWwpFB7FaTr8SPft9TsGn/FLFj0FlUt7tejIJzO+DtANY1s6X1H
THsZsnyWTyn308qp0SF5cBddkU5XGTnVuvHT1g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 58960)
f1kqH1F+4qjeFPgM6UC3B2hzoRqX5KufL4pRNJv07QIcZJzNz/e9ZlbydANItP8Kw2vIyJKw9oLe
uiIQnmfLaRadxlqwv2/PVFlji0FXS/Au7QD4btFH3E3c6dl+wEGe6ZPbnaLvMg6igMJN0swxr1Xd
np/dGmxjqlMwMiziQb+Sz/U6q6DDccE/8ckhAVC99w7Cf29gy/QtJld4qfv0lNMIKNNOKkP5rcMl
ALQKhRM7k/fUonxO3UTMW/urRm5CE3z27U5N/lX97wH57sDpkjJHcwweHmvSsRb7QJDd9kp0FcpW
jAitn9q21HvHwG+yS9+akMDsmtSObwYrwiaYE422hH+uXcMijRX+KMAf/HqzVV0mGScSQhwliBD8
ADbgvs8zzgIhbTEilU1fGmwwGTbtoeZgERD4PPw1DQHKWFYNFYMihV1v7zKsi5u2sRbpdweKE16j
9IBjZ7zS2JdtwEywS7hLZe54gSQL7k51TiuefBAThUmnTaFk9J5/1+7PR8H0GnF/gTNDtbGtXmpL
I0ojWwq6QGFNwRMkhrB9sF0PDF8YT9/E9VKc1jdjOnlLorG8HE6A4j8gBxi4BCJ8fVwYOf470b09
Y94Q2mrttMDobITvw1kRRi1tT7of/cVBTiTW8xKr7XLFvHPBPFLk8y8v4KXzZMIyQ+xNCmgan/OK
hZF33C4/hIS8h/fTIwZw+JARC4Ege4qbBRIQympFO+VKos5dqki1HaVgIDKcuKNTpy6cja+dAPsB
6q/bUEncQeALtuyHERtJuGbdFkTMrlaT3kb5mHEgQorNWOmNXSQKUgN8Mip+hLOyhZfBqfUS1asx
OA79GyCtLM2Xt6AieK+WyyzgPkUvu9mIdVbkXCa5AhyYuRMMHiK+o+StuAq4x6mpreC0bhBxemoL
xcWVY5fN+1OstdT/2i1Q++zz1MHKGUKq9LkNZz+mB0yVwLys+73DKnbg94kV+etmBiIv8Oj1PqOm
k55LxFRUOtdXz0IzlBdOQJKpp8Xl0NoY0iaOBceZDe91OM2chScIxFXoKlV9+9J/QWRxdvq384rf
1RDkJ92JXqQnN+BRUmTVu2q+VA3ZSFRRT2BgZBDyzHd2LzO6j0HsqOrAPZ958hMqMdIC+0VBy4LC
iY1EjYoWyIt1jeeQmG5XPNuC1bVjSqrQHYqXzLAKnIekSH5cHmmUnwVqUd3TDrKxifWIJ2nLzWRT
FWmSchagJjQLV8Os1SxBEmhOG84m7/p628+fcJtpqRFxVLClQRhTXY0YB6AAW9oOy3sUMLyT88hC
oC0szz2V7d/beTGZQIKVma7AHSWuPwKT/aplu4Mo+0YeHWavA3Twxp42UJtnp3hhya+exxuhoPEX
tlLM1jyBr4UadB8pxyFuuNOpXH8r1bguEfLLi//v6Iuvmr+dtU3eOgr1FfKdLV5R+oGOC/X+9jy4
CHf3x8pqxGi6DOUo0qESxseOMyD+GVwVhoqjjtVpw0vX4SJjWGUfLGexYImJM+Zsx5uOeYqhwIDE
WXCqr8a8h4eQE5Q29fWs+bBhchGnQssdx6LPDeTR8jVy9APttFs4W6zeA7NniJkmwiZvWSf/eQUB
FZALdgpGRWgNFYW13eTXR9ieNXW3QT0kSwNOMfnZEFK21BJSDOx2te+rHuagVgCAie6Flk2Kcgv0
1N0iGOBqp25baX+Hiqe8IwaqFbeKx5yuudEkEfqJAKQkC7NPeeid2FpbX/kOxIBkNMfYmGzW72H7
UPPj9QDJe3k8QgF8kv/J3e/K3AfmudlG1VBgzqJ4IF0nosck4wmOsjtpEWsk32ivlfiiWRM7EU46
EfkTjQVD+T6kRgrvQEkMswTVGdnA5qQiILbjKeqmVCwZmj3EJ44SjmnQH5nYIHMiKWv5/5Qk9fFX
RxQdAKaHvunjvRWBSDZyzIvIqsyBglKX2z1VMd/2wiTS5JR0H1tvFufdov4Q9CFpYt7Sr2Ti26E+
SCAQNG4rcmd//Sfx4VuDxaCPDB+1f22UQH9Wc2tuNERom9r5bnMdmFL/CC4x3XHVSEX3qENW2ytS
/HWQwfRrrN2+eUJSfELAkhuEa9jBsjIfSuX4fK0Zk0I/twzGlIawomj9p5ZoF4ORCWpBvcfWNulr
jK5AUxLSFTi9llmQu2dwQsUDOkrG5Agg3kx2kl1vCJfB3vBLucUC885TN5XAJV0AXvsNWVSAf56X
Gej/Qqdeb4NfdH9ch9tYCOZOjBTBtMRiXu44Ri6UnC8CN1+e77o0AiDgXLDhrhxM8g5zBUHpAlXA
eQrNTmtnIWJ6NeirPFqoyuUHELl4ia9bGSvu4ryAmVsI9TTEsY4FaZdURy7m5xJCJRD97epxAu4O
O1Qz9oNSbFijq3cg80H1JOdFI4IAuJ2pFf5T6tpOMRP926GUBk2nXMFrznwlWg3klmMYmFq6eycC
BwV0FNPOQ7dXmGUbgDoRUoDLKNEdavBnlJbAar7G2c6G/X4fxuFMnqylA4IiINPQJFViuKkwXtJp
ceMs8N88mdc2MAQoAfBDITu/jriF3tucWJCiP5iezgYp+FvBK7n55u21m9nAxM9yLY1ues0csEGJ
rUUwY4x1TKD/ZgM1LFQIx6HAu74iNosqJJ0Ea0nJw6j4OAzGItaF4mfOneJf8b72vtMALLfY4Wh0
7EnqoxXqvHcXo6bZCy0FXQenZREKVy81KqYrr8hjZIr3IV8sTzU1DjbY9fw1y7F44iqCT+hxw9Xx
jQt16rMzsP0q9DBZU3anUsf2V1rqHHnzBTepPioat8UyeA8vEyVTYt035qql9KTumNBiAzadRjjJ
ajQT6m4gOoUPgvQupEKSOl+qBHSogV9Q2TNW70AGgs50YXU41cl1aLS7emF0gM53l9MVgSbOKYtz
+wp1yUPkPgCREBiXxC7O/1ig7D8T+3xh47xdiMT4A0kRqOPecspADoltyzPXP70QiJM255eKh5/7
Cy3AnfqIrVnZSd7/sq7R2NwA2wNV56TmMKt6iw/FOblRgZiZfok/bYhSfPMyfUmUClaGDCN5SFEK
69wV1bgA3qpkmAVB/aUHpsANjdi7O1g26RRiRZ8H6gNfZqm9WiEIIXI7bOq6LKwEaErl4JbWtppk
y8jhNLXveeb8E/bsqBSBAWj89343BgxEVnHO1iXZNsovqJz45nP2kNAXUGXqvTX1tMlS7K1mozjz
QMJzUCEH8vVcBJxQMIOzo5zvg8GHTn0Unyvs5AQ17mD+86T0DaB/DDTK0avADQk1mvOjo+U6/Mz2
4BH57SXt3sm0WFjge609G19A6oBBC5fwemgVGv5+DQCGtvZgK2uZJqvTszCn5LFk3lbPjdFOMYS/
4RDMeYD5VA3RH462J0xZwxjuJYHePS0M548PLllvJgvgv3j8mB3OvWPVdTe0EjWsCpsgXoCPNiJg
hdFiUPINIZRreyPWxHSSQqAru3s0QMrPPkZzirDumrSIyioJH2x2wPBTjW5Z1p9luLhFL/Eb3rT9
shHjjYC/L5C2rNPCpZPwIyVQ/T2UamoCLhGX1kvEVKvvwtK7HDjrEK3D21yNdxb30dmg/wI60gWt
B/WvJLK2X42CFxL8KUIbJoUejldM4LaSWIt15dcQS85zxQLZ/hs9KWIxCvUXPSmGwvXTRqyRN+Gh
Oh0RLWDrPe1pYwB5lF298cEY8oa8a9CtzbAqp8sMa5eLY556RbChRsD+7oKkik3hYtiWb/ACdUu3
zPuHXPk/eSruhxwc+EMmTxRdH0rkcNKMezBTvfWb+MZ5n2twednBt5TzK3AHx4YsccKWC4Ph1gse
Jg3hnnW80gCa2Qb2LAcjkOnnR81/IlT4odPzxzefOpxH04TYdbD2NuBqI3NW64UHbTfkxzX9pPJD
slWt8o5FLhr5B91A2pk+eBIgp121bKoJB9+8200oDoRt0+KJdeAgVAd9BWJ8ZO4kIW4zxfW6frX3
Ug5LUO6f4yp1UHGYS+WweQIbEbdnnCa13vR0YcZUb3HZpPOG0f2zZWJa1Spof7Ck/RNyRBFjcTPJ
8tB9dr2lmzDA5cAVJMwquDMaDmo5K0DSrnxqEjkHeXVcZIGaUcDyNueGaHd5H3qG8369zN2gbUhQ
40fjgm3Vwr4V9sqhlLMXWp08nDKI1jUUZ6p/UDRaZPcti0TV132d7+Rvoi7QNO1IDTvMCmdni+Gy
o4xrOm/JhubDgRMmmKRYi3cV6YyeToWmz6mjUQ0Nkm+gXtdBq9QPSmB6hz/aikRfQCHp9+ez2SYm
4Q9HMtMdDdoiRTM2sSF8c0VOcWPr0jUEWKsqkiU4rTglC2dhwf4/9U2Xo+VdONIDqHaysIuOM4pR
I/sYJ4To3IAoqk3Xi0/SZus32MahbqZrmTQOhzM07EpZgooAjisccVEN7klDqXg8QmG0StGyhE63
xJ2KJluD8DNOf7z7Xqo6klYN4i3DkHXZlEO6g2xoTOrWdmJWPn/ujy/KdTeaHVd2+u71zCIa0omp
VbzKJX2VEWjB64qQPVFfpAHNUWowTIgt+hoWcZifHBQ7SuNJpf5Q6RDkKmzUSSw7UZa/ropgxnTC
MISHjV3v8DzfMh3Cw3IiDVsVevrWsAvpm0B/9eW0j8a+swGIuu7fL4Lk83FS6RQOHw28BzZumJ0D
NerakAhljLnvXfxahn3LMzZMCWIdzg3e9aj8/neQA7TD6dQDi4rWuScpKwFtF9+BUIeWg5lpDqMx
GPS+Hai6vQSl6/h6EhMWnw9AL+C+7MuPRc7NDLPXpRWfZRCMbFEeMjDG84IxDTlCkb03w8orNblw
OXZuyqMCLyennouhFqN+aP+rpntZuqWcuE1EAbdPLrSI1HcEMrUSMMRl0DaKNkLH8pstsq9ld7nU
UU4bTTlRXY8wGiuYxSsFJDAimTIJKuQb6IwAPs3VcgSRWTJEE8s50TiCPakqZtAK8t6CxwGXesRf
KVw6tPcEWAl9/IWUUnOhOE4sOrd3NPwX+StUIi+nVeTn1YzOiUZnEEmhyxZJDZEaK0V6ByWWEkDy
ap+Osrb0aokdIUYvVqGw2C2u7gRLehEMG4iA2XrzS9BMStxI4MicUjfMeVeINikLkwlyHD0zRU5P
f65YRD2Wq2mLgRPS5yW1QGRnIkVHBNpJOZOMX64bUvCF526hNIwTYG8DD8E1wwL4nJ/GExMe9Jd3
mPbqWLmuP9HVbZVmduwUn60QvG+Mle0ZeW6cWr8L6hTuPen13cDmrpa+V5bdEXNlfoYjhidy0AdT
3sRDQwJ1CLXdSZh7aKIZvS4YpF5d8sfNXbTlueXR+8WOPN3lHbMw4cEFUIuEdH6qVN3TfYsgCYZN
Xs0XTJVqnShDNIImwNLo+u+19Ix10GVcwT1zQ5uOQUhwcSwPpt8/NhqHw9b+EdIxzQieVFpz+q43
IDNCDaOUwFdVchY6jW+g3+C878YFGVSwv+VIQ2hb8TvMjtKUADL+KM8X2bcHg/D/JT5s4AqwNmuS
Amky9hTydm8KseDK6hTtaDtP1pBEHqU6/QjWyBIoeIGJ60JYfjocucVQgNlBFGifxILO4Jc6Oh4k
Wr4cJsznNuYgTwjuk9yVeXlUxqUQmeb+s0Z6fVymWU55Wz+wpBqG77gf6bQ88aLRF0dsqOYs6gsF
kjJQlC8pYb9uMO/XoHx7oKb5CPK+rjq06n3oalJoPDBavOOOd2dp/EgZglWu/DcbAu7bwEL7aVZ0
PnVxn2Gs99hZomOkgycFRFXIG7DeSHX9wP5VWjtwjAgrteH1qN2afYkGl9vLzYaWkO6dUoZhFQXF
ycqs0LboFWALRmk8Rc2gUgaDYmGADNxA0jtz+eMj2mQs8xxWuBwSZbuMLxKkuwvi38E3hppQlDdt
5kA/wAAnXRn34ivs+Ws/PahbJeOwkf72VwW3L+Zf1wssMXoh6XtJjXQsP8PtTG3Be/bzYhHxg5uM
9xOK25ncSfFlncFvHdfAhuMT5a+EiKF7ZOvmWh2+0ZxKy/ZoUzZqlfDC4yykJxvTrRe+dvXDkHNU
sdz/s07vnkhomHWs7HSYXKHeNoXkieSgvDwNzVUd1vLJ3kGb746ONKthC/ZyqqUkigH4achNtSyF
P8Bk8lzhwV13sSxpy4BQ+tivb+XNFhZTlZHwDyK5jCR1XLurPrsbLEkxW3ePg9T47qkrZK9VvWcP
pycKFI8jYXJvKwzk389m8si7bu1aDrnfIRjQ5R3/rKURCmCCrTjgGeO33zantl53l/c7cmF8/Ovi
lIcCh46kkt4TzfT847v6+hdZ2m86F8f9KnhXxApZdwi0jLLxt3veJYqY2CobxfBjZeeX6tvLwVgf
R26Om6upX9nPII3RXAINYMkvGjqRat0XC4+MykN6df0UeinzSXR31GmeShM26YMPBWx5jAOuKLeS
Iz+K7F0/tFKHfovT4hf6jxMNeQ0sEQFCzBNqpPQtUoKVJuKC/04Oe9672PqGImcK7XIKl/nNBk2O
dO+tIsR1iwPdCUJzAWMsmq1SDnB4ywJjVHreTF/O6sfjMiAj0+A2cg9IsWiJ2654Bo17ozFs2NDH
J5I0hL9v10cO90d5ItAe4XAZSHn7kUri2lIdkdgkgTdU777X+uVrBci6wDKBdLDtMbL0Q3n5q0/h
vUP8OE9Brr8zyVLSc93vLNU8DlGAkOxLC2yfAy2KDzqMfayZ8OdykUDe225Giyu0ABruTbiB4Emr
9ro3DEnpKrBLjrDGdnQeIPUkNj8BXmjUg+gfyGJ1Egca7vcnl8/OpcngkB6+wnRt5EpCea5gI/G0
Pjhbk0/L0yKe9U1eOixk/hdBnRDFARvIv01iwXoIBnpAqInjcY4I41Oda43UApFFpAZfujJn8uHG
HoDsRdDOmB+SDEbtBtLxKu8VuGYqX1CJgoZYWry4a+HuBbNO/AICUnqJA8Z3Q/cDJ22nzf967Cy+
779pbO9D56JpvBzcDYc+7R0uetMD7QdptxCbu1vOwBt7d53Yx7wp5d1J8vSKA72/0J+gvDMbNvIg
mtgK93K1v/wtOQ8YJyHnQXvK7QVGEWFNfBHVP5WMu0sNSL4Yb9jeEaiCfnayGhvCtul2p/wmGlOL
yW8sxPnWgWVlutE1X923hstOuhwcwkHG//0fGFxOv2ymIdBFhc+c8zWcsfN1dhpmgqFy8S7ZuhC3
ZjxNwXb4TNAeXajQFXfsdfGm9L5pMpPZNgeX6gg/BM/suSopIxst7Czzje5sg4uWKO2T9NTZk1Xk
q/Fk8Yxoe+3t3XLvgYBsQmAorNmzT9OLEkEGehG9Nzsg/Ljz2DUyWLMEy+8IoJygSj4cJBrScUzR
OgGWK2uLruQSRa2azab+dyKOEcNy2YwjIOjHTmrrSC8UtsmtWQ1iQGg+xz53b8R6rj4C54FBWLYq
LmxiyoJY2a3dgP2wl+d4eLNzuaox3Q7D3UPvHZRxIibILNlRW+9ioUJJnOloeTwRgqhYbgT+sHVC
a0P9jPMw1xylQPvA4W3ITrm9BlkGQJwgJh+Aibr4AZXHMAjfpB+0sNJsF7Zi2gLYnBuw2Ru2H/RZ
dgGwY/GGl4AkZlgA/Y0o4rnnLthbgizjrk5XInSJNhSy3zjHxPfP1xANmaTz/7zP/i7KISdeStxJ
yCv157RQQuSHuT+fv3PbrRPDQ0T89Fztaq5fT/FEfj1XsI+oNjXEuxx3Mc58ydCsAUKFPE2zp7A2
skA7c/g0qUcY9U8TFB4w1GFppOVi5AXDbqYuxenxgGea8IYQLcfuRafuTZ40J9goEDgBm/Rs7/98
m/2VUUyi3QfYVY4Sh/cpqHjlpWy8e3nltYtFizGL6sL2nHikk7DZ5Yj62n4wzW7bK7BVsjr9nsVn
I5+LZSfzWNP5WzSQSbroK+ooEFROBz4ISso6Li+UswjLRuYPihkul0YSe8UaquSPAz4Mc1OLoSKz
u8LPozyC4ZF8Zpv8l/9OowGhjw4aMuHZ66Y1SJ6zqCcTOxhRcJGuPZfVKVY12btBxCMz5k/CHlR8
PmrmGCEnWNgQkEEvV6gX+sm5NgUjLup7v713xku9uJBCIAZ1Kx7z/kunF9zT9y1h699Ph/XLU027
t949mMkivZK4Mnx2eEgfO4VjGsAqlcLhNphy2rTpBR2CewgvY9OnAJOtzP5HCoaRw7J7Qff5bkh+
km9Hu8CVBZO3xlpMXYA8EsMkdYmDk7IcRhD/UObagNWQqDUyy/r8xjGd1YV898qgzXes2lnGiBvP
T34xSDqf98BiwKM3omp9qhw0Sk2Pcbo4HiPtYKl+kmyZAcHXF/NGAS9UqqtbXXUdkR3hP+L5pl9g
Qy9R+jXXQFeH7hH7Vr+QVer/2N6+MKJVfi4aTQvcbKSewvfn7eps4oL4L8CF9Kln/+CFWO/j/Awh
KIQBJi78bJTYn02ltKcKmCaSWrtqq3hKIvj9t8ZLlwcc52Hr+FY++JKNznJ8qXznFFqQlhg21nAD
cUx7xGl/zAlgyssVRvPJeG6GZoK9LbxQg5/f6HwaSxgRiEs+bYs72dBNqn4NoOE53UoSWUZyuqGV
epmn1GKP4KhKwrsPnhPf1zoUF+eNI78UKRnoSZNkjEUJbKkAYj0Mu1TRwLU7LfVN8NETVmU/PW5U
SAMFHplMyi3y58FYRGJvYJBv68Iuk0A+tzXRwzukgeZrKP+IxPCEhZHEC3S5qB23xf9s0QGWXn7N
e2fioaoe3wlfL4AGZ8iMyKAOuOhp6p0ATj2L2klGJE+LCiOBB4GuCN9XOli2xGUynA2QuVsK1TLz
37g/nzlMZreRsELjcsIK3ibnknT5WsDl0aFQXTCyVLxxHs9XU9dBTuvL6vUrSOBa8HRqY9+9zex7
Whu1KGt8slrfZl8zCpq6BOn5ZUD/lsQIVpdHu0GJmtm81rrjOO92lpcvjV5F8P6HsZuxv+B4Ld4F
UAT1UTjAoqSATCSgziARA+BzHOezwOtmodhwikCREnfH5QfKFC1uCcSIqxkb8WajWNB1KjcXIBhS
lT3Eci6Wk0y4PdWmXfVuiGjbhwimaw+jPUFjqZvNBpulY2plrIQPsK6RNA2GdvOv76Sxjlk6jD1n
DwLLpPoW8Szv5PijdAP0ohn1GzjE3Th2dglTuFD0LF3C9ZFyc6LfQ/A4HNqIY9uBbbHoPUdPY1QN
gXANDMwPMLb4H6ci4Go5eGQ7tSUBLw2YQ8aHM7/IesAgt2ZsIEl+Ku+AGcZ8RJ4lP8HzKjlHFqF1
Qgx5lfzR1jWqxsUrsQghLMg4XyuZlmt86jYA8wK+QgjUIyMY2/DCokuqxYpuFp8T9rOPykRJxVC5
0VbfMstOTLpzJI+EUuJsMPMq23UyGStWyKyHuBLBOzRlRtP6csZlIInue45NOWYT49tpMgr1BXOI
MYoL91m8VSRwdsyL05I0ZdAtz0Obi1gTvxiNuX1aJjt+UQA2jgH7iVoR3A4hJ/hw6F6stEyO+BF2
Rj023gSldjKwxFUKEC60jHg5hI4xsX1fnFfwZ2PtiWCAR2diHVG5zhOMBqB47UcHT/gF2XarzI5l
FpDcd2dMCDpdyduWVOjexCf4++m9NucPlg6LK2T5M5fdPzELnmo/HbVwWAT2giOkwKNoZ8zl+D9s
uKuQ/d8HkJfnmxQUGWeT3xE0M3FNTGnzRfwfKAzUj3GWQj5h8LxHZvisEOd2xs34fRvqp9Lec6Q1
GvIjGfavUoJImf3fFTQdmEPAYncn5kKY3WRu83InwICO2RJpNMD612ZxXtsI1b5XejKINWqZCuN/
sCe/1JpZp6owrVpJH7mqlPxXc/7ZPm8YPZxgFvAhfmFM+15kafo01ZA8Wx9aT31DVBsTpPLQQhLN
ga+bRxnkXTpUsV7yt8FT+FYZDiRaW8JCjgNlZhAJ2vA9eMgzJ6niJD02jPqFGFQkuwWYyXEh+gxl
V//XI4uGh9gEOTfC9CL6fFLYWNE53PFYwbANp+wI5FO7wfuiR9cVP9CSbmX/JJMuuWyA8BnTiMSI
js69HTpfGEVGta0hZAUAyerQBFpsFAyCde83QQLa82n+ZMTRLfTjz7g0G+IVZYJLuYgYwYK/fagT
UHnqlEGRe6NZSlrwJ5TyMBpkG8gXvut0tlqZXos5WWV+HiZS0IliQ/Y6adjfWn7vhRiSS6LRDIa4
NcugnBnEYLK4vhLP0iTB5BSxPdNRP27oMLdn9YjLudtIEkeBup5BSoN2jJrHc65zSpMO2rN7PniR
CD+AZIyoc7tEDgcJBLdd+B7ZEkuZKwnvf5/drwAxPhdbN2j1UZsSqNv46Q5NJxiZiMFdfhupQZdi
YpetLfPZMAxAfUY6OoLt/AuzHcpim0qeQzEtmiKhfEqA/rFXLFzv6jQMge1Ik/EG8UsFMz0p19Pt
7MAXG8OdZybOYfmfEVb6B2rXEDv9sgMIbHdvv8z43fbi4GM4k+ao/o+tD/o8UcM4HZz0akrekIg/
KT2Y8oOBvgCtHZawpgsXsZwnoDnR4PZWuYI8Vhfr7+V8fj10hnzuCXNLfperGM0I+Yrz4yeR2VnY
hOA9JTjr/yZL8ptiTnd3POcaLBfSbjRiKJ8c5R8gjBb9NvQLkWwHhd6ehF0IhCwgVlgoRXlY9oHK
TFstXMTTfQ6NUIVN6L7csJkLitiGIIeXmRMPL2ZwECm1OlZwYPhcTTj5OemvM/DMDWIawFrcd3YJ
mCShLsz+fw+lRfdc7UMEgtRzl2433FJQta2/7C9OHYtVy7AhUOLRkokK0PI/rP8+zlEWjvqX9stU
Nx7vG8gvnKwSBAPWrm56nmDeqsKIdjQJj8wHPRiqpZTvRLLJ6TkIoeYGgak0Cchr9ZqENTWb43FY
vTlpRZxyvNjRnNlfAhArTbHg7LvYoOA+MeCR6xcECmvQ5aenTXKGOgD3XLfABheS2KO8bo9spnRr
1IoRaGEOl0g8z43ttLKBE9iGO2iqStakrXn6RPrKKgEVJXIsh1MkP1fWpFgBLgNKYGsWukJoFtxq
jk2+6qhQhpuKqp5TQHYkS/w7jTEH71nY9kDRR2IgfiIaYX9Vyq5Hr8Ik6kIPJtrcAR6TTRAbiHw0
6PbUYinD0CHGEhIZNRSw31QTyTjnvdSYxEdcwJrPmarwljXAQX/VfWDi+cddrNPd5gQaXOLN1lb5
PIpyZeq+PLp2PfSxcAqeD6c0nnIE8yN1RM2qxo+/SkVjHsAWJIhsJRvPX7rS2kNmVuM+cgofQOSB
sig9a/lI2A2aYC2gFGS2uVhOeo1OkzRUZXc/uNh5yO+W4icg4Y89U1F+EPOZizvPN9muS0Quim1h
wEoBJUXIvKq1xUDwqwJ59xN1Os6IL4zLiw5DuRmvAmo2rZo1HGDzmjxLq4LbMVKpsY0JTNvb9UYO
XwEHRGSSc2TGb+zA/t63kOnabbpMwvyXbI4KhrsSzXQO9x0RdHWdD2gYOnnQg3MCkd+eLuj68SaB
X+cxOMCWR6KBX2OxprHNkUQae9BfqGX9BLjNdPsaCI6VJkSHesznmQIbsvM/0+gVIY+xUoTA75EQ
gz9G2ABlyXgCGb8tBc85PexGCkq8+HQ6px/Yr9xCZp8vRrT2duW0NFJDaAzfOZhzpov+pnYWjE+D
+IjQfgEMpVLPm4+nAh0r6sKt5zUwRoW9CkkLCs8ILrmqjNk5a12NUuQ6H2IwsIX4PfDrl31XLGDn
6p0lapobjXIyPpm2lLHbV129hCcGknLRQrCeMeeGn2PfPGJBZtbejf1R6T6iZJM/URiGEuiFHai9
J6vZi72rehUgQaL5pHMP3BNcP11fsXKt8wBCPPemSk7nPT1gpiq1vmUFj7w6p0oHONLRrkTwO7dx
6ic7uCgIRRLbAbW6RjoG28V2K+U+tHbrFc+EPc3Z9GpQDn4G6aLqkcc7cfjJqEfyD1sfJ06SdKOF
M7OPlne3/+xovE/baXOc1mRIm5DnsitCvP8sqcHmmGM7esE0yWHexrOBdn+w+tTCc+Ksd4/bsK77
h96uJVAz+RE8b5CmRm4y3cCCgZEovejnIsfM1AWN5cPx/GZ5NX5PmDVm8WxIE3ilzqOX8P4sUNhF
E6AoV61rSGO2YDTWX3+XFg0uYnlY3/CNqkp7gsqjkXvO+bYOujGWuP3MDT/AOwJZ31cfHBS7m2Nd
ZMPk+P6gK5ld1f8XjAR3EH1rc24MVNxmPLIym7QkX39aygxPCfp96FyHpH4UBR86bdILB+N9RsZ3
/F0U1rdxnNzMsLwA8xfqkLqBRkaxa0SOyg7Abjnpq05T1wXl4zWnZxmRNSBWEl/ihR6RZ51Ti/Vs
VEQ3BvQGMKrODkSVbduwN2l+dS5FMp19A7ruVqwR3z8dlo+KCNuzHt1UH8S8e18W400ybRq9wj7x
JM+WO1JQIZtubS8SlCmqJbRf5qIlqsp+vqu0N6lc9Qtp1uIrGv5VmPj5MsHYoKgAZA3S9N16y0eG
NBzt3Q/lGgSn6svXQ+S887yA33U5dhksyIW/1H99VRVoUEVBpcY1qcY57ycFN2mfgHrH/ECvNdZB
/jQZKzcpdbXUgJB+hKmoa0haHRW+ug/K0czJzKQM3hPz99UxFmHgyngkT62/syBUVk7+XvDAgb/q
q/elcn9ynvpQp9kOEm/SGw/NjNALe/Vp/57Q8N/7lcNLRwTG0iG54fTpS4BReMfx5PZ2tlRr5VP8
FhBb6wjZbvqAIpxnAFXDUINSvNVoHDpGTjn7eYIgCDsNyiyhJioJ5pyHS+Wr2e2mhH5WK0Mj5YjF
6N39mcIVIh9wdkkyfQXq4iEvqfWQNVFKO7BYuKuxJTWAGaynbJwDuSylqxRQTrrj7gzSwjosh5Z4
AAAfC+I4L2THhhFuVlguJTOb1JQaKkTmO7GaPmccE2b42hDeYPuv7VwMbwm/8LtCpM5IJtM6v8gI
Dv83hDQ8rSCJglH78pRAi30RNcpI3mKpA1g4uyGaSQYuQ75ql2uoPYfm1h0KNTAa7BrCk4xPRifj
mdTiEqHQfuA9jaKc13uLJjhP4+j2F8eMV3gcmvZySvPfgx4Ql6tfdiISZvbnoPocZOK3mRhvfIq/
ZlgSnVtPX9hDS8/BO4rXca4lSXM6e+c4IG38wfcL02KKm6DXrHUPLtpAKri9qmD8XbUP8EfcXDS+
Y0OM3BmtyuVmPHp673S23SchV/EqH4G9uh7MtfDZwgKYPqarN3V39ODAt2+pHu3KviKjvEQXrZ4U
dA9tREfd/AEcMSr2UmMoaXsRKMsJrp6D+vCBlZZBAHsetiwqt71jvj8ybq67wT2vR5/VcDsfY+3o
XY1L3OGiEQU2GbZQvO/S2yBmu2bnKd5qkF0ejqBQCma9U2LStgyqhwBiYE95UoferEpwDCrQz6R4
200LUYY4brKTxP53QmC4GHY5gGbXj8sjm6ov+DcvjI930B0KarFb6lD5nrcweU+qG4NonWEKK/AP
PlLZOqQsEjyLm/ShIyRX6hq9hcgrZMOUPJPLNw2SYnfbGmu33AuyIIVDzsQcQ6SfxUwIlM6AkYhi
Lo05bQBfQwDpGees+YB7byaN/gEocES5I/vuNxX4C5LMIpFv9C1qPf6JtFpR8cu1Niot+FgopP6F
BufSoTsyzQc1AHgtbKQ5thtL/emiIrMe+aVj/30FKDw/nyaTODf3jYy07wO6Ucag9ntCyZWQI+dR
k341Jozvsw3LRf3MwO7M6HgqK7TbSayzB25iV2QKxOqkm4Fw02sQV5HI/rVlSaQo3xlyhVqmAQqS
wXS3LRqiZt/TmmP2Wj62vE9EXJElSZyIomzQI3Q3+8bEjis/vNdcgnR2L7aF1IY6j+kgn63+g31h
EsV7IMQi9W4L4YW3lS5CBoNgcMIKh6YUdrCsXPwacqg52vVqpRhti+vLmM2R4Ddwe3g4Ed4SYlDj
o70/Slgy7oDk4DsJk38XWfqlZn6wn+Hk8Xkpef4twTeFu8sZcVH7khFZrn1Lp4NJscjY/OtU0YFi
PqoLi9h4uIynsBGGIpXqCgajFS8yNpwvV+DJHxpdBZVQPp2w2WK9UsyVKFMAIMTJDh4l1yHvAxOp
L6kT+3uwyW/FQaAERCz4Ug66MeZiSkidirL8mzWc62dx+5+Qrg9XJ/u+e79pPEoAdA8RxREub9Tp
QdFnIfEE0f29GVCmpLUTW22pTcoZste8VeBrYgsADzDGb9A0w9bYrcZ7szP2PCK+QdWc69djFUPs
5ZRHsPQ2j+tnNU+4m2yYVkVB0YJYNIB10YNYxi6FIabgpvaI1BlRJrOntpA8pmBTyD33iN8AMuG4
1ff2+Oz3bJN5Yw+bs5Hd+CF07ZS0V2XSAd2+pkso2VHFtF1V0bZdCoLIT5z3j53ya7dr3nevaEA9
4l2ifguf6DME3b2M1KT+k+r4RMZHrCjcAVHIjDFEvcr9OVc2xcrsWeNbFHjUGqiXQcZ5yIh2yUXM
BG6dlScRadUYhAslMkoRCcu32HEdqje1u6ZHdQx3wDNJFRLwESu7meK//l/gJax0f7TFcvHDBnk4
f5v6GiHqp1dTwB14XPWN6fFk94FJK2ICX3dOOcxgHa2T9oNzGrhKTQGEC4RAe8rLcSuyKh+88mBc
uADLz3DT8LFU6S1pOIdi6Inv6LZDa159bBP8UI3msY0R901Zc6Nxh8YTH5YdNcHlDdcWfzfgWcCY
kIomJrqSJzqnmNhIZ0sILIbb/CCqKvwm7VAycYrBZtBwAlAmKJK+uaMXs7LPVojkXnXtzCg1GqTv
f0jE8X9Qiwsk4rQ/FXgBKluYGMH2N8ET8mGvhEZfdqr5ocbDulDNTA5e5RrUyX1jdieeT9tbxoyc
V2SZz0BCTXpGiAKnH62NU4hHKvqfeQCsGphw322OblYTfjAGS2lu8C2Tovpy/UTrnIpgRuIS8E2x
GSM/psM2nZWKuM5l4R8Qp3xDgSQm+bufCVNz21i2vs5M/XJEChrtTkFYbq+UrnoW2Ii9oadYix/X
FqGaF/Be4Kjd6LyT8n0zbMQy2x9fr8l/7Mp82zFT80iPU8STxdM3Zgyg+wikp7YB7tiAoGg3PZtf
upYlzvbbrIyXoxw+JqRpP2GRkIFK+z+65uRDEInmAGA7ioS9YvWCT1xJ8eUI9WCM02h6vH7swHA1
7KcRHllEIsEi2sjrR4hh/WBo7Eww8i/lcXvHvk+lc6NBmEjAGAXcZk26ZczvJk61mLCsBulCv8xP
YxXgTmXaqWwAS3qguHFli3TWvz6OkHF7oRihRxmkT1aZ42UYHwqSk9uGoHvQvY9H9G5KQ+G5VkCg
ooxV4/ip2eOPYSZC3UHhgPFnG8qBkcNiB3lO94FwIY53JYTCC4Luv6Y83hWghD0NV7hB9hnNU7/X
U4ysl0jK2bMYAfsT7QmHjPaHi6w5haDVF5u6OXCQvRys4cNLBHLgEzmreS1moJAP4etGfaM68zTh
AD4FYayE1SUCQnq+4Th+Bpxr51juRNPyYr8IFUCrdFHdYwFtjo8tVFvcD3G/2GklRZNhQjQcfT66
lWuOnfKKwMG0LTAnRHTaAJAsC1RArYNFcGOgiSKgC4y5LB43DjS6DDmVdelR70UZ3w+J5qQ3siz8
h0HSO9yOv7JqZJv9dISiTFfLBgYWNyZuXQTlfbDG+2bz9IEpLdFUu8e/f7POH9IyYyE9n62TQi/Y
udBGeBpOa03hJjqg8t8Wfv8CNO1p9u0M9zMLZmUnDBEOynXhyNQWwz9sJz3ibH/MCqr1N9AVjOoA
CAhTcMot5Z10L0X/JVShsk0iSZ1+Xk522gLcgCwN3Ap7K+XtpNuyaWbQTtF087rbrprBIM2EadmL
3YR0T7yrkSM2/0XG5uQwlVkjRymmSTr/89zNs+bgAwRaJvcgtD6tzq+8C3NSAU+0ZEFg+5vMIR42
FNS8Ed5SXU7B32o39U1J8V8hU77s4aNS8Pp9nso5HIdz6+ct4pikvqLTaNabm/aj4ttA7IrRa2kI
JvpZRHZQoMb9NydOeQy7pgYHCae/dOYd8KyOLkS02q5b3xAWV/tH6I0uoRf1dXxXuMjyKpSvFM90
Z22+TTXiGDIC02kFATbKHY3MTeZcRodGGGSWHZt32/8iTTo9E8ReiCDOLDmrdQJWuZ0yzcN8rlwM
+hS4wOwlgI9RXMuhwZF0NRhbwoFP2JdjgOwi80AAN3VGXgRUQ/wEpypV+bXDNJ6LbV1XyTZFAFGA
dEXLw4YB/oafnilNW002FmxizMyP05wGQlpjUg2ESkVItPAlW+H36XJ03LPd4T9drstdZgKY5aqq
fW/An0xABp0fB4A/j+xP8y8QNGDn+4wyIxieZgGJbzlYjUHKHIif8QW0thSx522CgTtjdza8+0Mn
fy0NgzakiXq5+v7y6wBJAa8gT0yJzIhKVc2RUK0amdzjNON4s9yGi3pmXoP0pixVI1Xrjg4ST5c0
fMG+iXie+v3cR9wSZtWie6vWshamzRxakNM76/dThyroCqw+bSipTcCv3q/CUV3fch6P827QMZtL
L5oW7hztsltRV8Cb5janGYv5CT3ErIxZmt62WulGjHeVtfL3mI1k2fbcHsrp0LzvSc0RHNFI0znZ
Zl3CzCYKuGOVH2TLy2kmx2xvKocqcgXZYr8NWFh80ty7byNWhDXveWxHYgXd5EJNost3SHaj7AbR
RBVGAkbWYsyIoHtOoYtGuISvBFv1BuZ2F0Bi73TdXptwiJucpnqP3YIwjL0GQFgRJF4bi9eYsKrP
0uO6fMdItEv1g1AcUYoelEMw3nEZ2R9PiBWAR1WSS2UJXderZvphL83vWUyWmMenuhjz8aXDIn0x
lKSIGm1yEcn6RKkkIAEJh76g6Yn6/sdCD7qSa5qyCXKkKUlkfxD0idoC0tktsnpGqVtCkJg6Tuu6
kuev2jmu3Ei4ipw40YOyKDQ4DhOpqQt0GdGIkNH9p1bwn8vZ5ywBwc3CjGbEpEDHIYK5DKmN0pI9
f0mHYqTYHwgDvrsu5KimEf1cd4s+9O3SDLH3P0lbzGsOcXXl/pol3tUf5RMC41c/nyF3+hpFMeAB
UOfy5NG9XvuNFWex+Yt5DQSWYHMpDxxBaqt7EY8AcWcJtaBeV1MReWN12U9Kq/vL1g0JgttdMX3D
7Q6Wh54wLsjwMXzHecC/9JINTtZiwmE82Ldie3f+O8q1003Nry3qwNOS2HpMmi/5YKPtwvPbzpWo
AregL5KxUL3kumrNHAjwp7ukeHPuJcGshigUYpNirPbeMrr5gleAdppsVHznwnS3NG62z24rFTcW
TT4oNDKwKpiMC3NZNGlxxJp3EgtJruLeZjV0pi2dh4F7XL9s09OvvOEomCgKagKjmxZN6i+FiJvl
sUPdh5h0kpx9rH6A1QqrP72keQ+c+tH8yqOQfuW81TduJkHpU/7aOzQq0+BgK5zMf4ILThwT+rzh
puO0GpUEKElTDVPCUxzF5cU6Dg7Dlm8dqnRZHnuUp2H9Cva+laFSF7KglcEDauQ5mabo8xJrjrtL
sShbLe10e1ugedb7FrlNZNjR9Bo8AyyMm68DqKIh/YXOFHbR296onVkXOm1QCa7ygVAU+FYv1IKH
wEPkJ4TkeRBIeXf1PXQUd2zwKRVOJsZSGA58wHLPmL4p1XATHEN9Fi4DZyszgOKj0BwbEtIqTOr/
RBJRlZtVcEPAJ6/oopNpkcWJsYCHYLlJ+i22covmroxNDc/WjXXMdIjzrUpQenzlyVgr8hobtoGL
k3ThRml3mEpKB+MVQj10ZoT/M/7IgrbnlDxsq/jg11JjNGGDCIIiauX6bPSFhNCoKYW0oQjkqsD/
KaINDjmOvL9w8G5W+nv9BpycJUgCp1Du3JecN7DBnpcle+w9CBhPcWbiDVkQULOJnF1TLWjxDQ2P
NJKPzufs+Lu9B78lni4inlPbUDUTjRvpEgCfFKxfYkpXhsLVjPazagco5tL1qATDAH184oPeENbg
U5zN6wqK388RTnVMsAuOvJGs7QK5nBqKYRSpfYTzFFvx61fA2bJRyjAgiNbwWGapX2lEQc6fOa9Q
RaAShLYC1QHVlOAaf5XA/KETH2Piau+jNzVgu0OVxOxlkANLtk7x58iJORtMhD/DpWljzKAEqsxZ
PfygSZE/B4AcodCIm+/Dluh/316bV/fUp4b+9T6z7tkmQOA0DrH82OM3CtFbYwWiwbVRonkBhXsw
P1yE6NVZ1YSRV4GB6+KF/OLO9uLXJpQ0UmdWhjUHBpGAVBfotghq2wB13siZ2pdda1WhuAzFq7h/
TA2e47EhxoOn6sqmMPxnYgX36uqmyzpEhRYY6Lg5DfQjzyNuMEdr5KPNcWXZSUYhvE0nH6qco75n
a2uk8vfSiMyLUgArXjvCyF9OxuctBVKrhFCvS/3H4GPQde2pHKRQ0n+yR6mVSfvOr1CLYRytOzRo
6tKCyVW1FpUzOEw2f8EATpiMyqq2PiOjyPxpQtoSL+v+wSiKO1UkZ6FADR41/ojEdnYjfAeeMO+N
Nqz6UjXaBuPDHLBwQ5g0o/Btt7l3/bswmhOOtp8aQMQbjZd4DhtoH7zUqbwVV/ojBd8/5KS+ddK7
kPpZCi7a2yF5plE+m0vrp2lhn8bXlyPtnuasji2FRgYSIM+s7mVpY+Y2tLgIItnsIDykYUqjbKaD
9zdo+VXrZeZHITEiQ3+Iconhk6KjmTpb8/EuBJG9bOXUjYdyUmbXJnqacPqn8PtL89llmhKuAxtX
xN0+RULPSoS9ta9wS/qC5Cj3iBImksWZuzW/FTS+RZCrpZMfg97bxFfoPSRG6dBsIdgtUcBQv5ff
ftyn1g6DSGPkUXELqi6uDbPPFcP0VgRCgCcMUEDb7qcp8foCoZicljHanUlNLkEFDa7oF757seIc
EBe7M25oE7p2cMXtFEixwaVOf25P8JG7nHr4r+70CtSgvUJfPuFxy83vvmuZ23scL5H9NExzEO3b
/fMAnV1SHI/XEk+jgAUA/rCwVUxDOsEYeyY7LCbe7pxwsHIu4mSMCkaMXIQfQQzrG3YJ5A0iHQPt
KeKPjoyVJpDzt1jRGdZtFRpY2NTH1rRuL6JzQHxoX77dXpf8WjFnCOJfsfXYMGX96c+fPStNHSlh
YaVlVTcfPDu0hHL0UJTY2ADMEumwI5yOxxh0ntfsrTj+aEVBtAHjEgLS2xIk4W37fs6gcbBmciau
TdRRIXcffrpsgxMFVQhhFyrCVwXJFR+KH/Jz7Mn0KWdSW+c3WZSxsddIBvKo2rdiLIHx8zM0yl9+
5FpAgzZMfxpH8NxF6eHHALozPYkhp6qnmlAncsInOIb8LJZqhdCdUSS6gLRWwgS6QRRwaGFE5ZyN
77TlPCFK/9MwidGE3yYBafeMNvsb5pY78mkMf8ktcqDOzpMzZ+ZAEIsQUyqhW109R5/BZww/KfQn
vKx6YyvkRUwZvJr+K/sICrNQBro86//U+8+Rr16wYz8i9PcdBQGktAVar8QCRphL3k0KRC0P2ZaO
TFGWSH/QchsBrphF+a2IxQ2hfN+Hf9S84ic4udRqOZ2BZBV7zKUygPuW4Keagazi6rvhyhKEZKy5
Kj8O+IekDH4u7RcB7DiqqsXQxgpj4KG3uvsnAg0UqcKKadecq1KKa0CBcHBWT4PGIf+1QYnpMlZ4
I+DKgAFdrxGUtS+iB5k/rfzWcrQUeh2Y/YzkWxLcsqC7I9QRWZN2rCdu/THTkyN8mih90eHjG9yj
2FulQm0p5/MM/xgGgQBuRwlIBAaEe09Dz5S1y8EII4GZUEH/+rJZUA57AKENvQ85ZntdD1mRH5Tt
e7cmYH/BRF12f+TXcxCDDHHHpp7MNPvnVFC09MP7XktVig6l72aIry996KLyl8C0pZy/m688Fm5h
VQ2UFeH38+/Nu4+oHK6SUHNfYbzYDRcfNPgrKl+d+FjJTpwmXH//m8tSAC4EohkExGTeYNrMZwCc
l23unQkgid7XK05oUUWW3Bl25ZmMNy4vCx4jgotiX+ntUh3jyttcYz6CK0dYT7W60dAPvyFusAKl
xFx6fujebw0xwTWIQarRnwo1guTwHBP4MVxco1YWhf64f+u6yPOuXO5NHKfDsjWYYBF23jg9j2B/
FJ0S//Sm/5raatzUCP4UqjzEjEWUl4CtjizZzBoguQ9k6AN92zIYK+VRvNqTwlCRbdU/xpncThsL
EVzAkvi6OG0ObiPscLTsYMoVmHlJmJI7gTPizIf5TBgzOVAEWcEETT7KBJ9T46s60eT3D4p9uaIX
DyTVdKHASsnvDYhseZU79UQnVkLuao1rzLC8sbf6Cmu7ky1xr3Gw5KFeeDKg/97Hee2eFZxbufnX
yPl6NLLAKCnGDIlQ5/xsdegKsMkzYX6ZsI1syi2eVHXIaQklHElJK8YdBo6lHldzGb67l/lsQvi3
vqiNMnVD/unWAJdd3C1j5UB0b4Gi6owLB5OF19KO0tzWnc6RCIgWK090+Z3eaX1bKdN20TFAthpZ
SFkPEb+VRFGWRkJ2XOIrTzOaHjYID3A2Rm9ED6czX/IHMWOu3nhq4ltJuONXWY1vdyYcaJg0fCgW
FFdZRntiQ99Yzp6jUE7MEPVafKIOCm5P0SqilQ8jnrb4fDVHG1k2LtDHh8IFLMCJzWtPAau4BJfL
90g99IdeHAZDbAwypwqeXHGNBb0yGp/5+8YJwlC3fdm3ghgztPu+0V8PPrtTN9t/I57MiMVbEceu
HJQE64pQhdRFdjqr5K0DFHP2gGfJmoIczzjEs4PjBGV8r3D8aAcB5hNxYsvCBE8nlaB4aKvYCvZk
mlQiJXdC9lQEvaqaSL0IJL3zVTjZjLr7Vos1P1XT1vlc7gOOGiSNOjuQ6et40DQM4bWvwnY4X8oU
4HMXomL7mmWt0WqCzLKeqx1P1FlAWa4+kujHlZjbCxF5YYlsgmlHXOBPgeO6Fem7nZdbl3QQt9/Z
jilCaJw1O/1aCUoZ4AwWN0X6jIJj6KHYPsoTOFmJIByt719vd9imQ3gVJYccK0UXbhO5B4xIGvjS
HGF80y3ctJDbQF2npUgY0M5YcgGVJ7y0leWQNFdgcc4RywnqXPi5WXCzSOJTZrbZRPsuJXGUYFSq
Rl5lR30rMZ2FWTnMr8SdmRvOAZ0NjJm0FbYnEKCGo2nG4BlHbokNw8Nc+CWLjSd+eQbBx3yyJ8EB
13vv3lBwwdFHBwWWxlYRPe8DTdZWTHuuR9eaBqrURRYgyUFykqBQOhc1EFrwV/kkscXD5uA89rwL
aJmPqwCHBmeBDdXIOOEM+H25CqnXcGbTLzYOY4ZkxHuSRsNi5fV8JK/6hIXDhmjSjcm5Yw84etYX
ZSC10l4ZoCxPhfNgp2nV3w/THUMJUqhDns0m9hU7CiDrvavK0GtapnW0FWd8bPfnygq+W7Ai3Ndu
xonGM/aT/cmLKBwBb6rYae6wfQpMAbmLDwL6LlE9rhjTQtSkZLnlwcmwENtgWp5dtqc8VhEswn8h
b87tfUPIhxe54x6pdTRFaZ97qJ1DhmmJKqn0F/2GiRkqNWvs4fpijDo7dpQLQoD4qiwvIZtiuDhk
Yo1Yv/dkvKMnRlPydeFQOEOIgwVHkhLXBtJPBrKDz/OGVh53NPomp0QmV282Au1drmTxS4JF84QU
ps4ocrczKtSTfEOKcTVnRTSr1+cBK3VuO5cBfP9ikuux7FowiVLLutvVi50bJKDGmC0Ia7tSo5Na
KU6+MAKR7MnwL9VVqLhSgRKf/Lh1jQk4TlaxpPQuNWNIgY1axdfCxfdQ9fpG2n1waynVMtRM3t2f
t8iDxvvF8AjdNEZe1xR7FCPn0hWYf3ZoQVdqrzEYgKPt1qEse5xiXjQHPAS+LsGRtImqmoPhcY0Z
rty4CY2oSOI9GUo9m5g2BMVyra1KsvaBoMfFLooOfaEklJOnk6FMXrz7GYgJQfjC7bFQdYhUFOm3
/HYBQKfd3YhJVvtNq5uDNTXHfUBK/WBESEI0S17a0saGAeHpg9hLPqPXXfnXi7Paf/pSD53Nv+6V
yJ79a+747U/wdlnArvLWX5o6JfhM0CXErI9yuLDzqJwmhIGNw3uX0HkPiBLopxZVfHh7/TGuUa0t
37dpBMTJnSlFWLntr7Ct5Fbh3CVOWfnaR8ILwQ02XyACByn9r8TomuemJ0R9cbDGEm4O1RDhBJoG
RmJxZZeXA3v+20FM1J5VyiGq+CSCAg9G2Wkw7ZgDXNRQEftV9p8hw2TnSpXFM0UTMscVsJCQC+A9
ZTQ/ZAf8AO0W7IMWfWlaGfK0HrO55QR1tmvVHc4X3rDu6BtZfIemGsjd/2hS/11FCVmFRVDzZyGS
ETPT/uTU5rcx/4/72MEWB61s8QHUqZ7rzVcEsPXBuPdfU7If8ZE3eCjaJi9lwCil1sNsbvGRhViu
GYX+4NZkIcDjGaf2lvYM3Xiwn7gX9562eTWLxwLrCf6FV6yujtfip7iqjrRenA7PahNRtfVJhfvW
F4MmU9lzwTD9dl3mMf9aUqxeR6yL06bGyLaN7txzbotooGcIExa1olS5F2nu/Nc9JuIqNYlPpVge
l+z8/r0FgJi2BzItauWBGbym9cfe2EjyiZUEFUX0OYwb2YR03FdYOiOSxLBXRbH0gm+T7D3CTyWl
icFs4tn60wyYZ6KIgKDRCU1AEkOa8t0X8eHYVUvxU6o5Vzp01JJZ0EI7tfxGukCZ3dQKneuavc6q
+Lg6Wxz+G/TPoJ9MCdI0y1BLal8EJazTKBdak26OtL5w/ypuFKgganLiRxfakVRrjiBk2mSE+6B/
H8fAogqKvTCgrtUcTTYK4kzuxSjbjMCMl7MFJJCg9XUUw/XoO+wKpv+0TjDZdZ9Xdl4nI5jOPRzs
UQHJIVto3YeOg2pFYHhw10SWLi43onhClpOXoRGShtwIALKBxu04YNeaiUIIdkF66N/yFwSjDH1T
1kXitOPzHP7ofwbdUyTGTqlYh0vml+kOqbmujs8MzCpBY+lQGrWgMuT8eZ65ycyAm1sQObql2OKO
m4VynBRMQ6YvPNUHuQPxNVs9YFxnSqsLUDxCrJbyNL1nHEamhbD7JlBhfpPlzdDZJ2K/YCCOW4yw
ENXheGNLfZODyLqeTdTgBXFmUAAD/c4/LashjS/hVjcWy3uGHnAN2ojOAit6nKp+zsnAcOw8bwGo
M0rXBB8h5kRqQETG6/EwYhTHdGF60Tw+MECx7Bg5wMHDZqCWsw0cT/088S0RQH2VK+2Kj/jdm4AO
rPbz3YF45FSnC6rUt0CSPC3W91lsgn2v3yw6k4iobCzNOSXsjAYihoHfkLQBGE6KxIrPxtRAGT8D
ydOcSD+XS+3+xyBZZNpCp7/zRytcJiZ6mTLNU4k3kzGIfh8eyrrqOBtL1jPoSsiKcWuvVpZQSDuY
aoPHRYhtDrsK6EgPqwMxTSt+z2PXgX3IxLKo5ZFcpc36gIW2lP437o5NZPBYqwQXLTfluvVE55j2
vqHvv4bjOr+3u4gxunifK4FAoLvWs+u90+zJfRbu2VQUReNmm18FPQSb7onpWBQRwmAPmG6zpErK
N2O6t1Klw9RngsVEJwYFN9T+aG2t70Lj4iTBSokix+0VcAQxQo6+F/z25SEkztIpaX8pGARlwpT4
dD1SLp/MKhpO0gIp9wPWIdDrhbzmBSD7Q6Wfh3sRGdZie8G2Cp8VH30ngN17Z6i+pxiqbuHg8LTX
YPnlfov4GivzIRIZrFquxg7ToAFgEGQppug5b9uHks2mgY50LBmNy0e+FxodGaX3XjdDueB1kFpN
GNcRitnS9RNZD/P9Ltu1gGUshbTff2bUSsQztvfDw7ImyobnVFLujVJoH7yNTDb+rMzQ1EVva5In
DjmygNV6tKwmyQ8gNs2c43Ah0a6r42sF1fNSfQaVIl/ej5A31ErDQ1FbK5UiA7vkOHaOm9CPqAOZ
PBV35N9fSIwyhgsUBDSGqacu28Sbl25fHO2D/LxOOw90+U01vvFrDwJlZhiF/UnpPOBkaXD6RlO5
seOarX0W1wkblMp51DMDkzExu07CHcsO0dRFC3BUkWeCV1GrGN47+nTlM6nnEUj5uzZqKxQjbsyS
Qfs57aa1vmbbaKI66mVLIHE2YL1II/4M8aaS9CSPAtLr0Pbr1LaHQn4xkflQZGIGaXHy+I760xdU
DmaBy/K7+Vm1U1MdEmAMuH39picidDAsOA1ZjmbanCZ0E5gNG177DkbUfncOTEPllp/6ZF6WEu/W
qtiY8iXLPiYqHwH7v+PDcBl5jPuS4uhPOp3ubCX0snsg0X4NAu5NOT+BHOMK1dPy2kBeHQAe/Xak
EroOHXAlOMUiefLOBlipGK5eYHtVJQx1nAPpOgPcgyMBI4ouH6c4wsTYrItfriV4KhowsubXGDBp
fcktQ/HTNs0fLsI+CcEYe6RdDHzcr04BqFAWt4rO+xYxGP5eUH/MeZOy7yBT3l68l0yCtYVHM1ue
X4eFVyeLkvvoFw5Hb30/KUMTXUJ0xtiTXN0g+QMkMnSRboQF9Bb5LLQhni2fDG7lRnOdv26YK0lp
9tO/A5g726XrHGUaW0Y8EZlMbKUWS5tKOHLt9A5BIfEgnCjP51/VDuwpteWuTlJcja4Ya/XLSUCZ
K5x3IrWp/WJFl0v444iWNjWIuFIGjl+kAuP+I3RKDn13vPLlFJ1sU6wmtpO8Arre67O0NQmfjPzI
bbBxxrT+bMVPLVqNqOQ6xhQfC6CmFw55viLtdVt3h7cyRwSu/CDVYzu/dRh/jfmNoz70K+ISZ011
JhmrycUJwXz0pPj1DzAxGvBoPNjYgFvpDgIpiPCMOmdlnT/IJYwuw/Y78WrFlCGZLH0vz2Avao0w
/0OTP6ele9xIhdy2jHYkcJBeqWbN4lxbaPGH3/NU3U++H4YxyGxu69P6+kuuUlB25EiDMvCCPgQ8
PI/dXpvQcu5JPwfC7F9uwPgGAWQ1Tqs+BbDQKN7UO07A9v9Zfks58B6wHevKKqb0sKGIB21R8tdE
61UES5xvGRhGiKOOHBxfEFuaa5y/W+a7xpSw6NxZuKIMT2nSn741v5iaJ7S+UesUoCsOXL9573to
NV032JGQX0+DbTITzfjBcf5eCgkjDSEqkLtuGo53Dmhs8u/e3F90y2MZUejV5AMpsthutffjE0GO
IZVlLJlb3Jq6L+9zzCjPD8A+RDmcgJrVrvy/avHFu2fhRJ+zl2oXFhDL8soVzmissc2YzzgC4RhW
Vyfv3ngj2Fq7DCqPPyC8p7Ul3wCfHfH5z81I6dwcF9qBM+Z+uUkFpIOxmyklQsBHekDDrsvb6OeL
aw/SxQxZSGA+TKeuFPDvkM/GOXEGtexFzmskN8uu+PtCEKoBm9H1IpvYiijwDHXmh3c5Uq4/IoG8
ylkHSCsdgyIOuMNd5nmWGCjHKtjWZtXMMA0rew/QQrfMVA9xx3ROPeUS5MGQ0SF/RSyLeCkz1rnc
65Zkln1E2ubWi0jSxu8dHd+rboR602Dm2/qvYU6kz6g0O+qXILMRMsIikXKUbEFGcpVzFSLudG7a
EEzU5L+i3yowBmgi3m+HrOc1WfVrsvj8w5NpJb6U8vCbf5S7yJG0VTaob11FFxYuAc8e3Fq7J4Ni
J3ZnGl+qTHWhEUuskb+gKnqfyDscyllmiWc93hpgJG6svz+0td1mCP69m5joc+E6JTmFyH/SyMEL
1Q6Hs2wa2+BqlC1OjMGq2CDPQXdjRsSHQRrzhCTUHbdm+RK0div58n+ud1B9L7upvXrqztXAa7s+
2+aE6yiJOQRUthCouCy4Aq4PC/aRQzt0usfQjDxMvy/TLXe2R0MvsTMHacmJF4TKvCityehMUJUK
4EMIxuvb60I+QoECVSDOJFzmFnNojHhcORpyatLcW9GMld2gBs7oLnr8Ir/ziJD4SvnoRNt9xnzp
Kx1NwK0bw7hEAONeN9djdzgyT5pqPL09td0z09lTdcriHxlQFhIqF9PInHhq3MhnB53ijq+119Dx
r+kR6F/DN40duhh9MoouymLpSjARIyobFOZFfPJf+S0EVsMXlg+rqy4sfp0r7bxIy5gZnctDmEM+
E7ZKcbdXjjlxtFApV7rUM+5HqkPXKYBn3N3Cll2V+hdTMI5JQJsgpi9g/GSHy3JPsN4lKovulFKl
hCvFe+Xd0afcoXXuZcmY+sPt1Ex/Nr0rL7bySCVWtMt+zZhUlfL6S1yPID/IBCHAi9xgrnhcfjUq
dGv1Bq1DXYVny7y1ML2CSYjQU49QuMNB3bqdYcW/3fJ5+gat9+CXq2/viaBsiKPIsCllHsTbo6Q0
7ZksdOi7bzzG8R7KqSDQtthPXuh5FQ3kUorM4x4TEKmPAUENz57XTB1zcLEpawj6taSOvuYthwzL
Kdn5EzTLwPqaKHI7UgthNG6WJzXOD3m0wcBCbfKNYs5wqkc3G3j0MwkvfoRKqr+zt7dF0aZdjWP/
qPJqb9Zro4XFlWN7LuuLKBTJRX65KcO39fA5kBPxTATwWKltT4VHhJaXMBtQI9lvS7vXMRdYWmqs
b5Gnqf3SVv1cJLBvj14vx3QQJj2CxQSoaYmT+MXbcskDvtNL4CDvDR+TOoRi28zIIr5wa7HodUIl
YJ8DqEOsbXjSZIny/Ycr6qWvrUJLz2y6pEL+cqGBhJfj/Qx4dOLhnPzaoDJ5GA3GBAQ9xYjNWA82
Q7FBR8GHGkssiEnHSnS4uyL3YnuzlNwHUaVjx0jrTDUeqX+YE8AdKXCHyp3rWPLC/AV0V+0FBwcY
OcGTsy8sEsR6Iz2guz17OHbhNmStx+2rAepJCzHTWzY1M90rxClDvN76+j20+a+aaHBSRL+T2WyC
FjoH/hzffwXqTLGfLbhVG/oq36NY8lr92n/McLe9jTHcXRCf7hc9S9Q1N+TyljTEY4ugtQHM8w+F
mYoz/uD2iGFppqcC1Si4CKoH0oEpd42Q4jsShcFJg10hZC+OX5QePuUwfb1YqAb48MmMsZKwQ5UV
2xEgwWPtPrOBt5vA8LpE5hp6qotM0e7DPAoIK3vCH1MFHPyqqlSP6Y9NZwpfgBzicULrGtnVGcKw
MUtTQJVJJpDgSRlEPhlww3HD9pSu2nLQUvEoEi2IDfupNsGt80TvJ+VwBAZXm+0ucpxVMXTagWRi
cMnCPm/D14EQSrj4dx5TgBGwXtk/Zwhx76fPT8AIxHoUIu8mvXBIVnQ/H9+RQJ+Gj4XGF4KcYJ/V
R95glq86vCZ0kh6Ju55NRfXUAMavEoYvQNmYZe6qE35Ax3d2ikJpShZHTlwYntoLrOhumdt9l28k
VcKfCAu8h0QFzNAU6tsrrn7s4RvwWJmr4imN/umAHZLp9BvnagEYcoydkWJ41Kqi2FhhvRcHiAgq
i3q76/kgMyssYZIMkRU5nhOR/85MC85c5xA2AR9c+OLxJMBYdWDLYA3hBRXsscJiQUG7FOo9PLlT
WLljZHGFeUBF92AQIlz8y/O2FNyoliljwy72jYHTk4AoPRbig2A/lqSOLASXTrFjq6CMp3Q1s+Ho
yJah11yUkHYH0pdwScmOeDR+4QYjAfcI1En/ZM4JcPWAiBiNJhvoodlZ8HxsCGhcmhER18u0Ruwn
grQRIGeOXEDOTlMpjUONrWSS/QWZBgpa7vtrpXlRNpuUpWcfZcCgpuVl19knN4Ymefnr9SMy9hTR
ogC8kXPGk4I7kV5YD+N6IApf+GKsCJIxa5suNLYQ0RKB/ftdp9XtQEWpjWWGc0H9xjPUxiIxZdSq
gFuHltd9trVNGdcvBQngFv7nFPyhiEQU5qvWBe02ELY/6UNL3EFpH+sA1gihUy1s4BY0j7qTFnfX
G12vPTRRo0c1GDewGKofT2pdQNJGZkmgPSOcJTMMfTIlhOK5Iflwak1mQHeuqUe+v8GktLKRUVD9
jpGNVF2x4WGxmj/tl7aQxYByYbs1mYoXM5xiveD/d1stTSfLVReAD/s5uZEt9wXnSMwlHPRMIfjm
xVdF3U4QsLO5HPphQMh5wTlo/5u4OUDQEZNdD3akwvHvbThwYX2tH2JpSzsbo96q32DLReRNrqv/
L2/NfdBEjZg+Du8Gq9WuDSMPMDSPgv8YuLHQf3r/sb2uY/CfSTJEbueVAY8Z5+wKGl+DWYCEL8cb
UQGSK3lQiNP3fsRjBEOnh6FPrI/Lbkme8Yr31aZnr7++E+XkoideWpUWgT9hi0CP1qUirmnzqYo/
8zdMSxHyf0ktavlOwxoCFlbn/nVczLlVXUxQ6o7Qy7Y/7rUcXXOv8T7xF7TbZITufml/wHAn4mew
IrmNp5/u0o5ZfvKzO97fhArRrebjjnBUg4bbGgTDr75u9D/nCZq6xHi0WgMzDnnUy8F4mEuEyXdh
lfn5PGYM1ng3/9TKYHSrvgPf7Oj9/q7sbquRRXmpo0sitRcBeOL9XtuwR61Qyg57bMZi1at/iTNn
Jlvi4mMpqOPvRUXWG3b2svtI/M/QZhRoOm9sNRA3Z8sSShYRjtH9vzxuFWwL4peQmCnBaWy3mBkb
8I/24TNFgX4vpwZKCO+TDilXlAwGdc2RDMpEu+2io2X213gR0uTXp+17ZCldk1r8M8Si0HxzAGwk
0jwlTweeNMu+vr6NeyfCnMkqaJwzAw2EQxQvmIjMHPMO1JkjbjTe5Kv2ZKgS1aB7CDXPvxDZTA1A
CE3PfN6Xao+ihE5LDjF+OhWIn+kadO1wap+W0IjuJH+vmzmsx5a7hQFGjDrCv/ojFXNuLHa17jdU
2URkKRQzMqIUV0o3y2whslBBg/Dgbu/MHUYYZ1kb8ZF9DZ6lSLhBdhcOSFRcnYhX7jFwQuz0C3tY
A7eMReUFu2ag/y42R7hXrw/64Ld4fPakzJrDk3TrW2SKOzGQi6n+/d+lvYLU2QHjCcN8IxCY9VkT
saj7Xlqwug9DH6jh3BfKoaHA6ShOt5f9vB969QCTyIUScW27w92BiqwpHIVR5xig5giDcVYPEw4f
/aGmBHAmzzEF5qFy9JXiEoBxxUXb5fHRwONfmhyjFQVJ/n8UIEbkqyeBNl8/0Oc6qRQQXzNauX8y
DOKWfmJ4FiJ16y82DQLALeGozNj4rA3num5irGQdM4iJUrelxQatQRGrHWTyJ7EjovFWlMVRx3Rk
JCMkDDvpt1k1g4HKuTXEVQAFZk3Sd/nUrOJk+wSrOq+w9XSojg0RKtfjLP1faCoEb5kNDz+5+C+h
1eGq9oeT0qoxWzCZYZMYMB/7ZNNgguD3Zd0Ko/DvtSUQY6phxJn/2umXno9jKhrTcsN0kiVux7BZ
vFHxFyah/XdE2Ny4c5gfjDtyYM+gi6xQ4jZTWA/TD1xDF5gLfjC51VHrgl82V9ZXqyFMzbOm5cJU
ug+d7izhKroq6xHtsvwjz7L5OYqc/aHMFlMNV33rB+v3CukyBtuAogQqvuuWeUgYjMQnZLLyRJXq
XwakFV+tN3JAzkuZ6cERDblceOZsttw4all+Xegw9wgj/ARa/PksipwL5OxlblKp6Sno8Nw29CaE
Gsf/lllARrwy3sBg1LMYgpHxVgUnLzAJzWTsRVSP2VjbfwOSzv2le8vU5xCHpIGGduOvGowj5Sl9
0GxT+LZbn++PE/B2R1uNuk5w/ny3V5u35QSF7YeMS4t6kRZrQXnuU2UgaCYg/yfUUpczqVe0TsoN
eoXiY/j9HNs+hAU+EtqRZSMc1kaMvSu70SLdk69y066k+73P5tj4IORYaOuzWS8HBtPbMytvABcu
3IkjWaG2k8q8euyluNmFDuxMItbm+KNI1TqhYW0OG5EJ7Izz1b2TyEFknxLes87K4k+3Opbjrp1J
TxnKsEMPJlUhPU5jJAvWkn74JnEmYv0hP9LRehVQFRl6WBGtfxbXs74sEreYpv33uuaC/VdibUpS
AJMrWRwBQwCIpnJ2Aw9ma1crNUhpAQ//f05RTWR4LTAPQuK5W+e3cQKk93bzYftVkTOeDo7cGUuh
hOTnnxhQgGtOqYdMjocBe3got0SPBRArNHQtMgAehvb1FtTz4nnrZJOYspx7E8S+6M6oHnQg/k0Y
Eyp3u4VJmcEjL2t/ABYgppVWc0Tje7CEXv9rbtq9awTvqQnsB53HmKJxAe+rzpNCQuRFVdrqy0Z9
8vmO1opkeV6mGNU16hXc7K7j7SqsS2f4jtpHKG1ZfmFGpNZ9u0vLYlEgmOWVuQJ8S4O102KYctMT
iT75I2HrTCWqkkpIoc5zlrBMEuYPIfz1kdgEAOUeIi5fjGmZU2XA4k3HLOVUW/pp9g4bo66vxkUm
eoOcyORdQTxarucMXhWbLV/t1zn5TQ3BFe10tmIAPWyJmLatB6wXO585JgAWm00xRnr76pdJjXj3
awarBoA3iFF9e3egknwLC1nNxLz8FLCSOQDcCwv0OfU5+QOKVPsAuBl1HZmkpacfNmfCBAarznJD
KzwLuDSj37hQHyvmA2oYYgU2qqwixdA1/dyORP7vBoUDBUKvWgxucmtKm2Ea7z2AwXKA2Z95TAAk
H7lcjZWZGxblXEE2+c8IOw4KIWnhG06AorzjKgiiOFic99TanlTmw2pffqKW7e1MlG2FC5KOE+sd
8rVqoePpo6kYNeQ3v5sYKC79q8QsCFG7IHY9rMqOkrbCnHIvb8M0Zp38M3YteFPlVuyE1Gkdv0pC
VbTA0Em6HFsJxZhaP55mNo1KwTM+/W96Gl2ZnKrKkdgAcycMUFve6qSCzjpn9xcv8vDdn+dIW+mM
HW3NvCzXo6t+3Y6+1DsWW0FUOraKIE1U+3q7R5ddEBduabOKXXrkcnXgxFWP3i7tSFUgqVeqHkJo
5au3rMvmOnlM+RqS7CpxvLEDG7O5teIv2efZxKbgdXk3gYW3iPf9ZLXm/jVjTh317+6X2q1MPMFk
JJWqFlwtDrrn6S0Qrf4ji73TT/gLmBe5Rm1UAe96jzIZSAjlOy3m1rRKSr9gMCgPzcOuHw5T1OjX
EoRNyGgVbnLtWBEDB8FpvhXKMCxEOtJPaTtZ6c8bmfYrYhk+JV/1qBxjF/OqyhbATi+OoYvxRepm
igfIHZdrWWabkJPtffS3y74lMzS2K1a7CUiY5ae2MB9qPwrgzUrE4k+0ql9SunVrcUOMRSkOG5rV
FvRO11094Au78QOx5oehDHDKEBycSML4PKN6sa4b+UO5/3XhnQeiLC201RBDIsUlgjdaiqHyLeOk
Hdme3EKW1F7vU6QPOKOTpslC04nOiCWrfuzlSLda/WLA6Swvx4P3cLHlPiKwRK2OLkj0PebkxLHg
9kXim63rAATYlyGFUUJrCAwTxoQxotEe4RiKSKbr/wtyDJcWo+gvo3I+hUi83Ejrph3ZvlOlnnD6
QezWnpSIGEXLpwE0nVAeiTYeOnssdaYdzFZG7BK+/B6+2JHGLpz1YJPqeZzf9aD6GhTb7KHgfuEw
44KBe0exlgzsPTK9MEvzH6AHkItVqFpWC9NhVyAG8BsrinNmywrzUwndIIJxUfisuFln1Niu3Cdx
ce/HrHTkfgRO4QlMz9ShjldGWSKHiDFwrnArjFQ6v1HXYdVxlhtZesUF1OsdsFvM6VpeWOjYVHX6
HWT9KtTdlbQO+Q4CNg2/weLY6r2tPs41l6mloZVqo/3Oa1wfuoEGcIWFWDDDGj7L6ybd+v7ECLBX
zcBMGyPczTisQWFxxafdMX+KcWCXDiRJmz0GJZPSHJDRTbKM7PK/tvYoVXccl1CUMAY2Nl4q+OyO
PB5dhHgRnKClOAGVsa62DGh1HdwZ5FfbY1xgDkmmUp2IPzvV1jUKoMFV5u8q71oZYhB7zzbXqKW7
v3MX4wOhuHWuYtuo3xAwgOkTCddM+aN7TY/ges/OQxQhmrDf5u8QlnahrqVJnnE+Wu3JkCrznbeE
z/4DLNplYIB2zm97Na2lMiVa6nBbDV7MR1eHlb6VlZBP3S2LKAEk6TRp7aqPcklNJGsiNs1zb/jy
nZTAvoVssfrMUcgpyIJap9bTDz6+oCKX5MLermsKX7vJJcZAYkv/mZJHxQKKYgfva5i1DU5xkOMU
Imu4QmwCvYjliTQDIKhiNR8aV5OKsn/yyUF6bA2snfnjlDZPp6CjSSUSNF2msLk8KkUAD277LsV2
MC7dJTv8ksjX6emZTsqm/UwbiBGD0hWakkc3W84QZUADG7LvgJUkroe/L+b80L0N+4Li7hJmpd5Z
N8pgEH54vAjwlaowYcqDRlIJddmkDLXNfraPKg4f6WAxCzTJIzoM56ZsUy9tH3HzOoqyfHH0FzSj
jugAW84d4VhoeyFA85RbRoWZX1BDJdV//4nORB9gQ5i6hSawdsEi+GJMazcgsK0UEWh5glOtTwAK
RdUirVIkn2wnJYQU6ux9zrvs5nKjtUQX3kmUaf7Mh1TZvtGDbDqNVSMpnKZ0y4j6aXhcxRji6nXf
PiNoFQfbfnh0yE0oqorLQFftRbcMXU4U3I8QHrNIymB92eU6/OgxrpxEC2nxKlardZRWaksqy8yn
DZ6Srs0XBh6J0Mo8N5o3qmRZ/67THbOnTdIbs8pfgBX5g2/rACBtYJ1AWeZzVbJ7oHqifajVM3Xr
mskDBR1flQNBvcQ39wzYp0aPHBOA77vWJMPGH8lu5FCzh5jamKrC6GrXFm5G7SHdnA+ZvQ+1fzR9
CA07g7eFMAkN5TPsKcO5A/NY8/oDBEUpVxfLi+U1YnQ30r5CpQAuI7IizsFoEUgS1HMC8Wk6NSZP
ZfaNBlPa8N1WVLDVd+kct2BOjH6PelKGMmOIjrzWQPun1ZqaQUwu3sxusoPWFR52KZgZlQIz6MZs
vvoykTi61bu5sD4CSLOPwIdGmL5PX1Og1PIKwegddgMCkTU2bUq+imqcUQhjEUxuBageen34LA3K
Dq0vDCOEoenZP5d/STPlT9rLqm9lo20OIGLiGJ3utU7hscfQvjFHb3z1Cn7QcdVhUdgJJ+3OHVF6
auYHbyNnKv2vS9q3Uyy+6fO7yWbeKfLjYv+4yphNifwS6LX5zOsfr8oEateLLti7a3Ezsb8IB9c5
DXpgZSCRlf/7s1prRBlGscuEd4Jc3ArwjgPR1gTJDel7iJ7N2a7lmgihdkUKdUuPp153zlmCpEY2
gzkMkCAKsIeyX7a7zNaxUasrSt99CkeycSmCqhknE0ppfNiyiRKbm5SOn9Iwr239X1yzFqmMjnap
gDncP38COWzAfYGLElQgstXs2MGEddamEaPv22jgiW3H1BZ4CASpeUOQUo3H4uBRSpFe2Te0SZF/
UVdZhU2+/HgJL+vcbTnRM4DZby71o8SK6xRdPEEJuijlJAMF4F6EcvTYSAIF+6F29KfBxLdiRrQz
eCo7F2Dxx7CE1ONW/DdezqdvT75MPA6Wlg9RPvypClmPE/KcsxkB3ZBQPd0L2YnWywuexD0FW9tB
GzSI8t8Qvia3HEquAgxRYtrsu8UyxubQB0LUR3i2ENZC1V6WD85x8NW9haWsXNy9Yc+AA4tMsUFp
5U9unWS6ixfkFqKodrUwisWl1MDX2Ehg3RgS1vbRaK7LQ358jnguKB+4ofxLwHkI+nnjpLOWjfg4
YCS78HFwTkUKucTOT4VgM6dIuogRd62xUppbmH+mFZNYb6zyj6zhwnaLCCXcrcLPy0atcql7HMgD
llgyAWFcSOW8B7iqBMNmi1baBdLtDZEcH+8qTcIqPCvp/vc3JO8U/IFYnA+McpqllpLsH+ggffrE
5NQ+QI8qgOHMbSTZCQgLVbgKFmExWOObT/VVUJCmiOxv2CN3pHScPiCQ51syh7HOSIXeS4Ejlrrb
Ad5MPaJgzoaEsEb8j4X+04Zjnlu/xRyT/bpYCcNI1SY2JzMI6WKdEoNbcyMBRiD03Y8QHI/YWMNY
wNMSu8Zn3g1vMj+4o7tNXAfYkcENRYv+7g9XCcAG4oAN4Je664NCftthPx99b4RKQGxWe78FB14L
cWQOsxDeKYYYIXTN8UrporSTXIFav6acFLX0TwLoNZ80WxNv1aAeqy7ysfQLtqwPV1Qao/FkHrcE
e5cwCvAAHxcycIcsMMzlWNPd/sBv+ELe9fcPib69Ih7X6HkKfL+gYAeXfCd8EMUEmrS5tzWObZ8x
Fs4wQ5TN8CcGsPpBQKF1AHtv1eJXiBntQt9CXsTinqjHBa66qXm2hw1sukD7ohqp4zsKHPOm6PS4
aeLJwjafiJeB5TJ8Gse2Ct+wH2D1uaGEpl30SdVYZhLJnBnMjZ8ugq4lDY3Gbf6q8nFd9d5zNupC
hH98Wxb1hSKgxT+YmeVz9gLIKvZTo4X14mqZojqueoGPO9QgyG3OClxGzpEBIoqXmaIl4wwUqTHG
xvfAftyeGj/HltnihrwG5kZG1VWrwxxRNK8xs5Kr9Fsl/K3dlHT14SdPX9VZVJa5CJBTzrSFjG2Y
g52lKypL3L6ZMjvkkG6HnsXpegHaF7Eqz7gVeGRQFnvrhtWXT6vkDj/vKWSDl0BG4wJc4HJVBA+C
iJUgCiZ2LArz/PN7aPlEvrPKEBYHanbz7jptzHOuhyRsqUaT6stwpI7Iyx/gyvtuqD4Zx0lQ9jT2
GqfUZr5svZqHoe4MeDOqybzEV+HmklROyOQgJnGP0sX1ARvLbQAJpFT8BoCQcsJ/ZGHUOPQWh2Bj
rngwvQ3ducvRivfRFD1DbAO5DEzjcj6X00Nc21NUh4WP8msM0jSwr5Y8WFpg5AsuIQR0sXelgmr+
Y4iDKeiOjQi3GtqsofjpRP0sy++gPvh3TSi72yaTb7aSF+hJw5jaVz3VkxdFOvQKF6ab16Sgq2L7
R7jirw53UrOG4X80vcoODM1JSXRbO+vMlbHgo76Qr8KwaFb5Fz0OqkGNrkgvJcnuD73LWdoGZN3j
5cCBmzXnJ9t/fS8Bcib9pSUN20ehH+NSdWHN09zoorfigRJ9yweqcxLHvOHnkOxp98t+UlFy1Ex5
P0WzPtZoheO4DAxZZA77HfjQ0xWwumSjCelx7/t9VdxG3b0LaWSXp0dWA9CLj/RhGWjFjed3XAwi
plGA3ohwyaYoFFONLsDlJtjY9vIkkEmlV47T/ExiP6Hpu9+WRscdKPZdpwxNrvKZ5QAdy8jArRdz
hSQQ2q9S+0i/jO0l6EQ1waCDbMGbFevFJj0X7ww7IYtl6ZbOXle2a5PsuHJX1Y+I168msok6P2oT
D0r560I5PTbgcB6I5+7KQCKv6J8u2skzO2Lz4CDHSkNkYoSLPk8M6bWDM4oh1hMwbzqEQc6b0f4/
ojoMHZpVk+J++Vm+pddWk/HQtzgqoIpco6qAGdtYuytPnsve+Gaj2r3/jfHCM9b0h7soD7/c8gaC
44Y7wZ0DvrbWGmo3KzWZjxuf/Z7yDkF7/FuRAs7I6mfNA1kb7YIbtHW6fW4YwhaQdiYfv8lXuXnj
Ud1XrfzcEaOxQ2zOZAV526TC137o3tf5M2ySehovlQukXbsvu5LciSLZWdnqNrCJGkpi14pt1zsE
fU0wIAnWr6alG/cVy/LU+vKskJkY2CU8hajkteRcYRVlj6KAGJGV3AAsj8RuI59wC34hXKzaEWd5
GaHf8CxvpWviezD0i3ck6nToMIB8AryhlxeH/z2U1zS+ZPpw4N0FcwwthIa+/YDkL5vqGnRTiYTa
KY1AZVu1AUCGeSkJyWnod7bs24W3d/RbAgiWrDpcubFiyQY6imqTCvemWFoAPAf7mz2suXSIBZDc
0AtfJDKoREBQFuxvw7X21QW93X/LX8dl5b4nJL692xYy0YKCCcAnN3SKbmAUH7leH52UuQPTr0yL
dH7tah0sXV4olNChGkPbt8dOVw+AiOg+AlViKbemN/PGZm8jqb8D1G0E0Djz9l8J66VsEOIsjcl9
8Te2Jv9DrNEriCRjdKZ0PqZXOV/7A1h1XWT2TC+XFHmpkDhwRRn5YyhevYXLf5T6X9FV7aKiAVCl
syp9OApMjkNMw7y8djUJNy3uLnfkh2PKLGNgV3r9/mmdCTPhE2gua7y5wAsCyAUCTRvOmOfyy4oI
io+TQhHE/QVc/UMDh/dNQF2k2gRUHIAYl5qiZY0RgGhn6cpTZewtjegq+9/iSBqhyBhPZJslyKmf
d1ufgTccWRRLkz2ZmCw0v/87bnq1JdQ7y4ExvpgFNr/eRb5PxztOgIm4B0DNfQZ95q8D9StsiNH8
2xuavNzECQ1J28dKjUIU7kXGYcjXjjjoN66cDTTuM2vNYpiUX68uwiAKJ4QyYQshr/UR0YA/ydkb
jRPKuzLBlxzHpiKFIZ7UkUXUAb03yVNQnn63L6975agfCiqDZeVF+qYQJkvetk2RQgJTBBIeb8FL
gBMUaawjWvaK5nB0kcK3xuDFcgcuIo6ih24gbcDBD80lbJcIwsFNuN6wDcCJpRvZEL6v4gOS6Fao
M8j/csVH5hpUtMVbPJ6GGhsp+DyBIgh94ENaj1smTLgR6GFGrt65m5FnyPGxuOH1odtvuFevIFJH
ERd7c3eZgsYkYmtZTNoMotn5JiG55NsK7FVXy449EGgdLiTzJbpmFx1YSOSJuX/u3TsX84Tl+eiS
8hnxQHdTWtitwJ4JDaOs7OUuuKt4wZXlxLeosHamSki1bkLrnqDvUKgO9Vnv/HAaMmBuKX4Bc2nz
HZKzBP8dsQP+arPOnNXL6zg3Nhzwkjz1yaNLCxsm7vpQ1h7r8NByUl9LvMRlpF4zeLDldhHd/CIK
3fsO8YpWE1+BXaxbOC49mL+GHgZ6CbogiQYNAtDBi+ln3w5491FAR19HhTh0zy4m1GPV+73tu1r6
On6Hf5SJ5ss2O1zbTRAY0/FGuh6ZdWjDbyLF88Eq/M+MYCkRDCvGw/4Dul4fGWDyXiC/eRE5DS5L
dxS3L8JJLgTSzXzMo2Umzb6tnRYfM3Wxu8zuyc7+rgCJLTHldW1Gt/fQEm90gHVipg/k29bJJE5m
ykgKbGor4yE7mcZ14d3lG6OeXRSZLZt7nWJfL1qc8k+p+ItgumuX9quw4v7Ckt0GQmaxgXtO1u4s
73b42oUHTCZ3aNBydjFGUMwxKg17ovOIAcd2iSGT8r2EQdhItpVxLEKwByHNft7VCCWSZyngXX9x
RtEwIyUdxIGo03HBgtlMVWmZcKLDUBgMezla6JPZ5yEHYWkIg0ODKn6KpKVC33oIzKX8nHyUI7Qr
aZZ/Blq8O9AwmCFsBTKb6lBSFb1SM6gRydyZxTKH+5lfBC0dhxw5djp7ueB+/s9dwYqI4p0+2iT4
L5EuyaPGfmsM29upv6A5qY9KX7Xut0alQQDkB+o8kzUQ2SVZaHk+RGSowKmx+2aTKOvQX0vEBIUt
CXyxl+wxw0vvl33erZZwm72sKC8Rr0wujV9+gLInzC4owe+jO/p0X6BUgMLrTCVBMz7VdaNKUDCi
YE2w/wLt9++CoIQwA7tUXq+CIEG4q0mArkbEzm2TvIyeXkIUrPZp6lpNbjuSB9lia6hEiCVP/NtH
VYsgaidxdm/yA/0TWlezHgsrYgvvFKnoMkR9khnx1RFzye4pMdIAX7cDEEHbGW/2c/Ad4sC1Q+I5
FBrLb/MVfcF/k+2QyO3w5/ZNwBF5B540VQIpWfZGerVveFtbL0KSoQ/8Vk4ELww5QQVAphh0u6zk
EToSXvxv02VD4u//xnxyn8WBHQ+9FA5wkpGjTwfeTptIQPbE6DV6NbhJnjgpM5X7auCwm3fWIMPI
dRLpHE7PlB/f7XeGQBpasnEobo1nb1MGTJsVjurdY7JAxxegdwZzOV5T2YjCwTvdK6hFc2dYlRaH
VCT357uAzlilAEM7tQ+h5tCtf7xMiZecvzDhyqQRWUuKsiBYuSwrSt05sLM3yipgPfg2Qty3QcsO
ZwbsAFa+ZcgaIMV8ropCKAUj5Ws1QSVf+nxFNliH7ztQhEK7EWXeRGqtvWJkQzzXrd4waFC8fljp
M+KIfErr9eeAD7ILwYBdOGyU0l5n0wu2Jtr5zQVpjYysVP4PbeXyqHu1A/LI2YU+btfEcIvXjqoy
G71Ud5+94qhAbcWgYJVvnL/SyIx2wm+pNtkKAh715YyogatzBfc5xkPSeuDd2yuycAIaEnC6YnIa
udVLnuPGmin70jp2OuIPXY5fMcLOB9Ewt8Gga5M8eO0JE+7iFfa2Dq9mH25HUOS8UU6S23jdW7Fo
+ys/RLnOu68lJH4ruB5SzepxrLqdQV7SbtOx1YQz/16a4y5yFOcPaI5LWZdo/1uWak4HXsxki55w
1ZEXPF77l+A8//QF4ds5X9SUXxG5eThQRM2t2sruJ+fzYrX9fF4Vr6+UXeVNnyySdn+h2EXLgTjl
tdQGChBihbG46wIuw89CYm+6INSKuPXQNceyZRpvbol0IA5EflBU4XacFhTeK8eymuoxaqS6Omb8
BCIY+gAg+Sn0SfrWLWnoCqSsDmBjlMmaAplygLM1bQ4+4BnrqKVjxYhHwkwnxY29vLK1rMcf/+Jl
1muAXapOZb1cXD0L5NTr4sI135rSCpasY0UN/U84TtOsMl/1CQ0UsJt7vO1VhNSh5Qrmz+9H1+mq
y7DCKHMDBixsts+t1H6CLN+DRABPhH5tQGkmhCY9hD3gElsnsBRm0F7DAL2EpGVBSupn4OXWQymf
hzugtGmWce1+QLDDWAZNSP8WIzDwUvk5wf6dwS5GBFGkW1ipmJjwA/ckxJjD6lV4yUs4j24/Xush
mSYPgr09MBuQ80ff+7gGOglUeCo3Vw6UP/a9Tub0Z3Xjb2UnJAkCbwogvQ9zb4Yxke4buve3o3IR
200Fx8uGhZn6LsC0HXYwLhe1vH77nX2hf2BFLQeZbu2wWgvjxvS8w8Ob3MCKS2ZC0Eql92raPeQk
tgcbAyeGt1JPmzR4k7iZvp103kS/cIOibB1ZRQCoqWwR98Q5z5pgzbabGXh8coVWW1fI93kHeV3D
DpCqFa/eEl7Xl1kjwwtjwhkoBYOrHkhMCFh3mOpSZPC2sv06nX8gNnhWa1qwWOxAeEteJu/N1Ogn
fqKwsawlMXzbxLufyw1hLHcpkVsYM3qWhr1yvqcQFAuYHI1NH7UKUN1vtiKcEsKbx6Qul5+6Jw8S
aiPKhTnC7baVb7nwUiZPILK/vzT32w66JOpzY2KBXxHBswzsq8VrbuLFBfDI2H9PFbSkid6PID06
5HTT80FPfsZcAkjm6YMmnugAOn1/H65j4dUfKnuvWJ41/38ZsdsP1Dp/40oMaNAdTePFwAl5zzCB
t0IE3QIlCCDN5hOPm1Ew5jhRxQ926+B8rP/Ncj545ZlETE9gRqsYtWEuZHMgLn6TG7aY6DIZmKOu
az0vqXj9zPjinL+wDizOHgH1wxGXSRMQ+8HYSoJ6CRtxVdQpvHCmKFUuoLJCm01MzuF07P1DpU/u
j4O/ahJZdmliOYdlU8zrO31UxhG17LJPqqdQ5bUa2rYe1h6FOs1LMwycBCQPQRzKaRxMPA5XUjnb
c4HXywVyMTmDh1aZ2xsU6epu4qkRPCdSzUf1P/86R0pb3/kRdfkRnPd6mMPqOb4TJW/0W2l6+B8Z
G8IVaUHy1BOUBJKf8uDJLmX29vi8vO4U6rC/r8FwvBX0gZCOoCbpaTHluQB3/VXMPgXVfT0p4h3T
a+W28R0OmMY9qjnxZCGy93GtV3p7PRQUtv4RpHe1c1bhuKI9RmQZcFpwXFdsOTZC1jJnyw1RpJvf
B5UyLTcKQ5OsoeE0/HUCKCjqEyuzK9D0Lfs3dpOw7VXt3aYpUyP5uWzjuEGZ2e5oTK9qrUBpTqVv
JCq1gvKf1yuLpjUX/dnzp4Et/N8rSx/r4sS2ZYFECaZgoaQfyH+URWp1mK0CDaq0fUW39D3H8IZD
CTCpdGhlk9dFZ6ObwSxFtvBN2ZdraEMPwTEw1r2IB4MQxKZpOlnOm3eHEf3RRPhVzz4WLcNzFYuK
TT0w3SFDFEI3JQ4yziUrfg4z0EMbGRqlF1IZFLxG09gSEoS9s2JpmdtVOM0lGsG3tyFcEOIFnBO6
eV0m54iHfONKZu+675Va4HtvUs0sidPS2h0/TLneH8vpk+ldGHO3/+8ObM+yelA/nGmL8PucpAyM
bnqV7nR9C+ayWD3UDxeEX/ckHv/f+Te5mXO8j9nCCN/SXYGBHk/w0/rirTrdGxKgbuYBPzUoVXMr
KxR+ZU/5uIDmfWEGb3DY0rJ0KoveqP+kmrqXjGKo1UrI0k9hR7Etn5cPkLZWtQZefJF0BhYr+vT1
DlJgphik2FHhLkGKoY1ADa4Bgid+45PpYs+sSMeKPKC5h9f6pwA973dKAuE5cytKY9YIHZF8SmeF
P/FV02PRwliYjPv/X1KdZRYPPcrzxehy8fqut9EVInRgsENJvxh1Xwg7BKordcQtAUBPG9h3ru2X
HSW/wiZmo5ZRihToAQOfGHFZ7BpXs6wW/6WRfoXe1dX+dMiugfRqrRTO1uUPu9MNbidknSZP7e4y
7mMVwBWQ5hTThti5IfWvlTRPswCtWo1YEhGt0HXxqcAGAhZMFoRS/5k7j8AAZPsJlO1Tu9WDoD/0
BuMYxHZMOO11SUhPQMKOuBstAl+q8h/LLu9zuPWew2Q/BS76p4Dv1RhtcAo19T5QDmtyx0qfxemX
vRxEM6PVBLbelaCWc0DfCKiKHdzLOmwEHLF/Ck/phw1NMV6McCp5QfzCV9bhJ0qvR2xh9Ucl1bGK
Su5qVkDXkCfoT/VsozWNyevC+seuejVEHDEDF7rS4NSoU1kEiO0upUkyts2KUatwF4VR1tkPQAFn
5OmAAlMNpBC0BdXvGaL/s825VVKiWf1utpxaN5BWmHl1IEQXSj8lSzQNhwBQRwywHbwnuRBwYT3I
IPWdxqXH8VVIJn6pocCiN+/aZbw7NPvBz0S+IqTt6T7aC67P1XMutYLmzluALllkuKwqMfJFnrzg
CUhdiCESmNL+QkQMEf4mUWDQHzwntFppkcvkSUAa+oY+FAHB4UT8q32NsVvPY9XMD7D+8I6R0aYw
imMsUY7dn6v1KzYAf//pNX7KSoubDKgD3/fCCFoIZaLO6aMTjRZRfgC/GDSHxA6Yf/5a+KamuaJn
ckJ/O4Ve3U66hfpkwUntF/amCRRvRY3q82Ot0JK2ony+HgDZc3EuuKDDuZuQHqQlDxEnpw04Hb0h
j25k8ImYIIEJvvO1LFoYnSuQBhYxJn40j/rROA2zh/TJkTM8n0rP66xMEv7m28JYu3Ti3GN4+xqI
exsQBMmMlAiiy7FG8E17gaRQ3rlwAqFyZaFGs3SYyoQgv9mpa5U7z1+OV5DMYrXf2JJNJhXHP9II
dLtRArSrMyGYPk2PAPQaNgzJ59vah/C0A9wrx4fsUkbf2z9fjEvZ8gC4ZOIxn8o5T4xNyD/bKIqg
04LZGSwl8X/u6ICjj3O6cqa2HccXXatEiOHdKQhiS6bTtyyrrsjRjw9yB+QJ9urU4FoKkDwR5YT9
9iyGdH7OXpHD+qvw3dagBx7n6QmR5CHrvb7y8mlmMFrfr/MyXjRg8uJzkK0NtjWa2gZsBChcBGgU
C1vwhvKfiLlwFd+f9Ak6OYv0iU00CBvKawJXWZxaMOcXDeE0x5sZs2hbP5J49plTqXX6i8aW2Zsa
0JwRs624RXJCkgSMpuQkh7RuF7UXdJfkBKv2ep82IqzyPpfgV6zSc/YN7xCLJePp/IejfMkTRlRO
ZtXPHUxTRjl79ufVKGptyRSWXW55fnmdawbY5tJIadeaLR0TyW/bojcffvnAm/NG/pBJB8hzQ7A3
yE9LRmjoiw25QUTqJC02JMGIhnR2meJjxQWTWxlKWvHHXGlbQEQYLj98pYIADEstMtvjW6YwoJcC
WYU2tGPUJtII/YbXVZAB85xGeszSTFIl5ykwI2wPf818hMK6OMf7POSbA9x+zBnGXc45lCFC67fF
zkARkHB7oYo5/CHvYIODIk0zXkvACv6y4TeBVxc+8MlsE95rPgAxE6PPf9SWNjnhhhbsjnm4DPyH
RBNzCcVwAejne7O8cbd1d6JHwoJiFYWfRqN1YNZ7yMn1lG6Vh+njQ+uRToxCS0PVX/pkfHfsm9im
8paCdtkIARBpWTc3kDzndf9VbqM6pwtTb5fp+iy/bYWALwfoRfdlxiUVxJ1LiTOCcUBIRMJmz+ls
sQNK3rxz04AmMozy0/PNSASzYx9wSiMLnTTt5PUB1dIrbiFfgHxU+6U9nPq+xGhKcXiGGrfC+rA2
oKiFVp0v0GXrOvRLuiyQ6G1cwpZa7kHzJaki3ZdlQLhI6eVV6iFwZeKMxuueELZ2oEzV8JMYpZkF
XjapUTyuafF6yKRxFp7K4pdVzRdGiieoradtGAOFLIMZGtycC9EJOxYLNtjyz1fpGhbbaWdg4o6X
uoAwkha8mdIxY4gUL4K/ct0G/07du1OgOmd31ybMr4wMdIOnU2j7v5ghKZIjMsYWrz8dXLE068Kw
p5AN/fHAY4iE37meQ2h/7RToZrEZ1QRc6IrAbx6BG8102NeStqqH1j1XAcGbgfiMqjP2cxEt/Qvu
5+TWXOosidSLzI29CHTzk8ZWCHypCvSDdBOk0rRpKXsnI0WB3+i17oCMF18sxJBOxb6R+9y/mEKh
2FFrXKiN5sAYRrQVUdyXAh22Yu/URyLF8dZYhBhUfxruZIztoOLQV21/rn54Eoj6TSgl1uypqsaI
QTLEFsyIeoWVws0jqTweAGv8RHk5WCChlXKkfYsnYA8S5DHi0vinmfCS50HoCafMuH/VzBrDRDHd
YDU7+aBOnVEV3NYxUD3Si4di4BvuaHThVjn+emJLGCPoxnkvGH5h1VGUdPtzWq1OcrOCzr15Z3ky
GHykFJawGxRrLHRdmAIKr8Aj/NoUJE3fZGL5WLxVD0Hch0CBY6yB7fVAuwgfJ6r+fAeuBiIpzyUE
ZEuxzK+hMDOqGhL/FB3vDUHqea6wTiHh+pTMOIuZmu0iYZx9Z++Z9R0e5MST5GISFebLLduhoeFj
cVrTLfjl+DCCa2F4Nv9iXsKv9Q9NPAkdp6NjGQbOp/CB3g7DXmmyu/95MDHYlH0los7c+2NiznLo
IvW8UWecvXNzNEHdWLUdSRC9xXzzM7bXejDC1BgA5JWt1RcqNN01/H3nAsLS8bmxG4DtVwoqZOco
GX16xzjeLCP9MUWrueQEYCP0tro7oEmJ+SIprv+tL2zwALj6FVZbctnnfj2dcRd/JZt+vZeKqhgG
l/ZpB/MxkjHfQ49P/KqzriVBJ9RVOivBgrvz7nrOYsb8hS6H0x1KRgcNYkeLHA3qe3/hJHj97zhF
KhgbJzAyEZ9VknYmzLhhpsimeajdlPhXE1dmAnfbTY2c0bbPG1B9XSaIGwvJqguWoY1XHMb/DnCd
GvaMVN5scj9lN4cUTUn5pcnRKP189AbU2LKsCSncAQPri3NCX2AWrPdEmaFYHEGA83nMBmMcMd9U
6nItBwM2+QOcE5jJz7PYzcyVCXzhmGuQ7CV8TOgWMl4pdd/d+n7vs3Fdwwa1qa8itBAKLypVic68
iItKlaGkq2cYX5Qv9oU+FIjvERTl5JbERoiXR1p3arlck2G2I/+6+vG2buOCD4uyeH60qJ4noEwx
wBOzykzL/P39xv3PfjBmTilvxbM8OzWGjcrJhol/Tq6UaXenwK5M+fdV11gx3CVfZSfTRUUW3jcX
1NgiqizwuUhJejZNDuw7BYMWHAqftlncd4h2hCppGhyKAvIW43etZF751+VY3hI1v1drRXDm+YK8
dmvvrlSMJDAeY/bAnf9UWVVF0m6uCZgkvXUGqggP3RpJKFXKfR2pxn8qk56DcliJRn7Oy7M6+Qpm
YCgleLQwi3u4HvuvmvdRz5bXK51lR/Mk9SfgLYtZXwpav/d44hqsHRsjtzBP4uCwfiIdkNIkA4LV
SPmJ/dE2cBvdqGMSz/2XtSPqE/SVxro/9EeBxM20AWLpM+Rt/iWHE+BTnaOTarvR0NYO95HunL2Q
2/slWjkH6yzOPbnZgLhCEFD2aLOISCBYvIIVzzix3N4cWW+mgbYs9KYjw4DmxIC3gRWeQS5mZZEB
ToVLVkRb+z7QJ3jiaxYtVV2tZ97Eo7dcnl1UT7uXKOB2AfaPTcKeBhl0E/pvMRDBq5RAvfuLubft
DFJramy0sTYNT9bVEDCAtT+xSmF5f0OCf/ZSiH/4AsxZrCIbNMtbMCLCP6Bn8rl1X72SfR7Fi5Bk
YyRsnLcEr2E8iRh+/oPcCoMn4jLjC1qAy4sB5vpUG6mdKtRPt5WUE3jDejc1GFyZ3CP0fs1R0zLj
q2SfqDuZAZY5nqEVfvxFT0DwroY8TGsPWPR/KvyasF/UYQiEgCnBN9TrarLlJSMrxidp2eIVprbj
cfngxFe0vrr1xrQ6bcE6o4w0hCePXhugcpATSdUEywGI/UhzxGNQEaxl8fwO9r35SP80dJauxyyE
ocMfSiljkrwvye1JbuLlt8+2JQCUvR6PQJboHx9NgUuc1Y85RcySjTblE0Ziw1f8ZWx6SH4TZbSc
ApKv52TH18Jue9czZKx2ttZ2qy1PIHCHOcWKu9eLaCg7KhMwXaTdcd62s5fPFOuk839sJ+aIVMe/
0AHEeT+dN8GyIEXsmwdY5dERbqgoSrTMgeMEP0UhGftMM24sULBWMtZrGkRh0y8auesgywiMTcj0
rH6kWw8DzZMm7ZyowWnsvYb91kXrgr4Qr3oBUq4iJeMj+vGHaZzI51hp2fcsBMbBsKkEDKT6kCnA
OxFOPiBTMZ9MYFrehCKRYtTjaSz6w2HEnrhHAn9KsRrFP4ZNryxmkk6Vr3qQ5VQYIUR4l7A5wrzx
9/Pl02Hf5gJJfaiKfB+o6WXb/Cjo3lCaSrChwRUAvV3lMB8zeArHa4DUbf8BqT2+upIZuCh8G00A
7mJ59XZFuOzjJiiv1a6DOVOZPDz1i8E2VqH1ZGzCjjtpgYkQzyjMpXDi2YYjxGM1mW1tzpMzgzAL
6lnYbBwwVpe2M8DevMmik3/aTA2uGgJaiqt2f6MyTYVUxfPqsbhsxd7wEIxJu4IE7y7YF9JKaacP
oL8+cq1Pw0cyOnHHwQ/XEzuDLNHBke1POgB6CZJXgOerG/5b05Pn7/O4nGKc4sVpOiXWcP5qMVtO
y1z25NVOda/FFzDvmzqwvGHGsc9+3FsLtL5+NxaMHeiYz13ClfqeWmvWX4Kc6YM6DkSFYrdVczdp
sORxiCmj+FJT2XsacemPQpeiiPxitaKxomM+pmAfuHl/eOl6CX6W10PPJUoXuvEUHVho4+dX/jSe
px6+gthJK6hnygwSaXZRpzC/6ZVjqLKd2MVv7m5oeRdXy+Ylf56+wekUg5xmOksPgf5Tla/lTa92
EdNEJgccCunKezUT2VxG6n42dLQ+RggpJAlOoj+ohB6kmPPkV9hwj2EhLlTNCwTrWnrXOf00MQ6W
EKKcnVbfKCz7c5ujMo8RxEVngyNj1O9C74va7NFUM921466+jHAutB9a33ksIu5SGUtBVcvFiUBV
PMaLAtVFqwmdxEcl64rMDEgPnE0vtvi7LRWxf28Vk44TGmzTfvrgeR1K7JXkQZGrCBE9rin9Djja
RNyi+wer7yBsKG4jVndirqSSIzqrBDzLJs25OZB84DPGDs4dCDxc+FgB+PNNwSi+IFP2xQ4XAguS
4P02+ZVnLEcqF2WMYFs3okE1M+eweTJwjLrCdC7MPQ5I2yO8tMdIEz8bqtsJGDcvAAIe1BqmbU4x
CYH3SgteVKF6v00GRPZfGxTRYW0jfupzax7LFdz+4xC03+wuRQFArWwlRu/epI1/70gyFiOc1+yy
3dqJHjed81cU9ag5+58EjA2jQb8IBiHUeudMat/MGIAjSceihnmjG91auzmx78B6ph7CgaozyYIF
H/Lkpc54HI9nQtpnUacVFs5ttCj82lgAVB83G9MzaTe7FnMP/3DGTkpHG/I5Xu/oZ6FsrIAFj/BM
bWJU0sC/lpR5WWan5NCYN7KoLs48izKYArlHa+i+wIiAwrRVP8lRpAOQlonQPNuxAsTLQ2iRLvZC
WoueWXv/kwW2TsAZ8+YKtt/NRR2L6jzA9r96OUoZOLRqQm06JOxnYld8+X71HBRlXH6uW4pX+qhU
YAPuN433FH8IIZd8RlZHjEJ0iSVMMKWE3UD7Y43QHOuiZcuv7gm8dzJwdX3Aen7ZTNVNfzeAd9Cc
/TrPa15Wwz+cItXa2lBpXbTT2DJrlaJdCaEZtEp/qQWrXLhNeMNm6zvmN4sZgcLObnIwrUX6mqme
6rbwMg+PLzCLEGtYzuVb3EaRMo6/DvdwfNHZwCIrcquXkmdiUCYdcbSqOlJ7sa1viVCnIsGxded3
yNKvzUCopGv+MHkqBjoyN87Vz4gSEyB/wsblpWsW1rQRpbsbd2DK5+iMkHEkklLdRiWIm0c0aUHN
4t7XrzoNx0rhZMYaEihD5qQHZVm1LgLeDelGKn5YaL9PGQgZnyYnT3R5URtNXeTtsqytAKMihwG+
ffz8WdciYlVUDYvwYAtRqH7BBzdprTyveWwEiwggOv3wWFUtzD/cEqsVrHbQFoWkarCXpCJSP1cS
6xdJKT6fMz29o4mHIsBRH27xez4K2pci6HfpdsqV8oYNBouDGuNW7Wv1G/2VSQT+HKLYj8SSsX1u
2IuhjXubwAM9GBhfyB436Gn5j/hNTi/2YVc7eJBUiuRVKieJhTM+oqCo7a1iFCsQANaedP8M714c
YxUzGgkoNzmrKszmqO/3b5pLL+azMOh+qTLBPY0KVT/1lMz2wkQE+9By7fYmSDEQ2+jdDtXWvxDg
Re5j1LpruXoOLRcalq0Hiik0vhyxa0lRb+rDO7JXAUf1OM1bHRV4RITLH8gFzbfIkm0wjm3/KTCm
UH+22r/GrJAYJjtwfoxBVp+JBVD4vJM8FQ869YlroX3K61ON65j7/7lX41z72JQbabaipWsC1BhU
lyfC8wfzqm9Vs6eUuKpU98brCRVALRxiYYYsKiUAfUKKONx3lS9WuF4pd94GzwEVwv/Oaf9GaUMg
nArbLXYh4RuCdLnhVuHL8+PAv4RV3YgIVo1rS6VpWDARGEdzHUc5CzZUC8f7pNt+OrU/LO32NswH
n3Xl31WkWsexYgbt2G7u3JkmLRly7VOYP/tmKHZ/X0O8ZaYRl4KzjdDYhR7lTSEK37DFaD2120oa
AqRUouuu7NzjU7znCmOM6QbN8OxWmsakVB21QX1E9ZXUHGcMj5xM4ueVfPh81HmB7FVpbTsTI9uu
I75ksRyUrCJZxPNkXK1DRLnVxwp5P65qwx2HsVPKKTkOLN+LrwUuqwvEzoF+mwkq55MOsdilSiVs
yrpJa/rUt1VCIOVlqpuSZElYnEIB8IjLPHLtxnN02SPqMsP+CTBCQ29g7U4hx9xyL0uEZhYumwwB
i7eNsZF4tyAT+Fei0MGAa08PCJ1bx+9ZA6jQCvWXQ5Y9w8rI7l3GDowkE02d4maEeK1jtQlfRCzT
o8PkWhp31qgqz4Xo2qcdDMiGRTme8eURHBsgCj3dvfMk9lyOATnbpqPiXU7dQCT2kZVfgDyN6iKG
Vn5REuxOEDojPjXjofj7DXBiXqXVNvaOGX5rTkpGAsu8QnBZvLy5TDj9ttG+qxcRNezydWNIk96F
O1xfRLwUCZJU8XcOZANpirWiReiZrwmgTldNKvPA+cP0XHLPL/TIfjuugq3q7G5jzovDSbZMDRPa
E+MIhmvZ/HezWd7DmRjm8gQ2vUH5tpZvoGprHJqI9i9eBM/1MajeqO6rrpoR5m+gvuPKl8GwIZih
blsnNV6QbE3v+zZke75iVydmZetjpPEq7R9+6jhQevNbktnEnu7X2YbsPWipFssl5V7YO+Azynym
jAw6z8DC3TCqbBDGw3hJt0aKbVWqClFGaCM0HSoeWj8HbIrtBnumm4QuCE/juej4xGtckV4FAhkE
bCsQYHYpIZvO9LoeUefbF/eFu5IN051KBgCKpluaALLLzEpVkBa5bBtgBOffefalw3OfYyKxK9X/
qGoFyKiQ+V3glZxAE5jC6GTQ3+5zFfcTUq1No0eRc8ubyu/rA83FfzqMBmF0aWULHYwda+mLsHW0
gI+0kYoTfvivZOP+Hgg2oMSzuC8XfScHuZDqaTmaRaQGP82eQba0ysmLv1xDY9wIDYNG9OkFaEit
o4hxcR8bjQrwglTfXpAR4CVbN56yuXLa/ucFO2bHW8FUMTGzGZzosXO4Bf0rH/H6EgPb/YZlduQt
YeHwO6befvowXkEY/5svKBJMejc7i7g6wwZnDcP/heawtWCoVBsTXldeVWB4m4/R9Lri2N8/BZT5
sLiy5um/7EDSk27kcZ+F5d70vucByoCxeJwwHgJRMI2q8M8J5sicgCagfXicQDWgEtPDyRTUCayT
a5Z4jpaVTjJSIaLl1NfBFlacT7laKrvbxddQX+Adfb4LPFjQAPwYjTO4NfuYApP2nLflL17AuzRS
PlbyNvM7mSEmWX4//0l/pUxn0BffPGkAwUyGtry9l/HDRQolQkcCRoiiVIRh6dkjCjiU+ixUER2i
Mquk0Rm7mDjNJlDJbfS+4Ee9Gi/AIJnD02+sZ//n2G7JorUZJGjSwtJm7/5d2WaqpRpNbs3pJ70R
jNkbtbWXwswpAjKKRtql/JEcqAE/EY79IpwalyuWgE4OiqZuQl0vtf+tKz2w0sRKjqvrrn9WNn7Z
29Nf+9Dyh3EVgtNHmUln13DovUU4wEUC1YVt3ARREX3N91jLatDWLCVe9H7Do5WmQEXpsBKEnhO5
mnFaWC8LOfNln+aMGGY7n4t6gkZRHOEZ5L7DZMbdZ8/mQl0fzzIi6LmkjomxBF05hQQQDjyNkqrS
0jzWNZXGOBLVA7/+1DxDm/baRe9UI0BH2xtpz/25hc0i0KR/v18RliYEsVsYZZKdpGZvAXa5tMTf
6oN1uwRJ3Iu/OMeBO6+H7ne7p3bKbptAHANNVjJrYwUtiVtyfrgfGJipiN+w1w1fgiEjww6PF0D5
GlT+WzoA/oBJUx8lgREI7/ioTd41GiynJAGeA7G1sUW1x1lgpdERvr6Frqrof2kSYIxjKfUqG0RL
yd+mcfPAh9EwH5ie03+Z64bVRp7+u0FBsPR95Dv2XzUOi2eUakaDJVh5oNHuKTVfBWJiU0Wb0BPZ
xMIMjyQ36Mp3YYmCU4o+RNJJvGsikK1xxa0jAMiOpCzTRtp78c+rVzEfC3izkpCREdr9iKhqeTMn
gmHSfqIQir+NwksmxOwV9k9mXwVefLrVfN/YBlZWZ3GLrBYu+FNdcnfVV4mRWFchkux/BT/4EPeX
dDQ0NpSOjN7BQrSKXpLQK2QK+WeU1BScv6dCV9MdgUXFVJwNF47a4By8ae9yXe511K7ynP+h0P7N
INoSgpmj8LbusJ/xuZmj/kRMkS59hOKRG5TJ/5nKoNdAOPnDThFeg1Ofy6BixF8VLQIdWBIUnINq
tZLaIvuIdR71fFf/WZvl3cTIgFQLhmV0iGWbdA0eHJ77Ul8iJVcIvjOtNkTh+ifkh0kDPMygQZ8o
quu5GSffHkEQEaS8kEtCrizE9mGqMlyDi0Xh4wc/a6Tuj7cGcKY57XkQaozCa2g9AnAbYRihojZj
jlHk6gs9oDcB1zZvrmBiujXMy7+3YS3cM5EiPcRcH3YpRTlAJfhtXqpmVC/yDe5S/VLjma9cbVor
zxVCfPWpNUbf0xKK2sNuM0QL32p4ao+L3BEFOsLq+kNDWr2g6ciSgRvAAVH8sjGWw/c+3dZ6aklH
vUxTQ2m0kupkeIXd8V34xFgK2B1XJZI8A9yRHip8omNGtirLlytjHIZhZKdNi0oumTGOsKkEP4zY
biJ7kA58TyY7cznLYrecoeBPwBv1lESayTiEMm5yihjxdcI1nFL5kSc5Wrfg8Noxjg7X9aRJ7plr
z+XS737cXfLPFMU1d3cYfY2OmToFePCeL7L3Uf/GTRzY0Lxpm+uEu9/T4jZv/xwnuH3xxpYb8oZS
nZoMphhH7u59YcGoMWIB7dtWFUmjgRF/IqUqBVTZ1X6lB+L+Wlc5oI1F/RCsasR5vYm/QXVxX+zo
CfbUBdwhM6KpovLN8uBBRyBlpqSvBoJCtsZd6PC1u2GkQt1CHxkwpBiq+Kvcng5IDXmovBe6POlT
HAvT5OwwUVSnBzXhgxjVxa+STKTDLSsv7NtNvVF/18u47fdk50UhscQDRAMD5xTYZDtFEIfeqgwj
e6ykfDfYKMKFqbHQd7J226tpyP8mmG/sCDoWYNXCNIe520z6HJJzhVTWi7QgtsbzcG0POarPhEMK
fafyvLvYoFr3cQpBrZ0Lswj2PbzBO2nr+Rna+Onr8mlrk8MVqdjwZg2jZwOcrvDMu91XB399HkuT
eFyeavg/v+SNypiHCpSNu+iAqNPJMPmHOMbs60KuCKfibyUeCgxThaF8/7cxz9RSCqW/6gtBm8Ph
1xnU8JAwUpdb/6YmdtBk99590patq2PpAMVzmmJF5ZB6yatD31sg0StU9hUaTWNXkI9eYv3RLSWT
eS7jbRM1utTOpEBFngFiSS9OT1Nhs6erNj7pPuVRBDexZ1g1SirYlOeK3bHsMvYaoao/bcvG/5MZ
sYNx5m/8vj/aVb8zXr8c4+fWpm49yE3/C1bKTqGBqNPhBcR9HVn8KHB5wh7sCzf1rdEkBcmQh75h
3bCvopZRMwLJVF9T5amqRu8Gmdtj3nSNkd1LR66DzRoZxBdBb7dvizWMhg7/DRNub1QkVtzBkgXn
c4D0ezoQWpO9qUkzvIqdywr2HXYWkCJ9/1TQT2XDR1QV1N8t1cGJDoylNeOCiISfxPdn/T/ixCXo
5sMar/E31CJJ7FT11PgZjKfZ7FQo3Bm/dRDnU6MsulaKPB53gTiYDq7+BzAwIJET66ELUAXRt54h
hju1NEJNgVzZ86bHu4XSQdisBLg68/T5gglK7EwuqnFBwRDAZ5sgPMd4oACQZMNx30+hryzixlzf
ZXC/+c/cdJRFSmX+K3YuRGXnS/RDBUjspQ2Fojh1HM8R5SrPZ+JoX+Zad2Ouhwor/jHAa8zyn32G
ahn09i7oswuVvZkNVby576agJKJrbMrGoUMoAbn60jvf/mq3H0ijdhnkiDnUWykf62hOFUmt97Yy
ZyGnM6ybPByXLlQr5qYO2h9eA2SBu9v1T6XqGFHHJTadP0ScdFYYfmBq95T5JmM5mmO1acs6e/3p
i8PGitCoVRFYnlnVWLBZrgrjJRwu9NSrBg8OmxXBTBWyLkD1R3HTx7vq2Xxp1t6wapy9xJk0qaD2
c7z+Kzt2VxOFaJwPmdVgcu84og7eOScuAajw1BOnitMIt07Rz5Az+9Cx3SuSzRjByGpRuahDaOcX
4rC3Sn5fGHOkq4aQsy5ueuHdg3BODVDJzJHWkRjAsb0Tex8DmuoWE7dnTcX9omL17C8+zDs6I0mV
B4/aWathxVcrKlD3YQmYa4ks5R8x/PrWM6bV7XrkfuUcJp6nd7vzT17//mdRNT7r5iFO8D3+pE5k
a4IfcXbJtzmFn+g1n/tkqyTW77BgP1I7A2kFjm+5/A+hHa1zdp3diV9jNdZR10LeYsac0WOqW0xg
y2FJ6qsy7a1yhhXBk/yaXyksSbAeoNc1I2e5HxjBXg6Tl8epeXv4juXBTp9OCTM2XEGKcs38A9R6
QOXRJqMruBeayzLe1JfMqtUWdosA2ypCM+UGK4wFVAoqmspiMIwVSkiMpPF0ZDod+W8ZBHMAOo2+
yngDxlHrAgPC+SZz85PdlzGqZG/fdNP7dHX9DpH82BSjmLLXM4kk6FohJuGTqNajwHyEIGP9hM4P
nJeGzBvaKlmvWAN8N1HPl/k4lbYTQ3WMKe/C59uJItUZa7HrUIxTxB0UDKebkVdX4oIePBmaSl4t
DxVvW8p9NEtGBNSj9KWA27TOVYpADaTPj8wKzbLMBdpEjEIbu/XfVajTt2S+7EVjwVSqcze3Liyq
P4yR4paqKGf+pkUKbeOSiEPE8qT7WA2kVuVk+AxV8q++qVlhO8iCj8Cu2nDaJ851V7FSTrPRuCAo
mx1pElVOyudA3O4L2a2akaqlBsjLZjA19Fg4cPSg+f3lphai2lJJ8NfyDiqLMZ+hJJU88yVkRvQv
FmmZnFK5FP+iF0GMMKSnGYLso9mVX6davyJQYI2JnR/d+NAQn+qV7wNsW/a9wqiDJw6BI27hhBVK
uPXZctsVsFXN+I7aal+4NFKsjn/cNQzioKpnuAbMiXtO/zkM6V81IMAbxDHfoOrdpGkRnX8z+wPN
bWXNV/5LLwX/ZXa3e7vhPahd00u7ppdlPl4cJ4Ccel+yeqMFY21A6hkXI9DO096ZiTFmJ3Shiyuk
ccJ15X0rvAE3TlE8OcGFKAPPd8H/fT3bJAfraNXi8vCs7Pqj6tUeyrVhkWzyE9nALyympb6akjIa
mw+vatq1AXSY3v2aMm5JxDNwD8FV8FMu6qE7uCLp7edf0yQeL2wu5NWJeRQdkuzsIYdRpjSbfSK7
Q18o9tmksmMB2tELbSf4iMZp1XVT9r7awY2RK3O3buuFjCjiE1HZJwoRZXUEbLL/lGRkmTnRKwGu
nmqqOwc1RF/9bxFuP+oTrgLl25DMQW7fqYImfyaYkzh9xRSa71pGJSZrl4lQre2C9ZpKTtqQh9Vo
pkB5xUgCy0TXjuToaaTy0ikbdgkBaTpP3/dyBDh4267+IHQmnKMY/zyuWkRd2dfKBHCE1FQ8nf0a
d2BkH8Ei+PyIg3KDmCX8ANj9PCHdmbHMUvf8xNvTD7E7P7hva2Tf0wibdRupsM16+PrznjPcqLdE
u7oL/TeBTNhKYSC3Tt7cKWkTgKyPVA732RbfHXbJ7TsEHsoTwxqSXQIZCYfc81M27bn8PGwizzWq
s5eBaTpaPnN67HIg+btWCGvDihWumNQbfj9LJkJwsFS5Oc/w0tHAzHYW7Y44Sx0yjzHV3HoeNpVF
jUqoM7y5h4O+M+05VW0hECtGrybFPiMAYsB0PcVBPnxANRAnTNAv35tvZODlyvgOBpWpMTYwEf1S
IcpAHJ31VziuV4Kx9VGoAisyRHPpTk/1BaoV/wNPNRpyYNhkOe+sUHaMUQV9n92P8W/Aj9RgMMYR
e/AGhGAufehw18i898ZlRaWPIU7PMwkp5WWwnyFs4y3Vv2y/CVU+uVm302nSjaCv/VZuwrC235o2
IozxfZu7y+x1ClKBBcukQV/5NmJuLY3DNwUDDlVfekRQ8fCHtLQTWuibJBG4HMYxFjM3aPn+Lbi+
0LOyJDgwLJEDiKovM9PSyTcjt1b/YdH2IKiDaA5eGc/kctSW0S9THsA1QASuQZ/pqfGW0rj4vjho
oK3WhkTCUwwrY7stIobu4FAoxR8Biygm70al1+C4A4tDzGwkMog6vlEmQKmne+6hIM2HkZAxfXTT
ajOklz9Ys9dIQmti7wndySoZZ0adOo/U1YkyEuKihVpTH0kHaL0MvnQxfVJ/Y3gGxulzFpb0clOK
98U8mlW5a6dWMl1vEdCIVj43WeSg/NYg69qAttacsxp/tSJ0xChArI+9fTsP82WDHnqgI6SxuiJh
HjzQcneedq9+5a3bVKknPopcVZ1qZsTK0r/6uLfrcu3LdT7jV69eDZj3DCCi9ZhJtRNr9X2q7isP
3ETwi7gl617BajAwaPRB/uBziZUpGq5Kdj3FKx+Uq+tewCY0KRe0URBiw/rZRf+keh2wZSBcCHoW
gZdwUoYavRP8yaYqqy+XdMnUpT47gvL+qyuj/254k9rFaFH2BJrjU2whIuqV+vUqed/UWTM24nD6
XJXc9hr3OSJuNf77Ku0OosilsoEOIfu62eZzuoxBzqPxhquodyJEZYZTKr2NYR5PVoEfc+afon9v
seuzSG0Zcveb25SWjWfDGwi9nvRPPMqjLe+L1cEW2gbYTsx9hl9se+Vj1/UzhNIPXYTNU5dfEQuE
tpqSn3FXB4yQpYnWGp7lAYr9Vubr1keFkTQt5f2Gr/D4GZ3WRKzGf3drsxVhFRw7H2S+zYzjjS91
1yD17ZXe4zDiKIqcQDPSg9AV5bJud5udvGD4f5Htsx6KwXWpOUCJPit4Om5TIR3Mmqp38y3wSawz
t+A/LHvAFXCrpA5Jm75SsLG/6U5yTgStNvvswshJ7UaIzF3H4oDCO9SqYTHe/XF8IV6t7fY/ZH3W
m+iif7ecS2BHz7g6TVy/6YHkmdCl04OzKxEaqUeDzC32qled/3mHDFCfhEqyBv4TCpEMyit1R6/F
p1tVZVDRhEeoz8eQMj7WS3BfpXRbS7igCrzEEAflG3ewQeWx9pcoLmCRIWRsyj8M4dzYzshcTRtl
X1wJ3TvKUciXzmkKHazVo/Ts/xCyxUkEknc8rzB84+m3ft6RIUxmkCkuM7kKdKES8tWB+LbrQGlE
heQyybIa85uCSQ3s0ix94zKnThMBP4sS3N3DTx7mFhhxeBOS083jExWCz3a6MHaqgGUnQ+pPaoD+
XY1AoOgNKBYaS8QoT2wHF8cAN+MFs+hTvyCukQzD7ftqGZzRx4Tpr7P6PQDMPQPrzxm1hbvWWbhA
7+1b3S95QuGcqYPtrfFj6Nb8qq3lybPtFCVLtm3PgNbKINPf0b62NrSA4TwdKdbBr533o9PdXJen
EDN9xHDzk1M+BpTUqQF39VxK2PPBFYK3CdqELD8nEJn8AyXbKuNtEkjH8L3/4OYoNbcR0AT3I7RE
IZc0G3mGFTRRQvAy97Opa7yXOFitOiu5/bkEGndQqjiAdx+GWDkWKfqMc/FxJMDugo39J8QiHZ8x
5uTb/IZ6RsmARSFqbPzok5ehsVtre9TEkIAJeUMdEOkSEcLEJV+tTy3j0bFVG1gauoYuSmUxldX+
9JJmKWShfxv3dRaUyMm9r2kjz/Lq5kjD+jrgmxdVaXPHbjXnOoSL+Y7fTqf1/g2habdlVmO0QAtr
1xm2/K8Frw+6on1ZPCMZKzK1SKKJWDbaQaNXDskWGDvnP9Kq2nvSmlqDourLJz1BTRwyOstzcNWB
14y41DQ/7wBznjk5dfMVDnIB16LHtdJltzo+O+GQcnbYv4VUzcXRm8GaYY/DAdklGmeSqPWcbDUB
rTL9hfNjUvYUwyBBm6a4Zy9lXbmPUPNT9jzKXxN8+ysxPPjWMtsrNSpCFHVbSn2IsClaho01lb17
dfXMQscvEhNzyEPmF5fizPWCdI3gGkxvJ/AcHgnfiSh1bxgKw0alZIC0bNwFpf40xG08ZPBr+anV
WYgLhgdyghtyslNDlVZCSopGtjitwoFmXsQ0wdFAhRfPbqGe//5Y+rRyffSJR50uylRwSL+z+BC8
5OxnBs4/zT5uJAPsQyW2z06yd1bEKLoJj30biWDWgtCWnKZQqBczwqvXmP0Uzvb6KyqXVWuve0Iv
VeuMIhrah8lnt+807GmYOwrBh3fn7xYBvb9JqOD7jUSIxh+2f50D41E9WNPt4a/m+STiKs/Bq/xU
6Os2VGtpyrFO8NhMwKOzycOm+hh0vdTelsmkTXviVeiSGqDCy22Xr0+1dbxQ6KdWO5t+c5Z2Tuvq
y3CSvE5H9xzSPCi8StAtcCps0/8H9ujZXZRLvlxDo8USdez8TCu/nVCrFuVx+VA4E3qsFcqtY3db
5pqJZLpNOqITwvE80VHYhGMKuo+Z4DBH+Z94K6TyFJWYT2SSYvv5ltXLuqIgn+CNiDLQ1bZ0fln5
jKosnJFSRAe8g69EtsyHxx2aOPxvZWimHkqu7CLTShYk5cQb45poruW2I/29UuAtg1pN4ehOwxXp
AwYEQGM1l1DcWxR6gHSQvC7r0MX8NFzRvhhG9+vwD+N5UyDBf2Fpjyofy5zBpQJ+M3dxRxjQcYIb
sxIK1nuX7c7tbL6+GYcdxw3B3wh6sUlRk0+vffQmM9A/lwHx1KxTMqR/KQplvJZnr37mZ83hM9o6
kUv1OeHo+Rs5OABp9Sq+KpKkLvKEpDmuQ+/RRfvBAwxHdCsHdcDKdYgPgJ78j8he/o+YrPPQ8sE0
eoI4FlSvoZVa/R1uCsgT6+etTTuKJlQF2KLFo1926lPVGfrFb11O/RJTBAY5+9OEwGvYQq1osYun
nSFxxGZ2S7o/LGpJVaRs/BCo8D37LPouQJ+znNqYP6DwEBKtKeOwKuXCHLaovgEkv/vwkUS/UQda
Gv7ARbLxoBYkKTeXU/p9brcWXSMO6L2UdphyHmfgtYkUL129kHkxJuULZyybd0yvvo3zN4d5VMkK
8wEXJPQ8mE7h3cieaIAHH6/bE/cS3XQe4iXXakLs8M8bMx1c5GxhHzSqmlxRTlhwiFPE8XwDlFTW
ilhJ6X4mkKA+4m8zjX6O0c/xVPgWuBWaWhVDgawVpyK92insmUtStZyTJdJRgca19Vs+vUmvGLvo
fX2XT/nV5p9m0JD043c6gcNnEfdTgwrRLKjqdysoRMaR24NV1kgVpddeIjZ9NkbJhRn72/qzQD/K
5pN/syCXleNId4KOYbQ6F8on2+TL9xEgGb8vnSxJFJeDVwUJ8iXv6C3nBOnFVVRWgAKgSdtQqOSG
c10mELvizxkjfh+n2xHH9wIHaNn9gZnK90RwWagri81g8Srjr13cIlC8Bm5iIK0Q5woqZs1+tTdu
3bFE7rBr12X74YL4et5ueCcGzWoMOgkCAow39xx7SCrWdHYNVjEdrbbRIpn97vvgcEnTdwZsnR32
2PW48PlMLFCydsyBt2Xq5CssP90W8eCVMMA58UG2/Wl70uESev1Ytyk7ce85uzS24RzP6KBhklqS
4my0IFGd1U0YmxxEREtcnst2xuB54yb7I8VYvC+1vlWFugnHHI7UV36b44V0fwNSkjoQo9yDwRU6
ggiO/BtDkvwvywiDmTlULf/w4vpqWuydv0mrVJyY0wcrM2UeNZRq6XusmvIb76mJX39xZSmkx5kB
N09bqlCtuypm4+2uOgC88fdNMEftyNLS1lCjbesbnUMG26HcMEMZ7ybHj1MeQOLwZYvUJfH03eBT
aH8qw0Y+3xqawl7W56yNUprX09wDHy+Zlam51QupVSDN5QH98UUINF4kE/mlY5OglJT4cGsLC8e+
FQe1jhcUSm4lvNBdiOMnj6xXnOf/Zehp3XHkJGtndGnFSt5wF4VP4qEEwwnbcAVtmHOdNnZ7/cPn
nJ1KYQJ0vP417aUsQlTYoNPxqkREJwGpCYlPxnpWbt/C27YlxWacvdsEvKrQSExSkfQaN4PzkoBl
eJ33qzjjRmLAM0SlUhHTsQ7s5DgtyyAX91pcSLnRB+CSya0jxC+dUoId2n/2HvxRVSHEdqDRFWz/
zsoya2vZjtPYk5bYsws/wGnH689U/C/tODWV63lQn+tDyFcKgwm9FZi9rh1jLaTdo32vHDB8AGfu
nVgLM+obtPU/KlPBZgiGTYdT0czUCLnoiD27RJpOi8EObd7YiPPSuMluJmt368DDVNRt9P4QnzCh
7Gw2ZuJr+7K7QwHsgFoLZqhQ8IFOSr9JLeGwme5syc2GXRYnzgVFlFDBLOtatTg4Mx6E1XY8IW4I
TGalwKzGaRYV7y1QnQqV5TVClLkeihcRFgPtHfJWYc15ZnebrUg3xuAubwy1GCR+Vg7JkeEdr3X3
i8AopyB+a4df0iIIvQuI4Wgzn8GMBMyOi1OMI9KL7onlqfHcr6EKGEYgXDsgNRDu3B+sJu/b9l67
DRNJmPX5hJZpRDz67EQGRv40MmJj83HytM/LKcDyRBQgQctjavJrNj7/lvqngB1Rnmer35x3S0Cd
hK3XaffXgGxs3VHTNjdL7gAh3YNJOMERyijTHkWQ5zlsspGyqa9Wk0vf0uh1NUoZWU8ed0ZGoM4x
knQC7yAbcHMzzDcsiaRacuiXg7VopL/mhHyupYmv8D5d53nmcTTTDCZxSUJEBA0Fp6txZJBZneZ+
9nq0cj+Mn0ZcIbocfW3dF78w+w0lfnP4T5SIAUMOwSGg1bhlOVuoNLyXfPBAXJRtaNKXQFjHiW05
JLsfHGJhWsckAlXIME6iR//fAbdIm8zDpUQKvTTJMpbtkRavPJGXOdIlsv5pPiqX0HuvAC1Fg2nE
zYo0WkCmBfa/C9wdcQ9HfFu6iagwQz3IBmtXRae3xdz2BCjw2+P/aVzuMLyNmeX1cIsMkaqHLdzs
kxwbjXGOFKFpE0R3btdMTafmXJjSrQ5B5DevrYowsoPAexENsspCHrz60LcVJqXUu0BWz1l8z0Z3
8GZ0/cZRUS9SMR6UfYu08Hn4uulW9euHKnV1+9n7MRP1+przC2/AQHzQI8EOL5Rkr23bdNwxS7H+
rKwsyBmZmeF0D8DqfHeuOhM87dL8ccAs01A4DkUIyvNvyQIPBo55f/7QKOwD4zgb+pMeRHzUgodY
aja5KlsZ2Yq+5YHZN4GWd0o8DNfFDxVckChD0mk36uZ4c7JC+dsQxPvhqbY9m79ZKoMPy2LIaqSi
XQvEQ/Fi3aj0AIGo/wqdjUMM6Bc4daFTOF/HPxSjU/Qgi+0U+C2iEBWKM5DrX8bgCbNnmav4wgTO
M58x7RdpPseI1FvtumqpogxJBGiopmMfs/jRRgN6s0mkWBS2CBRRUQVDVvQWudbp0Xp4giobBgnG
nqEJVMiRIm2tTmnuMphGhfuitHgOCYsj3mj+S71lVlGQEzzfzL0ZFDHqnkJZXCcRkPniCQAhsfQe
HZCbHjy0vvH2RxQai6wo6gNpwC1uLeQTiSFYj+p+9xUlKVqnR2RBE2Nc/bBKOT7rmzOeGj4mr4cB
2Wk/wXnaStXYmQviCjJXMbWM9scnBEEq5fI0hVIAC9QBjgsA7LEB+8t0ChUTVVuV4gJtt8tvl0WC
Il1QbbdDgN1kulzFPIPuXyx3zgMFMRszNe8ToOsbp1OmiLweSmSg+S8iK0yLxJl8+jnFqxPUvFyT
cfgbmcTH1G3VjZYlq0RcAxg9ZbqCsGhu/JHvdKmljv6Jxr6BzEucJvwTinoGjIzeBpdBIjw6tSwy
cnCFMP1i9Xt0kqoJfVoebxYelIG8xdo/PkreCLWjDokBTz4cb9GVhkL06lKB61TE0SBYNfVR0Qy6
t/95YdQgIyEXxHB8qiXk7uhsy5WmtD27oU1be9F7gwniGClH4OloGSrNGdTjuY8SBGIWHy8RnINr
bQfBEZ7Cs1PWjzmjZx7W2hnHnAZFvt4cQXidIwF3l6nzNo6Uzfdk20gs5MngUs/jhbHJT2HYBDvH
PW5c1NZnrVSfXHs3DTadqm7GI3ZC2RyAyPYJGZOwhl2zlwY3xuS7ko+Aa7ApOus/IJptwzdSsxe/
LD/ckIlxD21B+fBEBFhR2UNUFCEXdlMFlTfeCsouhMrNX+78TE1tBQqtJd6p9L7ZF9F1JOh76e6F
ga+0ycHj51/4E0ic8sjUYYdzMIvSW+DR64dFfnj5R61F9/d1fM8Haig3/N2sau5PPwKVnvmpoL0i
5pWAIF4zrZaiiC0cNQwYCdavxM9XipgYJwyQpAPlZ2aWWeOCnTmy3PSPcG2tLAapbS4noS0ZPRK7
zCSErwgoYsntYwxS8UWnyOFB5wTigh4aWDMvpEhlb6umWGaDlg9i4AZ9dAlDz056sTVMa4Xw7BmJ
NEDYEvhGxlOaXrKzRD0NwEBlsFn9m9Vmb5dp+gk7egSKli7A3+tAOAJmzyMa6eD5B7kXRuDK5c8n
f9pEm0YF2yyirT1kUFNyDfJxDD/yHKEitHarYynRW7cgkCLLLR0UBe00LSsLBLoapxwJCmH8xjk6
dPxUiblF26d59LFKV9Pr1OKovvTjuft3ieW0B9ZeCqvwgu1KtMOFJvtCD/5JHt4CzZQBz10yinTh
04/Gg1vrsab5kK5Ic9UquiPfNWwDMIfzZRfMLGXH/eGZLavU2qPXMSTXRxE8ZW/2fCm8xJ+JWyw0
dzx8InqSyqLr6zzk5LYLNEGuYVY2xOfuREoFnTFOdiVhZzlMq47nDui8q8/zZcZ/8F+bMP6nslpZ
8PmQHi7mJ7Y1SZQAB6eT/LqXUwwBk9ExyDfIK5yE2dZ6uv5aaAk4+T6Ntd5+i3JaQX/d2j0p7d9m
wk3a3S+SCKDNt4IilJ9JOLFNgrKbKm6CFo3LEEz4aebPmrhe9djoKTW9rJRwxjgiFwQuBHPCK2wl
DyHslFI7CzF8t9zoA4jxYTKQVfZKK9R3Gz4cYQsYoK9Xdy2bpM0TCb1Fc78ctCRMbI2zDMYh0GIm
O/zTSTuRGJRF7zC5dcAtaEd5FhHaIu5/bMiabEXoXXWEH+/S+S1tWHl/Ndn1WoBoefhv3W0mZgWM
/y9loVDHBZirUOOBwQ40z8A8ElqUTp+C/zLF9LP4dB3iz226LE3Ze19WHBnXHlTqSkL1tklkmyoh
mzDvjvGagryQUNJfCP9987YNiG74csAprSv6wlxbfTBYnmVEALhqCnk/2XNwSbW+I+ib644Y1UJP
apLMF0xA7qXnbX9gG0pThntP1luszWOtnpHjEWXlUzGMq1HSZiX/ADymFJ8jVoxlR/+lnW0vE6yL
WA0nueXUiYxE/lG/pz+QM1vVRZP06p4ov54pOs00DT50UeMku8/j4fxbc3w3z9nRvN2yqOWWN3u5
CjDz8/J3Yt0v6p9+wQXCa8OEqTtkCwDQPOL0RM8NZUykxVh8YgsCTEgoO+YbnUQEtImBY96pNsTh
UqpHBeGLA3PTi+d5Rrhwwqtoywx3YQE2eXISh1rhOyDURoQbLKXwcGlw/WCyNXj6QVWw0owjpCZ3
7gFn+2/QaZIDUK7CuV5VdedfRCPeWGS9KvPZEC8weloJCKVwCLS6kROMHWaFbwY9yZKyebocpdjq
uI550wTEV2ZkfyuGlQm2G1oU+JIiziIBMsJHRfRIZArQVNO6+1sTPAoeQx7kwOSwTbq31jXFE6vU
YMAl/QJhzXqObeEBBavQr2yxYJ/0TYfJPcOC3ym3iwggp+qqM5cxbsYKxZQRGEugcjy25uJAS+IS
XOLXOCDjAMXaSWWh4+KSBGYtTJyf6+Bp4qinTEOxYIiKdnq21Q8xMZ1oHgp+3oC9c2YYp0aSm4L6
0m+PHJ63NFurtmmpOeHHqa6AfMzN6lhaomPu3cAyvk4e7GwJI7P7Nm3IWbqUnrSSsc8biJVJl0qi
3RKHRGcj0oViqk1kr43S1vb8hGjqMakkc0ixf8CZa51n8pAsfJHQ5kVnmBeE4pZo0Vmt8ZbMQJMv
Zzyf/hIbOxi8VY+coONe/nQS88qmRvIEWH/WnyA4hp56qxprPNVS8TJ1+sUXQx0z7KpzifMH0xtx
x0tcv4Ui1zPPnEZn3DuqNI0zhBFatwwnkISkbiGuS8L0Pl9LGnu8hOpnkC/zXBfx7OyyMQxQBnF+
q7AF4Kmx1VgYa6VqYQjWiQQiCWQIuo/njtEQi5W4CN5QnGN2IB7Ima8B59Q5jhwfB+IjdvsdwS5l
WZ1c2VpYeGB/Qq0hvZCxex8kOCRrhX9Vy2qwJb63Psi6QBHsWsiPnNd/y3tIt6OyAN95lXUSPKk6
lSZZkMlDF9OeslYi+raH0j4SSLQlqVglhzNjAim5DxoNjMmSbj1NaQDuJotvX9RsBpz0HhShdHWG
xE3ruOh1Ai+HGa58B4fM06TsRGcWQFWHq1lCdtHmh4IK1MKelJpK3ZcI/PzPi11H3TyBn4IHe/9Z
KI4RHUxshDWP91/HBiiN1Wv7fPQMuHwuct6n6MopgBZSGbCwFrq41UAPde3B3l8D2z5AT8MKFVP9
BvlscE3IuWsWBM6WH2pu0aD65GtE/8Q6fHo06wXisnzswFBAagQ6yBjBW2sOyiXzMzqGjkVJYMIo
wGoZ8TZNAldSCILTFcEIYUvOQv+TWDhsKq1i7nL1bxog/bKgNsw0NTQa6Ii0QHmD8HSKSUE/liym
vnBGnPDZrw6naPzvSTTTouh0R5HJIOXjviBK4swMVdJAGeWjcSV0K4QgIePZ6I2sLXi0zflKa9Kg
+gov8es0ydCrW7HF5KtH4X5uV+KNL6RS9Pzvx1xgc7aTKKOq2d7lcdCqnWiKINQcpUHsKlQYTDO0
+U2FKuKMIrXu8tTDsxVTvLI2izhL6ntoLOA4udq6esze7F4r+deU0TXXcWFEoP0bvSb6khjRxutm
MIyXz0Kefe0UNzyXB6DgVsbPKr4kXY2xwrPvUq6CjBimiAzUFl42ibUqgOFrmSg1ydJ8FyvOKHU0
acQDwv+qdDRszSKC3CaeXa4uxcM8YSuapesuXoB4up1RFO0pZXW5R7+lPty3Guz2nCULCB4nCz68
n1OEAmvNYtES7TCYM6lERUSext5prziCIBjWSD3osbxOOLzrA5mFLs+VrDgQwY2Ms5ODSaDZvr4/
tdVxxgNRoB3c6p5nFTmUUqaZZUoim8Ak7VLAsb7vBT6ttnj+490so0Qk/k6MBmpC2KLQ5cVa458P
ABeGLi53hiM3tOn349ISdZHz8O4seQ5hW6aDamXERtrQH8Pil2GMTjG3I5t2Wch2vDjWxZAfCedq
FJspvy3c8CLkLfIysny/s/FDlrwrMaTx+M0p4xgP7EMBNBO6yAakr8kwUMuH+CwjGqtAP4wih3Nx
idjjPjb71bkrN4Xkt0KenwXsPh2wZnUmssk8iUYLNwXdiwcgIxVk7oD5pEaIvuGsVH4iHxRndYDF
TAlNqsbZjIc9+KbWxgG4hfA3oaxP0K5rrH65q/2F/9jTLhWdRFCBh2inoR2N+NaMNg+I2rLPZjM9
S0jJHEDBC0+mFF/X8eIZ4y2GRHvO1ogA/jjsk750ejrFVwF4N6bHbR4TCu+Sh44jhaKf3wFmW91X
T2P3nu3DbaYAidYI4y1UvK4aFUFzk4XbFwO9tF6hNE80KWP1pLeEVePtKCHL21Ua+8NgaXOiiSRg
pSe6tnnQ0YS3WPjYrzYSzhNKvGsDkgJ3QA2AQU+i1ht+J+lSIpf5vUmZWBhBDSC5Pgkfl8oiiKN/
K+9HLkomemU04nbmpP4ZTvL9l276Kz7qfEQS2Ng4D9C8zZgHO9PVsthxzfPrNupwGK3WQVAKnQm6
czu5b94UzU20wcaT+CWRjuDQCOSdJgy0RcsCbk2qPrHGrN9aDLQRfsdlah7RJnWxRMjGkxJYRvxC
/oGlX5DrDZmV+bN5bU39RFXlhW/u0ckA0B80ddPQeHlJQwvViNaRkJDd/ffT7bk93azU0j4FR2Vt
keqgoQOA0b6dMVy2Q92M98jDtZ+5LxKt2RUuibjnOt2m67SqVx3VU9FoE65bFTfK00MT/dlRDEwK
vCd9pc+ZyDegodIYyWjUU6jBPN3LeXVtL7I1D3aRqMs30OWvF5gI0+RxavXaTyBMMDN1HSoT3+yD
agqdq+g5/SQUbeOQajtPQO41FYhprhE6kyyUuA+nUUJb2FJpJUD1+WyMjx2SHshMRsIn37RTeIk1
7nUSgTOM1nwPNCaY1yBjHM+MLVV86SEM/A/hewhPhQqnOjhQnKccKPqAKaiaY1OYITFcoNeFwh6t
BrI1iJhUZLlLVA4YbvwN/CEZuye2LOZCIhAIL+MckXdfTAxQ/0GFdAqS1W12a46LemNk/nXFu9yP
w66sgDp/EuAyz6lS27fjg10SlQr5XE2+P7VpmhQ0g5UjiKFIYZqKyRL5gDr1ZVOhdpfCpBBkGNb2
0A4V7vISzWsV/YV/rx/sVoddJZ/6uhDdw8F/k7pKhZALeqCoxNYNJVjRqwkMrXKrfzECCdZz93yk
NgdwYLFeEaG3WTwywn/L6D6Ixdzf59aYAO0YQ+vB3p7JLx9yLMxT1IHrAkcFn0Faexj/YKl70sv1
iOOgt52JBo2DalGVKB5vnd60Wa+B2ra+zHwNWxvFJJ57NFnvLg9E1G+K/ZFO4nDxarPSlPT6pqnG
yy2HUjQ811yDqBBE5PG/FaUm8d9icJJWJDV/yD5Sr/JTy1jeYtQcxBqo7sLdiQB1nZkz9ENvTMPU
OEeFdJHmjFgPk8zRAgIaQjMETRkREZxOmNS0oPQA/3uCvnHp1wuu1t4vdpftyDEEPSQIvuohkHzv
PnPw83Yh1eDIZFuIE3ZBKQCx6HkEYxV4Sa5Uy8oTF7uGix0btZHC7hWz2kARsZZ+T57keWJQaCBt
ZEqePKFsnIu2xQCm6RJfOoMkfYq+EsMCZjAsOaYBCLuceFFXYIbnE+cpsna4wYQ/Ja/DLpyYmkG7
O1CAwdUpmJ6Qg99lhz0zvYKnXI4q1YLpWTxH/Nt03cgyJhOutiSc948Vn9ThPBkRZXgV6xyW7J2c
ggTH4IxhlwGNDFjoZDsxov9aWzLi2Psr+I6A0R5bapPtM67ZSCC/IwpnmuAXDNVJLZarHH0pbDDB
AYs5PwWKrARPGqZrZMiQLNuSDNt7fwE/dS+Ja+cDyMEAaykOcCYYrkRNCpF2BHdfzjEIcpaRN68f
11IU5/MQHQkDX+mvfvx5f1Vn7fi3YWXpuAMJnNVAh4I7OU+lE5ndI1V8/wHIbhLo8ZND895t0IHt
F23YNlzuOaoxVx2raHguGDjAIvgPXINQcAnYnkcicvC4PeQllpbzHVjqI/1ld//R22mbSDjFUzZq
k21zsP3Icv/HY0vUARmO4Z9F2SsFDjJKEfD+vcageuEJNz7XLtF/1PJseEuvxbaksiM1dFfN2k0i
a/Q96rYJ+hWJekjf3rSOqveBM/XxNZ1HGNautqaqcMaGLnVUDjrVEsGaVhqBv4TlgWVg7UJZugyC
pJF+HleTIxa9CyVnfyru2iGewAV/ZNLU2bcmx0+0cdCufj3/FBaFzmTYJZRHtra1BMer5pK3vCY1
VQaJlAb1JL/z50ZIcIPvhN8J+l6Uw9eJzUJZjaCxdlYrgZiM+JGOTfkmm9qmq31r12/9EJ2d0pf4
AI+mhDyyeP6Edi6sg1qEbYS9zK49detjiC1UhEDv/+PFN2q71WSmF2iU8Qoh7ffHKj2RDnOkfwPI
OndGWCVdRAdKGbIWIM7BccmGuxOkfSC8kxW99b5V67zOlDGad7kH7JX5TNsTSO7q+MavVlJxdD/b
oYiraPkqxILvTXDoO121T87ROk5w2I+twcVgNunVTpIOPDcLLlGW3i3XmDAGUVMn84G3VOt3HOeW
pbcqZdDoV6z4vFOZZ59vqviZBRRXWlGzRLRgTnNv6ZlpG5dkXLGRx7oEGVPxsxQxinVKYZpR3ADt
mgJaA0QEvVBCZIfami/oYdVOhNAUak+jDDjOC8F1ZnGazUg2P/R01Mp4avPxujigLGu1+ucOp++p
XURk2wKq+Wkh4G2alcZD+TPzI7q+Du1LB0GZjHltEzGZj0D8OP2X2M6XUpMZnoqNY/gFRqO6GlAa
4xcgzqjME+0P0X1+AOIqSvghoeXRglOXZ6yuumtvAbL4FQorgVvYB4tuI79xj8ik7Fc47F1bXcMM
XhKYEk5alCAZygnQwzSzAQks9EGVjJx7XSnpUboGrUMq8IAyZQXlq0pmcgYOvMayQoAuMlK+36/p
n+vqzmwr5W//vWLhFHtUfzfLRYGzg2pSXLkzmWD4RAHoQexuCyltgtoHtn7OVR79YtzoT8bWbOHC
fW2H+bJDqCYPHi3WbvbYDzqBROIxilb2ufRA+UnvFqLIkKLHZ2VGBLRtyIbZFP0abtk/snfC630V
TMVO4VxeT8SPHOmP6+XzEFHd79HYH70o9bntJ4V/GyKm5tnXTlI00jLkdFPHO35pL0gRR/9nI/mS
zxbgeX7jbsz5PIJfDAFYFDg1oDWwQdOypggzaVI9e0l1hjubgm6eHR+tS201BOCP4EyXn/l/lWNJ
/aaahjEGEVYZdFzIcwgZAkvesC7hvkwQK9YKWrFwl5co/tZlGn4dlXOhB+aR30QliN15o+zUzyQV
JTlJfjT0xg0FwYuqQviG4MELwV25VRFuehwfyYiB1RJavBEcZMxtIwmVBppcT1IW304tqPEsuGZC
QPVR4jh+Q/TuKjXdScoxcVDphQoW2VzzqsIKK1EeIPEvCa/LphLoFHngz+tAO2zFlZlLVnWGGs8h
Z1uPLkCkny0iGE3ZTLM60aIfy8mvCLfy79IiTJhm/zwSIXtOMplm6wfNKzoWGCIr4KrQZSzHbvY/
ohFhrXjDXMXolMQ+NTh5jpv3v1oPRB2ub+94JFsvHTC1xaHvvsSY7nyJroZrMeIVfOGUxVSdhnGj
1Eq9BplYOLBtzVvjyb28YGg21OAAKzbt8JrmZawaZCxxnAEitfh6cDDPvXH8OOY5bQnrT/E5NN+O
GQcZ1+wVYR9TAi1XKFdFZW4faEkwDl1RS6y5hcXZUGj2PtlNcrsLDBiG1PRyBPdyNyTxc2/5B9oA
x1hhu3niEkPQagAOJHV6ea4HTIjcyucYSjauwsEyFek7fOqGQgIytAW/zyoLn9vFMOBNgiSA2K2M
LQaeTFXIZaxFQMuDS3nBU/BXpdp8Rsgf6R3ojGMDnqY5I2e9W1/NzYAIxup7reeVJcwT1jpc5Tih
/YWCHsz8qaTZPN2sBt5bxu5jkrwIhu4HTemoyejBPZBr7pNn8mWwaShLHUQsppIVRp5zDEcVkw/+
zWO8Tfu6sQbjgN4VT4Q6rYWK5yXIkZgIu18XA2pvpeNAk7amtNPp81aCeA7+iGinLX5LKhiZkP96
cxzRGYwmD4V5gfh2TcEdHOrElWwIuuJk1NtCx/4AVC/tXtuTb7os8jlfThbBL9w9nOoWAWpyZOKZ
N3S0oM7DXa6boMh1/DB5LYkH2PE+N+/boDuD8KJhtIuDKyZ4NjsogkA9MW/zJ+AHK/vok4Wa7t2p
TOs68jA0b6fYX/33EVq5h+N+NkDr5LPmrZSO+ue0GBSGPjFVX9PToS3CcXqTT9mwOtPheVRaMbuP
aE6IairSiKxD5BOGMYXojNadZ5GAluPsPtE7W0I2Iglj1rl9+UoPaY0XZSGKqh2+vK3/9XufZFqj
mtxNDTojaft6Kp/yKpahE1FNeKa/XkDBmgheyMLOZ3bid2m/RWqP7Q6+xhdZ8PT3mMGRKccWN+6R
E2blyiKqk98BfFrrubbFJXt1xGNtSdQDK1JbR6flu0HkElQzrK5U6MXH6X/PZIJPBvfK6g0x3GbP
M/JgMpK9dFeq+dj/02/RJsqU5HMB4LidKbgo2r/reybIWX4o0ZAlpGfR1Y82ACUMpUVB6PZIBKRB
nYZIMI4kUFnBqRdjWrVkNQ266EQ+KSS5cu80IE/Zcr2aHLRTC8Ik611TcnXiY/ks9tQVJ1AJG5Da
8SlLn6BqUO2KD9KsluizbEDW0eAp7r91eudcXJ58FDcsMGFjP3MY/bMDRNfCydaHpEUQC2a5BrI/
tpo9CB+5M5vQ5wyB+3xvmFfr4coVLMpLqFJ7V2BK2VjOTkfPuXrXLuUQ8fqWqMWFbllQimQgz4CE
lcEjInbDJsqDrMlezXf6A6jov9htmeH6ktqdtFjFadZt/pN0gEmrsylhoqvq3MqTwvMMh2dtfUDs
aQBqBAmjrldGxNlpCYFEhjEl6sBo5eSDcym5wRE6calHkYClp+VBmYECqaDCz0ryVVSMgkg8ywi4
cK1JbdiHBZ6/1XZNURGO4CGQa+Wjfh5fnn0akiGXDJkS2pHgBfLFpRmwGroHweFooOkSJXC8dbDg
rd6Vu2UUJIfUoMljq0NM/TDXx+5tknn2BP+cbyR+C3t99jE++ivuvKNadVQpGQDcBfZXVbFWqT1H
1FO8OixGsi5hj/HGwZ8cXqsGoeHRcAZRm1NOfugd91hYNAL5bbUXoX7aheowKXQ1f16tI8/KIU9l
XpSb6x+pQtfUrWbjsHaPzebVKWJAmUJN+dKvtJFfUIJ0c5ahRhuSREDIoeGjgjIZbI68mG1EwSrb
ND3dP3FEqFeueyYi0P+oSyHIhElYw8Xs4lwwA17W35W6lS6JxJQk+rzYZDLBOTnp2DTmvr2btIvf
VN6dxI+P+aGZpD6wn/j5Gay28aCcQpRs/gNflWL96vqbNuRP5OD90TZdBiiUFAbjXUrL5p2TvwC4
1tzFzRwS1YCX6Zj22od0MdELm71Z+vpSCZG2YA+e1rwmThj/1uLwYlo0o282nKITfQHoIvfru0oU
TPhHeC+6YHH3FjDkv/NnDgA/Jf4ropo0ZrEb2OvJLAHoJqybUDA5kUvrqNgEyofzsNFlv8HxSyRw
PM+06pR3cij6jmHkFn08/Zz/jIF3CuVWnZwjVaDwA/GnnX8XYxj55iCjLfwOnKDIH1tEZAMz5zpU
ooj8L9DZ0OCnNHPAfpSOIYyBZYMnaMfCrLf7V2u3fH3QLitl7OQvR+4cDa/9hzxTgV+1mdkI/QTH
l0Wu30oNfrK+8vZs+uw2RIvlMi8tVOPUQ+EOLb3nhSDKeZ2sS1N0l++xAfU7xvFabGS5cC/1fK/A
ER2yr5xEUhqGNDZiacsoMFye41LisVWd0S9mX+tzxwIMWQpLQIBiGcd5QAY9qiv73AhXL728uctU
RkF6kKC8weHyiQBaKRGkWnp0GTn0JT3G9ONjgUEQFQh8VExPCmcitbrLjWMKR+UlYOIZ2uiTBpmn
UNDAz81aIKXrzjDadqy9kC7CPSdgkE8nggmCcvuV0v4ibNpwTdOEvpualVGM4ZUUKFJlKQ5neD7b
eR8wKX4pqtPYqW3AVeFbQ15iP4PnDSFYpxnDmQwd5F4sGSd658qvChNMeNuQiiR4AghtXNs3SAV5
AYN+wY0ddunFsmdz8mF5NqWbI0nHOYkllbxNaYF+5uIh0VandVjKtlCw8D5k2Z0v4JDsTvsrMWOJ
KKVORaXigTjPo1nRIer0X48JV/woQUIbCCngz+emoskc1Nv5+bJRNoTWRd9p4uDrls1/wl/6T2b0
GUPStDglHrXPvNCb0cS5iwuFijYU33H+cKiYcdIHJCLPNXLtczIo35uRmxmo6WdLTTnyqtkmiHE3
8+06XVrt3M9BeVFa/zoToEuDKRyxK24FLrtmQzQDj/LFCtYz6oLliwbI1zqVhuHXt61xGhDE2tpw
z7KzWV3ViUgEx2FDe0dDvbiC5LIcKsC3ZVNJu0KgrQpMyORMAXd++zO/M2sLuVE7RY5xcL+i3Fa8
RBdnPToMEs4LvJ9E3OjqR8Cjx5uL0REZA/b+gRW5RWUyP8x9LicpShx66MO16Vu0FqXel/fKOBvn
nP5GlWwsV3m9a1FwHfFkFRmkKIoJDEz642EHM3xRb4PcT8eqZWGb58YaWmj2mKU7AW4CIifg2wWw
t0u8MgEAO8GmeiPUs9Sj+fZIEPJ6Y4D2BRkf6ednGs5KRLOF1TLAatHzU4vS1m5p4/M984GDvPyt
iFr5BIRZURlvAm+zeMugt0e9RBdBV4ExCxqhDYHCYnCqDtdIv4bJLzPRuY6nyuKh//QXXeKoE3f3
v9ioMKkmV1U+W3UbcVflg/nNpd4BHYvzDFJM99pe70+6cF9dR/iIW8CYCi/ptPm/jKlN7HlmzfFm
8J87ZhkliC18qhnNZWmBdF9T5ahxYKE7wYqwXLmr5CFBLDATfjcDMXyFLm+pPuGnbckWPtinHgiZ
vaYUnzJrdGMgx/lHplRxXjPlSStW7wU1dI5wHAgTVBLGCEIAU6LDNzF6nZm5wbpD7ii44XMTO4Bi
AJCByMLfMDTmWiOxOcZjgSupOyRdgc2yqtv+44fIdxf4MXzvzoPWZNz9tY6ocU/3WtqxV/DnoAIS
yx86HedgQ8JQE5sfC5NW32dq7+L+EVP1ZakEQOEax4Q3coOqlCFyceYOaELDD80R0lTMZUwHkdRX
9c+LQZT46UCyyjgkd0NI4mgO1UElPty4dEqY+o2l/+Ltt6j6X0OZiz3Lg2RRAW9S4iOG4UHEeeTa
rMHX6Ko0ezz6AFPnvExtk2pIYlr2jle5LgySd8fzEGB9L47gM7oxhxqD6tmYclKObD4A2Jplv1HZ
5hhF4u20wXyRG2Wjl6VRNtVmgP05Kz4wE6cpBlukQRzypYUtFjzuAbk0eVQdybv6L3jH57noajdB
Nzn9hn4IDI9QeEHulzLhyVGwSgWsZthl7aaZvsLtNqLyKmRmhNBiQWeqkteIiXuTUEWFVPVglxkP
sLQOGLkA66byUr36Nizg3nbang5GOpM4rapUBV1Ytxk+mJ+CJzryM8mclwpmmF110WrCiFhn9Os3
m+Dn6CSKVBDoyj81cYg64DF3sddhhIiC7YNF9ztVHiN6LX+e7Sv/WW0bdMTbjhnnCreOXTKxu4We
efzcbiUvY6LL7qbGVB1QxTFXkiV6zKwGzboUuuGlNCi+EbguiOM/6ZMqOXolVrTWY2uJzbJjSE0P
BVkvA/3qsl61Z5Hdkbk5AoZygDlkqgjRQ3RT1qUsey6OEsk6gb9/4mCPfhsjpD5jNoBS0eiLhIan
2wiSBrl+Bb0Lv3tiGH0AHYLVFyNjZIWkEg4GZDzRc0Nf/0uLTBPZnjmqh/zSU3PMw+6S3sJKserH
68eRcKKJRcI431yaaeGjNiQ6mH0BWMA7tGSnvdGD2WShakWPdSGCMHPOym5JkaMxyOFl2KoaQx/0
vtoHi0X7nDlLWeLs67PqdFRIXFHxaemEK3dV1ORydMOe5rOj5EathVAH2l0xFUnsdbjLb/wlrDUC
3d5ypeN55+VQelOzNN+lWT3BsVFQ1kTzO4c0TvoY0aZxUHGh1H6fn87w7yrNfxZAZ0HmnQudmkVh
12u8d25jhDk+wItmWrJHTv2Myztipy+gj9KSJ7EPAS1RGHEUww/vZ56I/dtitVY7aoh2c2o2BoVv
63DPFkubS2E5ziCpO60HVV8Dx/7aDgvoM9FrfgY09OwpJyIZFeOMKugM3HmX2GBMzOJBbNNfDp5M
kiUZ3m/X61d4R2pz+fd2qKz8IAEKOYV+48j9VFaEQTfW4Ky6pW9l+U1aZkQuxXwBXs+wkgg9wDqW
CpyzNlGyz+4yE5k0Td05Aea55fQzhczFCcMCk4G34A71wDUsCYsnqnv9h+MSfZ4nM9Hsx7bAjmNs
0ioC0LVLZoHdJm4j1VHRNnT0HzkUvUOfQfRVOZsmxhT7yAnsBdmQ3JZnQuCkCTDdIhXrXrTF2t1G
/IR26yKjEmI8E6N1hMvo/qGML/PP0M3Pdaivt+vlyYGvwtE0UynjitF4cWb7OydF1tl/whgl+DCN
1RDbQY1nXVZL4wNe17gSEgi6uHP4Z4X+UiDtdaAkBVQSmrIrAMqMBLeKI9Ifz3gUn7XX18cxr9aB
JJJdczUG76yQqk8+1+AJ6elOY9DOfEsPQbKw4HqNVYs0cGClmt5tJUAhV3bUZ5llZU1DFF9ZJAWp
jOOpjfKGcDhue2Yfy8SaQcgU3XpXVRdzx44npFfmASQi78OZS1mROWkNkMUuyTUzmFqmXhT5O+Zw
ACNQdr9FXhwPq6YlGYHtwOa38ZURz7bMmIUUP7SnqecV0sH/yjNQwYTox4UmSFhhgOnwN3iKalSC
pew2Nj3lADoy5P3QqQWPpuzXiDNpJSHRNartWtjvt1okAkSYyFdT9Kt7ecsmP8aE8t98smXy2nXl
BURzf8ICWfPcy+GLGCLPCb3wa4ElJXQMGTTHiTUdJqOhCxuISkq4ZTxSoKTb6VqpL8mhQAr70a9t
ZYhDU7lDN0W5/bPcrCUPpQD3Th0CA34VFDUtaWFGOFO8aYERL1jTNEWxi6IHriWdVja4ESlWwi8Q
qukwfQpQKS3cA+maBqDU60IcXXMuTswbtaqe7j2XTgbOfODzVd+2UzUBaJKnTOXOcz8b79GgNtax
r3TgV6JAVly59NrV6ldlKNpIO6Mg9AZZVWNorXIfQg0NaybBa5fO5YehT9v2SYQzHJHrdeAQ04i9
i01cPwYzuTarrU9Z6vhQ2a6ZVcjSzK25Ee2gggXHxWcU8cg66rDwNNj/fNPpItbjWDXid+64knnC
1bHLbQ0QsazDvGiPaYL68jOqS7MMfCICV20qyDuecTPdSjxUsRGNVy89w07mNFIXg/IiF6f6byau
K752DadVt3hKQZa07X3S6XjT3BK8mBJwzrjWQiPRGbYzJKUa0aXhsJUF2lvFSM94Nf6MmSwttwhi
sQmPx6lhpts97pwjrxdqloLUqn5o0FjBA9S/wxBvsQcA0wdoPGJdEZHd3GFqypMqRHPMgJ1RpJFi
+wW3HOxBYEk2WCZSnqE6KtsrszAk+VnVW4pFtt7uxe+yEYob35jt7MB3WyTc+3evG4P0T57TqH+A
0/Xqti2Yhz2PsIujMDbQoaIPNyrkNKUgx0uuEL9ecvxTAEhHCUdKAvPlstG4WmXFR+F27L4wPYS2
e95Z98gRvaUPcwkc00iudl/sKiCCSZgs5qbBXls9fkmq//X3W2UmE2y+P+9pRWvh0XRNj05Dj9H8
Hrp56ViXgmyMgu0usp7ToLiYbBOPB0hWWfSqBt7eBGKUaKWeQck/JrBxz8OP7fntPpdL45fbnv9C
2b3pMViJlFlyHTUApGepZ1BmcglGHR7MOKbWXla85wArRRDwJ5Gpzj/n8RkNxxY5ApMXvYYtfxdi
Nf3B3sayXgp+Z476kCIgLNgfyESw4r/WdEw4edCXYiu9Nak9k4ucRDJNd0KvZ+h3oPOO3D5VwdTk
turQBrw9Il/5/fCsTQH9HquUd3tjf5bHJPpNx/r2FKsw4MPidyfgYYf4X1tSQWgh+Fr+FJfIpCo2
xkh3OvCWgyHMUa8Md5Rt+3kaZDLJ8W/N+8evugx0wWdR2wiVeNH6D4kiQf183JB7JqK/zkh8UkeO
6R8i5rcyKhSgEkypt6ZqN4JbnRUQ8rYmUO/ieiOz+mK/KsdUsEN2Qn2wDjhHGV9Ed2qnb+BK3Sbo
MRl/ry48rJxrbM15OWapQ7CTaCHrDl2ax2zR42saab67LNb3uJt5WU0zVUKgKrOFVX5CWbOpCssE
gE44vSbRo9CfbwyY/DPbBpK3eyS2NNPl0fwvrEYEcLIK3W05LhGD7cvuweUaO0Wxu7xPquI0IyuS
DmyJsnvYIB+DQ5N8/uUnZShpMEDfC2UkOG6kp7pT1dyChfYQMvEy+7TCjU4jid9IGLSxLvGoNyP0
4U7CALu5hu1XuCcRcfk4AUTPnXytIaa4BLfcRdUA+0KCELL94tC1oTc71Zic3zKQLkqNpqSl/fWv
Dfq2gyV17WdYM7Qki2bRIxKwfJ5/7+piYc+t0r9O4C8L95//wSbIFym1MD3AfW1XoWXurJ8zbFzO
KtYB46naXNGQeKts6h1RUwZ346PXsH6k6ck4tf0Q6yjqnV+l/+f5uXiJlAYLAeUyU6eV1UmeUKfN
R5h5scbuilrEfiVt80Y+rEGd1l7QzvDJW3/owbyYMA0sWzW5UqMSjYApDY1AyrFfJFtMwy1ZyTEw
xUp5K6wOhkn7NRxCSYKTiYqz3xlQFRWPy5d/XvfvFCtjmS3Cks5E3BtC9ZbKup/vu8mAcammwnE3
Jd4Bo5k8ZUxDtJMl88m5e9RbcQCF3T/6tWSq1hLspjD/ysic2Q5/Gaqc0rkqkWTE5FAjOIvt2w1E
mr8Pgbs/ReMV+WdWcpG2gQHYdHS7A4Bs++c4qWAPJJNphO8OncNMqadmgFaSHkdLmpb7uGXXa3HX
3cfaoLTdI7KeWgwrMwuKW6dBTB1xHzm1Rm/PRE056NlHGznx0joZ/yZn+2iYMjjbFvyGVmaIdXdq
WjM8ktni20R3CkEKIzPAwqSExQdRDeB1zJ72GLfWxirtfDqTGgWhGe5NJTvbFDFFIQhrVY89nQ3v
XMlX93WBUszazGpUfFX4BzBItJKKtPHff/fdyAjzKvMVqAq+nb2o4MQD6MT2l+4fzvg8BkFDOqh+
f6a5T51GRLF7ULfLs2nF2OWSQeuDFEbxU4cbOb4/ZHo3zhcvKYNIn897+tpSYv/W1QCZJADX8NYH
uH8abMZXyniWsNd1VgJqzQ+VXNzpWi7rYEULK5fSUTVui8nr+7F2Vz4jkF2DtLjzuH7RBuulJD3m
i4PJ9yWEikBZpsLJy7WzGYZYb9ORRfX9Vzj7tFLu38FFP5TI+DUO60w192ATOWL1GwtEap1qq5wW
54TwsL74y6x5LPTpFOGb2QGseWUupvsxzmdf5YfLnySSulo2tzEqAJpjwaQp5SnN/v1onY9qQ326
ttlJtNfZuLNO08DdAradh6cOpgEMbx/qyKlG/oXnqwSFsfs7yWv0EuqI0YfLbP0U2yZv1LVtRL0o
1iPr3N4Hi58e0+BbrWP1uwPVO/N/RD1eS0OIMlyuNCT8O1oVHRB5GEgWdfaAY9bzKj97IPil+Xip
64YOTbF8DB0RI5UDQA5nsubGD4NAUm/10Fl1RjgJ7cqxD0mU9QcmGaJRT9pn2AFRloknxXaHf+4Z
nTuVxRmmijLjnj4AWDP2l0j7nqj7d582TX1+a2WlXH+bHj90oXXlD4seNOjqOT7mPzI57qeKGVfJ
RcGVSlPn/2mgRfYXukfUqOoOC7SDW01c3Xkgiv4XDfCmGCkBNRkgyxE4SI9xmYvQ2FIMYPFgq2vv
08mtuub3SfJxAsx2wsXAbxrsLRwzNU2Jvfd1h2R6aeXgHRjJhy4g+wakmw9QyUpY8RE5qWd3zaU3
rP4GyFhcvFmUcgs/KfdNF3j7A2eXAHcxuMZjvmTONMRUqavJF27/KtENdiFeGFuQHH+7iZMolfdL
Qid2S0lgTFtkketuyufP+jqdmRoBV4dYsjM3GE2wbVOfHhy2HXna/FPjJqVbo/qgG0qF04vsQ+23
0vP1cVHBrlZ2Lr2o5xv1vEQs7HfCpxNt8SBONwHuYxLM+xihC35Pt6etYZF5S9GkzbSRPn73OcdM
0bNzpBD2B91N/TaQf/pkB++IMrZvJ9xbPMJxFtlJOTzKe7r4o1b8Cytq8KQ34y43iSLP6nQ+CTTH
+jHZ1OoGOOo3eSbbM7kFhBIzJ1Mg9LmBBZTgfoAAK811dsaYNsVsS73/rcmbW3mw9uk4MczqCv1x
FJ+zoDktLSsKoY7mUHHrKxhZm1aS8kTvm48ZVw+DzDfkC25GTTQ5uXioiNSVOMoPQn0NpsjE9ST0
1mEEviSBNira0IoT47wmmLhJEQy8dhK1/RzXWmyz057HxF4Gvbk06uyTEq0PWa2lxiWkCFABm+AG
JJU0H/ALr+G4kpDXsV9FldkzpFESNCUw5obs9hnQo55UbRxKZlKExv6ZDnMVDjADymanaM3ogScw
qabdVJRyvX0er9ZRKMf8KPWJwO+HvG3nST2oRGmEK++sNKQ2IrYwCDjUgGGpsRdFGETYb5khEfyV
M5vdjXdY4J50s1Mz3r4F8/tZe0boaCaSw+bvVD89Uhml8UY2XSw1qWvfaDkpWEX3Gh1FbECZe8PV
YPRung/8meR1SzuTWYhh0YLtp/fVMt0s3EYrhsxQiMnURiUn+63QG6vbrJR4iz4oif6l+rrB7fc7
xsRIU2PqMhPON9LqLiYRcTFfKovme/OtkucQXnPlT2FYcNVxPhqpR4L4Ho9lT9zyBmtfgZwt/k9p
rebDCUTEWBuiq7l3JFCN6ebeDGs4ChtDbxCjoZLAtejV3HZaTR9VA/HnZ7/8WXaxnsTYTW7SEJEl
9IpOyB9vTv1WRptk91YKR6S0r5S1O4+6Y8oH4PxPWAhgMi8h4XoQ9K2WZxt2w61+0F4OomxTzrap
s/J+pJ82c2mvzeUkHQr3XgFIv6oHg6w0POz+873tHS9WX3JQfxOsW8BjOM5hQiXwJRPlQM+HB2eQ
6by20BDE5OcDDd5hUg9Z26614zVBSdYtaFxdMwG3Bugkk6tOoVjhIjx5jUmeebjdfyu5yH2gepqB
/9XvdQUC6a1WnvgTqZFvrr1fB6GWjvYz39URN5qNvkfbiM4nnTqkBoM2dM09B/j4MCZqpO18Xv++
sbKXHZsA1LBWbiQHsWlQbTGPl0FkmWP3J0f3Y8HV+jK39NTMyiSygvWTzukeLt3hH9v4ZId/8p1x
991+zYI0kK029KhDjiUu5nn/il1Q86HZaIYML89JYVffm+uwAMGksF8jHyCE5DxkhAmRB1K7in3T
2/HgiugbVR3OAEjFwrbk1A1C2aTekAbo9IFEUrpnobBIGljy/kyf5b5Ylf6xOyopyNY/IgoBmRuB
bg6MADN1ujkzDSxzs+07SgbNuVozizeuNKgJWVQ5ADO3kk/ULVhcvk6foldBXNZgkwcxEafZ7VMT
T0ljR9q+7LHOnme1TrQx2pWDgkYp9E57SQJCNLfpTSNIiXuOtJZthHgf2CNVBZhwc826L22UwNdt
HHFgjRYk1ojBekn9ODqw7yurPfOf4VQ8cuA1dkC/mQnZqwNzK0wgNvkkxWKr+vunlK0lLm3v/Kut
vK8nloG7jC8HXcRVwRLyODaOrSGKEo+rwwH2SsS7yI0wWZJfXpmd0s241RyaxDbGzGJ03FiojsY7
DOaO+3zdp6PWCRpkcMQszVVT6QMJ0uWixKsKN6LeEr7PcXT+uQuwDXY8SHdvG6aobM36mytw9WSd
hSq7GiRmegwGFcSxuvKTQeHD7Qn1DOOgX/B74+xie8xPCPsWW+Tz84OqDITCsZP8Syc4HkSANDE4
76hGQeP8tBd7L98WusAs7F5BEP11Tuz4sVww3b3gpzXNEy7akJfi5RwdVocxCkHdDyUWnT9ZnJqX
9esQKKvkYIySJYFtmu9uYOc3eHdhJliOxEhcGRiGk77ZcmiAib71CK9bi5GFK3gyTCyALJOfAMjG
1N9w3FmFZcCA6UpuSCfBhoFXi5RsZk5cvRsK1UuMGfV8xEIC4lXIggBS1DYZiKYJQ9desX1maJjq
hHdUbeoH9DCDiO0PvocEgvcsTdH9brvDiQgCzerFpw6d+b1M4gpatOb+CFRs40AJBopRysUD69xx
kai4zBjprbnLD4o4IowUsNsOKG24zJpEkrDkdxNPiQ8049nrbphceW8tUDBA4U5ABVkW/8w2wlkG
QOtnwOWgqcRQDmmkkymjmJ6gOOBnHpNwT6NGuVYIl0OTE4yGaV33ILL6AdNAE03sYET7fMmpY+SV
lPZw2iVUd7xlAg0Zh5DQ5vVOqiM3t9kcmk4rOuKK/z1ZbllsjmdWWQD24lr5BGuahLu1xH9fnPNF
yx5wQbs0kk4XJDrXrKmANzww3aQAczIHL1QqxvRSLMeKClJ/JndeElXsQLrL+jagbSZHVjEfWD96
iMM6xI/lMtzbsepv5Q2qUIbQoC0clm8TQOwIXr+Jdi5o/MHpWYmEnBKn9TWfW+0ImJXi+WHZy6i2
iWsznuF+nV4dI5ojjs6qaqjLIiGP+rLGOoB7d4QmjH7zyUbgIHv6qnzv23TjMJKj69EWsZN/52mJ
uu3tkTcDOXqIcFh8Yh+3I78+Yi54oJ6iweQq3flCKHjsltU1EiJDjgvxyfbv6wsJBvVgRUDH7EgT
t+hRoB6Fz/xNC9ZM/EkDrAIWZGPUz73Aj0Vm8ryfyoyum2+ZONAQwPaVL7bnUKhZeeQUnmrMpP3/
v+DZYRjkgsNdl/Ad6JDo8BCaFU7QnLYazDLpmNZVVvUHhZOkQpVANXaYz/2jzd7Hk3ftNXqrQmyV
7Si6Qj5fwlAFL9AQ90QrEbiVFqPx8LSxFGbwDYTQjhB2qklOX1Rf/ofoY7cMn4WmzT8SHtdv9+pm
EQIE2ggeS2u7SV4mHSV9MzQ+ZSwLjZY6omLcHC4AKAcR8VsN7FdQLNw5UshHpvBGQ8tK+tKs5W0x
WLlR0EKKuSKC6A/h3dt6e8rHBBRnBVACQDvnQluZWAvjp249RQJ4YmryhkJfGQQbwoZ+Uho2jqPk
pn56g8psbnpwpRVht9LbI/VOSxqVxfcG3L/h1xg2YoJlu4fVXaRPh8F2DnUk0NlgmSWzmyFLZtHd
/ijMZUfIQvoZwhFKQzGUMQ7CkTS4Z5iV8M4e7e2KGDOP/RymK1Ng+/hsRqHpFn1z4vXcxugbwdkf
TGKCWeZ4Yv26I8T/IFppinRGthc6OxC6KB/lFFybUyq1z+IA4eJ0G38yRpqamzvxkmSFeeRzvCdP
3gagv/L/JP2q/4SszjWsUkeR9P+uqdFoO6/F+lH7cCgMZRhBLBo7ia0eWD98u4IZzgvtWTkNfXJ7
IVBnRSE0Ru5753x5oSKS56G3VglHt0s13jMa9ht9MM0ukKNueR8onR26oSHpGyIJiipFcmrbLh4B
uQq9kDjjt/JIVyk4uSYkIT9zFOw7tn0smsq09mZ4tTFKOuOaXcMEOWfnYmIiGIDtRil5y8tKu4wS
tiBj8gHu9zTRCuGcpOK6CfMPVKGgLEljtYRlv0vjbO+UmfLjQtezntpEtA1uShB1ch6JxIlCPHvn
NzQr3yt4H7vMXpTpABAWYPHmuAsWqMZpc6p33/RrniCacVmqttXPu+v8+NqYI+9LdvE+bhntuKY3
vgeLYNSSF9k/LyxWEl6kDWAHbeC0cuMj6FAdZg7mH5xiu9iDi0rj98QCPYHV0xZPQJ+hiWR2zkv9
XVCVa61k/5fIjNYCINtFiR6QD0F4ZyZtkbAvWIL8P0YiZ4flN38aZ1CQwW8WrhvRu+7iiJzuxdQY
nrRtFVXNBNm5acAtwB//rZKnXyfxnzmsUbqTE+ux8oXLBArKhmcmbSTWW5PfoomdluMZEGMqVYq0
2fEoc9yM+aexHCRSZLLxteyjPlHnuIv6zeRq9KFg6VATb+0Ttok3MweeLsaa+TCwC8lECJqxuQuu
sCk7ZWHGuH24PvGzdlR1ml7YLplQ0o0Lz2vGJGeAizjMx2B8GcSodwb2F/09BlfKmhq/4ctDDjfH
vm0roJZvT3bFjkmG4BsNLDgp+hZXz+tt4cBiAkrqSSXoW/8LlsIkXl5dg7EYvLw+j2+XI//Yc5n3
wSbDbiYEIq7Pr2fsMGhUElxVxfVsv7H2CNZnEuGS4KeQS/KJsRcvs2fjIrtj0Kg5DKYK/2/YAOvf
NcTuloQofv4exn2KlJCDtL82YYd/jc5cm3mHtWxUa4mqNicNSXmbAnBdRivrjwy1WeWcYYHeSfBT
o2jAkfgbmhVvcySz8lEHY732SnNzEw==
`pragma protect end_protected
