// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:09 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FkRBRAAEZtGaky+YuZr7X9FKG+8Uoor6kkM3JDS7o4xLKpJnFhJLBxLXBqmyLUm1
CUFb8oO8JpmHTmcATmvlYVhJEYS2HAgxlRK7PwlHR3uIt+qOFVG1jIhW/YkaghSA
Ik4vc9+Yprnzu6Pw1wMoYNOTAMRgzsq9zwmxrK8d1fQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15952)
CJPvPJLLA+dRQXgSqMCdWM69+Xpp6pj8gkf1RdBxNaeEs39ta2G+4DhfxfqfcCv8
pCunvzUs+6PcV+MDHNFccK9tYziThYIdCT7kTWlpDh/VY9RrYr7xTvOzkeR4PJsY
7K70H9Yzwc9dJlTgPBrT1jyAZxxwDVg42RPYNyFIRxCU/ONKkiE1ikqVdBJssBIQ
ym/JbQjYhxDh4d556+wYbf8I8LXL7DgeAi5WnXOSpQLlXNK2A3MfZ1d83teAf7DC
BY6chmhGn4+f1L+kIh4NlDU10QtAYpf7POhaMkMzqfqiaofkv44ec+5e1L+aarwu
n5PHgHekA10Mchr2tCvmBmy+54XeviBb4OOKnL0kHITmrRJPle5WqNoHNzGLZUei
feuxHJ2MHtvL1R2nUsh1qvaZ7+68h4I1Vr45iAf0i81p95cT/AyaZ13v2N7GY8fa
hPyH1c+O9eWlQKUXsiHRILVwhRDWN2oPUHw3tE+l1kL2CQBa2FEgHH6KUU3AuBix
2qymZPhILTdyxWrtdahZN8gmFq02Z1Avmxn5FIeCqS9B7TtT5cNhBw/i3muDw5OR
VKSHEG1FevTmAISoSjlhJRKcRS8+TJ1y9cbkPesjLgBKls8bYKDe79PsO1TwB9t1
o4CuSoPkFCK0982uFWRWiLFKqCxWmkRWUXPBMDIjHZP2OZJ7298D3FO9DZB4qyp+
GzUPIdUH0+64AwNRIIP/n4jecdEAC0psypMBRA6WXyqBhLUO37YIhSYf6GNKgJ/7
wOd2odCIjic1HfbcPEpXlg14l6cxqDS+CjYhtXVrB5H3D0tK4uHxcj3fI0W2HDPB
AciK+EYt9B80buvROif7KV64NMnlLUvDh0XWiMtu+brtGOSuLnmnRbFrMpsp4UOu
IPcqT35ReDJRkGaPrsFJ1ExFk0b6AjqBqHd5sJHEmS77VhhsjgvvyOf+C0A3tSeJ
77O0lfTanyvXbA9Blzgs55dCCv2DcXptGCbXNOvJb7ubhMUO6MZw/105CpwrOQ3r
L636fWiIail2syA3BjxLQbIq7fDLal/jQo0UDCgml+mtV8v3AKMfYbGKv+K9ibbV
PJfu4xh7qB94PnNBmPDNHruhgOeYPPV0SzZlE7EVjV5l5P7HxjXQwPpw9Jx3eeNG
jslr+H9/cSORI3YMrot0dhdsW9EmIJenyQpcbF0sDG+Jzv4rCpVNgNlRpsBsBBpm
HFIu3+GZwh9H78F6ei7L3wPMqJM0dZXhEl2EERq/xYBgolzYdWQebMJLZSJELX4J
cvXrqVvd5QaMY9+X4Hvmu+ZSBm3D+w+p7ZtRDHhEOoy123tNpt/DI2A0fUWsdSUi
HdMqb/2gJ63HnyZw8PTWn3IuM/p3jlBHI0dOAWjtGpkXYv0EOEiqDOY57FoeULS1
gW812xyzKGTd8PYldlLGldl7FxHHa3W41xAYw4MAx1H5EXJBNjAATw5EU1bmAjtV
hlZv4hGWsulWt/kiEhhup3J267X+tKx1wrRUx2FswIFE74tcZHQDB3cDSjs2n7L/
sUa+4UIlUsPEjOmm6kXRLVNQj2pGFEJTg2O6gmV/o8gl7gCUcP1VWomqWEIGycVI
cI9VIBmjHBciAc9ksKhzrnaEKUFyjTEq5SLaocL9dvl0rEs9mnBIlqbL90SkfWk8
d4BGMNs1EcsMT8HUaRYVQSVsmf8wewinPHvaMUnTZTqxvkCyAzRHwUJExtp7K7LE
T5TM8fhymMFDbyfuBMqr/5FTTqOWECKCANUJObE6wu6nuAMzrScxY0Vz3v4Nwmit
NUL+P7aFD6BupytGz+5yc9/KF/1e5JISYYcE2Ha1v0oWguO0gW3LNpNwJSwzw2QR
XM6BCh5bgNU93IJ1TAVK6G1nKl23D2skCWPDugu8GzYHuhTfIhm6S4iBsklz9rex
k1nkxe1Q7brXDhlAaDNb8iYO5bj3M2u9C04R+cgflVQhvNqPtX/y7g6/dWNzrzg8
B1bp9VokfX5mZGGT0iuYezY6EXSrwdORSM8jL5AY3Wn9Y7cIyK4RhtDjpFoisIf2
mP5o8VNi/pd7+uwHsn1oPG5Gy9JAj2UeD6NXoHyVqcr8urlSec8KdvMnc0RjTh/y
OstBsYzxE7qcTor8mWZ5nFb5K273lZ+VAU7ZYTTS3owEko/RtZid15vD7EAfskka
P+YBztKHFVrNla5+2FXo5Mo7SnNE1/EoIjN8EQeqbMg6DsssEphoeptLOBTDg1Xp
6jIqfZrhP/bXjcZ4CUGzHp/ukg9ovgiV1aZb4tAlOmIirJSLJKIbb+b6OKg5/RNe
6x88pKSO/L5MPM9/RwlUPjgPPqNptqj835PXVSTl+S7cD88EJiLL6RxuRyGWjE2m
383eZ8w9j7X6SPI/zGdwYDBJJHs8BR3npJqJzioEpK3oNTpIG81VKVsY0oHOXy30
h+r3zSTHvV/9jVtApF5jXCd8dWq1yNu5/8zct3Oei3a0+aNEc/Z+S2nZW2kCKUYM
YDABPHGdflXlt+WDMTq3BDsLa4raWoHReIQzkULlHR+RLFrC2zWt2/8nPx+lMIZI
nM7ChuZhJFEXpnUzlz0HaQO2vkBBs318WqRtxbDL3LCJlG0DhOiFEAv3UzAl3Kxb
Iv5rFtTGqENIDtWkFTq2mDIcXqkxta2PP9uzOMJ2ncFwZHhHdiAeNN0hbefIcAgg
HK5cnh2/ge2mO6QUG88MniX2KlWx8bVueLPw9qQnXPOtzn/dqCqQp7K0p2Lfs8kt
22PFC4/9nx+b7CXT2yJT4xoyESZhXVYorqAFAjGrF9ZEQq7JRyd4CWf8a/swXhx+
6VEoEaUX/b+d2Snd1yk69vuCoHhilTvA6k/lvzYG4IZih3QC97UoWJGrGjuMUPQG
JQR5rBGbHb18nT5eWw8w4pT4y2DhoRoIAm/H4V07a9nDmk9cU+BA0DV0nCX6dEg4
4tS2jRwn5AFUFw3gL+56or8OLOJIddLCJuF+++IvHX6kf5KH/mYj6UFpOLilaiMN
RfUvycsqLsRJsG2bQ+hZD7wOqbw+fahMvGTScBpTNKjbrYGAYP9H6OP8LKybg5r+
5bc0sLlovLGlXCgu78BfzjQyTzEZD9nszrKa5gXBnpBe9mbJTN6rgq1mXDgbw4Y4
KcVPQyvQYtyytRQfuPKKGnpeFP9kmaW4JhmpbjMLXvPRBW4FYdFwfZB+444gzdhr
AhcO70zNIdjaEZA13hfRHlMU2hxPyoe4L7YhG8XXmUaJ8JRxKfOtEmWIalJcFcR/
TfK++GXX8EIu/n9OouRP2THQ2s8aTSkXOgt3wrBsFFoD0uDfpUxEkL/GwQLr4qZ9
69Ej8EiOdaaxrf6daYjr7Gpfzg3Hf6J+I1aWc179vtyoPLiO3JsDq7p2r1gaHd05
aein/UWW/FHmqIKfwFz5IFi0URBjfhXKHmYXGB0NtzxJY2TutedLi3HDSKg3Tjvo
4zH2VZFkIL8bohmghFDC6SSHOa4r3F9z8wOP4w4L6C79LvGkEq+Gr2hYGXFoXoZC
r4VAZ5BkJ/ljpYCcbFzgRUdF4Mn/NYSbxnAh2lc4sadCaYhs4WB46q6P5UTcY0+W
lR4IwxSaswgH0rinu1fPmnRnrMWvSwAMwVPNF7FadagurQHTH/p7BzFtFZgJ69Tr
iGGjddcC6MriqnTxAX3U7p7fgb6c70BSI+lz6fSofiS4IyNvs0ZdXtazZPmGNmNi
jUF8soBpr298a943YHMWacRU5kOzNZkhMWElbaDe2Jon3n3h4aoxR1u3BVzuVqjl
a45EsdgidWiwf57ZOGpY51xkV3F9cktt3MoHOn7ainVQv+IpaY9KkF0W/Z7dP3S+
o65rb9UXZX0m2jKqJGSh5eUtIrFDOqg5ozdRI4mwRaQ/DxhbMMkKV2UYFAPHCfn1
md6IyvutdTFRcbZ1LM7hv9Z/y73ZnfE0VVoXDv3clPPaQ4fQuPmqLXwx3v/3z5np
y2I8xNyrYaC6Ze8ZAnaVT9prByV6SQUucoGJ7rL4zchRNhJpEbpI4l3Zdi+kRT3v
S2Pt3avLSxdsXQKSNirojwEfl0TzFRVlzINGUn8bT5zfe2U9kqXRMsQEX7KfKI5j
EL4+4mEYVXO0lvQbyK9iTDgLWzS2jb7G1AV+Kvks7XMx/YpcyTfC7QRhPFqaFR4c
YuCrbrNw0URCFyA3M2efFvkcGorkwzQgj/Afr5sNYmTMIZhxHX2JA1F3rvWit70l
n0SPgd5fW+CZdrbz5Ib8NqkYfB34crIHMRli8VxUiXCHab6QEOTWLrCiUB5y/eom
DlnNk75wM38c5v9ixHfsGlRU0qiYpzN9I1ablVOXDMS7rgT4dqbygjAcDpnsoy8A
plAvJN/IpZJJRL0/vscBNB6+adiVrF/jpWOdyRETyyBEjOoqUw6Kwm9jKitdblsg
TP0mj2GapvIf85u/1StqKY6ur4ZPNkyYKUCVBpt9ZzK9Zou1a7v2nCyURS4BYjKP
sccksp7q3Nwy3J4tbeYAu43PgtfdnCzHbXd5dvEpw/oTCNhZOxqp86cE/EhFxjaT
3E0OrrFvMIJrrPeT67QTRYAoMxdKsFtHDFafUlL4AUUHA7Q7u1xpqAhpYWK8K/xs
yWbw+S3EdaY/uZcTCWKIHoe7/TU9NDYPXZlXwpNc4dH2X+Oq3JSPnlGuaHxmcwA2
4cxNDedXgddkM4pu7c5xP2FNATQYlJ6DNpY+CYdPY5vKQ7SkmyTQk/zD/IyPdHm1
FO9Vv85jPJLgUFrXfzvdZENY1Mr/ia5tDQ2uG2qW1wrLSqjb23MEPzXW/sb54liN
tHn1wUBcpX3DA/cJM7MAOc1BGTg0NFfmWnakjiL7TjTAcvPGZ87Ft1pKauDJGomb
6BThjArut3MfL79Ds26stHh6y4k/9d/wVRTHaLnbZI9CON1s8IWrZZPbEuLUFHYa
4hCIm9pXuuDA+itKXM3Y/KiQrlYrD/YEwWChjHIbsuJKVI1Xayq7QlnyXCuQjUvB
AijrIOo0ZF7V/jhT+3xuZniP2GjbY4owyCTJ606YIqiEDl/tOEHGNvtZh/4h0OgA
OSgvVXqeTILg7leDu8IShXfu+L0ZHMMmfnv/uyYeYEn85r7gQ+HdLe+mzf8qF/ry
HgffKkh/AawqeH7PHIycNhRz23KT9NhOcMRCjKYg5T53NTXcgGBn6k0ugreqaGHw
GJT3+KE9GlTnr/INiNGxmdUzwbNAhMSeOzK7h0iQqHs3hHmiu6hGuo780UVEM5vZ
XzMcoMgiLpmBmVXceKdEVUCBxLvyjOvAr2QzCoEN16MGxNLHAIJhyTM+RFXNRtQB
6KfC2TskAi5d76Pya0cOr8cHvOBNx5n8VISehAuIBxr5OKQlyqsPJQDFJbEt8GGt
g3mz3NVbAESzMprJlDQVZQw7pIl+V35e6n0/3pi8VRX9oRyN37JKtbl3kfyUlnIK
Joc/9Xg9j3CgATItxD3rpBFRSBKwKJaodqWOx2d2svk6U5CipPC2bnHXRCdYbHZ7
0anCttSy/rnPOWpoeUHLBlLuKk3FCmcLpCJ+3K122mx8UaW6ZmLouT3SJ0WzhsSs
UdgvRKwOBshexGj90ydPIsQYzfIvT+H5n8+Pqi4r0dl0vdlq3hYsIj61R+RMdv9W
4Oj6XvufaLrva45oGZSRbPGwNhRbe4FqgOYqPqYOrxOO1N2DJ1x13HqP9y67/ugb
C53NBvHXxQQnMrMFyJ8RHpkIYiXPG07GXa9x0ChEME6NCKliDk0v2honIz3lxeUR
ktFLhBJMFPwPHzLtEaVKcaKtV8cyatQP68dWpURE5z8NxLED9te/prgJEQTBmyw6
ea3EfN+IzLPCLm91I1wzpSrj4QAtRChKD06sqBxULubAqE0isvUXlf1xx9IStOZW
84uc4U1BlAII9dm1oDWG1qwBb1sXhx8JR1FSr0gsEQKW46lc1im/P7Pw/08+sq6o
0Esipq45wOJ3RL8VLxxxDucDFB1PRxPviadmhlZDZR0GrADkj3i2MzEub5c1R6PQ
gj6c0oAQvdB8hc/gwwtDdW5G1d5g+KihbZFG+ieA/SWIZLs+1JblEAXqag75Zcod
Z9R5tT8YTXJrSKQu0dXkX1Zvq13HvzzhhVQkwLmBzqskh2jfitTJLwCUMUKnlvlb
le6wIuNgQs/2/XT/4ZNBHChGL2SuiDkV+Qe6nu+chbeAFP7HeTKEnJJmhQHRMmam
efu2R2g01Yf5kGsZPWukgncWRtZGOCq6zNCtF7wsi9qkqYRDJKYKvM8HIkvaqKVu
PfyQsJFWGisXkBclFhdBf/fk/TtT00qWT20eb28+REkmJvItDlzW6VOVw9zDX5pE
96Fl/krvfxuqjU9xYH90V5jzZnWtSQvn54G5zsiLpx9o3hE1O/7lHjpsF5/uu10L
B6jneEaOOYX+ZaZPTcrAbDaG+87hwsdZzr0ukdANa6SzZ8vKEuM3MMIVaoB1dNqu
XACdwT3GuAg26LTaq9b/jGuLRtorAUSigw2ULa6y2IHbImJs1/uu33i8/RgfiU8x
u3Uw7rfwiYZpjCHGXuAc/DqLYN9imdrRhJii7QeIhaTSJVZJkLNrBo+EJ4o1/VTc
01ihWtKsxAuaMnY2QxKGq0mr7DKbY0GDAshOSpe2FJX6K2UrHDnwzGihoRXcHlK/
PAnG58L10NSI7lDMFUSDz2G6e9J7QhyxxzwP3GupA8FE4/NQosmtb5tU0x930kOB
JHElnJ6tXZnYEnkb2cvz/E7d8ChuvuMKKzU5cOUMpg/z4G0lWNcV0DgoufqexR4h
P49Y92uAOcmx+5UpSXS3wnCrS+xLPwNuaRK5uZHEcLf4AjV1Rl4dTxM/MEOnZ4fz
2BH6QjTmt/wH8Pn/AZlN3JQxY0PhcKh92lyAfsypmOAR7rTjaHHZx8SO+FS8arj4
w0Z+fh1szSPlrg3AffYuJOHpWNzpAWdCM+/YeP5eN1vbaZj2IezHrMQbiN33ZGyN
oFmC2Tt6+DwrgQKpZTHqCOdRmCs7fgf4ugyAKuSFQsQVCAyvq22UolCx7f+5tuIA
pT7MBh1pq9ew31Z6rBZkH/7Jm3J8O6Dfgt3Vn+01nvOsFT+MqANjpIpXpL9sJyIb
NSeNe6I9/qZegShgJ5dTZL/Vsvq9lNih0qjM6WTjls2zi2VM6vQqGIrBs8Etpo9N
JJktsBqqJHEM23yfUNqGdMD8L53pga0afjI25WS6C7iu8oe8ZJPZ388LrrTocD1y
H2/37F9412DcnGZMw5nKhFkxRIb+EnkLk+skoRl90KcsGQc0iG5Q/pYmNFvq3+ox
pA/Y8aK074YNV2H9BXG/RTWEhvlSGfkVve+hs2VM+S7T0VKL7I2oPoNDZrJzGKEv
xO7VVBftLCKYOZVqhC2tbOh2Psg3oOjHXQhLvgyiAvvgnlJnVsto1Y2nwx1DFU9a
wZuMOsUk3sFV4tiGrJ7JL0497uCZfQfdDY/bJ8Pakxxu6gJtb+daa3vr7REkB9NR
laZ+gfCLBIC9W5EZDuh26P1dN1Qb9Y5wUlJ1U9i84brl3syJ4v0UjifeV+PzW6Mh
CvVSRueKLBxVmE29eZeftGFEb3r1qwL5Tx1I/Ueb58Z537T0uKAZaHpaSw8AHYVA
c5MP0sqWybX6F0p3HeSEWmtMDjK/55zOsbLHgD4B+P8RlhMPAfBXZxfwOCVbhhes
p2wvzxCuGz8Y4h8qHIAnj1HehpWvuo9aFHdNnhzT6jdJF8Az0gjwCIXVrCvY/h45
usHgiN7nmqZ7acPVg+ejpLS6QNsfGVh9hy8L62FT2B+hIHiupg8/Bc+pe+MHYG58
NIdcJb6O30VzlOAVoW+20obmevGOjChVsL3Ay9yFaRdY92ueHl54ctA7ExQviQ6z
Fy2fIZZUPX7pev/CWC+wn/jCtHLOBMVTkfeXveuo82KPOR4wIsDMrLeB26ew0oCG
d8iADjVUPdNiOZjnxKuYVb+M8R1gFQMh1+apYW+IAabTctPi844ZQVb1/4XNRphu
caunP+QTZnp7qAj9u+mq6cm0e7FUT7V+mhNJTaUAWtw1X1o6zybCwCIbOBEY9bhf
6ozUiQofER/+eISOM816eg555CE+PzQI/RgkueAI+CiSjSriRWXug2N+ZEBQiw9l
8ehwAFWmYGhX27y1RcTU7qOhiIddtsvWnTIuEdHAPmWPTZ75+gB6c/nt05izGf9/
6Rfx1YTweTdXv9GJEuwjMhwx7IwIC74lCuvn7SXeCZBHvG/p0/5G434ddzFXtISm
bkIA6v+r5fa0JYBJjPVIHbZ8Bfu9DjuDju5RHsSIRiPHoxW22hdDlZNY6hHKekwT
OnIQIn258neMBy7bZb9twSuGyKhOYNIauSl/ItSyWGZ45sqdzUF2la5mCIgj39R/
QM83jxHLsBtTbBxtmFkc1u5TMOAi7fIahQ8w6D/LqbBZkatNNoGBHZJfpaRgP/55
JwtIa2u27nE918PYU9sydzLz0ic4HiHzwmb2cQEGUl9A1qaO/MrVq6Y1bGP1NyaV
9BQnhDywCDDHNaxy/CQk+Zd5wufIbrMwF8YZyMRhr7qUY7wJw0CA5YIlcaGw6MMv
eo429vaKpHFb4eMMgEgLYh2K4sUAirD8AVE5jjImsyDwrMv0NRpZZarU+rz5SHUT
MF5zagy7u61F4eOKz+JezxMJwOR8c8oqghTaTKHMQvy1KJubGS+cjqbbxI4TnCdQ
xFdcIXBlgnRP1+JekVe853hUO4sbOnyWTOk7NL6hnbcYPiKvaeRXIOgzMGGyEnYP
DtSgN3+yI4b9DvvWFawlrexIfwtcq8LXfN4uiWuCy+zKtejUO3x7KOqw5UIE6abM
iUrzMmWF+wpDXI1X23HP3CEN7E2aFBOGUVufiSLg6r86I6slRPjvkvK6Z7z/ND4k
gl4YuxKneLa0aoeeeOdnlAwn3SjWTDTKRxDEetBiXVGz/3VxkTOjp2HtrTogSKqG
WCBlWMz4I70OUQK06UAl866xsrIcyZUCeeg6eV0kik26518tkVFWiJWn06u9OtDk
suun2xqMAHVpff/ki6KxjpFQ9xWhzswNlyqdm4cBfXZxqJdHrUyKla2VuILFeEhz
WxQ7fWg4Hb5G09aIcm1dgUMPIJlXwGirJlXovO0CjAQhlBKqHrG3xRaFytnYd5wL
BgV90S92ByXB5BvdKn8/91gMLsLDmHLryQjJF/vxoTceMSXE4wvP2ePgclaULea5
XpHlnI5WOf+u1Nk/n1U20smCIeLo4Td/Xq+V/szr+HznT94lNHbFTQfpYJpJG0MF
u32DHF9l6ZQmI1oebHCneuDaWm6MUppn1UOKZxUJIKJyG1T92ZpkMtzqreLl7aUn
Ibz4cZRutoLDg+xGMqSbBVJJHA+ZQdhAVUAljDIITkrzOVy2ZA07t/jEROfVfoA+
LU7ve/mRbz5vogu8WFc3rADa+hm94FV/diLtOTHEaI1LJI5v9cgSfm9R55QstfZw
4f0KXVqRo3yEbTcm4e5KTAx/FEfr7M30afGi0/ysXaR+ys+yHi0yFIKZW1El3Mcy
CVHX6r+wZVOPePQoybuLLz34daLJbJOyoVGqSpz1yqzwlrJTN3YcKpZIayXwLBzh
XgiVpqWXqoOTkKuzistjTgbbRtq16vS3RULGpH037WLI5SKYLjiG3CejA7UFEIBK
5d28W5Y4ApEM6zvBSv5VI1wKwdFzIrupwVI8xc4uWk5maz58nWBafVV+K571kH4Z
Xq9XJ0+NAiTURnqNLfvykOtLawhurGdBBLDKTZvGyPOz8EgrXcahhOgUKgb87jkc
P5rOFIHGTvhcZPBYQObMZ6SsHpm1ImK9Hdjwg8iQ2/J+Y8LmTgqNrfpuD7GG63ML
5L1j1ZBw5VSP1Do8HtOGXviKC/jF0RgrIw+ZLLGM3dJ8R9pEHz5YHgD8BBQrQ/wF
xHJVS0KLYbt1KV7KfjbZoJdwApJRh1ejYwL6WeXMKtIVxnbrn+HPzzYFcY8HboOX
tAjnyfI5IACqvkjM0ZsU1w5Nxiemp6NUR4FOrWzYQkZS33bQV9M7wxve3xibHPHv
ySIfkuTEPVDjTcI8h29ImaVE+lUs62LMPIdp+5Bma+hZ0z2ALquyDekxw13ui0VZ
+nza+1b7bH9mttn5eufY48dpLA61AexrGxmb4KW/Bf6ZRe1td7kP+SeY9VLoBdPx
/C1Vzq0LKJ2Qx+hrPa2fo6WGe/8tgfWlDPBHAqPzXoWpSx2FHhOCzNwtxxugiLV9
OSTKFZ6y75m04UGleX/+SmlYLnPjwZjCQst+1DCb9I2jAg4/bLBT4yKMM/f9zyxa
7g1mCb1Ddz3yeqdFM4Xo8/U0o7bvrr5bYk013d278NmxM7zyRgV7+ulHJqBeEhGl
wWLS1TSQvfG+49JbcH/dyUH6S+TWjZiAC0xgZm48/E3I8vjuNjKMhP2i6AN7CIDd
rAi4CPO8tparGZ9wHyfePJkKJOlHWfVhdBcxubO4z93lnBYYbyvO5k/8h/5nAOZH
gwQuW2jlgPak/CYYTdi/3iVSl/FBExNhN+Lr62xgeKZl9D6g+auUnwcqrn9GKDPJ
GUS3XYanKQLYUgfdyUJ04F9pcSFgTMUNzU2kuY7TUIPsFktT8IodA/tJYs/7tQno
fekeUAnMKYRPei8Qk7qmjxSoGWwH+5k758CZh+K2wZv06Z+lLhoSGp0IT3L0Ch9d
zkETnPKtRU5nLPPziZQGBPpDoJX26Pn0mbkmufdhbgdnmaI8AA6BDModZVG5BicB
L1jr0F993iKgcrRK7c1YmN/BleqAK8Xs/OKcvEbKBpo4abOekUon+YtDhOjhXfY7
v8Y5B/85digtRIix8+EI3kcblZKbrP5cKKspwUApNSFYxfmE3TMsEwxUQD6KcPUd
bVcuurbnJdm9yU7vJM8PEUYcqDkKfDZGfj7V+IZNhADseh84Z+C6jsdrI5xXu9NB
F+8zld12TF1I60fLyEqlkwzhK8o4zhTYaQxbLFWiCyPu4shovH+zPPGZm7oj6NhY
XYrY2IwfKTzQKHyI26zeprhvtZtY5oOLmBsLvhzu9hNnTxysbiX8opoIWTEVI3Cy
+8Rw5n+YcEFb3fvEVHpw1IoFj2rgKEOeG6NWM6oR2o1B51ZEAEENQTM0bOHpUmhj
BPvkvUB7LRPG7n2tfoFW9k6Gt5hBA7A0HbY5XeRDYoFqVZu5ntwivgCzVT8q0ut/
EY1UrVIeGvr3VFRRwWI1tMFEAMJLdsEOdRww53VIXjEIsSOXeV56nJn/bRT290WX
D0ZCNCMnbCKbfSfegEV2Q+m7MkBj4zhVpBRYfKy0fCIkX2k3YrcifnNyqWtISYN9
y8DMdunU2IohkEJ7u5IQDsQ1ouhQBanuZwRkYR7gyDOWmMEzUXw3zwj0mjvlD/60
2z9IUMiAv8tf9itfSrD96APcn41KOyOg5yViS/vB76zkS5/Lv/+hs2PwiL/38Ini
ZPmlZQpAZm1E2iVBBW2LT+TC77HtE1gEu2rKu3D1BtTJ8v0rvDZ8oHVG2RJU1I18
EKUP3ReAKxG1Bj5aMtosSBhpukAlYQRwo1shJhel5cGHFx+mJxtbBZiM57PTgKbP
Wgx1B22hTKYscZKJWHejxZdEZuVaBBqmsOJedMPM8e6fjddmRVUi4u/W30uviEnv
offseeUuX1R9oUNBxYUJRdHaZkGjetlvRuVSCu5QLrX+K59oUOO9IXZBi/koq4xd
rxfu0765zxa1uqSGvNXd2hdgwZYCmZg7Aoq9DpFPPnfXxunZs/rau2QnUxabI54J
q86qI+Pb7YggjHEId6LcUEsRZrF1tF2Pls6QabLBl1zTlypLzZMrUlvP8ZcXW9eZ
Wh+9Xdz/fU8m31SPTFX+XBIrBoG3GrQgsN+tndhDcWbW1bCA5KF+8xrDz9e01oK3
4FyEwcLnIa3evUgXplNFPOVbE5olZ/0Ozu/regivkeD0AjqBV+MIia9QQMXQEw8r
424/N/4/W9aSUXDcf3eSb49Z9OxgY4BHjecG9mwyuqBy2gREhItLVQCMfATg9wfp
cgX9IgCyp5rpsf/iMuRstknWKsr75lS8EcDOD3cyqrdLireknBXs+qILvN7HDyxY
9YRrNkr1Ulf3nK0dSzxIRLfHxRNa411hX0d/8lqI04f2dwjDAGaSvYvtpCET28k/
yiFu6Oe13QYCPEaoIx7dKs+YZS3u7BQcNh6EShOHvIkqHVxP59iN33+NRo/dyC9b
V6eN4rWOLDlHrKgXzCHqEGxcU6zshaZJ0hd1OKQylGoQ6q3RTn/4cbHinZf9GFAn
vq/0AyUYZtKmNJqed5efIF0z4AdD4xcXCqZWNhbsnYt+/B2rXJgGmwKNkfCTGCNh
AT5sNQHfRhvY+h4JIOXs63BGOOYUCVVKx+lo6AD3Z7k45bR4j+jubsHIkRt2/rzQ
e1GhscGhH2RErDCwBQ41q3pPnV6MBFuUfcIDJ4RIP5/9i/EyoOrLkasU4yymnLsN
lzr9dLj31qJRW6YAQDoW379AMsbfTXlZ5RB3Hg9vszR1wgLH7/Nnt0SyVmcX/gA+
MXsIUwr/iNl5nxzLHxBN+m38C5SA8T4v8wTdryy+WbXPMY1w3PGehWDzLVZs/0CL
Io9TFJay0ljLcirAR2oroi5F2tNIUPnPdGqxCFeQZG1Xf85esyFUY9xS0S4MNzrk
u7SoUnMQjCvgXnJvJsC4jsGehjkOCc5+73fhpnfIAfb+PlocsHYDPQxm5ciJ8D+c
PBfi+QWFWESO4MA0RHJ1LqeUHJ3xRpjIiGeUWif/2eRzMjfIEwNxJFMHVF26bmCI
mXO0aJnvylMD/yBWwTpRP1f66zPLFwODVhlXAyjETHcPZ7sre6wnSIgPfY7KE9CX
3jwTWsm0ISGLdjJPYNIpmpfUES5ftQx11b2og7CdbFHjYoY9KPm+ASqc6bpxeRnL
8mk4FMlFh0EwfLJcFymOGdeksvxWv+HBt3eU2qJU5Nic0+zqhKul7mi6Sd2Jj1sW
MWYB78KLALetKCpKEQqvOAbW+XNtHocEnLXDbUdJsKqfR1ZC4hybNpr2IAuUQInU
/K6jU1JL11aPSjWqOEbXnDzoazJAdBzuknDw9vnWU6BZkgD8oH/a2MN+6CyHxNk2
0VRpUC1bpL4sJKr/k5QUq/tVXsk0kST7QHN2h+M+vGvKsAcbnDKfcyHzenHnAGkT
IHzxHrFFxObFUYKyDhkw80aGNIDbXXJSE3Ifyu60BuwH8CNI4/MSIGU46hgAC01a
GQdiYpcPabLXRztIjcjlahq44EpnL27p+mz5i2wDDi3m4GRpkQQHfR43sKw1LOR1
UZ7D9LPxPne2h2WpRadjOnJ13LTdXEIHcwGVvVIXsc4UvK/mFfS9NhVO+3DhU8Cd
BnoZdftCt6m4yf6w1smqVYSQ12njaTDfYPGWGksIR3auhkEYEwxaUq8jI/CQnF9i
cN1uK8OtY0idpfWDcZPvcFFShDmbghVfVhP5yqnhYp/phEBp9e8P76wtp46Ao/0q
H6JFyZOV9XocJZPUfvzHZP9PkJgD9fYlYaQx7kxmWIwqJ2vR0S+VWGFBVY+bFyea
aHJstJP3DSczpkA9fo9ZaDDDm3sn5nk6Uh6KyY8DPekdbopBKOvn86y+tjmGKt3/
3QrvdOA1qxWyO10wLP8GsVWh5wxK/2TuYTH7ayWVtSDgD9P2bUt5pzzYlRyiptCR
fmqn+qOYRmRkJQy2kWeAJDUZElWES+YBE6P0XVVowiAoKJvyWJXFJvMa6DGo2ayO
ipNpDsINmUj2pEUEjIJf3R0GNoI4BzxbSvUev5xdSwUCWOqL9BXK6Ao9lWqVADD2
luOW47a7WONU8FO6mbBhkChV8BHZl5cGPoJ9ZtAvYq4HiY0BHQ9MjTi08RkWjvxo
zpOSmPLQaPPwW4xoU0UtzGEMipuPqA9DbvvPcg48FcjscEfDsS3yx4yVRpnkkI/I
bPNfPuMiu8uy0Oo24AFQHh8yNEy74mYZ8f7c4Usqlc2tJaSVHnT4tjmnA0UWCVe5
NJ54BL5exQr7uECxsAn/cwEZfQT9kgvhCmhoZ1TFp0itEN7iHz5aoL6ayUOKp400
R4ppaQnB5oGu/qLOXVx59xmrd93ShgmILJfPVKBUaAGhbTlTSvravoMnqJ8VFMUy
l1R69I9xffPRX/7dbE+rRcdIKU71FLDH8meu2/SSARsJHtxfs2iM60tu1C9zqv+c
JNahOsu+9qVR+gQ629wW27Npj/JGotBsBdn4KABpbZHNY3yUpHTKeeDsiCSRZi0F
yo/01rFAWn78x80OMqLMXI6PD9l00aXsPc2fzcXPtXw6trOURiGDHJY4fCMdhofg
xRxnN13Ek1dwc1TAvPjIlpV9zSo9oRX7eayC8ciwwtEbqy9AU3w1A8B5o1QmQnzy
QBWulzqrMXKZOZNyFbNW6PNo4sMHDXDtFu3PMtHCIl20yw7QqKuhlu2TNw+LP4ss
0KTMc5srgameY6neVRuMptvbwle1u6cXMcVhbIpz7i8kGdr3B7qSc+HiNxeLnAf4
Agd6vyoPV1oy4FEWxnu1YwPyiMR9T3PdR7RHF4qBL3rvQnsFMLMPzWKDApiq30vf
UC4aDBU3VT1yDip2xJlEhFPcpC/mLnQRYD7mc540VN+aGtlcScNwdO4xBL55I+Hw
Ri7+f/xXUeAoNSI9B/h2uBwrbwRLbZoQq5Tpli8gt8lM5I/LFawn2ylOjhEdZ0Tq
rf1OjNgdUHWlZcnyLUr7mO+A9F1LKtqqn+3rYI87T8492PwUdaAqHNaSI+b2G7/E
vC+jbXj0+iwLbCflMbikp5YF3rEdcI6jc9iKKYRmtD2paqRFqx1bMNgDBpg3VLKt
/wedlvxhEwk4T0cL2DWeOw7/s62l59iceY2qfpZxL1U/1Zd4Pj18StGRIUESb5kX
+guzXLg5lLN54KJGeui5vJ0RIsFRNtuSTPwdGRWT6amydbpN0El4cs9w0Wleeda7
RfNGoKS4pfJ1YxY4RC/480dLI0D0Gb38uZoOZP8aXJZNxrfWSesMwdUlZldItWk9
pwbHzCXjtWB9yXQtDE2v6f8ohnxwx+dZ4Zh7HEfgCz15nuUOoqu2b+VyPJlG/7+R
TsymkXjjFGUNfM2IKRaMC4CsYPSJl1gnEdYJuq+JBVS/vqgVQ450dkvdqTyA11yS
+OUcyWAzezI4aULT3Gg+Zs1kU9CY+dr83eF9LizhZ2DSEdVhEJbC2eWpganv5oYN
RVBtehvnKchyTsuCamWWagU1Cyh3rwTdPJxb9AVbVkvZPnstBaLvVNhsaLKjj0kS
TAUeVW6E5MAzpPAQ5gezuIHIddm49R/9rk5M3Vf+cI3ivewrgL4NtXTUb4nCF0BW
cDrnFKFN8xxnFOo+Qmhb2zCt7/AMksPNJGM55OiCvqRkJbWIBfNbV1m8W46rZiiY
J65ysos/+DkPvkeaiUZNgk8lJG8H18b0EdOSha0sUP+MSF5dwE0KtB3S8XFWLWRE
A5C2a2pCFdX5m5tjU1ffd+zBXrVTZ/R3GOPxlI3mjEi5Du4qYqzcs5HzTdQMFRWS
7sg69YJP+Yw6qk6UD3znkSe4JRRb/te92pvAdekiwaNTE0qPwYU6+kGokvflFsmX
jYKE162ZstOSscApJTeTQTmUmZ1clPmEkJR94sODYsMhi7GiHFSZO0Xh7mgWpM60
ph1FUoLQoIlaZcW6TPsYFtAijC37FLBxhmvisCQXvSTh+/y+B5x1IR8uwj4o765j
1J9WoLNPW6s/oeJxcPmDIR9h8IepfML3ylUCLNw45t4wfiDYsOwoUh+FX5VfpEWT
MmvfiX7m/4d2GNEFQtNGOojXe8VSrcOQFCXN6JWNwqNhk0qt221qPfqF5J7VKEVa
Gxm7LypWQL1mwzA4/ArgFKqtHej8/TlZYq77HM1D5uN15pOgN6r9A7Yd0GRCPTdX
FgKT5Y6MUHHNZDNIzAsqBwBTArXGTBRPF/A5NNKsr0ZzWdYJItAVzZRs0zivRNTq
Imk7DWQ3N494BRRkhODHEX13n3kjrnkR13NexdgWKTwatqaZHjpuSdm1Iz+GKqJJ
ncFdL4khWxvMTG832FePj64A7dy+wIX7ZFksCQbwx39g7z8nV3rjcaKvrMOJfsBh
+a4NoCFSNxo9TG9ZFLWmrZtGSgYg1f/qyB3vUWwLpjCr70dJAMiLapDw2gVl2ODs
mKdGPD9ExkoVkOJ3yCO1I+MEeerfrZaNNwCEEAspjnf21jXwlpJs9TBdo2cJex0U
Dy6nKmOCNUL1cfDavz9zD2bjKY0cYOVOzyOmGiBc7BoOq44DzfOfI9mIZU273gxX
HypyqrytORErJUk4QCjfT/j5CAZcIPa6tIR9UtDu1vOOiuhsy1Xwiq0Hk2UfCdRg
RfVpIoYPUVQcu9Gy61fKW4OA40xBK8q0iqlsAxtEVoABs8W+dVfExjdrF9+MdHPf
WQikb2QepeMsu0Kx8Xbzm86QNNdp3J8NQJo6H36FfYgSevtIUa0taMA6U7esxIWl
A7tRuh5BCQwhr3A3KJlhqhJJDNTmNvETFDPSsAJMJjCu4vSD0OAS6hc3H+ZKt+B/
G5OvTVb9zAP7QiLCoEmi7RBhf+vAZB1FazOy4fr2n5s92iP6DMtQXWrnbUVscPQV
VUQKHXhAtymzoVkMIGp4nVCW9HDdtY4PPZTOmSb5lEeZ/YeyPDpHp3AphrXq4fuL
2N9PcRTvJ2Y4uJCpM3iBkRdsloOiRu8Syw0gEtNG2AJlOZZ0f9wH7BwS9yj9Wz3v
Eo7thhT87exWT4x7m6Gj7NVPu2tcdxfvH6OFkprbgjkTqQWP5t66TpQd2o5/ZEu/
/dkMsWZU3Rani52wy0KacOBobv9uO9M1W+zSUyBPqmVYNyV6oiYgON8kWnRMkmyt
e+lc2CdgOarf5uUv7O5V/rKdsUa2kTJPqJSKMJVbRwCBxm/n6XSp0AcsphfrvkxN
WmDdGG7z/nkalNUE9hxGdseXOLHryZ1N8pjoeMBs6FODCxqQWuRcjnSfgnlAS5IB
BQBU56JAbwJJneBqVMhwcN/2dxeSY+9JX5x7Okek21pJcDxlKjylGgwep17kolog
6m/EJUjDPMyaIRo9sphHBflmzOJ1diOdN0R1FE6Jfy6kxct4QMsP/ZaIWs+9pKpo
An2RZ8qTm4Q9rCcGFD2dVtvbZJr6EMjPx1ZkTMiEGejOctswXnDjuM2K9H9ihdOC
CfwjyCbsKlBF8ID7unp4zdwee+6WhqOWXXdVkFI1OyVqm5SusnLAX8nRCR95klI2
CKtiVBSqYfIHZi8l8FQyBmlt2bbR4OKCA4GA6Y/eHDJEjPonBD+5uB6s9YDxG6bT
XuYrEladUYsyv4SsNAcwl7Dd/VwbNVFtN15yAN/kuGMJQWejQNFQuGwmXWpHQKge
IYZl5uj1PL4+kFX99ueCgRgaVmNjS8oeqwXXXOHMXYY4EndlWP/4GU41VElxshD5
plShxf3A70poNPPumlXivbGw6UYiokhIKES2NQcCOt7Vu2MGEdkJOay0wxEYW/ST
EOSQZqWIxoznBJegHP38+Yj899MzxHn/NuVI8f+QpmwTHezyXkzMCdWuhCvuukxS
60jis2KX9Q5uwervhOxQEMnjDxPyYsz68Jry9e5/QRiaH0rmUcZdROEVg+3kq+ZV
lykdpV/n9D7hKG1F0sl8aRBX6gIHJg4M+EFxp/wRT9yYMjLrGbuGn9+Rj9JYlV31
JaGpPbZc8g9Q14oPDqXcqMp09REnxcYjbZLNWRo4WSnH75w2wlSyhmfEt6mcWtOj
2puFZ+p2FNiiTE78YS/PoIKp9p5bOfjMOnGy0d9yBx4tNCp228gx/A2n9K/JP2A+
N2LWIyRtguGupqW1mXuLBhcpk37XGViNY2ITST3dCVYK+RnaDVbYozn7FQ0jOL6j
ysSA/+8qR2WBMjCVCGNEq2iu1F+OmuJ/PHWLz+AhOyCA+SzC+j6zWcuBvpWo3Wd+
3cuIKkRKFTYO38ino7+6uYEW9TNlWX5ug/TjXmNFEKHoVQxTZC/MUX2mEllKrfcx
EI/9rtcZA//cOU8eMJ2185JiUif+kIqVvW5bFykykJH860xveF4/+nlmjXdEk/H6
ND2ik7pUnh527q4N86SNjwdK1zifwaI3L+j31fBbdUVNtBGjY4gtW3Y+wvTuTES1
IcTuhxrZSyHeCS+AgVCT4CCF6/FbkTKsQ0oCZ4f0JIyzy0IjCO83B4EYkd5s7D7E
0gNSjJn+arB/JBr37mj36FxHLd4+ufkOyLyY/PtDtn8us4PfGMeJiqy2zkylYOsN
YYirRWzKOfkEscylm0kmZsveRVqxHt91e1WhBljsjp/8Cxe87Awq7cTRoqsUMH79
wPNAR5tQ15rqKY03Zs9GHZy6nQsSVC84amtNhkQvsxBPiBD8W41sz+sTVX+PGBOt
G4kSd8Fl88zkB96wv7yu/noBG4eRk6tE6w76o8G+mTlDdrpxARGaG9oanxJjZTG8
RSnQwqVVZE9XV/jhtjU6ftudJqEQPgeLjdpXg6jjxiG+AvXrQpokFfZdouSiWaEi
9hH1SGhzgxvK+hPj+HNXCmiE3/fAyu/D3FHhwVv1oe76stOU/huMo+eeZj6SlRh4
MD4tiEb2SGGSE5tfjq/71wT5Re8PsXmojO1h0rMvxxm5t7cyQlU15wLYAxCqlQYx
QSCa+DKqeWFNbeX3bTVE3/+ELlTxcXOruc1qK5ZqBVibJn9Y7TCOgM8Men3lXd4v
a7NM9Th4XUG9Un8mySJB7wJtFjROOQYZJaTHNnxPr6Jk33QKPKQ4TbX/wkINySoX
QMSMJ6k0zDZ4Inp4oJAOIlfFxXUGRjnEcv40I74PIpS3pS3ijppTsFrFSMTeLYIX
MvYeGpNsrgAC3af+I5ymFWRTXhcmCnWEFu0nW4KlZtgGh7d57hjYhjgWeqS4sIIc
3EzVI6+VfMK/mQEcMBpjQKE2Nj5aI4iT3aqI/F/ZhrCPk0Y2Fdim8kvhkg+usOOm
ikSMhxyF7soPLkBiGvRjeI8p5dN9RGQ9cMdnprTioZ0Wz9UEdHg+RTqA2JZmtyWR
amDqwaJenJugxW7qAAax8AWDeuZYZ0P4OmuowQCa7N28ACEkVBu0dQWs9qxM90nQ
uttxzM1AElL1ym+H1nu6F2KRQJpIwTogZ05nR+G8qETRyr4W6pKSIcLASnW79Yf8
BDp+L5CgLdzvX9KTOHa2hKEHP9mQEi8ZGxDLIueeX7hQQRVoroSqYt0JzUzSP7SB
MTOK2DGHTUVxIMqai8buNH8xK8/5B+AYdcUf2iUwf7iZrc5mS3piKtDr1PHkKxgo
dVe39yYPO8W9j2ufFuGUd2hTK02BCTauIENb512OYQtKrfM3VZbl+Qy/KckOAS0I
MQ2ol+6GxtiQ+5RvKQUujN4oGJSmppKDjeNtYzB9vdbr/cCNlUjeG9N5YE8Q2JMM
m7pVMlziDOamKyTwUZBsYWaNA0eiaQMT9e4fyEH5C6d3Nb1CZ6YtwThedpzWb0jK
yr38hbyVC2JzHwpafLM/TyxpSAn2Ld8X8m1wfGoXjrN17RJXfg2EnaYqd6Cy2gc2
ia2bDL4AJTSmARJnpARTfn28s1zZ+9gm73cRnhqeuneV5qA/+Nwu4eaR2JkpNoK/
dtxlmSocJ09NFCT8hmeDyaR7WUr8c8lSs0GvT8SAPSIr39ENAiD14+d+49aroYvJ
tzGbLsPKQOwlbQJ7S6/AnUHRuiZ7/eqtkDv12WmsHbxAiU1SDq8eCfO3EQNVxl2o
tXeeqb7lcPOyC2XdU83TM9XiAuV8bUg3BqQrh2pxIUW+IPuDzC76K2oIlHQ+prH9
e5BokRrQwhaaTvWRfkEggPQsT48Xe/6KONJcMuVf/T/buZ8QKH0tHTubahdTp5/W
pQPGOXK7NbNdCvE3FQttHWZKdULx9RGZSVlPYEUIPOT0Cz5YtEsVcrQ3r2Atgfj5
mt1CNGUyFD4icOIPC22pyf3HKQrNFaaen3KeNyggimBP/n10WppZS7O19qrK1RGb
bhjb6GcZrt5k3DODTT901XmQKu/6A4Gmlrx9v+G2ctEmNdN1pEied+wfa1tErx7z
JKogpBsCpW9JonJM5TEjV57+qPf0IbJddgoFKWwdyhu5f4UKZ5jQ1IJI9gGv0pC4
Kplc1HSRDmip6mK9UeiMUoUQsP1un3l+ALFOXWuqM6PDdlVyHndRBBXdRjozhBPq
0Skd6SWj1hGnsLmO29THpXo0YV1p+hDFa3JwP/aIhonFEbSXFsWrSKnqNpNgZKyt
PGs1RR/CiJxULogGQADFT2yhNksjGUEqsrrkdxx4D03d2Qb57/O/Bns3wUsIJoJK
qr3L63Swdom9jsQ7fsNGxOIE9RR8b/eBbotTTkAbKni4az2SVrA2ueWMpo9KGWoh
vODVz+tVQkUeqc9eFQ0VGNHge+932FKGvTehS2P6W0IeUPFQ+dN9TGwxuwHa88EZ
1VeJpyuiPIJ5Ghcmix9I8sv6IbnSyeyzLjJGTwQIimlBdGA766Fu9uT9/FWd/Dtk
LeGcbJmomrvoIg63oCphLLNT9F19FiAfAnAo7a9vPQuKFTUvxj5ohtj5g0I9pkeH
848b/hDjOjasNFBa1qxyfKNNq6okoX2bR1IuUp9p3ZQBNv0yl8sCCEFMR4Visq84
J6gCg4XIg4NKYdeUX8sBk9DlG6XYaU+otPMzsRmdqcive2RQQsRFTElp1htq1maz
Eqz1T0hQINS8fsPtxZ7v28UsbNjy6wOiN9DHfB++OqIHNtoODMdSWd3wvVp6QCXg
5TF8j2pXRBfjSXkikgxQxFsZbd4sPXz95fBNt0QQNVU2x+sgVhAFLHwS8bC47rnk
SXyJC8bZ69aUEcCs7RI8mOAEQrbgjUPPrhg0pcd0kGVKwDXgUB/r16VzWyULgUJY
Ko1n0UojNKqtWvt4kqaWOQlE3AHbnxDztdoAeF0iTwkKkDRwRDVz4WHMJhdrst6H
CEDCMM8QOgvCly9JPSZAO61zUMqwAV3v2a/VsCUckZZ7HXxHHmOp7hIY/wf5hPsd
QMdlzEAjVY7BLFEmnjTuhHX2j8DFOajN8+GgGzuPQLra04SEbUMV5a8521aKOfVe
s6NJ/amDLBDdp0h3uFHgKhVwjNoJAktRyFHhI7WyMx3GnI8dMPeEnZUkG7e20BUj
tY6wUN1dPvgI9F959/1QWEprrn4Qw+wfQLHY98/1py7axlUFNzhusgyDJAwPXv5u
HSaJWu1EgTfM83Q69zcL8g==
`pragma protect end_protected
