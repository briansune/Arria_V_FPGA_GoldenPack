// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:21:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZoJjB7LJQxlln/isIDimVNfxkgpRIaSAAx/zVOZtJqmNmJyydeNVD8zxH7LVg0lc
VO4UEWKLkPAb20XVa6RWzREJIP6mjHwQefeZSfVGjGlxIgwj/Aonit2QPYvksuaU
RA6Fj9KpASxDNViAat2nNx1xXYLz49GNYbsLQHgpsvc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8960)
zGR3N1ebUV+hvJOlOj1chTMorKyYH/X/zeoJ0gjQu4FRiLmjl8ftMe1DFvjZnSWl
AlBk8FwVmFHKeoeLJIAOUOjqfRr28TxXmq3sFs8H1eY7ZQ5QbBEcMaILtVZcK3GR
FSV0LqJAq8oHzq1LjCcIQpJBKZQJ+tuQX2niTJpUSB+EoRgsRjAKBcnv3d0C8MYm
P8YBJODIAAGHfN/KqSOoPF+PudYPBleHOsPbGvMLNCpsZRYpOh9JxHtK1qx46dCn
hNduKNZZCER1MtXtBHLq3AYLJ/9jscmyzWw9THjkqIdLwWauandgNL3AkZj2zzYI
Xb1oopb7eH6HOxhfsBY7EOHp5wf+FDPY9qlV4dK5L3BzKvhKkwxuAkIUM5yhgqxf
Hwl7g+r/y26f1ux3PW5m0uIbpKveXl20IX2AWpR3GgSE6/XPWzgp90Ndu3h5PfXc
3NigsmhIJ47D2JYrSDQiOaEXLCIRLzxvq9YQ+6FZP2pHPWvDuWBGDSWVJ20gD7nM
f50jawpTS1tnRHz8X7e5Haq8tJ911evI8/KzqMIyMimUXR1kzC3zW09qFCzbACC+
FklA6JBA8jcqnxjJCzAyg6XMhbYlVLYgNHEkS6qQRkNPF3yIaPUkE112flz0VM5i
VCn+4FQvqOzVET8YSNenj6YDg3M3j6sY82ErzFjVxpA6jb8PwltDh7I2ukjo8p3L
1B0288yNwG1M655Tf5lVlCiK4LFnIweOhVOMEsSL6pgPe7eycbRtgC2AcP1tKsnF
S8DJjfaHdxbgWFtMlZ/A9ylpnXMs/HEwyniSZxOTitlV7beUDYEVeZbu0NcikEUD
XV4Fp2SzLnbhnEBDophW/0NQimE7SaiM314mKIjywEvoSqBYo8BfvFRB+1XFsruL
jkhIuYKe/skXpr0HfdPFVmR4MsYxQaQuubFgmq8ZtipspaoTvBeLPfox4Wg/jEMX
N5LQH+ubv0XjWtiYmsewsTNo+MDhLDf9/HMr05RYLmLp+FCb/TO43fn+MWrgS5F1
/Q0VJ/T/sLCfx0kSluPXK0eoFzJ01RtritkIdv77nHmfxdQjnxs/dUT3xu6IN8C4
Ekr/uWCHNOpto7lkCbwskDq5NPVo4Pq4Y4lmg2mZ+mvJZzuk+JcW+/moyVLmNKZe
Ntw24Bgk740MjQdG8/5iB54zL7ypd4WkADRlYyyAsLgos/erRxOM6KMcegMfvWwq
RjkShF7IFwZfS1UzqDfQcBn2VZjxNyVXPU010JjTXcP9D7UN0Z27Glab4CGk8Lsb
PKRrObSsCcCEVWx96jnE5PJPhk8H7AtG4jlK4bDyXYbycDdkOgSRbp8vhm+HcwID
MJNULEfcNuz5q6+M6442R7nDKklWxv2aAMpQZ3DyBrs1iSy0rp2J0w7TskThNBvh
zetSUPAja8FqEVINBpMUOmZIF6DA+x0Pmam8zk1nCIHHQsE6W/U8n/3Ldnm04pwU
TNsJdlRb4SBO9F+dzI/NO1UskgFnmP8mkQQmsQy6vbSC/YBUDx8aFQklV4/6kruu
H5Wq8tYIG4nunEUi3bl2QaAEMwqcjKD99cjH3iEwN0pR+RWhlqiJLXBFGZoxiGc3
hEC87I+tW4/w3ko7Il2qVSaxEvUjO0d9WFjUL5s7jODs1qG1+7CUbDwUS7SXtLl2
2cibMF7j1DnB0IqOBB0bZ8xzPn9e6M/Og1wPlKW61M28AtfTppb39usYgzVKEatr
y8dFFTN2pegGCBgpN9lNFKNwX4LieBo/LyRdyAfDUObl16oitu+4pT7UEHFP7NtM
k+c6QaAgkULN49fuGYKjiUZxVLxh2t5FgNhiEcWKWQRAH6OtZCuEzEWb7q+52JkI
KkFZ67X2w3THNv84JzcgkgfJdEmLFi6pjoQoIZQpzgToFXEDpYcfiTeuN54l/V+F
O1c4po58LpKeDcqPE0Z/kbGfRhiT/bpeU8WFWevI0MPFAG0PseLw+F7CM2Ho1e2N
E5UXUYC5sC8LjPnd3lkTCHqKOWFND62YK/HBkKt0QFMo/zDnV7FrMWY9EhrB5Xyk
DmqGv0uIHR/4TKgiCPGZMio2dDnzh7bu4Dod6pYYYQn3ctEqr3FdNfYJF+ifrka/
Q/Yv2A1xi+qo265H5izbX16+NlQiwUk4XA6h6jXRq3B2j2bxBcBhqnTESW1e3c1A
HUDt3d3WbHo8K82UIVUZeB1HpBkxxO1UuKRGs1xofSMARNTa2qzRe0ZiM5j7tPqk
UFodjFRj+ygUMCy+TBP8NXfaHMgCJ+rWwjnYhnfY+fAbwQ7E4VW5SiUQ0Td6JUxO
HOC6qQsL37YYowpJpEEsXUDDzmUWq45qU4qIE5h2UHeIXP4IZOL36Ju6QeNeErE3
rgTTY0sDQS+weFrMnmPMjiVP7Ngvfc02JsnHqJc9qXWsxY67HOLp8fKZNu7r7l0P
afWYAlsexhmH30InEN7vLzO8x44ZUY7O2HXg4DyPKP9qpfulShWZsl9jYfTZORnC
Ypm6+kCxZQQpPCeAhILsCDd0tWC0piQd4Ul1ehmOymf3EzXigUCzz1fF+DHnufHd
9SqQX26lVlmU+FBglte8j9UABRikmfGj6chymtIi08nVfBY2xxbtT00IKRVpRCEF
ZdhL/4Z2M1bgKLZi+qDPEZj7VDoWv0oJT+/xct4RGySi1pBOkjSVWsDVaUiPvQQ5
yXoJ2Ftlb3sUFvpUlDVpGbekQfhWeA6ga78NlmSE/wLY5zIEEAG8sfUbCP+DVyd4
PecRiOHYVZur8+E1DESMUmtnrICOEOT75TuuU/GV0QAMUdhjm5HxDw02R7XB2tT6
b6knKpNQXk4WLeKvNJXSosxD9JJ66h2AbH8owimeHvefKJ+qSW68xaO3otIk7FxB
0++oezFllJw4CCCUqLT7A4Eci6eJ1b3aMsg9t460VkbISp177RlIRvrXlqw7Kazh
LT6nUj/IQb2X33LmLOJ6mc8n57HNgPRQC3ch5WRPLDPzkW7sR1a2ih1Frz6W5mzI
RP7QSd9oYdjV3xuYzPFq4X2oaKlFPIg7tfga/KjFp2WnUN1wLcmU3O5h0UQVvFWR
FSEVv4+zrMnPys6dBZuZvwksDkTZzTa7ji7ziJ8vrVelWvlMXsm/Alp8AThkhE8n
l9PewPEsYLEUVprAll4MsZ8Ry0aMCSRAeijM/iduhnFiPUXYBwJyLuNxVAejns6n
5TJVCS+AfMR/v8RT5nQdBod8vOXCsI5FZu8rQnGjhwE0ZPAqQAwL9aEAa77rD0oe
5N9ET1AJ6pEq4/3y4JSeme7NYkBdnmaT3Y7mFZUhIAbLOqMfUwq7hQqMdY7N96yq
IIIDlgyCgxVRAZtEkUy0+/xBu6qSwubW5DOh6SgVok7ADqIw8x3372s9PS6aKnbW
sBuXzmb/IyPrPpeiCXXMpATPuTz/5JUR9QOsFxKeLQu1EPmEjDODRMLyFljfuY9h
3Qc7iFsOiMhLyKH+zfwvXT2gDGBmrq4SPk9c0DCNCN6nB+Jd68B0bE62h2p1Ipl7
vCG+Zu1KwWcH4XI22n4+CdsPcuhytBI4L9BLCBCEkylZUQt5V2Ba0yxb/veywChF
h/790S7KUmpR8P+pcNS7Li8kFyNz6P7Y8553Sk/pl66MHGUyEZ1VqqmLOFdqY4dk
bXqUIRt7QHgxlJ4CdrCZS8ujcSmvcxNZbyPXZSjj/9HFsMJWSSXncB3lPoI2sLaq
aepzywu7FSiI88mWBGH5GfXbK7NQwIe4wC5pl9vLy9qNl2Q9DyiOXtW/IiWrcGnj
FIgBuwpfhEpmk3VxCL+HCpiNB5Tzuwd3ghhUlEjpkDom2v7/0SMkFfuQOGOS6wJF
YOEQQN4eZ4KqvMYmsaVFmXfsR+R7hutoewOyUftFDKYW5CxUD094VNMDTUWDfq5R
IEn8CjP948F9JYxFtAd2208ns2tlwfTLb0EgARbBBz6potLh5KlhceWjma8IeLdg
eyeSvNIExux3aQ7pfOJ7eKwotm8QzzyiXjxkEAVtwyi1/zaqB8LiRnE8NK4PHL3u
mCNV6+stgcnL1YvVImAqGjFV8auXe07lzn4qbfrmznGQaS9CymoQJnRGLPITklHP
SVFbF47rqpFH2Wpql2GDl+yRv07a0tf7m3lg8ZIE/xwl8vlYdqLi9yAGJ87qNwpI
KUHabldqpH5QYXsHB6p6TZTLblQ04lZqAGzikhjknxl1TkSnbC4e9YBefSWIlc2w
U+zZwMizZoi4VuVUECd/itJF2jiLhc8W2B/kohBTa6DugdRelhT3Sh2yCwsezuP9
LM5Uo7jICDef4hFD/+fBWOBWOgzFe226YoZroV6xsUdNCok2ZlPy+GN1bDJJ1MSp
VSDbz/JpxMfodktQn5/wZJFpmZYrYKc+AyKRHtK0N5ZgR5CfFFRekobwCVV0fdeY
/pNV3yTRk3ast416YCNe1BPWvjWBFOSkwvk+ldDeiaDOlNnw49MxRd5xE4MOnJkI
GpKWbsfCPwE5WBbppgXwYEgiAHOwKCp0noE7JODGBuY1x+fAP5qkTkDAjrvzxchV
JHylx8mcFJakDUldt3LzkINvQn6/eBgm6d8EjBaQq/UGoclhi00IQZ3sfpMYldG7
3n0k16iciVGVrezPJAXnPy3nSCyenvRNsfyk+CsifSggxK47C2cEi2ytGWBqrTkY
cZmjQ8UOo/LqMpCkHH+KGPIviSsBpVIWAdlzg4h9qrhhy8HMH3NPb2oIomwWNAub
hrHS9gKeHlTI9ezAFLqh3FGOAQgf9cXYUG8pX6EKIwvNkg3K+sn2Yyq6iJS6sE8J
r0QV6aGmzGAkPM5Wi825JxRpILm7y/FFhppxpELanoFbpAzVbN169I0S8Y69fb3Q
q4ZJ7bYcRP2R4DdmYinB0pEmMyBaksqXEshVfDz/oAtgnTHG33ilIPuckd5Pw/5r
7rsiHQkxZNwSdgSnkW4/KxP5cMc5ibQapF7lE4AMQ1Gncmm0faN9aCKrBV9DiPsX
YKKgSqrGFnJrQJUABDeGhpv6Gu0lIORPtXNGbh/q/dfHefa1J/sEXVE1J7fr4/WE
oaw+uppEBSUPUWotCr5dYj76+bHTfFX6ALuncJK170bXf/zxAAym7JGdt20JbIAy
OjP+Hvmyh0+LAwc7H6LlSNeHbKgXFfP81yX0MffLAJKpnJD7dIcMaZ7fuzClCq9H
OZJawG8ksYyamuzBmGWHQQl2fymRGW/Ft5SiYkl2NellRoI/EUzWF1YhL9FoYTW0
fv4qQbqZxacW0Z2cT8jYdyRIb8eyXdo0PDq4KYP+duxshI89Uhlf+bVM5RLy/OtB
3JuqJz9zk1S8E2YkCuvzA51jTO11P/gK/vWvTC7vVJgsSYkJ3VrbO6BBRhNNvhRs
km8XlNfU7z0tXto/9wxr8BRJAYKgAybkmAHA92OfOc/NI1WKCciMLi/B+UAoXSTe
FhsqVxfYVFodWc/Wwn0XOK3KUEa2b5EUB8+O0ypkElX5iu3iak+bGv0yBBphWKKq
05nPD1x9ie/ayDyyyL9gGhaCsMO3/9hpovIOdZVlqcmXknX8yhvWexLnN9LYf1Gg
dqK+kljHaqghaUoUW5y2KyhDJA8g8sT3Bv8c7/OVsb8v3mDchzlVp+u/BWXF1e/2
iBW3bz3FQvhOdJkrIyRxrvkYYkrEOGxGwBSu0Q5aE6cmv79X6ABzX9zfbsgVmIpb
122sAk/S1lRMofH1HzLowOuQwsRSbtHVfdQUekE91NhfIlVOzjxACBmirQ6xb8+8
MysjnZXzPDY8UXzQd+itygjR5PK7SpKnk5Q48S0QDWoKAxSLdAJ/Q63HTHpBBlqI
dxn6dMYacuPSO+u3vO/JjVMlFMJm5MRFDIidN32a5KrQtMNMFQPt4xhZ8/xB/w9v
6DAk0RR2wMCQToNxvXmOh06i581rA97Unx10ccmhZbbY9RkaLqRzDp/OGmynjcBb
J0qbd7+NlfNUhMH1qKg9QZynHSe0GN0SO9q6B+6hvcXk1jUaQHQYRFZtKtRy8Fqo
Fym6BuAC+qF6LhijSCqHX7WVyq2dk0Ppy7A4s74s3iUj6ZiSG9oFqn1Zq1MCzCLr
XOBC3YweV61EI2aE5w3j8EP1Fe1fJNIuYIpCyUv9N41nCPvnY/2s2lxJNJc2+NZV
W4rjdEUDZgDnMbofOeNMSXfqzkoC8jvqZCRqa6cmCz9T+5OVmmYVTtxNZvl0hZkC
BDPA3UuvcSGTWisnPgmTsFAlcBx1hWMcmOMOGrDFisiz2c1jKrPGODsuTwkKtV54
QY6yF2sVvJhevD1USMnn/T1GqW5Xxr8mFXCHmw7fnnRjlyO8fIAaM6KdIiqH4TPL
alpvFdAcCkAFMAdCrmsERdfVty18KhHb0vSeJsR8G79x0KblwBOEqdlrEp5MI39N
WMUkpneidPa7OtddyIVYe5KwDBUOMp2hAt6Q1yjxart1QOpMLr28laiIkwaSoZgR
z1dBxhs/h2in0ZTgPruezAeAwWQ6vCu7Zv3GoVz4rPIsXFU7MM/Uvh0YayO/8+J0
L2la1Wz2TeMHh3FdVKEvpMx+Ryc0XFzRzsln5ML+aFvR0MBM983mrm/IOspSu6iF
QPhSp8Ozu114PkdskQvIDnTu1alflzxc1RQG5rwOuA2GWJ5Ifk/wvB/SNAEfFSmF
XzpRzQneOLatO0tKfG72mYOhRCQlITx1EY9Gm67qE3FciwXJiuBJMoFpODSn8hkD
PhQNPjywjgAiFk4WwVDmNFv1zHSiQzg22K0L9y4oBr4aoPq3WApk4KDDSOmqXIvq
50OU3z3xAr+ekFQJLr3TN18wzRIW5NQK78pzEd5h3LHsLpisl0dp0+B9zc7PcaYc
srkIetPteYjLosX58GBwTUsFEhGS/EHA8aVzDA+Ke1FRL4/lZ0DskYYEMN6u7x6S
bY65IXaIe3pXdkb3J6POM3MwfPdM32kOymP0Mi+eGJX0zw4A2WbAQCEr72SwRz72
tNBEajEXNJhRmDO30amz3sAu8GZwdgQejW8o8CWAsnzjqks5kPDoBn1JMEFiDhQe
px26ipHwrORHEi3uk0uxUdokztF+uYnvaz9CC52/ybLFu9YzTieAOKces+VcYG4E
VF/haGYEPIdp0/6az84vDTFUNJAmPg0nvvv0zz1/5o6uiJYNjOAFo0srWjBQJNAZ
6KH1Ua9CzuSefH+HCMfGmW8mmbRoh1UvHlK+zpHRTM5CR6UjdC9p0yH4AHIdXaxz
m1tKxPFCrRV96ljW8MOJefDXSFEeZcaur3VrE7taQjIPQJC3+N9FRosjqZR3nmDf
DCg+oyzJO5Eukmc1StCvP9oAZikyWk3XCe2X1cZ8EUZ0wkhDk1TqI1wPEpdPgV16
uBnEFS0xap8HmUFUNQ8esa2mNopkLZYNyMclXtSYwpgFIo3vcW1+zVicoj/Sstaz
8aBODFFaMvZXoeEzArXzses6tS3Y+tmsbL7O5EERkp3E8iLLltvYZjKRmAaY16LV
2tLlthLCd+nOpWr1ugS6vILqMFXg0/jvQu2g9j2saYCjybTVQ8xrZnZGreTcOzCX
dFOYNkpRolclBmhr1hMZN0XBvDgNw8Rio1e3tKS813F7gstHW+iRxvoNMmm6J3K9
XRX2J+mPnkqK3MtvhEh1IKircQFIIe0f3SAvseVC5tYi1NMELi6aJAMxJYKp2Vg5
vgVwpXYSa06GWzKR7iEiQeYkOejiQmjq2kbwNcUQObteGYL24LrkdE7lsj95rNtS
9pbtU0UaQROtYh1h+5zQkIb4iXUR6fnJImhqsXztoMxDcdyNTn62HO6v2cMHHCLr
mlw2ff7/2CoZQFb334bWupqDa+Du7xlJwaj9qXYOqOJLatPWBsQYO3awUmQVJIql
qEfMMiZZ+3tJOzEj06+4c9YMN/5GpM9biReMrjb1wneH1lJ4jrwN4pyWsn3TMUwz
lYjgxyqP9sbIdkIULl/2qOt2vmAJDc/6ylguyoGOcr2GetSHnjTl6QeVDX5uF0hO
LJjNNn76rZpWVAiKxirf2lRh3YVit2hKixeGNQCidQez9d7yu0Kf3SoP4WFzo6wS
35HVD0BAzwdOrxAHEx4h6cMi2e6JAIJj+7gmo55EWB1aBHVSRCVJWW/EXfC6nea9
f9zUvcJa8Xpx9kGfvkuB3ieP7SciG13Kjqs5vVdkfokMNjCPXsuyDrNrmdzzXQEk
7KMQw2/ElEEA623lFuyUYxfvurjXH8hRejvOvi93xiD5Gp3cnNSS5nJ8QQfpCNHI
6Utyuc6oGMKEMcLTqH7QrjrodlHib2g8o8WX5+CW+7v0mYGUbxfPy/S9Q8uo6D+d
aDbMLd1U+FP6S5e6mBzgVTsJHr6X7VyuQ4g0vLPFUtbVCPkGoZ6vPa+b79cIn6fi
KdWJ20l4SDGlCoYiJ9YkNFQgpALIGLgMMaK23x9HFItRfQ8LclqDxn2fXQ3QLDQ9
9YnPZ2mj03IbYTGzvwYVruxilDHs9baP1ezxAmFEoOlwm815HzDZcdizmq3HawZt
9m4MQO/DZ0NA3ovOngqD982EBmfId2wPXazCqc9MEgqE6EpqEqpO1momoMLCLL8k
pqFqMhYxc1K/li+z8rCGaMJWj4JoCX1jSk/ZDmm+LFScGrcDd08fBweSMufVbsXz
L53HGLSVO93fO1RHn+c4c04mW+C6LEUeO+Sw/EfLfKJaJkFcMcS3K/jQ7P7emfJU
6feNGx49We2e5Tsegv8rthrrye0x9p3btDYlFBB2qwoG02wEA2VURfowlKBYwP9Z
dPdOBcj5NnsHe62IUPrZzIpIazojMu5uSMN9MbTBfukTspWPpuYCNjD8QozTzywq
NseVkZJ3jOET3vg8APBQGrZTV0xMM8a7aFB2RA4bB/IS4YFfj5x2lRFDJoNLaN7L
AP+6jFY/8817Y5zmUzBh9rQ4gPuUhMbXMre/V6DfFjGaPR3c5BBtA54gM9MvWvXh
9BBBLANKx+hwsB4gp8h0GSwI3+az38piO+6u0FKKIGOPLCk2GGwlADdDarXgLxGU
szxJv6uGh1KFt8CxCq+NW8rAaMB3W668+bGTvoLrgOMdbY3J5XrZL0xBZ6frt20a
8vknMjtWAFfV6CQRmkxqg3SE6kBO/bM9Zg8H2EfwURB4Ql2Mv9WoDplaRmbYtHKc
KGEd/VEFTsCIye9lEjL35cZ8cG5FSkWdIE53tt6sYXW6gERdYtWhgEWRIt2LF7ye
jd/FP4k6MAvHdsoIcb0Bh7pZ6ar72kqCe4WPnRUk79EWTBAvwcWmwtnxj2cBT0LT
17ItcO6mqn6LhPLkvWdGuAzJazirgWIhfv1W5voggs7074GgRom3CAK24xJTIxN0
3zIXT/qn1VqCs4R0jV1gKEXNwRVRKCdmNGXNUQwCxvinqTYmnwrfC8uZd6OSo6Z0
NcsBuz2f8HBTRfQgpjgYf/rVspfKGAxwB9da/MQkuMTkN8+u8GNshJAIpZVlzac0
tHsRUSF50lTcxblLGfmouR3Z5j9Mpt4btEd+inllwXLp2ar8qGEG1hKJK2cDlZsH
KlNsmCXBsnKBmoM/7d+OZdb1dRHoXKi9fU8FCkwGpDvHDupyCSFhZIm1/8vp4zUZ
yNZxA/V3PLy+NuRyNZCK2i8Krvb5/eaVJRjp03Xj7LiLfsoLBc5FTdJYw14TgHhz
AVj2PYasxS+1MKnhQRVCNmru5wEInfwLxedfKr/cLHt2GkaE4rbJx76J8bKgiG5g
vAjouQVRRR0gWKOgboqBjwE3bpBpMtBAuC1938HYXuVSNUa+i9cy+iCaT9Jv2EVb
WoH/UeXnXvFlUrvRV0B8Zi+JfiREH6C7WYuhb5zOVQTmRai3KtNXBHBL+qZ6O10s
bwxi6vWpS4U1SWU6BPIVExYHnBh38P2wrSzg0ftNiSOOmxpvG4Q+AHF+xZeclR4E
ydy0yoQ+Ud4maMa/fmRvZVZq+VmcOK1TWYN1I+74BwSNcJoVKtds8xMgHwQX39g2
qsNQkXs1To5rDbhM0rxTm7ARxgDw7JftV2taAN1QrDCg1dnsmt/+uAIBmgpot4Rq
7Su9d5UVCN53kpObXegn/JwLycSeSLcVo0Dup7PLrxdXzDKggNnjaZppzb7MJtqw
gkkUY7foWxIQN76qbmmiozWiaU/VKUuTKvweaYdRrVZIeIfbkjS/rajrLQwL4kLC
FaUu3v/TyCTNeux+EvaWj3w1fL1GC2ZSRJELK6mz5PVkZCKxNiFyfPWSNLn/TEW1
riT++OXmxkKFa97y1QGBJCWYIpmmwOIbCeEAZZKSMjZW86XYC92BpaVLypDRdPXu
7YWVBJor9sdJ/o04/XJReqOCe2lTLpYuhv8Tt9eRvR9gIXro+zvMw7DIr5k/9cY9
ynh5tfF8wp25I5bgtR9jW3w1i3ikG1rn94sxlsP+ZY6BcpdiRlSu/uAzNP2YJZk1
05ZA06MqJf1tsENiS1ici4ZopNETl+IXzPpToTHOipEgeQlHXjMZjbmH7cSlFarm
rIVo/3cBzlaFGsPXzD8aEgBWNAtUusB/1uv8JO787C9MOv35pil1vbKKJLoBgztP
N4iw42S6yfnstPLqD7Rqc6qiUssISO8lDd2oJ0Rh8UdKnVEPc1adxMlPHE68BNz1
a2ZavLaTGtuXx8HAFhsX0tIRczlfuHxcm0MBEpGAJVw/gRat221suT29ml+SNyzg
NBPcTEL1ZChWh+kN2tBxgIpwRO4fbYxVZRNLpAIQq5YdgEblTDSp4ShrLbyNroN1
/urBNXkYwaymSpEIxT2bWBsip+9RP9emhVAlEZIZoCTlu3NTO3c5uGv+UIzSmdiU
DxuD5rAEBqOx7Ov0O1zJndTxC7Nkv0e4/iv2OMwdSMpWCydpBH50CH6QbAUH39UL
FuU1o4p+ogrXBWy1ErKvYIqKMC0NnttHaXEkU6BrtGOrKJS8oA8WFDjaeOvBAsPp
joZmIMR44abyMskG2Ah6rAjpAWSj87Tpu+vOyIvxb+7j1fm1kfMWR8FKlg1jOkY2
nqv54D5vFYPYbEtEhgl4Ppk9A96hjm4thqSfsz7fu9MgDJQ6YMB9tryQiMoNgb1k
A0I8cBaVAEkPbjh+IeBILRK9rOdWnNOc+JTsUgheAeLE1erzZzqjEwq9vJOxJ+8H
85cPCQdn7KuyA9Q5g91JdU3Ld70XaOTewWNLWsKf9k4Wn1fc+qa4P2480hjzvakj
VyatYxlAb2GI+n3CGPmerE3hS1hgcQLO6rbOViH7FxD/MBE9lDVwNp1eJdfKswSI
EoFB12BbkArsBdQb+XQgC7rL3OS9asLqiuBgBH5frbMf9+S5ubO9fG8dnDJskTYM
a9GocsN0rpUmunw+ew8LT0vgTUdzQpWY6mnxMrQHJSCA+I3kBfo5UA1tfrjI0+NF
ZqsBODU2iSIqquod1SV1eeXBkEmkHfwmn5FwLKqzPu77I71PtidcuzjUnIsleCxA
jhHhsXShhtYDlDJ9cwxUxC7fS87bIDoYEfloJyL5c7yKpdUGUlYNQYy6Mt4Nn40y
hw2o8rHQrcP0JOB7xhrjdm8aE9eS7a3xSI7M4uOS3bbWpzIBFgpiwhMe8hg5Zw3b
GBWZbejIHFvbcpaBFNJGo/s3yomQdBfNQLMZYG9zbr+DJFIWlBXyrzapJH70NdXM
Nw0uZfpaM+rGWjdzD7JU3dEGKMYEOFQ8Q3xx6neFDHga4nTojmmVj9WWRxqK/6Vy
AXTGZ3felGu17BE9AFjYB8L2xhlHeyUyYLGJ7758bClJr78Z54xT2OdFF1UW2GXN
PjeOyKBNSWImAzdqRKIWc/JEoTnccPexN5fUIjhMGiqVekWDTZWZyz7ID863PyV2
7y6MOfJmCG9kM5EdcE9GD9vsvgxQjK57h8Uimv7BA6EBkNCbPRAmSBZUiufideuJ
X0HW90N1yjnhFriuFBxw4QdHN12xG4d499HJJWlGNVA=
`pragma protect end_protected
