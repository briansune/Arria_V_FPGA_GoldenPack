// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:25:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F2ZkLrvOcl72gESdD6O6ssP2uvR1PKYRGjUGJ4ciqZLDFB6knAzGEMrW6XlW8F0B
JvRxGXCDqjoGIuutXQrJhdF2uczGZI2luIGBhcYFXKayXQ8VHAkt20gfGc6lI8FI
5Cdtgl/fSLcW7IRSW8xFL8XoJcS744l/Avsn1haJSb4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26400)
uJeTZ+dB4KKgp8Jw5HNXjZp4jFElOLzeRRwRPEACatxjUUaN6nKu8vIz1E6F9Nis
M3WKk4qJUFiGOPKz6qKk8uAk+9qqmJYpZjBlnKD/Zm53sQyWBxBw9K9MmlZ6GQHD
9tD3mA6wB0pLmZSEm/rTri/JzlRXiyo6aD+o1vnk7Lk+IvrVkttKZyyyDk6OPIJx
XXZOucNJ725sNEH6IT7dL3/bF7qdUeY8vahzffwznlvtv3/nJQjIRC6bnptD1QQ1
dujiC5J4MT8TCkAPKbgIEfhn/svjFzaU+Ma9pnYNi++rnQ2WNlf50d9UiBJVKGQS
slHVdjiwucFOHYHp7JR0MshHuhqUrbofMLHR0/HzyE4wWHq19M1A+JJKuZTrN3er
xkg5ikit7OO2pe0tiPvBxV+N4D05vWMyyl0yz+zMkN6PYreY8i8ogXu8qI6j6jSb
/rPj2qN6/Ow7R7nMA589m56JJwueyWWR174wbeSMX5Z4qyrrVJZiNIwjqA1cTPXN
LiiH1sWyZFY5k9hiOJxdtSSeJj7rH5psE7U5bylgGLnU/qF5QdkziReFDFSttDEQ
qsgjMdVag4LPWDD2oNUWvWizryhHLs3BtJAuE6pgYlnFoiIdBj6PEIadZeFNG2Zo
s99q/r/BJKsQosSbdzZMSmcZRmQ6K3xcyRX5qIV1f035TjWDLMNejrM5Qh/zJDck
5gZzYEwn4rNQ7lha87hDLydZVxRn948lhjo67kTs+n80gvLmGEqnQhQdCqaoAsaD
zvJ9CMLKS+RXdUCtODbru7G6s839+Q0fuaFWpgN2PHBPqjAjjE/F1K3dqMlbTWzh
Kb0zCuO9qO+IBqlGtLQDFkwmMnS5HUkWGtFG8VVu9NDxluNZMS4RIt1cKoGQz6VP
J7J5F+nRg7Kt5sgP3H2VsAVW2mVjyQLD10CKOXBgnrqlVbJqO0R+3wjSO9Hh8OT3
LlK/ZYNhpSiM7UTPcgoUv8+QaEAqmT9a5cRB6MH90MsrxGrp0n+RWvwO23ERnpL/
I3tvPcGpfM2tP3ppJ7HCY5eNyUlDIBM4xA0Zk7meXxGYK8IrEvEz1l1vcqsxJcOo
h0nIhlxmMCyHODS8BPo7pX7PhbXe3v6ii5m6yyeTwaEnUAPqWUyjYYhcANwDPYqZ
WH62+Nssz0hz4bAKuRfkZdMxPaapgc3d19U0LF9f2MZ/K5jZi1XHYGLGY8SolLvn
dnovjr1un1VryelgGcUxVjS5laUvTf/EbvnupTkxszoH8RWDyql2jApz3TRKhiaS
BFIj2xf2ExdMs1KBy+X26ptGpFuAJ3UaUu31EqwGz2BXnECgwL1/hQGTvWicwkmP
ibVbIhXzbVSW1uvvHus5TdMzd6OXRq4gcv2FT8jHscZORaBaqUS5O6KGZ1lzQdb5
h+HpdWeKAvpEpWiQXcRyq3NyAG9qmqxJ/KgVdusmv+XeECkhSvnarbydbi9FLmWQ
jPNTuYZBvYAdfoIS3S8EMv/xt0yFn0ZQqYJPAS2o2RglESHLemwX1Zy0KMiPi1hf
yKqtegPrCzJ1/WeI+udNnN9s88bRDdv0x+AOwR+ImYtwKWBI9vND8QAtfywsX1Ae
MsMcsQ3l38Uuu/ijvSps0niuIAOlhtE4E+OB9a7sr/ZVTL3CTBcPzbwThs+6fUfc
iIcxk5DOZNVvPeSbqR7i+aqUoiS3Q66RgxS51m8OeY63pRIxx/TYrZAtvRwKbVf5
89yZ3DR2D8F9IHcuG8tLi0SH7VAXWHOEMGprwN8h384rqaitvwel0+RUzNwqGtsr
p05WGFmx/xX1BvWaXifT/vuSEvw2+UmLkcy8UwEy+LduccUYv92N8Fi81BqNO4iF
eOV8du//jugpelQa1gf2OZXFXqTTd7wxQiuiPnERkxGy95OE1IZ832HMMrnFoEtK
F6zEBBb00oVKrbipp+GYGXBzYUH2KdJAiepJLwHq17/Gg8cT+UMFMFUOG9SvLpJf
4N2gBnnWqGjI8abyOjXSjEsZt5GgckiOSJpbn0oBwIla4TELNULKU6CMVr145Xmh
gNWmn80FFXuhLziVW031nyHCCEEu4mM2pfjJBi7Bhr9TxVp0uYlPjVdgTqLoJ6gj
H5AL6qF/iFsW1/nYjCCQpXQka1XlVfBmDLcTIzVnLnLNxYIyRZzF1Ocj1vLCNQlB
QbN1GBIa2TJarnFVKhiOgIU/UVlVAHYBuWKZmNSWU59mY9w4vuHQzuduZ+l9Orss
jFD1zLmD2ty1P8S3L0oTxvhvL1+Vapk5abQI/BUdtMJ1s9pIJIIKgwu6TVv6ZcKI
PxZG1q5AZnO6qAnOcXsNZgukOj9JrCBylbBGdCcBENA8z2eXXXI5pnYZK7Lg0LRy
g3pTbXQ0efPqvan9Kki0LaDeLLDE0z+769gX5TK5mlKTFME7Uw0+r59ro6BgM337
Bp1DuRrvqrCHsXH21iJlOx1RvLYltoiSmWS8ofyK9Zu7qpn6psWQg0b3vKyfMNb3
cWo3FNVhdqD/sU3GEpylMWcZukF5IqxADVwpBXaUFDsbfsDnqEUclnaqtRMfYvvr
sOpLCt0FEC49l60SHeBfQ8UJv4kyKPFbFVfDdBufQJ2wL8i8NVjE7p2oq1ODSufp
qT/JzBRdJpZT2BzIr5FqvBCunmF2iDzgPFAjxlcco4oohZx6TO9mRPdL3UfzILsj
MyBj5HZNK0BtvjzZtkX0JYY/EcOcVsNuolsQjYTE2MiilcAfuuOthGu0RDjaChIl
5jNAei26bUb67LQEafdK7dx+oSH+lmJDUK34Yl0phdM2kJTL4XWLZqhbI++z9VqY
z0+ONJHtE6RSn2mQe9ZO7/zsaggtESClsytgpqYr2af7wyYgIMBNTutZhFT5Kdnu
Rq2lcH+IQqHg1sZkFJN5vhKCVc73JJ23cfwrzUoNGg7c5GNdjLcWQTMysIb7Cwnj
VvR13iFSn14O8M8Q8/WX8BbABJeURNmmt+q4kdUAz1xGrFHHJZs27pkqyFQ8IeGH
eOXKuJ4zBkv1dCwYPwnhg+e2F4X4ElfcWKe+OiRr9Zsop3JEErZ0Pg4wXoMYHMLl
yoa6NbBxR7KJi8J5G3/LC36F/043ADQGOYEB4RJhVKVi5461Q6Jg+fL8Eq4PxXr9
PqYPqsbqLl/3NxoSA4OIV5tZ5px4aEcpNGv+Ht2YEEuZIStZVegRpJB42ldf9wNI
W1J8i0l1D9YtY4okX/GpvKBv2xZQNvSVMz/CWotWAdUVBjOidRHF7OrOJPeFCodd
Y+19+H3+fk5Y3jwvZxc44KDttgqeF3VD28Cq4aU+AHWvMEBirHdHClbw/BjjQvdJ
dSkVzuOmX+xHOx5lJWIVR+dz9o5/5GlSM+T9i4B5dynD5O1HjOfsYAE/FpsSxX2P
pcjFFKtl+mhldyCR+pJmgKk0qI5MVDcQdX6fclFgb5QQcrqqYJKDbbcbMoXpaR+t
6Q16LYlWN7osV3S0IfJL2WvSFGgoshBMjthPWtpzkWONtzfbbUbTezvawIGgqKxS
zO322yJ5FCglg29jZciuU7j+NlkktznWeEQ+6Hv+/Dz0HcjXgIEmDwhDodcjDJqQ
LCd9kAW3taq1Yr0N88i3z4zME0kn/tfBxSE45e7YT2bEhpGq554NwZ31EIlW0csz
PbXzqdRV1kyCDf6jhbW3vdZ/HqZF6vh4ge2SbzHUfSGeqmcc0VpQmrjuzP8p2Ny7
2hFEFPFkxa9ko6945/eKqHaEF2X19NMtuKl970mhhxOnPARp/aoWZpUj/g+LSpmV
gSiNzcuUQrj4ZfeMOoF/z8Q8qJrPwj36hDgqzX0PmcnIFxEKKaLBot5vYDvByyyU
LsQE87ela+8BYcdBU93KcONrgcR1+DHBLQfEWZ+6/Q44hqsB3qvmJbP1Zc/9igjK
KXQesKoRtubVI8neYntEsijwFTbpl9cznhu8w+D1SGrtfxJa/zVsMX/EhLPHhYJT
GVl04KSH5t2P6VCEddj836H0rP6+laMUEBy/Z1AXkim2JIbP1YO/GFXpT8FNMos0
JWEPXs2Az+jDetSZZL7f5LjSuQAfreqTK2Q832bdPtv0547U/+Lcr7DZmjOLsZzi
FnTat56u4FV0Ajt+Qg6f2tbm2kUzP3LIzq05/LIMXpsVqW3SZaRFqczq1mtqRY7c
Jlxgz8SQ+L4zmCpyMhR2Xqi1BV8JvLzaxCC1JeaeYhK1N7f+TIWHVZ4RNJRjoEwV
YJRnYwZjmN/+xKMqLWIfCKFQsIrqO5Myt7QPGcTHP9RhcoszssJfLaw8VZhvIiqk
VDjTF+zFOL0hIG6MIh2sMjEMEw0NlOXgrqDy5Wq6CRHsu7OxYg/eom+RYMdlUKUe
/k9qcobU3Duhv22aTY9VY+3W9LMH6yvbiKq5QZ4fFqOcrrfwPYTUQLJIO79S+Gey
HEsR8bTD67qY4xgV2DYPgS1U2uGnmB/Vv/bdEUDs5WuYRcXdYA358wXNFmMt99It
O7guX+pTYQ4BtDW+qI5W5Kcbpys34caD1+VppbZxf8gZfRT5xRA2M/VjyqU4+Kyh
11S/LTTLN2nFaMMSj8qB3o1A0Ueyfxs3rfEeyikn9cMtIQ1R54RdQvcW/Hqg9kNa
Exef1wusRF80qJJnSvU5VMW29511e7LbdfdEaBdPvswugf5wt3ZqiyHfsMbyymJj
L9kvE4NZ6QxUi3tpSSpzn0NujvF7ZgU4tTRglozYWZ/Hgwlvh6y4OZp1UzPYDL/0
livuhlAVdwD4BYICCHuW9RM3ncz2kVNx7BKWN3sciJy1iNUa9iQ0/14JEEv9Rf8x
RhR3FsyZbTlaeUv3eemD2GrJgvd8wXxBVHIeqxeHeL73gkiX/5o8OrzTxBo2uvbs
Tmzsk0XzNzTW/3R9Z+UAI7jVfohdb4w7gHiH3w5R3GC/owe7qcjjDoirkYJ9nTeg
iQxlOD3Y+FZrCcP4H123veN9mgV1hYFPS0bdjBcGVSKFHjGyoywMM2UYTONmh09D
s+RKPbk6heeFwuraCZLhrPzt6S2lmXTtyHv6gqlbsNe2taZmrkWfph8976oGwpIL
2YU+sVlts1NvUNnRzv0puxxHAGM2MtSpwbbyyLOUkva9s79D3obhDMVxegEPoPmh
i5NrIm/TbXbKIadcVQanvzM7HUrQUBotirceQ2lYknxG5BA0Vbcx6psPKGv70o9c
x695lQcOhnSlS51DGrQ33Y85ygDnfzZiq64EHAkqkIlKgvPEnhSj+oKtcLdlBlJr
iZQOM8ebcw8kRjddDBlVwWiL83YTND637XDDk4PCcqKxdMBAjrrKL4upbZ+Sej/c
Qp64u1+TdhVIKG/YjWcZag+yNcKNMgIlKCdTJBPSR1Bik+kVERQrq/EHJ1hFw9bf
EpFgs4cccEoo1jpptKCF1IJRMp4kZDTvQd29vnhbvwnQeDnWvh9N7tt+bKxL7r1a
AtTMGXXwwvJsDVPPH1UAsu7cx5ynsamBxT74m8lNc/ojWCKS0vtJBPfM+GQYyubo
FQhAz4lPEj/XZRhZ9aQQKa/3pAvtzLmPc8ICCwB0ZLh40ZrBE9GYAelHOUzS5vYB
1TrpTVDJGAf4ojBCNObWjwaYteAlDsfn5i1KZAbeNC5u1NjPAeyDZL55gDIMzglW
X8XucjNj7zDMyj6L7di5X+ID6d8Np0GDb6BAn1BgAmCMWeO3jyBWRn+WcVHGo4SB
eOt6iU92OTsYWt17CbmZ18YeZfur8tAV4eOh4XFnWJ/En69Lbt44ZPJcsIsmZ/34
nXJgwrwyWj4/9bAX7Hps6KoD8YmSZD2+DG5nBTqqU0HsOU/UY0y4AgE56fJ6wz2b
6UOlUwI6t7yPR0HvhifuJfDJ39HkJF/ltnyZMswBcl6QJPgTS1w++VwvS5/ih3Lh
oZDKfnH/slmiCjKy6pqJp4uiUcoG8D4BOvWTmXmg3eY2pBzCerfk/f/6X1srNWc+
eybbRbJeuh0eawrXYM7BPEdt02mJLPt2KHqlpBVo3K7dcvqY6tMxeaK1l4WCrIQL
OKEOeHwLQVns+86m/ubeMLM3sHsRc9Wu7BHObIZuDwNS5Y/v/hR2WIcRtGYa+3Fo
tpJyJ7+QhrJ9EmFCKVAUsdodIEZe2TjRGsy4vMIEKEeNKH7ho+cRyZ6MkVhEs3gd
uM4Y5Bpa1U79ZvJA0aNqMB15LtUDF9MeULA8bXq3n8JvKonzwNxK4vScp8F81nyx
87gr1QNmpxPk5Ecr1D3o/CT3GYqp8dtHo7BoIWRGkYZqPo+iiqQXfZwy0EjSbFD8
uOBoEnLORnZKQ/90AT2lA4BOBVAR9rYw7mt4IdocWw42Uj/s2F63UzZs6youCsB/
0zmRrx2VAf6aXtbmGmSlwffx8uLIcDeo+OLAYAlWvXEO3aTgjJINmBA98Nw1qbS3
lZf7jifhWNwSkGL/CdEJls5F0PVmdMmOBtyy4qh2wZVa2gD/bf1PG3w9m3aEnfF3
pzoGjLxfYRrSYPdEH1kjRBHgcMTMKE0r/70abLJuLojrC84LEUSCPYiZ/skeORkB
CeXpPCclKGoYUJJLzHI3AOAx0mWWlqeXqtcLGp9RVNK88OlYgMbILdyy41QVc6Nr
eEo82FSsU4ecqz36kDj9pzxvoScIAN4/QgWRe94aE01dWf66OZHU6zxPRWQtgUvw
EPoN9jbeJTVfMYaiaRLtR0CxhKps2/x/WgRa2i/IjjqLhMeL7CBWpaAl2SaNnRy6
wz7EcGr3i1aUFm+OeImV3ngrgOexnMfl9ovui9e7lxKEZh4Lrn34IBq5S7GH6ENU
G7NUzR24Rn/ekVSRcLNTHH3VqOUShKXf+Gakq7j1se2LNK7IOP30p+nIOb4t8PZP
7RLFuiguiM267N00J0zriuwDvfb/Qn5knTzJpuwPAA++0T3DCyXWfx50EN5S2VE2
Tfru98lIcevArkawcP74sJsa22KgfV1wqdQz9ixrKomn5h03NiamWs/cB5CmEw41
IUgDz2SB4K0Z27r4lT7KnMHSRcxv7+dWseP2hYJCEirodag6d5S6bu/8Wm6ByNxN
tyZWN8VsvSlviwXUKYU8xsqWexSWBlJ3gW9OJ1Ejm/2UZ25yVBHwLORlm8mDJn8i
wsuRdmsiwYTUn/CnVomx2VjQ71iWppzIGSAvwVSTQzDxtZcFdQiYaGq0ojgOtWgH
F7H3frjuffwOgu6KQmi3TBrhI9fzCBhhEStmlW5JD6cmxl2FtJa8M2wX0kTRXcmC
wqPmDJ+Lcvo3ucqzocD9z/WTwkSBuSYtdfI2C0RVcgReM1pZ8sXzJ5GFBYFy9SSf
JqTZkGfyPn7VYhOIKC2bpzYIptTCWleg56OTpQ47E6e7LFs35Oqtt5WQiJziTstc
7DKsrnXRbJUpBioZo2io8LnO0r8RQcTMDDZQfmqlkl/8XMyV+xJxM+32fsvVsszM
t64vbgGxa8GQhcHWfMJZbeFYdnCWEuCQ98MBNg4c99QIQCnLJTZ9uHBNsbPGL6i9
dbgVjcnKXQ2iTd+lGJcW2dXM7J7PEpJ2FiYkOm37sEtAqX26M6WhxcSD/w1JUQm5
NONL+oY06FxIBFfj9ha/CqE43/gpe/FFKXDHzQTV3Nj5F3HPLSUpVxzZVFLedmE9
viFSR5R7ew9m2AMgrR3lVNxstOL1vXxjwxUWTr7QkKPUkpqsBhlEuKoXA7l3p3gd
NaT+OqSHFnGWl5mCc+5MbaUTMe0k6eY80ks/rpC0ABBBv2MnDM54P3y2x0pHDaNF
NObHCDCwlO1GuGo/9ecnyI3xac6J9NLkZBwxFQjm9Y9mmTTM+ucncdPOJgjlIXR0
jbpU9JyTjefAtchdjmBVGGgjUDGf3uOlD8nDRHVGufX+z1/Q34J0JtQCDAY3Ni9v
SWhI3Fhkxgp6NiW95QqRlnyJKonlm3rBFNpzFR1vMwlOJUra0UD5duMA5HZu69U0
pmR1Ka8mhoaWzkt8SuifsfzeS6e38utCcl30pt+k/Tdv44c0GcFkx98egbRJMM2w
t4Cei7agDZQgHP1nfqAVrhNdPEsuqwX6Jji76OguxGP0ZRVsk445YAoke1CHFL9B
TZEvnay2MdY0FKCiSjWw5PH/v4w3sVX6fuMnqjT+OGJv9Al0iaFp12eDL9vfWo1R
xxGXxuteczSV9oxxeJdt8yAXvkHySnG5lpv/IA/gwmvNirtawxME1+pWupoPXAWP
lhfrQpokLa4v2NNSM9W9DrebvXhDQIyx5nhPTY7tmFsDKr1elwX5MD0SABn2rjqS
NDmk4HaK7GnqJfl539Dml3iqz2XBqnTRgACqjt4EI8vuEWGhIEdnAAx1qKzRbzvD
NSukW6zDVNMLTNvgk0TpnYctmhGiOs31LjY1px5BHcd0TntHg2krTQDlbIEptMhk
OkknLM6ql6eSMiiKx0hq1NlzLcJLmdKYi+t1TJOCldtjr/9KQVAvvSLyZBzPbKEQ
XttyQQErHbasrta9xcIwNcCkYSFg8cOxCS4rkdfKqgp14fIsDrZLKAU3kbZTGmBl
2ScWbp85ZHY9Y8Xd9ogpjC0LuP8tiJ1dS+zOsXfRzND1e6mvEyiEDNGWpWWxOPKk
L9PyVYLZyW2RBHuuPbfAMLh4FFNqbB2fZYJmWinulN8W5NiI4CNgBlpEa2X7T/lI
1OKMRAOPYVwbCtK7j3c9LeusJTiZsUJO+yMwXGtc68/86vG76IX69IusvlQNIYW2
fcs4F7hdhGss+v0MgSrPjSZyab48rrvvIx7P0BrT6LbNRbWu7moGmwQ4YByva2tE
p4CF37zEKvlxupFvUjVQGdmQeowblVnahAE3UUCT6GZYA3/BSixpY0V+Xf5zAHQv
wnTwl290XcJ9OswNPvl/y9bAswXxTeqszUWwrSaTp3svdLP/tJ7EBaKI6x9N1Amz
m4TB/MohFofSEulps+j6/VWgjSjTS3vSJOYDNEm3SpzyNxaNxptt+tW1C75p77qw
O0BsNssOa0HgOL977uqXZBPArYtIulVaKgaUjIUd7v4B2RxRiLo1J0JZM1fik6AC
O13YBxrrHKdvx3UhRzcfRFgdxSFVnwMHgsp4BVwmKx0TaquSWYUs+gUSUEQ0lRk2
XomPyxYavFhROl05PGK8TyuucBXBwm6FarduH30zcA+1zOAwPCVdg35xxfkrQO62
LiG1SYfHBLd1IlHirZHe2HENZSZ2mgO+d5IDDXgrP8mTEr/mKaHCcGsA2RQBxhwG
KbdJU3JO2LeF7EPOyzOwZatr7D3mJsDG4368Un5jKAWux5DAlYrm7jJ0ys+dnGSm
ixXL2G5T4KQt3MrMLZW4XW8N2MguwXVc+P4nNsE1QtWKweD5UvmongoXogXCtbYy
cLO6uA1reYBtDcdOuOI2W4AaCjZmpk/9044s3aCfPFbkvv2W4YTWMuIiejrq0cNT
HPyoMlc6ho12kS2OgKBPbB7VLnZuxZuNfyrEb1s7Ks6gY0Wy7iwFy2N7T8GLPaHx
mBROaksR4b2T1gVVI26usMYYjqOyFTYNoWZz2z0jlZ3qIcG1Fa6zaDc5U/a2F6sN
QCeqSnGHvKXm0M0pZlQoArTjhMWeMrgdttDDUPrQkwUT/FpyyNuBwyiCvTxOZ3z4
E/ENQPdlEOwEy83oQv6RB1oNVbliGZZqT+JPiq11+LSJIRx+THSZk6DhPHKsI7S+
RX3pfyhtYpITcN8NSHS8nZBSHoY0GIwZMr9TnPYbBelsLEw+SjN5nowR/QuocR2g
NXC8Sz1sxCFZZZb15Lmygzbtnh5jDPrNWluLa5SiBEcVHvnqn6EdzaG8AyQ5dfhl
bVJ78FynOu3NGggyizactKlxAXTUTqQFnqD2k4GWU4bKpKR/MfVVY6FizidRzBo7
lVo+hxLsgIgjevDgBhNYeN8/DViZ9ld4g75XAw9NRu/vzkGVo1fyq/8kXN66P8vs
lnQj84/UVLG6dZ69dy4ipi4WctEstyTSKtj/rXGzLSejviK3qppSFyPTKdUxIMPo
aepwgkh94ZBL89Ay9joVt3R1LY3A2Wb/nmEjxfESfL7o6rcR3bANuIA5Anq8fxmA
YdIy5f9BIIUsogdNsiiaFPhqnHwO5WgRgy8bQGIWRnzRsYioESnnpLiNqcEFYL0M
GZicYcFaabySzK/DUiewE98i5UdHW3DWv09USa9K0FOFPmHmc7bvDP20rSzcApIG
jf9QN3HUHVzYeKB6UsI83gL1ZMCu4Di+7yBPRqhJsILrDnd+DcOLYHNezkz0mSwr
Sjd54zMfL9ZTS4y0u7NoE9ioURpQtW0oDU0l980QS0wE9hQTJ3ttOQ0LnQsSHIbd
apRnGg4l20iRSIhZ2ZXChofB49SeuSZAna4jAEs9nKyZEKmppiNup2Ww7UVj7bux
QpsyGVBqafXv7F5iWm0AOGA4wuKdUwKHMmygDuOlCNFzRfd/W+inZPsyWcVSBusb
i16ornAQQmzOJIYRMC65dKGcrUdrJyh4rjHaB9px2iiIiCDJJT3jLIpX9QHvq5Ha
diuM3R67wPxRLy79oy4hCIFi/t+Cq1UKmxPdcvzLPEoJ3MjFj5S75lmm/EHWOQmT
8SneycNMO6HDtlC+1YGwcLKmJ6ZAWwsTPhMb6j5VtO4b09X1Eh36+8OpdYwc+lh+
sWJJhHs22gV+5+xjWNjDMKHJ9OuJ1z4AcWA7itpoIuk3dcJZzG/V2PLmkxtoqEgg
TaK4ix1DHMRztifbRTu9U9DIEdZhp9qNIoj26w+yOquSXEM9dvp6t33K4IXJgegt
uzG54yKKWyMsEjoueyv6kdTcqL6WfYuBrS+Q/21Y5CVOJdaIQcyaXauRAlX7xEWD
E/K18BkgUfvQqYirtQCMHktZabIeIpF9WeTBZXN6LlbP/YlxFmZ4YWpipBQU8mvb
KCs9uMidUbsmnwvKjWrlWkmJE0+6PjipWUqchcJtsJhydDekJUYqkywQ+94l3GkN
HHGlgOGBGvCZiw19Qu9ezvzwTfDLgMQAu8ryNNvZTsv/5+3F7VIbBpeHJOTKKZS8
xmHznhjWZWJdCry3dvSG7kTZmYdFP+/Rc/3Hh1kGcWSpH1+KpVgmVoT9BDm0jY27
eOLFSflD5hWXtY3g37SsAxjhvOlKpA3Afm3Y35RVS3Yi76DBYhgxJHXUxrYys2rX
z9AIKbs+pCeckeDYGrrVe7F0b1QaMSzKsu/98h7c82Oo/uKoaQZf9gL/YxwAR4rC
yQh0PclalymNFqYrzQlSu9ZPpiRz9Lz1yEeNe6gMeWMQ/OPs2fMWDtmovOK+lef0
4J4fwxC8XvTbecfnZ7qH/QbpMHpqkqQA1M7C5Xhi8SRLbq6KfV1Z3jTEchR6+r7Q
RgCHFV/FoaGZoguyd85ImgW3NR9Q5Fb6cKxWVMhjf+TaA0Eczx+8/UsrPhji/4EO
1ViDbU7G4VWmzuCRz1HskzdNAzl2RW62sl2KcmJwR/O4e1gsfNlXfQMKvzI97Ktw
Q6mh3vSwJG/+RZ2sadrOzhh7IMwUUlasn1vCAczL5GO5n8hKhOg0x18Kj+/AfD0H
2QGkGvA2p2LX/elX48PD9aqjB0HAcKFOURYgFCMLjdb6Cwt+prIHSKEvFvWxZpGm
25N57o/x+qZjndwDen07htu/AwH793HrjbVO+doGvBlloT2/1t8eYuM25yI48Q9J
PrwdPb1IvtauqFym5n2rgFubshUUQtDMloU1FGtlHwH1ezzX5S+RMiDt8JiY3Hmt
7McY616qe7jSb3sAA/2rSLwHyK5BKMn5/rJKnLcKAXSVEwGOa8QHeRzBU+BV4hfQ
6wOZhLQXv1vA7qOBuSow7t+w9pAj1cGSM6BbkV6fIm7hDMWBBRT0HD7yfPhc6vJt
b/cY+xU0NqPcsqSALhEV3jT74OsR5EnhkevwM4JtbRWkxKRHrKsWXlL7U4u/Uysm
NB/Za2IrbR/I4F3S6f6rlar9tvB0cYX22PwyV2VT2OpmvrsudQGTCnTy9kxAedjl
H2EIJ7XeDEiba4a7fdzBjlcJljGu6AZORPIVyA6NcNZLSapYTMnLdrRqq32YRFna
YeWavU+UpTAFV2JUhuUvJyQFP4KrptLz53GFCZR3zLKP8afR2MreebNrQHl4U5eI
VzTut8AwQAanUNo4OagKTPAo035UGjBipbA8AnVa7+GTSYloJ5Zo2TCVmWVKaj2N
drXJ1R24RHqGiPiO4bz/b/I4RNabVIEwZH784BVDTDkcX+AUya4a40Kx5DtrjML+
xTSPjPIsvQiW3X4wFgQLJkZnN0cgJBrLuW5Fps226ipjpSynLjhdql1GwfIrjo9O
msur8dxkOrrvKReuxF8cjeZkXq769itwwiv9c7eRts7c98tKqTjWtOF9mfbSoPgS
cuV8L1siv2bjNddZ+cy7u7xmcgSNaBsSh9NQ0gM8pyeoxRyUEr5T+8mVEMSQvKDx
Geqtla4q8W9nukK6wJjsP8A5l8GB5jwy7vUcbkT8jjDi14tkKhWEw9iZIIbmvvZI
hWhcRnCeqxck+nfw9wQ5a7tFff3pVDvuCVwoz7WkZtr0Zmz/hRh7b1UlihMb0ZC6
XGmnE3ZZuGR+JD+ZqjjgDmj+FOAsj9b/x2rpXpIAz1XFBpJKfYoyeQ31PTUGACS4
2YLq/vrr9J6MlXP9i8otEMoDCWe7m18q2PL3Qt0EY8ZO2ksj29SlQKK1PLL0vt2n
kSwAAT63FwScjSF3Aku4V8TuoAhpr2XlHzutRzYyuug3N+vpOpNIcjmpZwFYaeOd
7DfjxI8n2NGKVk2MQPGg/zX2TQGR5v82lHtKL64O+b+TSyKo5/21EaMedPdwK8Yn
MySdKsmnaNj+3mdwQGQwOZEdJc1ZAjEF3gY5jGR6ozyU0+FNKb4+7pJcKaDFlDzH
7HXAynZdejjMBJDMTMNtnAUF3AatiYdyrceDOaa8sAwnLdY4FFwFwkMhxpGU8hnL
hunvVgRmf8jAEVc3IyEWsoCTBJjWPZMfPox4559OOxyN6W6ZVdX59NwPUPASZnvn
MVLTbJc9xK7Rs4VgHE+8PY/gcVM53crSMhBUWzvarNa2VUQYEPqGUHZgi+o0Eg9m
hF3TZuDvRYH2xJmc6ch78piE+ldJjtWFa3zweveqKo2FlRWWl4bQEdDnoYrAyYas
dGh5cFB358WQ+mX0QGOrKXenYFLI1lavHKGAMxU4vj1c5Hmj3siXLMgjJEkMSiST
AMImnkC3jkEJBKAV2ck7Mh/2KiUg5N0ctkSii2eFgVcNNpWTY2tjDUQReKr3bWsS
avk1dpGkFIaPG+m9bz4U2uvJhKUUKE5nhx/6VHuDQb4kRSWerKsLYI/m8/rNQq3P
4rv+QUHhI97K1UUW0xvvtjCqHoCwOcofVX83JpTEQkOjlPMstyNufaE6W7JDUUDx
bB8OQSisUvMtY++LlUmzQLJid8i0aAGeFq+sY6gHWTUhifYVlx0RMEYF6qcwVCiW
A+0c3Uf2YRTQENaq+iFLGdtldNsFQa80rv3QtTjNjz60+UHdfFAnens5WpTHl4rd
hgqjyADnhG0lZXhLD/GUYrR2cUfXRdz6DxLhumiBxa6P0ox6vtSyvzguwCtW1U+N
ufY99XC6+NsSIKR8baerol4L+l2Ykgxtdw3Y//Q+WrNMqcG1e7sNCK+w015YtQ7D
N5DFM9oC9FUSRu48N7jqXugJh6tL+c8QPU6mKibRR0nU2jRrv9xBWwBbTxef0P27
DfKBsroEmrrtXwRHnJUMPzkzKKIEQ7fU0Yy9xqn3XTGWknQRD6rzoGg1jnsS1xqL
LY55h39Ukvustl7b45JDcirMGIcKRxR0SmjPkV7rqSgIGYQ8nf34XlcLkGPSuKfw
h0d3f74fvgsRyllHbBGEEwxoPEC+Lq11GDbSmoEmpLHJoi7rx9vCQ80llmJmySha
dyaBszmBoCd4f24ZZ9ePv0c7gi+SCHZIQfde31YwHRozkF4g0PdLfN20w0UAoIqb
jeyWtv207fZmIQL7m0RUxfFRUXhCgdQRJBcnj2xHJoeKs2H1xfWsjo3c31ta1adW
hb8Jg4tlT9HjJ02imwynlhK1BWcPZ0pMxhroR5bo3ysl5mniXYgVc/ArlW5dgpZz
GKoIkxmht+qJXCuCJIeaX9zaYcSy333SmQKXJbuAvO2YKNTcq4ErNwBwmzPZsGMY
XOoYu32OUaJ04dZbA41d8wQZDWw5v5WwhLB7FEdVb6YUVlfwqqEBpUwJr20ifXTR
XWmLWWT6jtMdtprs8xNhkbdCGN3wX/VVUfCdAG492GyTA9ta1CEIy+cwH5i3R9H/
eoOmIcr0L+MjHiYoNxMn7DCGsBjx02p+yCz0t0xELHJ3PIMcI8fkmg+pFS50Bq2S
JzsFtglD8o3f8qOs9IWg82i4MjtW0QttbAC6ZmC8DOAY2Ufcj0YIRRpqMncXlZi8
5VoKtU15xTJDA3ZMlT8bVJniKFUf0Zy90u0LfpVwNYpeNXTNVAI6fo7+ae0ZeAH/
XPowIEuh4ufQF309j9QA0ALT8P9i7ii6e+7y3FzhEMbMDdMMhK56vXkjzyT2okn0
HhWwXSoK1DpquDjkEIx7CYd9lD0509opPxdKh0OMsH0wYaYzNim29ONw4Dcv6c73
fBZxybyS31UgvC7zv8y21UrILZEQoIaRtsK//D3SwulRQh7DPssy8cGZqt2/SOSu
a1Mo6iDY1sNovueiUEBM44zeSnZ1IKq/QJrfhN+SZvR/8oQaT9hZHY78qIXBdtrE
W9mfE7w62WkDa/wxfDaHzC8ePCJ5khvSKsCiPZwb13naUAhb6wpPH4m4+6ZHtmCZ
BoTK3C6tknd/C9nYYDj1N3VWS+ByWrOygsTUYuIu31OpjnHLmcZQ7LwjZysWaNa2
AhlnadLdon8++quCWwFVd6qY85lmF6O1ZFC9+a3Sqam2Pe/LxCTM48ORgfGB3Qm3
kWyBpuXaz9GikooXkHumfwOS0wIwPEonDLk+v2VPtjsWH8shJ8Gi5dDm5Qra/NqH
lVkPGXk//HClrA02o2hYcT3HS0Qdz7VBR7WyTo5PPRktYBegA3NFu2+isgxnoJ+R
X0EsVR4wC6vfeiLbjlKYUbA0zuxvFVo3SwNnu9EB80zWTZ0q3dK2QZ5FxgD2C1Sw
Gs6bVbRlFA1RlQHPSn2cnwLhjkxZjBoT2EK7p83BQb6lGTu04vroajp7/I1zclPM
dT56bLeC5QB4FCz3KyeL/ZaUZ1tAmT+PD7zwY5XvPcDNAtGC0LExcVKIdRHn+tyU
/a6svO83kQsx3USE2muy3xecRotzIfsuvwkn45sSrOtwFEZKe4jWDwV22bCuXo8N
3u0LdTVk0BjsGoXk/BK8/kPFiKPn6LdUeutxZygw2d2zd/x85ddhXBpYBFhThT9n
D/mUjMp+2HD6vlx9oaOWaBNByOaRfS2oPMYz6l3/5agy3VWSFyGByMVg89m9Gh04
kuDQtr0ekpqyzshRuaw3nChVLXsYrD/Fm5MkA69YHumtwdnUxQ0TWUDbgLHzX5/f
iD5HJB9YOWQkuPReBJoNp+14k4a+I9S3FS1Js7kBqvi5DTnxFY+GixcgTFvLxUQO
/WBqB9hxgUmp6Fhm7WLJFcG3HcPptlWid68ep1Pi2+I89USukNYzOdYDcoRFbKOL
0FElx4N89i21YCtvf09M+fUDV9zmstLZ8ghym9IEraxWONJZy8azU0i3nIspWCfS
Z33giK5bjszvsXA/gZ27rvBfGs7JjmvVD3+OkB0WLy/78DGPdbZbonPGjS708xSw
QQ85cBVLhYcl7BsIo1h6vtNiuMIR7CbXoBYTzqhWx4HkTM3+yrat5dpdWQsrEi+T
BA+EOL8uhO02rJH4u23gH6Eq+zLFx3vVBsagKNkZ+qFvLTYV2rB5sORuSeBz8XlC
oeMSfN/lHgwVf9IndEmTYVpjQY++Uf0/Z0BPWiPJ9iOEYNcVsy3oLpcMqcAfnatH
qrwdZMfPUplaqAAqMMAZt1ZkHJhL46glnwNyJaKPoZk0O8nIKbLQfAvGMhGW6sRv
Bk1FC0qvni6PlNoVpARpfI0Bup5PqR+XOmXfHklN/X21XFGOMoL5z70RMmb2W4Sq
Ied+awtcLo4UjcG2LqPrg3JbL7YbyYo3PWZkoG6+098HrAslI5nJ+UU4fgdutvx7
X+gMVWncCRDG877GXdX0CN5QsvTHUzHLuxYyzsrwzpmirE0HORODwS2hjM1PWRqi
8QXdVz4BHTwiqn9/9jbREeEBe5hIIHrqDUKuRowtWS2tlMWlVNC6JDfgi9x7+Zic
5owcnDyPh9xP5mDU8zazNiUaY1I0Os6w3xRcRmWLIyrQkqp1twcCjsFq9Xl/yogd
T4PByL1dXdobXegaNppgUSxtK0fmPeUzP4AI3p7TL0/qzlertqdU/1nIwZlcbI1H
p8T4PCfhb3JiaXLw2Ti5kBgfOCRNu7NxHOPhIeK1v26TAvs70E9QPTuMF87LHOA1
TaJDKp3fjSLr9DdEZAVDoo5ATE+ra4DQX/vCC7lS6sy83Qyd3RVZurq42Vbp5ZNL
gZDRJIa1BA61c/DMKVs4pOCxVV3eKLnxWgSOxg8/FUYYpxfrgjqiPW88P41h5Nbt
3Z+nrZOzMQ90vBoX4W9WA/dAQUXgiQctDHr5W15O/whPSg1WBGhJ2uxas7lNpyTe
BP4GWdP8MOPw/xoWWJ08jXaFkIqUAzrUZbKLz8MlZjVDkkfRZTruD7dxJEbX72O2
IvNmRKbP4dCb81wrDPZ8UyuvbuKdnVN/wu0k0ogyQOsRR/OADkz1KPu0vL5mb1UD
TotzxwhHrY4GxD+6ZZq4JRwYFD2iblrMweHtUOmAcfosCd08pWq8nvGCSBWDNlp5
Q6v07oRy42v4EN9/sInZ1I3Hu6Mw8FOXrZoqZKUCajoEFis44KwNMPSOM7BrMMBR
BDXJz4LZb7ioYbNvZkT2B9VkvvSQBXo/Q4EwUi384qX1XgbTW9Ov6Io6LTdUaSjy
5iDzlhDZyxyi5jcmQRgm6LcaGUQ8E1aS4zYzsqN6TRIlTQWUN5ySjEqttDc0nFRa
BNvsi+DoCnBJ0Qk2985m6tRYdznzixw/vHUGxWMOnnA4SsMtm6cyza/ovXyH5uq2
6270+4b2Wq2QlSxP2HkruD97j4HWNx4Z47cKyyCgbWmK1dEe5svoJIIs95CF4y/m
NjN3YmLD2GPatta1RuL4QWbwf45zaf56i3Bk79nUvu4BTHp+XbT6G/JmbeLv+2Al
vYCEFZAkM93Blp8RTIsadbdDGZe5y9sRxQWa+CdJvdUuX1eZ/uDjAP3n5Da0rDOZ
SyfqBj0zENKjvsaS8QqLaTRGsf2VENjd9jiJw7Wc2PlPY77m0/IcN9g0opqcDTDj
aPdi0PMw5u+rgsNCYehBbmgNIOeilR1oYDkMASNaYr9RlwE6ndPi3m5WijW6PPhY
2bFr/63CQ4U5qItB34XOkQ4TmUGsGGgSjDwZM+9tcpcoEmoGkoy2ipBZSNsFjkSo
Y5QeG9BRWPIgsyCIo+iD8bhAJNntL4Q56gEpC3awBPzHynVKTH/0le8XAZ/GbqCv
fTvLDuZfwaajVSYXilx5ggzNCyxwC22KjOWBGfiE0qV3QE0yjjnkDhos0DaUap6k
L2uXbGmp+q0WgekA+JtIe8vJrg5wW/C4Y9773FqxfOo+r1g62h5zbzdEwJc3O6d2
H+Kn0EBliamlbnUi/juOqVd+ZGnz0yB9ZU0+GyUSYo0kZokeih5LcryZnYgMc5fA
L9SpZ183vBZkgS77ZI3HWsKTCmMmN7gyMtVBKxqw6escb6Vi1medQH5k1whjjQJj
Z8V9pDRODgHZkVZC1k5NOtMaYQBk2kSe7qGcLlhAG/X0ZU1Z8XBd5gOPT2xRXKox
nyRzyF9lZbwZFc0YV1Uw0zpp5+7fE0nhmWtLTzzDFAY6mytYroLB5jbCv2D7oqnO
YQdmtleD55aZ+HFJDfAPaCu37OdFq4jMGKkjSpjarWaJNtE4nSv00v0ZyunLiyb+
jk2CWqeIxr3G9lUq7iFRf2cL4NpA5iIokSnO3UFmHZYXmohzCBQlavAEQ8y0Em3u
EvB8wM7G5Z9nBMI6LvpHGjBnMWgVXffSc+EML62vkSrGJQOh/neKUDt+muY0Lsl7
8OykQVlspGzjUtdZgOj+bxWEkqDQTGL4PiDOnCd1iF9MKA+tnEB3dk0xFUFJmRhv
LQ/n9nw3gt15Z8Thk407UONQ8XwmM8dYRg4aKEUAjN5gFhKZegIqzHp6ME+Ew5ev
i6MyVWrjYPGFruAr6JL+Bm4Usyg0BJZl0grHPS//BGCnt7hGMHZWglsMgMBYAa3S
YNoHJ0emhLgY4uEOZtoORl8YVzW1GqJWVqOAM7qjyshwct2iLJFyjxcX0ickpiUT
J5lpbIV5ZtODYjuO6ebdzeN3v+69olB/memBK1+p96Z9z5zLmtB40NRzx8J+DJpK
3UDukbCJqX1hra7qF9eqJU0eoMnCRDBuSFooQFCT2eQwBnx87TYj7UJZCjVTaaZc
r5TOJUnpy74tSUQI68B/tRclEQOAr3BW6d1wRU3TBGlFhDZjKerND/KO/54LAUUI
xPGqM2Nkx/ywCBUj4onZYR6ZyhLOhPBSQxPm/i5kDYcmlZZuIGiGCDhId/04GewP
s8X0PeN2lCMSUKZnup0qUTEyBAe9KmeyjXtpAlNWa3yWXZS5Fz1UHSllMqQ3DYnH
D1DI5xfamcvjGYNUdR7AKS8b/0ObluOf04H+HIs68b0OBvKUuOiz9VfQ46rwOywi
foHQ3tnuwGAibvt5rmiMRAn1kmfHWZEzSMysJprgMqDSCMZFvS8PGCurnNnwUgeX
u2kbuCiSt1+Hb1O112jlToKFYIdNCpU73zQB0yL63uQKrol5nYOkbr/yCJAoeZ11
tDRe38BpJqY+SVvAvCNThVnyL3YGrWRvcHYr/e2M7CJ7eEqAdz5cxjrawoFZX1ok
ImWqruRG0muZK5UfugXpIe5bJlJoVVdB6pSJYhpDxPSWdjj1itWaTRcZUWyuc1a9
+qGTycO4Ci+glVe8RlCI6fOHUwfaADhfO2oTGmrLHp+Z9DFgoeCegp5EbRFSCdU7
mM3QC/UJqCp9uXlPe7i98QaH35LTFk61VtXZBEgDLLP8esyBvPpw4QuC5I6iRJEC
m41QXpv7sNgPc/0Jnv1fuOwaOhK1t2ooidQ0UNeCcVP8oEGYzDe7ubPdNBhAhGTr
mVNtwiquy3ga4Q5Ppw44798F9xxMOymi7Wpyl+HCh6ZYrzGjDf81u70cRJBPZVLy
Zq8/VZhYDDWGRcWRbxTa1XEWWbGwm3FwF5pCJK7akGLtkYWHEtgnkUpm1C1tnOt7
UuLudLEd+SFTyVk23lm9K2be0QgShW1Nh33skCESXImYmM3AXmOrnciGuoIF/T46
4FsUH9rVGgtsMG338qgKFiHwVYUqiBLBXYkGNiBI5cyCtk83n5iUcCyYEGaWI5mW
4vKvhg3DT/DH+gxxhenvxtD+RL3ST6gbbN5D3+Jk+q/mB/trK2mh3NX93JFUXgtI
Xqhu1QvQQj7tx1PcqY9zwHpYO+3yts03rJTYNBvyltNnZDQft5dmvI92tg2rCnAG
l3+/5g6sD03qrsRt28uLZ+B/cdpI2XUhIZcothjximvUbqPreAf17GqNPwVPZv5o
mww7Qd7gv13twhqfFQj/85R7iiEp1efeGX1BuhzK+zl2MsRBlTF5DDrChuJK/lSw
0rkvvJCyKWmIJO8QZx2zgjvzfkAa4IuJWaRPADPW4PvyZROiwCErjvYWrn/H6zs/
SDbWvFmAQYyzYpMI6SJIG9cPMVFtciIbINfouEehnFSsH08Km7YIOZgc/ip1vibK
3HJ2HE+K3DNDr6FLRNVZZ+0ck9pZfLnVR383bkpp3SGSOGn4AheUjPf2kDFZks05
gPwqJhDn8rCMCx239S07BhGr6TO2WiKS4ngA+t1z/96wNxkw+JJ0Fi8QpFfKUBEd
zj9Hs/zWf3QRGDqQ3Hpplw1UzduM2gs7aKyYMpaOqMpVaRoqLb0b2guVZXo8Q/LO
ZFj/KebwJyxj4/IpLmtuqvd13jdDdrF0f1SxB70B3oDRG+zA4WH5rPeRVEy2DmrW
5FDQMWAcTxGBWdcPfY29j302W7eBgRxrEyqUa7CicDaOyuve5/8TvbYd74OodNWk
QxkQi2oHmFXz1k4jMAexduJSGTnPPxgBUPt/GHICbFjBgYb1CGlSwiK0JE9R/d2s
4GB9b2Cx2ZuP0zN6UvZjeEGgwyiDJDqYyRPgBOnPrzZg+xEd07uAUhKypZfdsvWg
ojYCrdfoYSr4ZyyX37TFqIFMTy0VZ11hZUUDYXEN5TOnNez5MrEXRxh0OG9sw0zE
LWK+5VErKk6JOfC4vkRJCF9GtN/RLaJUt3eJB8vfQRNpgkX4+jT8UH1x8XiwuCwb
5PEn2MUBQWQEzJfbyonvOBLDeRBYF3bc6QqYnYS18hmo70+XEfrZ0o5yxpLiodi1
OiipbO+Osj8kLtaMXzb4H9SzvaBsdVfJg6vaCqwixryV1zvunPVLiGwalamoQXMQ
thTxs/NhCTfCmCWWqQAjd0ywr0VZAyQaPGVWGoUWR7Mf5bTVBniXLyTQ86l/Aruj
5TDTH4WFaME0YdFZYbc65y7TgsJvxi4BLjQJJWWo0yamTT3tp/cU/8iNpaWRGGSz
M6J1ZmSgXr8l/DvYAwm2q46zrFkBnZ9KZV81O0KsSFEOfm+MukAS5eyBJSX5JyEr
vbevgpP9+Pe1dSIpZwSU07rpZ79d2u0jFUqhLEF6xqUciXblczyDPQ4Fy99t4Lpk
NVbAwkZvlQAnSS8sFgoWd7ssE0DQRhkcJlPijSXNz4gamBOFCsF8OI37Pwm5RMJ+
4h8ezHFmFMp/71LvNzUmvcRRRejaeq/UiYUfR4p8V30u8y/7UkOta322QnzT9h7s
oUYbF5IsZ2utF8JGJmbZ4EwJlCCwY1PIvgwQR4QfXnU1IMwKkuYjz4VOYH5eJg4V
nYJDoHbojHGaulAJi93W1+oPmaJlTN+gZM8I/DjyYBGgTtf33yyJrZ1YqdZZTWy4
xVYUwIPdZJyEGfKc2va5X+/y4B2d+wS9JWH5SY0KI2wxDNZwy02+Ejw7W3JKFtHD
/ycozoptHOcTBHqS6MH4C1Ho2cZi/9sWlRojHeEWfV7HUQBLX6Ivsnkjmq95EsVj
Xij1WfWy7401LhuGMor26r4Zvmxz3erUYUe3MFXYcDBzO+8p7jlzlRD/RCpESQ4G
nKOYcr50Z9bXAHwIOVcwexLWNtowWGbU1DKwsEvxJiV8YHq1EE1oqFrr148DX4UW
61ietXYiZAIzScgIe72709rHqEUJMoJdN08dEnvhDVGQaGhviTxOHZ6ySeO2Xb+n
XiajInBIS9uDx6nQgZ3wBUy0PFyBpbuXVp/2O9I5X5RFnNvbZuQ3POf/aVvAckJM
q9CyBRfPSg0AALrJ0lEkBLjCei88n0whI+Tvmkj5vFvyN+XF8Y0VjxMdPfmHwV5k
DCpuHqb8MkkmdKrp+4xU5ZhTLhvuSvYUJMx83q8hdz9pYazBerF4asFJQrugoK0u
RYo+74yxSMrpSRvknyNQuTlR0KqZ/DG67AWlP8rj+uAqmPL/pwI5cce7zqJK+QOn
OVHO9pnVRMr93+RNKtV0Zg+aVLlBUlyUCvF6Pq7qmdz/dfWIkdW5WTEH+hnincFD
XyH5dkHt7gYR9Ne5nB3lSVwo/+kQ23Bn76vi60/VRyanoBSCEP+yXiJtOcPYTkU8
2RB20A17yXreTqJQWiXlkFGBTFlHTF3lgn3KfVdnEchbWndUhs4Rom8LdhamgiMB
vUnkrFdv2xn9Z7n7FizGYEtiQHak12QiHTmq8vai/i5wDfiSkbRsLZTrivTvUBUH
bR+2qA8o04lYvgtJoJ7Tny596uBVawhcyO6WqmdAC9qjiiYvVXzj277kRtn/G8PB
a4wdlizfuBSr2qoFNRf1OKb/BcdW8kkGHH47k904Pm0LEhOA3XClacxUDaxjDpPK
CGz1r7ZSxSB+eyP1/opzPlD8SBv41zN58tiXNC7Xj0a+MQGeWicWdT4qHlpKkJ3P
0syehlFSngaliiu2E1DW4u9T0NCcSgWCc0yZoWZ2NcwLK09udFyxQ8vZzyq+kasX
c7R8gVG+PAfuDdttluKu2HaEaqvtSK4qBmtKEqM5KNLZU724DBMFKs3G545LIRY1
2aMFj8/PCcdvDogtq9QdW3DJhcUOcYPZ79j90vu+Lr9+fPbKG3CGpX0dCxPrCDpt
5cwHRhPcmat/EL6O0qRVTCnMU8wLu0MCgE1/NiNv3lGzFSwoPyhmpdbUPw2rFzIy
C6glk8BZ8Q4/xMGNIv2Kv/HuIfwnt/uD52eO4QxwDuWb8MewnedSX5LRBIq/nIq5
Ceqs7yMQ0MsoYhmkxaXU+AAzJjMF7svJor6jgiQJuPBoBOqzKI8+FuCtIbZiR47e
raMqlMt00PcPXGh2PP1/GD5uauU5NpwRBY9A3O+BY7OKJRp7y6WSSE8EY37vow/Z
euO4tJ3tIRHmXTvk/XzCliSIjKi1gD+3CVhVcLxPMTFoGHyNt/zxTxSGY6qQkcog
dEMqhOFeGkj7DtdHxs3Za8shZ9GyqWusS7r6wRhksA4TwTFygGdSYuZpqkwZ97XT
Z4jvC2x9H03ZmWKiyrr8gjysld3fQZKffIHk+1F+JUo0q+uC1qy0yr4cCKfIsf/N
vkOIXaUvi9c/WCdA7TQ3X1mMMtqQiLDmbLxxEDDcL7EmYqbUSL+TMS2kIyCxjgwm
MuOOLS5ri8zPaTJgpDndy97p/RE+RwRXmF7i0OmTPdg9zfCqZf4IVqTuRjRIdMTy
WK0dHruws3rhVo2MYLUdG5eF57AIkvUBGc9Nv9UQiQwHpm/Fy7f40JYyYvIzp6LF
ZjQK44z6IaXB8qKyT2TspDA/x46OaN1H6Q+hW31AFaL7DCkSBNBQQYy++c8IfvRc
uk+PUT1TRL6ZVaXNKhKc6LnfEpqF5bxVbh8o67mEUoPEd11iryfwhrXoaa9aRHE+
GmmGW79bpN5X1mEe7h3gDxx3YiM9jKpss+5WZFzBbb+gaiiYD6rGI59Vo43DVOvb
Qnw/gnqAWIhlnDPp/Z/qPXePeb1m9Aqt/wa+0/FlKo3Y/8GL4R5WASAVNXo1pjdv
hx2PQG7eEJ5bJ7wBncNWJou5IiAExz5dDPqTAcEC14y6413JKFtbe4R91oxh9mhV
D7lxceD8hDL3hXP35B0uLC0SyqxxHieBocPknF55BUkqgTuMpXIHsytN431yYaKo
dASNmn/FJUNU2493M2jMj85+3VO1emYDWKFDZ/fl/Tr0fN2OlJafW+mRpCnxUMhq
3GoUGpzz6eQa7+o+cqUhIe4/A3kMg7YQ0/f1uDME4woGUA28w54k1q2dWkevfAC6
foCZ/uAmnZtwacak5mFcVKAejE25gIAO2TfjKolA6hqGGU4PrEpAIt0demlxr6nA
X70i/RUqQPCk7gwoaNE4ETCWoFHrSjUH0C/2bJ0S+WIDCpyKbXS4j/ckmlNkeEVI
5f2rocu06Ucg4BYxQsso6GwfhKDDILrsOHau0CbE27FBawfTslJLpbYSHOKpsWw6
Iu9BLfupPOXW2yVKqqyUj8OzVygDTu8X8lMtOI49A9w2vVYEnAROMJ7R8oOBBc+s
z5U8CEiE8ZBt7RcoSmUahF46qQVfMf6tMcbM4qPuiiiaxnsIjAx+c+ZY1KwiaPII
Q+yc1Uulid5WsbEt09/gmiDfzCXZM90sh0M6fL9HgpTGYeVg4fkKnDciaoHlB5NS
MRSr6tps5ZzDbGbxHE0mx76OySPFjUXVaOMcxfGSSY/qtTtXSpU9XB4SsndJ3sDK
fM980EcTT1W6c2H99Aci7fpuSI+lL8eQf/tCqOCn6jrmA4g3wcOBs/LJEVObmMy5
ysx8TjaouXdrg3uZ+djaqI0Ej+jkci+K8PlOELCgEPdwW3k1vIsZdg4VoQtZk3AK
tZjQV5IpL9bY/EFTnMz+L7s9auhl1gTmosPLjyu6kU85zJWCORc1PWEv9PTtTTfC
DaORUHZjCd5A8DrWskCUZyVQ5+7Wp/2pstSPXVZQqLt0K0eD4ZNM0dP0e3/SqjhJ
rHuym7HDqo1W4XJ1ORyXR8OtThYPS8AJx1V4/lD07sl9ISOw49bPwzLdayjSN6Jt
knYty+omokrdhM5VUZAEAl+d2atFYHI4oW1Ti4ineRRHgsLhc6AVGcoW44ccQEOu
ci5faJo2lylYu3Cotrss6PWaXGeUm7xxDyRBbxPVXIUu4Y9234iGACi7bHI0Gtti
cf/PCuUbLtd1wixyNBdjE6rMwOPHHtzg6J46VVU1Pzi04EMPh5GuejMNW3qdGiq9
eeEsIcBnzoRESxepkOgVGicePqYGn+Uy9DVh5rVTrr6FHosUw1plCO3J2pn4U1hW
t/ds7YfeAN4dhBAyc7oYd3wv6kQoO4POcwsWk52eDL46Rf0ppgiY2S+/Gb9677/d
rnbRO1wxehD78JLn662fAoLoiPyT5Px4Sxt/dGctr8u5iyhBb8DJeymDEEqGD2jo
tWvTdGpAZizydX+/gusWW0qSYnTWcrtHrYgZsgHYueejXZIj2zSxHN2/mihM4gl7
e0Yg7CwPCz2Xk0E5xaTuzoX0pheFA2lxTwkopsu4880eQhf3jdayz3vkFim/Qx2p
KeIb+Zhcel8+K+aUmjCKAyWcl56F9Qg1wP9EDNmvaOxoD7fZBvU7G1TCjophsclE
ccEIphBRZePuSDYwXDDaPUZxXLL1oiOuSywv/ZYxHqd+xQG3TpwFaqLe8j81tVWI
uWV+JpNS72qso6MSkgXbhulnwQyThJGosmOWcHI9Bi43FvJJx8o0c/mi6bXKCALc
q+5cRRJPv7UT87IitzTmlFBoPKVOcy74BvooJjh3doUH9wklkODqpd7m/b+AYpT9
lI6XjEDHN8wUI0z1O9hQmHT/pXm9iDckcDJxwh4B4gZo8ptIRJN+I6hH02yVJeq9
JemCiekTnqJK7gcAiMwBF2n8EyZ+cUzP4nCftWYsvFpzn8Mv3iFpr9NmQWHtVI+l
zCB8B0AGSIuvbuaKu7mvNS9+k7afQLPYsh/VpG23at1nLMonWVheO3jB7zFTzoLO
NpOuQtmyNcRBzWuQof7bk0qn/jl9HswCu/JnZdmt5BtnP9s3ayV0SdEuGRvEoYj3
WSPFemRpzveJBIPMGRiu6bHZAwLqQkObb+ecU90qe5l6K4QxkQXcl3vjuigHcATn
7IYufm7Otcfm4xfj/FJ1xfc1Y0AgtWPuhu/ybLHm15ONfeZoMku/9NT7CSwlQ6U/
DOz+llxD1Xz3nSY8CPYqkaxwNbdAyRxOT3bdrff181NUfuPip6aKv3megZbDoReK
75BPEjJgweBT1/Vyd0kNUfdDbwwdvoHf689bVYv4UtT/tcL2PNGtre+o/fbkxRgD
YAnNDq3rs+jP9c64KWDfKCWE6r2bEaVwwZiSfpWIupjTHYWQRzxglo3Lf9Oiet5U
/b3TaXanKxBflC7+wy6NPIVEkUhzFbvWQvyinBCLEIrx1MyN+ultoLCeh7YNUIaq
qAjqx9Og4aDNzKO8hz9k9ZKzuSr2AcwcAoOlQ4JESV5wsANwqjUHgjuqZMl6KVaU
Fu7/gKUGY0MESOIb7EnOE57fkBpcGDn/RSurBvAJl9fSvpyGnYKglNmBNmepIMHy
o56JxtdzqZ/tayLm7wP7++oOhF4F9vlu5//sJ2UoseJMWuPztS8+3vHA6EPXfzqB
xUf2orTa9W5Sw8M4RBHm+KWqOkbLagWu4VzUMaVENOeuHbDOJIunzRXbHvFwxd1R
/qX3XZJrUy3XZdBLs0PSUt7zUTbx/oMGmdCGlvzbSgBwSKrYljjK6ZQFCPxAnkhS
SFBfVIl+54ofHdbhBb57JWXvztr9pW00vI/YdJp8QUh1370plItxjVcUED6VR4HH
oLLyjjmT0e1dOopR3xEPG9l9EFF5IBVxGgf0RPVg00bO/CFecEC1e2jEGp91s8uW
y5/XuEmbrzb7QzM1oeg0XXqBHySwfnr/BWr+bT/n2Vn52j3dyGNdsBMrFq3+PWVY
QaDJsT7UqMPPS8Yg6QDrA62sN8Kat7lB1dSesS77l67k7+kFIkzNu87cdzRuMrA1
ahiV6/0rmwDZnIpz7SZdMDWRSPD6TMXYJkMQf7E4O+ZsZ7vnJAAOgUcwWKGQl6AZ
0WJ7ZRSWxdFgKxcsDbpHJy5d4ny6YSsAjvPIunnI8aA5KIkV/CPlcopze6sTXbu9
caFwPUX4NHuigNGRTcKtbfgwDTB/SaN1RASlvDB7paq/xgQBghJ2itKgHVEvCG87
PvZKKhCn2DWHeqSx39qTCtBxqSroq9Xy9Js2uIN3NsWZ2rcDeOUUh/Hj4F1YcU1I
5DbA4oOYsQJPCwpvPcflGlHYPCDOCOhzl6iwJ6zVIlu6r1qiP6K9UJOku+FOynid
xkUdzvKzNFZ/E6ySKCeZho29Pm+vkmJyvGfyQTwOrRu2gaatEC3ptmiaY/uPhjxF
2PhsO6+ekyTikDQMI8kCD6ieQMJbpdI0Y/KFW3mSpdbvHKyAupNGew1hUpkoFNHF
BvFipskwXvwOSTplL4Ow/WY/a+jY9f/HTj0QLm12SLU7us6iCvicFyWXm6BBVzDd
/1x1rPcfZFVqwGVviwpLZh81Kgvr+bPBvTJo4II9E4ksyZ0X8OUzQVi+G8HSDPKw
HN4rwymxjNd+UR9HFWjdp66oarA/UkHrTemugIFs9gpgvhJHXDJ/X9fnWo2lvzu1
OH6V2MV3NyYaSsIa15JjNxRqSc0nfUjq+Icq2LOnT1pbF4P7B4x9xNs7Uh6H82SA
4DPD+zFUab/fSqE/ptLk3P4WHw097L8NMuNbxPOnbhzFBIx0+s/bvlQehs1lILa1
bCDIjbMnG85Gg8xHNHcMAJB+zp5YPth4+OLLLJPbb/3H0wnYf/FvCd/Nag9ouguK
CkdWkuC9nkUuTRnvIr2Ofu0qz57Tp9cu5uCbSqb6Ac+9bre4QZXH9A4T4yJC6Ul9
mf0xzYmu6/HudvuH31oiefbKhA7cgmP5GyU1tkcsqNnm9hINwtEmfUa9S0b7u3rL
T8GWezFuPcuAlqVX/aZwhQQmeRUxapbWkN0VBWAgDJ5nZ46ldGsdv29GT0CLjDYM
X913dx9Dn5ZIhIH2W1WmfuG1/Xe3CJVsrtSBhzq08abgKIb6WmEzXEB/Xx+L1bvq
Zlo66yUeGJPFvz206OubCVw9kzZPToCPJNEsbpaPjCRs9uWAo9QujYbC4Nl+3PJW
OY7slXBe6uetse94fcTOrcybXb+6tQZUHmobuhjeqVmk0aNLtKx1b5ibKb/tXVoS
pPMVA1JZvHAThA77Jqi4H1D6F57dDBOLxlFy8pUA2SyHGvwz0GKWxeGwOYwxEGSF
Jsfy4EK5TqrLgI+BrhW1/3y0NXi7xpFvf7wlWWKwChPJgfPFGIo8M5c/nyHOGeW4
lRcjEQ4nXtgpjcStNtdt+54czYgS86LGbiEo9jkuLDTKSqtjj1bw49oHDm9JbN0Y
FTKtJ+F6GRBTFhdvU/voxIEuOAL/cVEFPUtA4t9bb7Mmke9s/DyOqsrAoEDGyt8D
alKx8tmXhYEk5AR9gw7s/B17XU3XmHbfxbWCisFraEx4+WvPp3qEI1cRmmGTjTmV
0kFhuWbLDsb0TbNnijJF3NSw1ViYPNhenS3NrEO+W7Dog4LQFBXL4X1XF172DOFN
9hDZVC+zndmCdVs9xlratYzFVy56PX7XiezRqmnsvOUeDclQ/w/Kbt6ZffmmCLdH
S77wNU79lKtD1muYdnfOWS5Ln0N+z6/e153e2C6A3XjNPOV3xMiLOgmxkoikW/1Z
xnO3OyX9WZ+E+5NlIzo09lAG6JOJTF5V/9ftVKkJzrpyDs2vsRo89KBEwrjZodsl
Qm0gnPQ2axXWDGVT23uSH77t4d/A7Yayxps3CzhF2VG1EnmfiwkThNh6VB0UCnFg
3ibx9LrAIhgYcbxSaf3yXrX63TzGFfMj53uAwyDMxu6MGerLeAU6/AgKxyRzIw2i
kT9CZbJBP9fnIA5od4/pwmMVPFt/niSgBHxX7bjySXEVs2ZylYu9SxTiJz7WSW3k
uPZBOy+zScpMwjFED1FC+t+t2hlMZ9M+IY+JpGWyMezTA7QbBu3R+mSPnl9YfG25
g5+Qwox3W9Qnp5O2AIzMrbaJVAjKD1wXq43I1gRn858Pmwt3R5I3j0pT2xe6sW24
WzTxMIdWyQKQeH3rPUzwHZYZuw+3hQGsEmsLd3PtVMXv1mHcW4P1kXraqF65qgCB
F/HqCjQMlpzXq1JSJ1O8oaO5Xr2Op9DNBvLpW2WXxpoZArXtodaAxkUreiAnKykD
SMBfVAPKnqdx/aF4CBmwWmWqaz2KshBhXXEMc1TzPxUoAvHIHv+QCl527J9/Yask
FRcAlzqVsKH47TmkxfQEJsNGKYqix+/HGha1hDzEiCwbfwEGQIOpziLCkqpDbYx3
TqFa/CrX5r+LP8tjAoAyMdGbHqFje+wN4lOR3LU/N87IYPL8log/PZv2o1IQWYX3
PIQ3cPQ2a72CRjwboOIYyeJOLnQ4sv9TD4YJG/fOXUY1klJjQn2zxj+aYc97Gtmd
MYxjB4Ig28Jdml1Bet1Eyhfzm7ahVr8ig0eyO3pkxyfQHR7siMtL5D7BG/g1Y4Vy
QAneWHUBMbnz23cxZtwot2CWe+4pp2mjroOFNrTOJDr3SDP1+WP9I0UdZtZELE8N
A4c+i+nnbdeClm9STQ2JpZ3lQaQ3xILux5qhh5c06/zfRnl/2mtIP447oniLZRx4
d/nUS/Q5dy/SZhn1J0BR1ceqMa1RHW94jdQHzQOsdqTcmfMldA0y88VVT+NwzCgO
m+ctDYo0YIH+fw96C0WWwhRtC5Baigirl/yJrhMNno/1KUaNkG8DeG4hH1S5jtLf
may8uo8ilwHKW9BvwSXgTF7AH2XyzykJuS5PtmoTS+HuiOznNIBMyX7s2E0dGOn5
tnGUw+3aAJLrRcBbTEtbfPSZS0/W6O3I6/pIx1fZ9gEcyn/FnFvbkAyDX3WCQ9YC
lLza64efsQPmPlcRraiKBE5/ZDulj4lLDV0UwiUs2qwjuCi+TWdNL0q3J6kVK1w2
tUGTpM/rKDMkMLNS1CdAnIamOOdy8g34lIZ+/OTrm0zgkufrrPc3vBN/EnR3hALv
rjn2oagsR6xP2OcXLvUrBi13R1jMKlViihY0wU5mGBHBGq9TLmzqhMw7iezWvVtt
ZokATwp+wkwIVM75c9DfXG9A/tT/uUW2FPeMZ5Bdm0OmEyvNJqfnvhDfZCk8ncbj
Rem951X8Xsfi3M9NqqCBJOsZY18xqzAIV38SE2GCj+Jb1DSPLbT5RHuL2Qeglje0
N1e53Z23n92vbyDxT6a/zriyOwfB2F35Wilfq7vut9YooYKzYJCaivhieM5eNG1G
70TJLf4/ogBLkJtLEpb7Snl++jFjAs42tOBPXBW42RA9IkMyFynjZWkGl6BrPUMc
5wWTSjidas3Pu5gP0BojjqXgZdux7WgEGU4J01BAQdQ8CRwXyuVpSYtj0TrQ/sZ/
aNIe4lhBkvq3D64jfUq7ek6vwY6gXoDvPjzi/ewalBvEfcCf5F1I66wx5bJztZdF
jmbBaeWF5eKORavBod9wlpaI3GuNJSsA531mH6Iire+AwzUw0KmRl1Tl6RaNMoDy
0ZhggvYuYM7h75ZQSBiGU16RxnGxfxb01v+RU6GtVpjXi0Em/9FmiQDFbPFRv4Mu
W0CYZHD8qTxzVPigfZWD3pHkX3fYsvaw+ftNh3wkwyBeT93oub3n3jMX89MsEFLK
xXLlWFYayO+g3k9bZTnHcVHetfawztB90FInOeDMfoqzJMuzLj7BCYyknPGBF4L3
gSRTD7uR2NPM3vKEMZx0hEZFGCA3nBrZJUS6OD+g+Z67Gbqf76bjoQp2aGw/m5cy
syNACQboZ0sXVLq0wZlRgG5yEPUNGmOKCfyxre9GKNovrb62k5VNb5UZmqcSDdYb
UgUXQOEmYV/5LkgJI8hDRrUQXId/72ldU2Ta1WZfN3ydLtPNoMMl8lKoDrBDHhlI
flJiYs6cBo68lQXHDIgLm2Gm2xlRp6YQYzUlthipJmq8jw3Oa71CnsrPZMY0nlaw
2m36ch+DqSMxNBBYTvztIGbA4MbYJaXjOGdh/YUbvS0LuG3Vb4iw7+ZgRvOpM9sL
atJaQCs+FmZYPyjFteme5fQQUihbk4clfjTswDFY12ySm/oK1igjIkr0Eg+nE33d
bay5fpsm6HQuxzIMf8unDAMQWfxX4fui0D79x1rW/X9wktycztAWzwFayB7GZNCJ
ZfG6l61zoCbh8MF6P7zWHU/g8paeFQLkPrXagLb3IycR+/xosfmWy3k65rFHfYM9
hhUtb6E7zcZcNmzcqw0qp7WT/rnZBudon3wTDC+hg0gne2J9fvLImEfoG99hSLCA
7sevx5bwhKGI1edCfWDf1vFBcNW1bBB7D+oLD1JA4kCxjjraygHplZ0jiW7z+Ssl
w5kH1dY5rUnJzU9uH4zQ62/oJmYsfK0yKXoz1Jrqk+dZnMWGsv/9nTBVXwI2enMv
sOxNkSmREorGXRoYUKf5dGjcbqyCCaiCdEVWrM+1qD9GpFIHABmIQO7uZdMA1eKy
A4KrE1CmuZ/4bAwJQYV67Y/WRbYZO0ofs9ewzQ7KDtFEdit3/Dh7HSN52mY6LUjo
N6Atdk4lsr/Y+4iM1zCU3LsTb1Todl5tNLxEUG8ZuRL7ZmhkVMA88H3GKFUsUioQ
L4+Sm1lsB1j+iGWgxGNbwEv0941+C5xk90X2I8dakggKXqdVZ2aZcRd9r176ZlEB
S12sU+Fk5NlC8auDeWpdKU5MVCHOMPeXEUfY9Exl1T3T2543UGpTOa7Pe1XtE6uf
lLFeQap6re45oikqvYabCXEB4yEPGOJ9b1SNtIppnxsO5q/Mxk3yigfwu5q6ObzQ
Bq6g50Iuryw5PBp30zoWg4T5V8eLpvQ83N/P9oOKJKajEdQbvJYK/2BtgIqxuKkd
qjKXBFef2FakTg84WGmvmBOp6wSMKE/V07U8PKvUdb7/56RcYCPwZfn0GKkDmahH
Y/kWNJ3toRnCTo5HBT3Go5sG62hkkmHjBk713wI4UXi7UBGPUNS0jZSAsKGbC/C2
mYFhMxgeXR+ELedA0TnQFX3atElyFgcletA1KBDxSU2wphVHTZZ0FVRQGR8GdQqt
cRrtDcVcoXQE6WKqONpP4zImEqI3iJe49EnFrsHq2Ljyvvp0AqtLPDbhjnl23GuV
pbAHQYXDPu2fVSGYG6DexFYAQ75qqM/fCOvVhWxpBQjX93ln3yQdZDaOipPlBUhS
AQYYWLykBfJ3STSLbpSBwh26KmYzkyscjXIIw5sqKoXSz5BpzDFZZAsjaoOALxpC
g7oSZYlrUg1SsjY82s/e4wPTr/0UCjVU3jAu+mZXeT1oOcpW1rzacTk/NIt/qf4d
DdF0DOVW07ZovAWGJwgKGBqgEZmfhzm/LQi/y87kIv8lHEsi2KVAIhCrETyfoX2J
Q1St1qYSt//xrhTLDvnpEACQlZVmgbngVKCsQlMv2lZwHGIiG83tTHP/nU0cBw+n
TfFru7IKkIlovTBi6POvGeNPLYzg7cqi9Y5fO2+gmnkLT6h98twg1TpxGzqz5SfV
Pzbkap0FszH58hbR7E+J8NdNPfBZD5pRndMvfMYuyH8e3Nhs4G0qhLGQPt6Z7hX3
I6ATaFKUYtyI0tC6fzKvkv+Nj8EflVVe/ii6IYMwEGXhBDStS9dSgmXK1TfhuCXQ
bGeFNN2xtiAQc08nArQfF5GEMtjrvq1e7sT5bnaUmYHjKjiTBDxCKUjINfG+kmMt
3U8MmwD4TRUVX27a8MIkoaVw0oJH7u83Opzm7u3DYZwuvqtV/OniLOFgfhMCptcX
MrMUxxUjTLbcFBmdsDPXhnmSpklf68POXUdFsUaHXIhPsAXZ0UkDud34DlLz/jHA
Wv1ZQzpPgTcDIKJ6giSIg8dNADkKTl/iyb3S5mA8EFaGgaq6n6PEOLuozXoRxXo0
TtJF59aYNkP7lFtmVBhCT3wsfMX6XbLd634JccZg3ee10c8RdyChi1jANQFt7lqo
EF3219HWSmJnFl2LhAsW45XhBjTyWVFkgfmUDxTGYRJC97watG+sJYKgFH8re8aa
AVxxY6LMDeiTI05xbOK+H31QP6xf5Iwu9m6qpEFW+7syrT2uyDCHrMOTpirKH2Pb
DTLK9ftyR1q2Lj/vUqh6tPgPjUqFlNHeuEiCCsqyo7RqIQ5iTaSeb4NjXZGe87ra
tytkshP/kIRg3gg9rMiWcXUo/xK+PW726HbKanVE/jlqTpnKCJ5HdzlEbRPaXGp8
e8pZod38HdBNSNHzZ7s7cGpCx/UoULOCda3RKs83ZVRCtfYHRB/ifDj7fHhONTsH
38mC6+94fjBOPyqLOI0Z5maT+cJxooxAHpWo5RrvrP6b7SV6IJlRRjI4MVw9xHb6
j6ctudhuMYeHpVsoYY9mh35OrooXGlL3r0G/kiZ1aAqofkQaSZuC83fb3rF5uLNr
NJSSLt2kYo2fr3PgxtiOrIa670firK5MLCfueo0rJaf83ybGn3xPT7vVr3MEcQKs
YwgniU/m88mSQ4+a7w08Epdpdox3t2NXYh7TObencFWdr/uCI3wkEMx+krZC/Tkm
gPKaF3upeX1X925WJIgtmE3V8Tgg2MuYj7P9SsuQIJdoPHBL/mz+0gjt0eNsQCDP
95guZAsnJTN18/khY8dFz3ZrhukP0oIQpFxMZj39DNyKDUU6vyLBuVsi1gC/28UP
3py6kP1CW6Spn1FEuM43RiddOxc2Z2OAuW7Tx+XHywu/oytlSnMJ7dx4aQjSyJef
eLUWfrcNiBwrtOCbTKSCJZq58m+IP4bv/ak7agTQTx6RvO/LkeuqraR/FNm3CPwB
DNKLPg9FlVD56W4rTKevddsX/jTdDHLuLb5emcyhqDRqbJAnJf5Re5gzkkipIiVx
TBqRAn/sUD1NwC8+HGLBC5UvNF/cY0FyRgZWs60+ktnTOjwTsDx+WkADlbXG9ud1
0GtPVY9xyY4IGKpZ4Z5b817NoENVIudlPZOCfBA16NBA2fbaRVP6qhD8hdrkGIGV
SbhYkC1Z0XeMOe4NAlJ59tUf1CgHLTWUPmvrSuvtInDeGoPQUH02IdJ8CbrsiWlf
omIjgBnShPk4a81mOMNtOuZY61miXutNRJKrwPZapMd17reMQHO7oyHOEWovyh9f
AuxizV4fDj5ipStoCh9m6ZZP07XrfOl8w0u2eh4ni0/owZjdlub28bdVUtMKvIem
xSKw41zr8rtNHy2Oo/6s7nLZ9Hh5qy9AFTLaKiFxMkHdME2itjySTEquU93e6Sjb
BTRU3GYOFkglGTs9XWsO3eiEbaUuanoj6qOXnGUDkz/3VSlK9V1ek+2gGkVDv5MM
B6a2AlNq+AUHS+A2JEg6HiEc4XXlND4V2VMon9PKJlKsFm8pbMHsvLxj++qaWCir
J3nQ4aIDflG39Nf/44SXWbC6QjKM5MrbJouoflegEOP1DxROS0sbzV+n/PBqRn8N
Gn4/uLzqbDXGBgoNTOKPL/yJ5hpUuNJ0oU7rPbtVwHH/rFccyhBDQywFFl0rL68U
/B80wyhmMAQaOGwO02xNrWl1k/qYTyGlrTpyY/RQUbrZnazkx8GP/tMmegyCjGl/
S/GiBCSUAtKB80CnHO+pkuOiVE9v/T6w5S3VbT51dqUxEJqfOI/MIWLN1/oRsVsL
baUmWO0j3i/GFnIiyw/eQsFlkg/lQAhHBaSRnK6ot1ypuSQ17qi+44As6No+3EQG
SMzlsZfMRNXSU3DvWO/vwmE7QXe3s9ThaElwRTmreBaFbtrzZyEIDIV7HEcsviDk
6dRVlETcNffDGxqxsex0+EUT0F4lFgX8dAdN3OrniA4GY95yW5aNEUQt22BHCU/c
RNJoujSCfkDqz5xnstnEcSNcbHkSFMkVVT7VCaskUNeYp+V2HFzG7TmNPgR/iLLr
JpX2HgP0exMOfkhTeaKW7YM9WuYFWFuF+d7ioN88utG4KGTcdIxa7/O33JEL4rf8
ZdLiS755l8kAOAkYCOU37vzajZx/niSYLhPC8sScABPURE28ElrZCWWqMrpFmCUG
7ot8AGiFUvD5RRoEgdQNwGqHY55AXUJAjnR3Ik8wx9A/rWTIxQMlumS6CrBXn8n4
JDeanYXtZr5QrGuPeR87oXJsr3fwgJurq/2owqLpo4lnggrQeN99unsbmo0ExV2y
LDBaQOJ5DcyTAnPrwPAlYU4Tu00tSSOmbi7xEX1Or2wAMBWj2z2NJipcpPw6YzDe
3cXo7KgAvUAcbjU+P9fo9U/DSONDWRDWUg/qgZLfcG8tCfLy9TygIjocnddPj+jN
/nQxYQhBKDmG1XEd3+dJGhkedBSrYUsNjZKud3aqanwZugt9izumMSE0E/fcPVsZ
tGT88yGShGUCCaRnyI8B2cFj3mFxfDy/dXb4oTbGzbEOXKii7XBZGDe7nrz4aK36
ZfmI3gTc/xPVH5by8rHkQSF9Ph3x/6dyulNq0MkWB2ORxRgDhNmHkIxsRX3pxuUC
maMb12czzgSPEXgzKHmhAkqPtoKELRaThMqFqOjOsrXk390KfTbW0L2nROy/IaqW
u6+MbfeeTw9Q3NzR4Lazx8Ja/Grq96PI75NDV3f+kvjRfBcIoLF/eDahugomKFyf
wUHpjOOTrEmU188QovY0oCjNyEsQMtaxRk6l/+0F7Y6XL3/DqaQ9WQaO0AfCNlI9
LI/734mlEbndJkKT71U+O/LaVZjX7bapwwGbxQD7g77WHdzcRcAxNQFlOk/pugtN
/cb8fDYsCsuKXTxf2YvWLXVpCrTs6TZESHu8TXQGQ7joW+DeWRgnNcYC61FEeIsC
Iat12b6IHPNfuoLQv6jbWwaWUb3p2Ajk5zWFaw8bmpJc7MUlVaSZU6jHmAExtx0N
3q5oEKbJpGf21hc3INOSgwihz7s35J1Kf5fXyzpo2p9o+UcGfAoQGz2az9/gbM5D
7GnR/n8w24gi9p1hk6ebLaV86f5rureM7CSGGEVTySfdWL/AJ9iEfafuAw4/3Zr0
`pragma protect end_protected
