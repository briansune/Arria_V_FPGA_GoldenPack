// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:27 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Sm5An0X+1lhAEqdZkpqq2Plb8dtEP58OhSVJXUHKr/b4Hji6sshnF8s/AMMAa3zg
WuQkLfgyeiuP+TrHSz/mX+sJuFG16CPcxiAkwoe3XFi+/6R37LPkYYgm5b4V7jcy
3Mly1j6zaQxNYwBI+DHov0LXEKE6xLSpe/1QDmvHmJQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
cpxyHyMiwQ7wCI4nu4QrHFIGVy3zqZOetUtJFz4G7/ShKqtKbkshptM2oYhQUDag
t3/ig466l/O88tkKIb9udI/x2Jmi3N38TjNZQnAjNjtFYU0P7+Dr8aXLKZfRQ2tp
n1TzdsVeYBYkXwYRai22Nfiq2WXH1WpEfm2mswuOGGaMuCFKJhZ7XbzbhZ/ejT7e
AzFnuBU4xM9oOXu0wC4NhTL5b3TXVYx8vR7X9lBQyFscu8EYo6D8N0IL63BaLZXB
Jj8BtwphR2+RxkDvc3wJTHmJdVNAV7iajwl/WuaXnUdNwbgs293UnpUwCZl0G2Jf
g+SqolGAZIP6dkbkIC3nagFxZX0lF2ejJnTSBmnrxMlB7KjEK47m86nN+WSxpDKA
lqjd7GifymedqqriQxF5X5HvNODWYpNEtSXa/fKK2xLHs8h9cx6vH+Ch+vikMiul
YoQoWhmkeR4e5JY6VdA+Cf8s6RGGuRlCg25mqyF5YnlMJnIn81HP/L1GE99499QJ
qKIjPJUX698ic0PriRV6pMj0Y8pR53bpxScLzhZ9Ai+TlX3Mj+8c6xnpUnfY7w2R
0R1WcC/ARzLwamfK5mmPEqWgqrETLSSsfsoqErREvZQTfkIn5QafJ34CIKvBGtGV
rao/aOlpbGE8xKSwYBvIJdrcsW5kFWjEUzQaH+DNdevUW4otx9vpiVSWgoTunXe6
sMsg4pbVE+o5F7IxVi+PsjEM4GztlqibCWxrQL/NNFwrrBk/7JmwL7nIF5BfsnNN
a5sx6WRo2CKP5seZ0y3TZ/2h3s3wsOI+7TlmCq51uQsmbwRcwYXxWsH72pQLCVqi
Cs0QZPDZ6KPUgFkMrPqP/CozN6kYCwq2waUGrKIqC0QX8jtZqNbe8SPosVUYMaOc
l5zVJf2QVUu1YL+Q3XsL+n/Irv9w+dN3CCcnkDuo3WkOQ5v4F+sVDh+T8rJXz2Nh
g6AyqP0kGcsohOsWU23+UHoKiod2o0iOeKMf8K6gMNblxBXCcN3beUDz9ScawL3t
nFXvZT1HWeuONiohMvAOsBHp+N+vvl0tCCK67KV/VQladsFNtkKGa4hg/Qj/ommN
bU+BkqfAjWmGPoyiLSk0IgBF3HPfuLaiWAGaW/Pwy3NCtcdLRypcTLu9YExiFK1N
nmudookzJv/gymos7NULV/0TlVFfbJOlMDfXpASAZhreZWXF9+hA3+QdlGd1RD9f
Sa3QRiFIJG2KppRgKGbXCN+yRlIpwSlF1ccx4Cww8tBYatTefyVVHE9469KZUOBV
cv4HyOBnBZm2esRAods+X8T/HmxykYeoLyRLzGK9qQniRqP0gpWD+Id0zt4zsIbv
ren6btR2swSHaVLy8cx/mSCu5IizrbWpp1nfKK1lYR1Zx7YnJYwIBcCRTvOvDSmE
ByKOl3ikSc9OikSSSGeRBBieUQBELODvbE3VRT2kCqj93QfuGT/HVRixmods8d4M
KFA2P6kOLzadqmHrpK9n/4W3qbOyN66uMhuw7tC3virhEuVlIjHUQoyXlhpr10QR
2GfSHTYOUHPFh7D0RAd9bO7iKyaCr9cVMryrsHyjN5TsOYymKG/zKv5GhmTbCBYq
pp7T9NNI4dM1ApjKXAHOkeglOuT7vsG7FKka/aJ3fuIGPs5lIADBl9nazvTLwYsi
Ys00TMPckDqTG+qoBsa/48+ilfPfMcPVqyJ8wd6MCQz9F3w1BfsK+Hpsw0934O/n
Ja7ygUguTFVIK5K7vPTbu/yqZfLC5CMYs5wctarnf8CpqORe3UeebsBy1wZQeOnP
+TLC41cvFaNs0mW1km/6CZMfyK1+/XfOSW+T7RloITcx/BniNBQ1aigV8PDKS1VA
y7cTuK8gFlV3S5RXBSOIAJH21q0gQ7Z79hEaPs/S/60uJyPvdrZBNSTbDdXr8Y4+
NMnlvPfrtXW3K4QJSVn+dwFaISxEMUMw/T3vCNnL83P2OCiZlxrdIjcK6+8wTY/e
xzIITh4FROiQAI6TIp7EuqDXolNwQ6tyQdIz0KTYrT/m1WPIG6lcM0CymIb06jex
C9f1CxGGUpJxMFvceikUQCeQEUODS5s5FCc0o1HNKlu0lmo0Y48vcQv7eDkxq2ZQ
T7gL7LTix7xOI5RuILQRI/qkYWaaCsLseZ9mAC150hXNT1WwLpdbw42G0g9E0L/1
P1ZVV2aJZIOd3d1dgCPrr7IVAdZGFpG4exGw8wiEoQJbpisNlguWHWGJvrYKGgpj
FA+uUPgFUuviJMwqI/+C77iZv82HVnqGdZtO2FqJ9LP07e8iW7rIjEt9DesP/1Gt
e/g0oXXjix6Gz51dpcwlnfuZJZ9Q+lf9pxGukr66y+q4TiUDQtAMi2OGKtULYr1n
MvfsUVqgKw7iMdC7M5VqTHZDZoNQiVPxOPOi/5s93z5fdTub4LOD7jo+T8Kwx1QC
0g4Kk2Etg5PHm1CF9au9H9Z9wj78yOLbfKu5R3EtIIB+HkQMAdU+ZsUjqPrMWbRK
SGAihd4w4EVyqMGPW0bFYHrWAO/vFGfwITrCNoovNUAvS8b6o79enuw66lZoJ6rw
E15osD+tMKYRpB4smpn1vjWzddSvz8677kYBO8jKp6C/29v87QV6YjUExqnrHEv1
R7ivc25Dyw/g8v8jYC5YsQemqx5UGSYsscvbRtG0/5HXU5Vay0zqzypqSQid+bFx
U95z38/mjDNYu6AdRXz1sXnlnN56b1xmhTlUGAE0cIoBD2TR+9gGSqolBG1rK9at
kUA5e+Tf5M+QH6tLji3v3rEscqha6NRRwa7V07rD/Emj6eM6mKoR5RxspFijx+c1
FzFBJjBV5mDnpyGVrE1vxEJ5ECINC8kS42XV3PlHySeQupJZ7gjNB7739Ifdo+ji
mjL9ZhHApusQEk00TBWe5TTHegasmsoXD/e9fPdm6sdNAH9YV7ghvZ5PBFn+/YJf
dMr7dlOZ15sKzri7zuT84+ZOQ5ZHUhyXH2Ds6DexZZeNHgoMnsg4Mu8zc2Y92PkP
9eHN7TmBXwQkMa4kYIJoFLRNYKafEvHWs15UawzTBl62sUtW4fZy6IfaL24AfDm3
RenI5m2u2fGkNMlMfCfQCTeq9OKLM7tc5OLBXKiyyP1AeNtnSFa/JK3N4PAHeOtz
ByM3cszcYUnqLF16phf+xhE7VO5S3Vq5c7jUegcb+vn2yIeGlIRSrSKQdqYHBvbY
AV0d1/VTbeJXikhaSL9r5hT65o52Dg5B3eDE4ehILKSz8nbold/VEfQR3dVy9LAS
HsGYKNnKYzL9rH43FAR78WvLLOdRYXCklIh/otqW/fV+WwVGz4F3+uuoOhRTVNi/
71/H4B+wJON/pCk8mLSszh/QNwCjy7N6sXZvbvUFbL8C+INLKQelaZaEUVf6KyfV
egHzdFliU5ZSd0GsecdDk4ZLEP4J/MNEiCWXDSOjjVBMcL8bkioYfxt23FIXXkHW
RrGsirHhkWMhs0sUlSy44eBh8Io8QY5yap+ixUwNBxl/aii8pbXLPmANR/ZW2gCJ
3DmtDXtPw/UWqHmx99Z0HYRNACjvpv/JnuCpBuqpmTnpLIt8cDEGi/SmfjylYAgH
kr7n8Z5stiwUKDfPnFN9lvz4HIxdiOZkPwTnclWlGz7jSiQdal3YQD9DD4+46Puw
10fs8a22JqYnaRupLplHmOJUHQvTk9AZb2u0QM3ZlAo36tX9tiy4pe92Y3TFG557
S5WD5xQuj4DhIH7vmUA4T6C68esmfT/aOFi3JiXi8T2U/G39dyNAI7EMRyG7lkS5
/1ZOFamSf/ahfLfgGky528A7IJlabO93PSOhhrTLX3D+kfOV6zwy6tMx1m4pIlED
Yp2tTe8/lFz01CT4Pu2vO0vce9DEzBGow1y8sLcC8eHydTaV7FGNecM294a0MT89
tciYlUwFQU4mM3Nfv3hMwNHcIw2v7vOfswEsedog7aZfoE4x/XOhgOL995cPFDZ6
Qj1Zf6+63Y/1X/jF8LdzKFAJkmE7e7xmrY89BgwEhvAG3iFItQ6d/2mnSGX2LQ+f
nmSfIhwGuE05vqZWIOCRUN5YcHbVPFuryZAt73Jk6z+RsV/t9nfupwT+EQMaNX6S
2uB4FCRUWX115JeDrt5KcJnLaMJxR0eNl9WTrE+FsqO8Odpx2QUEMaGH+pYGlDYm
uqBx0nwgs5UOP7nMnsNJYGAWm+h1gaykT6NdJ1ee54Q+87OmJA9VId7DU5ya7gMr
1xoYb/ATHT8OREyFHTiyoq8ZfWnvZVW2vYMg5dgAjE5zfVdP5m6wBSJV6eqMvIJ2
kMgz6GwxicynT2R8naLYBWACzbn6+2fZnjIwP4GALafP6C36xbiracCqwF2sgao6
Lok8GuzD7JnatWUaZpzRcMsKlKWMYo6VVHQMe3lewpj985EAEtzxt/fkG0cXKWd3
ahF3vT+pcbpuIMFnpd/l5nQYbW+jvPQeFDokJ+cxciKkg3d5s8BiCsc8cFohFij1
l207KgocffxR3n1PSPoN0CbF59zocU78F13jhTAbUHpRZm4OkVomGXvRJAs6nnD+
CBPFrXQa9b5K3pzboygpJ2VsxliauNTMjuPHuzkPLayIGdU9HAaiKRg58VkHJEbK
mX4CnVlPn0MxctdRagxSMyApWaxkNJf9dHIFNaSesDAuczK0KdeRvC9cV+XpVXvr
S+30YZ7L0ygC1ROi1niPjg0oujuFSVigFsJeqxU4Kar006u6/NMHC81GWRYTsybX
qZhX+MGL9nxM1oYsDZvehLFOwZ53cOm9UCvPRo624wc5m5RkP4bHaxGZg212+Wq9
968dqbCT2jhIfPTvDUsT+LYMniFqv88gh149chQIp4TxC2t3zi91nlJ0sj/F6ruv
69I4HSgOe66sJ2dcMjr+OiJA9BMv1hnWaiWlGDHJTtUYPm/mwUKbW4ansgsCruWp
ehbZZlRMfoJSNNGM6w5q3AjZmHJc5FP8EGCfEdlye1gKYPRHaqtz8uW66+5WI0gl
SgD0Ek5UiGn/EJkaUYux+UEmC1DPBOjK7+hAaaAj28qwZY9+2QHU/QUjNLiuMKim
r04tWSEBYX302ubQvBrvKDdP/CtkCBwuhrpwn29325W2OdHanW/OjVxImfW9eic0
cISpG78uWW8TdctRU+/jMQV5RKLkZ8IWKjCS156/tS9xwQ0UNWNHBNs8Y6uundWp
N8XlD1U8mFYHuk/7ov8ihwlZ9DsciIjCKoI9/AXCMckeYyLlTceowFvvym5QWWNy
QyeGpFMC14el90Q2V13kWKH7E141rV5pPDiWwv01tprJRSIxmkJLsSjl7MBTWKzh
Qqrkw4e57O73zTeu28C696TX8N3mMRvHmJM88Sj9w+++R2ciqh7D+PAAAvKfaZk7
JR79fpBOYOflbs06WCFhoY91waS3mkcv2RSDsH9oLlbWqBf31AYLmrDxPSAmF5mg
hM2+MNKhGVnLQOuuw6tXbpEGKgOn3p56fQ8U/q7fNJ87irayhYPQvTMs5hPTJjAe
GTa30d4eCEvOxAozqXFJcIgg8kjD4yi1nq4P0oCarx70skovDuHjWp+TkgI/Id3N
XPenDUAMn4EaKC6dZ8HOfNXHnkjK7eoR4f1QhoNuUobCxlxyC2JZ9Ij/2A+CLKSe
5vODzBZA+qzhGeCEFck/6Sw8U7qvRBCA/C7XybfU6a+4+KqW+fLax53PooQZbOIZ
+K3gMUekuSSedvKmKfqr6LCxu0Lln6IU5vSf7m7gEYLxDWLqVuIlfMmL+/wP0469
YFtxxuo+xJJW3+H+vv5NHWcxu7vrR1rEt+PqbbhMSgoNZI9/DeYR7CO3gc6wnMU2
va8tjRus0YbHV+qKhsNqeq7UnkgkwbzpKGzP0StOTjOvhGALkJdPO72j0Q4tW9U/
Z0S17nZz96LhVZRqhBrmP2qAB1Ae53UH22NSmmg1M9inyNUGWIYreEvwj/h1ZJ+R
gUc0EQYNJLY4xMF9azDaAueKKVxvdT2HOb5F80wuDHVCP4flmbcqX1okoB/3DvGS
aHYTnkzRFp51JTloo3CSdx6gPAfSiMp/m8VrrISKeOtpzG3c4OVDnY1ycCmBtO29
J3M14RCqcKJq2p12DCk6jDEbWQYzre9CQwvFfN3fpqZy3SWKRqPSuMee/18JoBWD
vi2nILpQxYvTtdYgu9jSO2ks5QqY4kqTbCEvgVo77FmAUnFB5DB05WCI9VPM3TI7
zuJVDBW6uGEG++PgME3K6B730YhmSNrb71CUo4bu8AAgio2YQnPv6o4KpEPw8o3L
BU3uhZkh5PbHsjizwff9nGxwPRi3/oDiX/4Zu9YbLdfyTxVB30TkYrYXCsvAlroF
ayUxNrAIvFtSoGUY5ormi1kmASfLiBSIXwY25Va1StTk8NXbTSD69NW8/v3C7GL9
VwUUb2vl26F6SuoiFj5/VyyUqNSIE54qYIAbyZaJ4NTN2PdyIhE5zb9+XKbxOm99
XQFnPouv9/Tjv+7J84h9EOgwGXvJ73stTiWsayEE04UqqHAWrMYdsan0Ze+oiYlV
WWSSgtjvnDJ8XiQcbESu9p8PxNqVJ5mXukZBH2f+1v+yhbR62OpvdRv6WYznCwfm
aixboBX1Ufqv5P7SCFbux9vz6ZgkxQW0GybflZAT1EuBWfqd8dnnZWJtj8/7GCmY
IdjB3kz28bisY3AuEJ0icT/1lBqeFvTz2+oXQLg1y+aSAN6YQHUCeUxWtlkBW8S0
pRPKFsYTmmIjSdASZTyvNJn5NUfv4Tmc60RnbOa1U+hEmxUDuAMhJXEkTlXsS/bY
4l+xutJeDWG2WpTN4jZ54E94pZbeCC02H4uG1Rdy4g9rSJaf200GC8ISXqSZvy3D
Zj2cFKuB+89SBk08Xkx+qbVm3aIRhcSRgRzd0AyR3lFQmrr6eA8xdAVli6fCv/cz
OZKb2bjVl5FgBHgiS2Xd4Xt3LRQppHZFIrBTSBNZLhPlR2pfawnkMyB8PwdNzNN+
UzQ8abtKyC6CjuiDkHPlzRUhbBz5wey2zDElU1+7EDQwEoZy/cYyO35TeQ3+VkNU
BaDjhxzaOnopT7UAxV0/ZaaeiM4PXwhdOOb9fog7Isd9HfLxvqOI0q0HO7MhPPhc
V5igtUtCIPhWKAIoniXeEoK6VtMBP2u2LIjj/vVlOf1zlVoFssnWlxMH2do6xGYP
nD6ZUz9ocmxcFH2TfqmfueYjxB2/LFgvNNPqwHQ8OmMlG74V8u6g9I5mRdLpPhJO
M7/a2yCOff1loI3Yo/i389f5rMuU4I/u5gHehakfSXkPOyyjPgTA06QBvMJ5Q2wh
4me74XgnnpOVSf+C7zqtlOZsHwwp739cDtF42DBJfW6f2wmR+J+kBH8b31CTTZio
OdhcRy95S1gkMxhx+czkqJUHq5C3V1tEwj10LFjug/+j8kwzK+rYwh9r4QxpheV3
mnsucFF0mIJedMkvTh6WRs0hSbnLY1IvlJCtKLQSwKIjt1r48FVOw3qkc83q/rgx
DXf7Ql+KOzQdm9SuYvo/mt2e3Qbo+Qk/Rymh2RD0aDR76pQibDkmi2c4QZ3sTpy2
BOTP7Ckrbdflu0eyd/3c1cf2Sthu35fSjxMcUd1RMM0jFowh/pkOrre71goEdqz4
T8lZCDPEFQZA8rdQieRJXMnlzcx+5qQFZ+ajYYoSuJVn51aewCOi7VPMlg4eBdmZ
T/yk+8CYKgJjw28PDt0Cl2cLpziL3SxvjePzwit4/GTiDRbfwe6KRUFqY25iIayq
jTHlvZjcSIQbKmIOP4eArJsOrxl8KjlGkjWTq/Tyj8KuKjGp96Z6m0WtGHm/nqii
Z1Z+in/N133Bu4UrUBuDWQQaPjEBg2LRLvzW3WSQUl2Gop6dC70XgV8T0s6/iTft
UmvllxI3JJqnqrK4+RxoxJ28bt6Spc/yQrJqJ+nvXOLJlMawGBzXmF+ZrXrJ5dEX
q2LNseT9RaybFSBIidQ8nbSfT9b+ptMP6rrXp4SJMVmErQrwkjiCjPlaIDi0j3Wa
Xj/kGvmnMlSA6PCSvbIwUaisjGAFFHoZcDzmUrNwCotGDnyHxVPSztlIJ1R2BAPH
xam0SMVaoy8R94agElkOwNWHW3XrO78oymoKVZG3io7OHca1OmnSVie64qSlfSiU
bLkMF+YEQARX8owT3ynVIE5GHWjPF8QrP3gMznhAi2fQyPifvET7giydA2t2qmAm
hnD8jl6ZRBGV5Nk/0eQn34xrswV7w3NZJnkm+dc/4/JR5OX4FG/FZDXiK2Uu7KA8
JL/vjqAspfzJNK25QQITYqAFNFUyXD13itkAyUNZutwi5/cvhMd+w299NJnFInrF
nexpzMmCV8JRkzvAUGcIGadDblVyO9skqQO8fFqDlJyNVItIfqDGBfdkAPT754gw
w9BHRBpEpteT/ScAql+uzvCKXEqAlLIAVlEau5NQfpb9/q/sOS/ZE33qiJV2Il2d
zGiIitccBM8JB93DiV+uL7T3EBAheI66Bsjb+G69MnjOrPxDuvpg1izpw5FHTK45
oOwcCHbuGLeUlBDistMqT3v5wTE4VJ754g34AUkaF4N7QfYFnLAq21u2JfjSy8HV
H40EAQ2UWO0CTk8tsiwSZU9sDFjrZXP3KeEuG3a0pDUgKnBw2fdFxOdIVhdOkva5
hDS1nTIcZWNkK1Oany4CqzkzyMUeumra28OW/jfg5rr4oBqFs4JcQ3hd9X55dQrU
DCA44RyVUtBmHEKndg++aew2XM2dPWKuci+OAuW9k+0ygiQtatX01eHkxOFSsfPn
eQqCVnXxSXkOkZYj6Zlq7BdPgwnYNMMORdqgJbE5z/eziutWcHdWuwLMqj/ykt4N
rIBtBtQGai62qgSyNqButRn9kosggVQZy0GgxF1wLbl7WF2xZ58VyT51W+CyALil
iLGBdvqZyPUpsCzz5oaoxblMdcQAIGTleVrLdmb31wgIQ3lTnFjFfi5lWDk14PFG
KNXf5hcoZWFgKayUP0SubP+uhMaVa6hbDHC6tOB1FO8/ocdXT4I1xlEt95lbPmB/
tppV1CWDgMZZymXbFjmWjVnE64xLc/s/NrN8AKgYxCBcieTTo9GXiOr1r2PPVF7g
zDUM1Mos3qkYdHAPeYr/68itJ0GZozgN8eOTfr1uWEmWO5lCiWTWK9A7VFqtHBnv
AEU4STGj9qkqGSvX/MSy1tQxV4gZSSLHO4LvqpU/ukSSiVNgM69N6pIFHB87EhTN
PQTKSjlK7axq6NqGP2wujHPZ8Rara7A1MFqc0LEbOX5YwbdzuKxwkMAwmVmdS6Fx
6Q8DhVmft7Qmvo2ICuxjQLe4r/PcQsQkz7u0e6DrfmmmoeQ/yDUhVZFkNLektT2e
KSIgL4l7pz3Kg+IutQ+ZWFmZZlFkaXfGrjZW/Tvc4y5GwT+RhqnjtATFnM5OOOaD
lwk+nSx1Dg7D5C5Xx4heoCGbCTz15NF2+dmdYlLtczKJL1X+vx32vcVPGmcimWQX
P517mjurNUAYU8EfBLW78LUBsOroHbzhcmBgM2leNMcN0JyT4zlACPdR3GQ9rgPW
qQklTu80V8wShUq2ov5hN+4bkKEtnQO+wgos6HiLO3wYV6ZXxpleDcPsdJwu1Erl
5QdPZfcgVV9k1bI8QE9+Muygr6RNqb3FMmcVDrqsKjClnDIMt5R73u5+AfdHALeu
luicv2oWSTrDp1ANVWUA9UF1gKZREH25qZ1Ybviv5rG/vTKaFflTFUThC1iA5o1Y
/sCwYRa4FLov6sIqVuokaoU3249MOLmcXAtY4Xzf3MEkjKbguBWUerDjnaDbrG6E
jVcTnaPg/+BxGs6BmMXiHp//9dlmTZFHHTolth8c25eAPhB35I3rdLWHIh67nBtD
dUddNg+VMFq2Yg7DHXCkMDsQ+m/E8uphK0Lt68wiYP/kg4dBtU+48IllmuKm5FRy
H307HGKEmGqxILBXKpDZ5HXKl7gUIB7G0nBDQETX1JfOxd+Ba0j6yqnZltczcRcw
anjQytCZlR9x+H1khrJ9q7quJBzMmzapRkne58S5+ThxtOxsdfF1CW0gg/PicM6h
FRfT+Ro/b7D/KmbU8dCXhVpcDYvoq2HgOuJ2jLGsJjksXkW7BT2n0SXc8E57BqpY
iV91aXvLndvh3sSqv5TnqwDuJLSvC/yznIYB1KUKjExxbYUz39cO8IGqRc6lQY1f
4Ny/KyezUzyiY2lwo2fxrCpOtDZ4v+cnajS+G8JPKpnoS9VfniWuZIOrX8GIwoRO
+FozyimHViORuJmN70sKx6kMy1/rch3UWpLapg3bB4DFffAMekD5HpD5m7R8Gv1Y
tDsTJJk3TilHSf1HmbZ0LsRPdpJP1HUt2zSeOWU92C87Wm6ANpe77fSnsOEt49+F
cY5nK9YNSCyy6xGvkjLuMh5vuThrIFeJx9nTr9j+fu0OMgIzE9dSBCwa8u6ZyUYP
dgGhFu/nZM2LWulzProrvwQcWUIc7i+Be/c5n+vw69y9n5xY4WxT6RxQViayzuyu
vwkpC0NMrN+BBEUI3xLIkfCvbilB7gyWJkbC6y8oHmekjsUntwc3SP2Ob2ywbxDo
JczGOY8zCWcHYGY/MKOl6YVboXhdUEB9j9uYPPz8PNhjTukotiUTXg6u3pIzVH/x
N7P/Qn8FyFQNC6RChTfdgBTX5k7IZvbPdrVsgmfoSLwv5AKlZssXHBhs4uJQDjJV
Y+i2blzM3PwPCrS09uwPSwESZaJIJYqHFYaqhxM088ZVpNShv95WQ01oV9i3qsJN
18mQwFxaPr7Oc/VaPkxgECEwyDdHv3G0aa9mEilxqCeQgjQXFoX0pgeFeWUPsO2c
nlBeR1zfGovPmS4mSulfWXGjcvOtLaOBAKcsf7FEAgO/aRQnOKI/dWeUK5zG2slU
8lc1OXnMQO27/nMa+C00yWjTsxc5Gg0Kw3BMxmipDhZ8Ibv0+vthAB4mLeXVyhWL
HChsCi5F8zPR6k4eCE+d2g0Zjz6jcGF2/drsvgV49o4fnN5HyqMbpn9alQskXvO6
t2CYG5rzGYjNsxh+PFwUTtrk2an7bdeIrSKc5BGaSOBq5iw4fsiUMrUZuuidlLTO
XUjwlShwrocQhg+uXUB31vdc2PIT1fdHcEAp9vuel4bX04gzMrozWfp9ZjpWAmGF
l0tRKTrdvyS7maBdXDlNIIjQtC1mYJhKDKRB8/nDh1fkGpAZEhK29w3UbeBo4srX
jMMbxi3cvWOW2Zki9f2S32aCotnmpNOjhVnvyY7yBJ//bzp4oqf3XzFl9+6Tb0s5
YqC8m9UKeAU+Fw4SmDdzImd419XW9CMe9KqEFBMT0A1rd4aDpjdV2vZS6cm/UwV9
3RX9zkGHYMwYbH89o1D3x1expe6AYKf3icbeNH73/bRgJjD2RPCgc14KYMDeDjvS
o8sxV7B6Iskn30UhmYCccFR51LjPVWHVrflxpNrUJpQjmLUlEqUeCeUaK90MfoFg
pk0nrwYm3HtBysS/Wo/iI1Vgq1fQqy6GrqvW8T3pbIaXtYnrNmpigZciDS60IqYJ
L/btDD4CyndBchmpaxYabS4I5ry+KjkuIoacyo95yDkiW3LFsvm6odPMW/s8XTzK
a2iVgxK3mZmy2MPEUxZWVW2tRvgUS6hEYmYJ+z7iYYWNa4pfxs+aJhBCAM6NFcOU
OTXZeA/zxveWCuAQB9i5iPDJiIe2sIeGqucPR8bxM2Yl+pJdcuWoxYOIiPmQbquY
Wy/eiUoSRNXAI7hN9UTLDPsFjkl7NW7yoYRMe6sj7E+ucwRms6teaVl88NP623g7
dyMS6uCPji6VYPfWTmu+AR/tEOXyUPkMMMjnM4QlHCCs9MOCh5Z1i2pNm5SGximO
cK5S1U8OVCTdmaEOZmZmwwxvdHvMlABPvawhZoc4HGayFBtu/FM3HGFkx1xl6VS2
19qxZ4LeSf0uEmyE2T7koT41nQe/E0RdvgEZhvIugOrslXBlzOCoTvUrpUQojJSL
qw3AGABijp0X1QBIF83xlmJm0P6fdmLGDs8tG1D2lyRORj9fZUsE2b6scIZIB+9N
xSEXUPWhw/Wykt3ipMrN9BzEbJDiLXLiGTOpIn10RU1ZtEG94NX4m9Vi17QDfD5h
lGesGEBn+WkaY6VYfxiA+ZDiAw4X/oN2DCZJ6mhzap4Luq/koFDPJ+IGB0H1KUe9
H8Pz8+4mstQwO5xmjJE00wKUUTkE4uA6+vGKxWheKtW+FMdvv4zibqAwk/YdG/rK
6OG9OjLcAMQJaUzo2EFlYRkYCokDnrcSW8Q3eGilia+q6Kj0eS2KCcG6GUNRP06u
K4mVozVFBbuHWuncB+UVWFF4Nw+PcxeYiSwr7FvnJD11bevC8vZOoD2ffn+KlCxg
RbtI851RYrqpr1gOlxrT2mMRtVeAXg4WLssn+c0RwDhqsiy/tjgUZG5j9Boqg7C2
tPzLNPNS39srbklHdczHXtZz/3nPsDxoUnfCzKf6EPNQYr24YR6zehxichviN6Ti
yr1o3m2ksLh8u8+Pc/hmmoKARt/D2jcREV9FI6SWM/J6zERlbA1dwe8bs39Iwnsr
nVcwUCTNegHCb43xhi1GbAKJ8zE0q7TfpTLHaWKZFwMOOANrwFYtjUZIaDwhYwgV
08qJIH8cexhEGkGqV41agOtSCJ4cXVj4rrShdwzXWbSX3Sxw7ZrmC7lJrCpFfwRF
iz2n46l/I34NgKwaWGFFezESZRbcCbaTPlqaMBoblL6wzlBKy+nMxyijrZjWYqoB
YM7CoVQEK/JtIq1oqAF/n8jCFZX11Hb4XtngB2kHkqUEj1ezti+QdjfVZDHQvwEP
uxaZFkXixWW+E4GC+WUyPmjc2uGrOvy8B6LYd63fFJqCchyCBNK3RtsnqHbY5SK9
EMMkne3N/mIAb1dAQy9C63GB6NLTonAmdWueR0CEt41xsGLhy5tSoSNKo7x1g5hD
kvNR3kAYftiwx/aNtAWF8OcrD8dyWQzvOhpPpF8uU7mr5AFnsgU76eh8u0PBy5US
ZX8LyZCESsFGpjgA1FpJgNo+yu2ywF4QKozMpj5SsqH1ZaA5cSofH7CXbSyE6Sol
H0VJmJntEX/wUGRMEsy8ftXO2MxdqOpYOnaxZg0RQk/NWgJd3LAgQyejSvryi7o4
elsBeG5MsIFjqoGtU3BSH/j2nzerVuITBUQEamzPXxUSiBWfUHQbpr49XHD3yVY4
4GGSenK1aUSsxj3TilzJ3Pe+7GE5ZwCJbkNoKSwilJX5gpD4+Xin4f0xsOiBxDry
EJdJJFP6PUzCrbqDvw+jED6+anIR++o0+crjzXuTkBjtkNkuyCrH3tk+oUNn/Rw9
QBPbGIzV1Bp1TnUlnZO2Q5Ae85GPuoXXpxczKDERIjv98Y1cs01HWDwi5L80UVQE
INPgOagfvXvjvFrQAA1FR0iH0ldx6kTE9uzgIHvyvzyS31kE8H3QhK8yvfujCfKe
IMCh/2MPMDZyyG2RCsiyXL5UufknoouCYYzH3fb/9kBgVj/6PMrZ8FNZGDu/QMyP
+dxYoC+mGkImnsVxkgbY2zOCXIzLWzz/zW6hINgANiOGjijnpLeTX/Jue/E6EhK6
XGNVEAxKlphrYYUT5J0yrNeqxppyOMElFotLzj1z4bVjaoP+voxS8xozXoa60AR4
T3Wdy4Cb8WkII43RGDpPk3aqVmHTJWxlrgXdX4c27dYXzOraIGYc2uL/SLmq/r4L
WlysT97uaOI/WWRmkKEwZRHe9ljOyb1IeZINU92RI7iMf4reLpH28aqhzywZKTME
xqFROafK5rZUzTtN5Lj/0vuBDttL5BvQwiYlkFSkPVHl92/IuFOQlPUTzYgPZZ+y
F5DlsZzl70IJmy41tNIH7zue0a0v8GdL1jQ51YR0O6IFDrlUZr/bXYZlSjzZ/WWc
XjS4+Td9L4z6gwvpTfX4XQ4lb746rXHJp5YqYqNgDJ2WwIPbRtFckpo5juVQ1e1l
ldw3GRS8XzBMfivPOGzKKSKd39/68kk3gu+yJMzKqvUiphZ3/ONzsbui3me/k3TW
dTdrFHUCD/iTjk4eYkNj5OIA4v/WRrorMFhGPyutgXlExJb86+I2usdhyornEV16
ozy1baw2ndiSNWOTKgu7RdTmf5CNmIm/Yd5+FayfR5J+Ioax+4iRViXYu3ZV11w8
/yPucuJHIx3tXqsiMpxHtPGAsZ6EMaMARSNnz84fS61DMSHcs1TsSfJslvZ+S8lS
naBWvnHE4wlVE9J3C/8xL4+bLaPbqJzkoT6hT9Ij3KCkai+Puc5OBIaANrFYF4VR
XvwrHnKRNze0ZYshJuOFkbWGtD9T/SQvkLbmj+mTJujJ0oaplApeu30hnPylpOqf
ziIi3uwaP7GNoXDzWOCCNCnjeg3sPfHGJMj/IgyD25Q1bv8nFt+J0pdN3OB8O3Zr
x6CvDsGba/0J/Z/wloFKZYVtrgADdiI+aamJF0xRKTRyyNk38IczJUsy6tUhFLJG
c6V71EICG3qjIxqTsDPYNAfWGcxA0Y3iNvwjM3T+JYXfAIuvm8t8z7NRA0EP7HJL
/eG1zf+7hrJ/F8U2OT++NE3yx4zBUFu3r20laKDfsu+OVFpren5FQ4wZ6kuO/VO5
EqobUPAdhJklj016upRLHEiZR4PHF3Ezqu6lMnU/wKejSSawfZJ9i4IbMZIZjoXk
iuRYUFGrTfr1Vg/05pzzWTVaWuyfe506F40b17Q0H+GdlO4aHPyUHzAsjIo+tBqL
xx5ePAyPfKAy4A3IfXMkMPjVgVKtY8W7GBS2/+V8RtntQ7aww+SsbFOmDPTIiOl6
hZ0QoyK/lFhoTzd3mR+5E0Qz8Q8QgMBMSpkjVvU3A1MfNSFfbwV10i+btkWRCZhl
VB70oijYsGYiu3rNvxazYN98hZ1QYKB4Ip+On9onsV2+lFbruyPZTW4KeidfccS/
QqSFho6/j+7wPGwqCoJyaHlbm/YlCtqzpiVmDBvrcI56tDbF3S0OliaaeAmSRIhU
xnru+DF8WYTcM5uqheAGhKf27zOPGPohWj8wLzusySmfENsTZ6DmFkxXeql92CJ9
AsFXDY/LrlqL3O6MABa3U1PZyQ5NR80d2cHVyEyzpBmyJOBv4w8o18CNf9Vgzxaa
3c8TxadjlPDItAGkKKcGt7c29Xi25THX/1wWhXyb1zU/GKCpucm787buJbEgNel+
VlqnRcyHwnIB8ykKunC0C70l1adSUpYGtCQys8PrvY1JqFZn6pYugTO5EZQ71r4c
HsnZUgKDZUQDBABzTWG6PIzcPbelT1sfmsRB1ycnn2WQO/h8rIzshK2drZ+5+Y2e
5tA/ZAydvHYP45QHj/ixlGrbf2wJR0CE/hpnuo4EO15UtZhL+RtHVf3w3njPMeaq
4cmfbpFlecckNY/4my1qoOcAckI9ogK3KF/Pd9Ls2xtkEGs8zaOoDS/NAG8WZWSv
x2VSb/ngf1uQN2QGHeHrdRbdAb2jLu+Rcfm2PrdxRMWBNZETGlCeFV009ikm5lNT
gVyS9qA0+SxsypzUFc8l+ykWpNH41ZnW6Kiq+jhabW6FjUlVId5qqivWsT6B3rtq
cPzSaXI8qZJh990A9uoddp7T3ufYIMDVBMOag4MhIqV3L677F2G6lvEBVgPW+ahC
zQVV2kSLz/mrLRvF27PzdGy+Fa/xNZ6pbxAaYg/HjxftgrndfbCygBEp4FPIat8y
yo32YqPZhR576eH7ETnic/fxXCHpZIJkZ1AFbLWUk7ksV+agfmDYr1rrDZb7fGx0
DrQDBj2iPacrPkCpKo89Ps5w3UJNMvcnWMXc8kcPebnUuNwoWxFmNI+uKdnwgVwO
y4PynR4XMN5RPZ00tvFRJsuNqIAm8U34j55A8mengm2l0O+b5TDTjEB9m4VnuGFc
PYZMCNRSJOAAO9x8okOGpKRvt9dpEy+AuokOzi1jPlsAR/sCATWoMATNsGQRPZc7
XoqcH9A4I5dm+tyzxvT3eW2bavbMWxE4SGf9JU7cM6YLrm2fRUAAylvAYnkQPJxH
a29GSJskZCF2EUb6VPjhyA6ajcznYqaScedoSJ1Cq6jWzKUlHBvv5+hg+A1ct6/v
thvYJQ+AocBx/2RVlHb1eGPMGYDGr5BYk/hAr+yHc3z2ZrpNn6bF7iNjPNaPnzYE
bDWWEe6wMDIj2oQn5iS4oLLzLywH7nq5CifrdV54TR5Olxr7QiIWjzzCZuC0Qhg8
YPBMrApJTythi01ZpQDTAt0qvivLgtiyK2Cp8bcg2Chz52y0yj/22lK7V2zdGoqQ
56TXDR3843TmOCrIGDN0F1Rd5kJsEtfuJSX0Xftq5U8XHLfQyRK5ffgjvPk8igga
ws3lB76vjfOL5P6W4PRVP6QRvP4vKABRh8CWswMfmbAaxARyTM5Dz2z23hijj3FO
RDfNe5UZUvg3DGF/xUzbyZp+QBOV+z2pbotZ68HcjzXwohiHPowt796DWqADnPYy
ZwfLHQKTUPts5/qxCtEfh4yrtwP93kqj+St0aZqs91wMfiOXV20v/Le6Bc1Us2YX
huAGMTycpV8ZroXWyLk2+d3h3peQbckQ/FwPYfBVa9lRxCc9I7PiKxepbj+ulk4j
hPubnxNk/dVxlFKMXfWJze5ABXMxi2uqqkny6g8WUqVBxtjAW24D383aqkQYGOIw
32jBN6AV8W8P90bA0fK5vMHiI6vPYyZVPMgc+qSBZ/AvdylWqmmBZYFVbxZ5jN+M
DTy4ay4Euc3JA3ro77wIaPh4XeSiFk7v2lpU2JZunRBFub5kBSES0+clVckCoVpo
RQ8sKHI3QL1ulmFmSFxmfKRSZpBAhNU2Ig6Qr7CIIBmmgxnKeqEN0Ak5thxQrmjo
D0iKWEl+xftM//JvBMhbsgRmwWteuF3SET4J/htPHr5kk8I34EfW0h6+P0IuNtN6
ow073TGbgK8t92IDyVqJclbC3wlhpa13IfrMK79XCTw+0mHWZuYnQg65QZak/A+5
K/x/zkoWiKoID9bT/BnsPCh2Yv2lpQrEIbNK+CODnacGT/v4/NlZZJq0ZFnIy87k
wQwl/1LzJwm3QpudKHeDBrtLxglAlDn+tBbObVONDVzIvQHD5Z6G4/SJdqXuU3AY
6bNKOXTCACMkmllbitG7CUUgb9SL8/Kzt7PVExqOs1GUGRmy8iDw0X1+yn4AGobm
DU1KB/qvsrXHAyGERAa1UR7iAl5na5vOL+0lKwdm/nWOa+xynMkF7o7AJ0WjozRW
cgvkNEnkp+7pqxlHZeEhKRVmsD4IkOBUGMB3kvaDsMMjY9mZTJUaB65QDeLKUgUb
cZloThHfM30bv5BcSHoeCiSos29RioX/FlMPwObDktQmgia/vvp1DZ1fvUM44nSL
I6qsceey3+Xd9wAey3DfEfPNYbXaswslJGTnHTUtAfN3fsEDSuKL5kWSJYPlUPgn
E9tX2/B2ovgFYvqz/Pye8MU+pu7RYoqqQL9BuQCBLeN882jMjDWmJRW3ulHCkDiM
H8ZsXQ4w2tdVGJK8Pzmp3eMk8nlW14ASbgnUJg2HfzdiBpP8hwuLz0w5a4IG4xmr
YeJlW+HIRl+1Fciysk8/lI3xZ6+NVhv6p5JlrCL43Bc2ERS3+N2sIPF7+8wLODzh
RyQFX0WzicBy5yyhWVL/LpNJWI3wVWwukjKumVjC++9yTgS6oMvWsNArsO+LkId5
xNRDwkXdkO5rT93uQtKMbrX7De/1Uk7075I+HSkbyw8M1zVJksPWE23tpftb+keH
8yoJU5JJkuP4marNLpCfumhBnAoSm3fBbGboodzI+wzetvAeX5CgKBhU3QJ9AScF
oZEuEmnBWcT8aAOrOJrdRoK2Jcc2iUnQZjdlyUyBdD8saFU9HnNtzonoTXqG84NI
xioayAwCA73hezJOAO2pDPN6guot5X0iiL7WyVTELhLbbtWe0TtehRn2GU42UsyF
+f4Ly9w9TeXhIa05Ezkn24OfLINcEfsVbtamyb4hFq0/7rpzojmuaqLERl4PrW15
+FYqbfkAtds3KGEe5PPXz7V3WNDfzcVp+f/VtTkw1Pv9z09EAa97gdEsVNsqiFl0
WjURO7QW3CNVac98Wt5AS1RcGhCMH6x7yTLvfOZtz32dxDvgkrKtnQ4MO7jl8Qo/
WJ6CD0T6OgJpcRR6PkacuAB6626hLbHRQuy5jBn6kdMcBWljJoLtiOkeDvLxpyb+
Fq3xLBJpsSIBadwnFuxxrNQfDwHD6MFqzZVV5GwGW+FvZdHcYdDfF1loTya+q2xa
kNyWB1aRTtMgsKaP2TxDa/pavx8h1bo0vbSmT6pynjwIqG3ipGcWG9wCJNhQJAKi
CsH6oAvmBWUYB4P3jcRb32wPqrDzHLtNko60QkxVipSaZSVxI4JXmPi1DcZQx8aT
6lErV77UvveP1J0BPeTaxviR1ZGP9457425d9MG8OzYdfKn+XjLk1W1IrYvAJ/yI
semb9IJ9gXCdjPOaA0/dVcknBVXIGtdJcN5hjT6GaF8vh/iCBcRi1SfRHchcUL3X
JyYC6P/noQKdMQ8cE6QnyrFE14u5UgJfwG4PJ7HNLbD+PTIcyOVJJaaX2ZaAhaz0
4crSSKZt20CHBapzX1e7J9xnCZ9Is+crEYxbg49Wf1ndh8jTnSftucacZOGt5PtO
C85Qm7Z6kBHhhMTlwUABg/3Z8cTf84r2pJqvEdevQCN5ZKLHoKlOQnU0bk3gaYt6
z9md5eFfknkunGNWKndQa9k8y2Co/WVWqjHQISZ4mk0Vd6Pif1NVUk0m6+kykvIP
wgxkOsPsHwDb+jLjAz8QEdEqhQGY8IJuIC+Db47xKeA6MNxnTsZ4h89H/rvct7sR
mxuWPTJyx8rr8UgzuUuJLIIAOa1t77W3HnZClSB62W52BeamJd+5AurmB+/JmCY/
r6Cu5wOunsfPY4lf3N0BZxo7ICEf8mrzZyfxesyDaSAXpx+awQ+nC9a/2sTwVEdK
7EjbJ5GwHR2rBB2QufU0qeZUimVspgONsBD8n1CUJkD2JkOgR0GIHrlmeC+oUCFi
G7OrpRQ237CzaDoudmuTzp5YArWd0w8O9lPszdaIoaoPWcv3J4aUIY+ORea3JLQ5
33kvb9ma4+2tHCQ2lLdTqd3+4BPYE1UpRXeXxU0Tq/2OY6+1E9PV8Ytqa+GN10rg
kBkMAo2ndvc0SmLOEo/w4qMKqJvqpUj3HTRMdRKW1WqIoGR10u3BRrIGck5MbT/I
0c0uM8iZ4fII961yIOgkhuDUsm8fLi4gte8UnIBmi0ZEn9nmFmU7+C4KtaDFKfbR
FQw9J72WVmwhhcsqs3Jw5OlO8+MrH3WL/O4W+Qcc2iLVcqODIwNrar+OUQO4FCbI
j6iSRHEzHLgYpD5AlBdCcQ9ccMeS5tR8iBvJTHJBOdGGuLbCTgyeb6VgPi3S7Z3/
/8D3Lz2hy6nTexSkhuHAu3ai7ctGk4ZOgw1cd5C+VqcCKJS2myGkTHvernb4FWJc
qsDQifanB7HM5ob/Q9v9cLFpZ95PMNpmP/V4rJMa2xOlVgSVUNGQWNFXEeM4Pdid
9E3odbF7XMpXPXc3fP5fIYpkq/W8QJEt7T3rYJ+wYjc/CUbAHNoJYRPW+FvF1f/c
7YFAD4qWdZOkC2hsjrFV9BTlw0GunOeV1F6R6rML12gF8sMUbEZ5SVX7R9oX3u6u
HofTwaRqZMnsigFNpV+GPOtoNps5Fm7smYtVDnF7yx1r8JaUEnlsJt+ZTv7qrz/5
mLaNiMx3Ws8n/xd+NnLnpKDTqQEwNFAwf0twN3S6AJ0munPk279a3OglwrkH4L4u
KnKlSS1F2tDUBF17lRq34CKI1evUOA4CM6MAb93cdZbZXbx3ebc9x7CBx9hPLxV8
tggBB/Pz/7vvCPBH7OzFchJYbRXfoUiU+U8RYFEgI2YbQFjn+3uLdlfTuz0MaeMz
lRQWYglLaMRM3yyv929nzX5zhbBzvyW3EySMinqmg83wikxA0VzFMSDUd7dEyGMG
FTPuwwi+dGidaY2gIxEIKdJO1bar835SZ3pUuoMmVvDGR0+Xfnp8E6k0hstrXVYZ
932ZZ29ZpocO+sbHkcWINV0XRMMcc+er4/986GzScjsNmzUwNwMyKHRCeZ4oYVtf
r+kPdDUkFaoWm2pVwtFjzQOto6fUqvuPSBVDAFzh1I5Yv2n7aiQB+Y+Uy1h73ePe
NleC2jHFhbgIpprx4fv+FfG2OtmTybSPC6NX0XpULvGDM57qkiVWDXxDLucMp8Jc
rBdog/VAnwC6A1nQ0gUC9YVz6Wuv7x+2R1r0oFR+rYlTn4a9SIkCzVBCDWwFNili
T7m+pcHBesOzi/yOXt36lMMj1r9Ax/EVdIPJnuyYpGpaIwWntjSzr+yqCIL24Otm
BKAwMj5ldFaDvbtRrVnHpUWp1zK0MI1HSXU3ttgS5QF0p+V0lwJWPiDxEjid+TPH
3pxZ9r49r8gmXrSXrjQn804L2n7Vrs4o7Jkoc4S/D7bLu0iC44w1W+NHAiD0KP8e
g5kkV8IF9kPBRQ7Kg8MFno3Kl6kR/CLuYhhn82lpLeX3ILWs5z1OPoBbCnoqWzNH
bPIvdTi3jtsTL/RkQryl12SIKe7yJC8265+0youh3BOGU+F7pcWPTBpPQ4qge9Rq
wRJRgiQCcno4MxKaS6fiwx1GJDasv385XoRADtNwTZ4Wq5r6NMBP1lYz4cYslcQG
Or2/X9e8/YNuF7DJAz5pZocsQ+SI7cHzw+YpYd719Gh4rynY38fU0OVVHmGW5EnA
9Aqypp/5AU/XDAVxIiR4ICnq9TiRo2+aciXiWH6ilI+1DJCkPN38ouYdR7Cs7qqp
L2Smpd7uPmdnn/mHQeBMIShdZxkNdh4UHTDwn8Sp6guLZYEMCyKmGeRreyCR1avD
vGtV5NuJXEeMI+tlv5Hvh/5WORFIq31FxsQAdmiGTGI5dgfHGIxOzJXQ8qQiYxG+
lO1fmTnZ8ttswCEfZ8xPLnJ929Mq3oVzJeWsuiFL1MWfa/nFTmgN7wB2C4CYqVCu
ZB9Y827PFHa1lWB6RkucjVsS/ZJAYDrjfGaClIXsHtiwBqa6uhOnKlLF1O5yXfDa
3TuFROjE8TAEsBydYMHXeGpWoDglk20X8ypA7B+Yo4N2BSxvLBZOkp3aawNPw+KI
hg7VS20859ud4tFSQO51ViK3T32S41izF0l4q7YLPWVxhXVZLTFUPPdmyeRI/t5n
8MLugnWNV5QqE6RZIUJ4trELOqS5JnJenQE9E+cy7/8nucdtLlU89xf8Gv0AuTDt
PG5agWqw93LB6HLXIrz1J0k3FhRDThnzrS2ixDqfhRutI3cnHZlD/n83PNw7CAk+
Ni0WhYImOh1bDYXm97WUDervVnXAa+ZyHR1alcuOKwliwwMCXT5vQ3HwE9PJah3q
0NS580bbzkcblkGg5PeCczXqqR358yaOaIHrFCGSx8L4y8XpUqwdP/R6fwTfF5Gm
iLeP7j6r14zO8KaM/urN90LVUAt+1I8cFMcZWvm5HaFuIhTquu6iRIraCcQV2NOc
KPYml2rNzw+uCJuwUuYbay2vFWXGxs2FM8PJ21t630MzRmD6XWmai1GxRE7gjh8D
6QklSIV5e4kKmY9UlLE2zUIuVrg8VUCqpSHOdfPR04Nj1RKRdysG/RY4F6zHw3hg
nii7AeV0mR2btXO0YcOhwiw5WGdc20RwcEa3ufbaFarjjUPSB0KzTqk78NbWgoih
DYq4BAVD+cGMG5K3DrkERKNmE4cWME+71ARjzmplFVqaDuxcbxaz2Tq/udzufWVc
V/xFTscjiz+azY7TdvG0cMKaEAvQnZmzroCgIWSUgIKQJvVa92+gBlPZnHfukk6V
lRmxflh23h9XKo+SXGgvbtkBwXMguWvob63tb4pQz+3qmWzq5sRU+xHPdMUuAHc/
L7WnWIhbEyWwTd75b7NzaZy86pNJg4BfX/3U4EwmRzP96GQ0347giicdbPlw8bnN
zkE3n+latsSwKmanSr5sYOY8vQ8avw6dSFt7C2ttUbxa96MQHbutyp+7il9SIF5r
c1iJ6FBXIAmMX8f/Pg9Bbjs0giGJ7HisUaL8dK+ZEbZkNt1ZBMeOw1rcIByx7XZ+
HzzPFhHYie/ku+NTUenMIUDloeXD0hS2jdHhcXIqg//nEqhJ9RoaRW0cT/xVguHv
zUsdN00stEeubfZjzIhIhW/dT147I6g7vtfJk8AAe3zoUQRea2VlsHFeyrRz1AFK
QCDDQHVm4ZyWCc03+PDHthsQ/pjRsHU9TuoDGIMhKyLqaCxKXes8FxophxnV0QTP
NfGD5ObtA2z2mkx/e0/V7qfRKlOX0uRYy1/YRvezJQChyRDrkhbztegfqUX3gvHm
tA5WF3bVwLSIQFprxMaYsGYSU3ngOfPG5OMVLnqTbLB4iQGHFi5FbFlmB8kSlmEF
KADhX4kMmzXl+NkWd2FX5TV2wwLec61JBxx5aA136llhPCw8whXE4hcQ9ihRd3dH
pZyGDasqNVuna07u2v6v0zCNjBuw4W0p9Sd1/UDE2PNeFgLYjdxnNFA2ueqc+bQS
s5dFCdWnKYUzzfLtbtB6SWg35LZtf6EXKWSnKSuNR4oHAPOe0XkRu1X+SLgeOvWp
mP3PGu11pT9VkaXNMT+SNhCvq97Gn1NX3CSYRbG12I1UM9IjCFLUI0yKi2Z/xybf
gVxyIuKuzL6ahlrfhiLx0PodmIhp2ee12wsje77+qyFsxTz3AAXkFii43oZr93qw
sURDzXMYpJM67nkmk8icMnE0sh1e4ZiiG5bf+o0mCautwAT4oftvAhT3BuABuFFM
/E4PCO0o8+N5nGybqur4Wwxe/y5yaLyD2LHk1zR2p+8F+N0cF0bOvhy51THhDNXM
Qw0V0KjkIMXIlgirMaT7B/nBEtPGxUa5FjLZz2D/iXPZMYyhj/v8MqYSa5R0/EXG
qd9iM4VP41DragsIGzdig99kBN4JoUzSi1hly298etImjAaQPKrHbPYFhNxEh5Ne
i/SWm1oqSEy/sP0yT6Isr+i+7cq5B+KsPgc8nlcx1bRPloF6b1GSQyD9itwYsqzW
4z5ffUzpQy7PFI5k0ifFSfF94dKfyWc/LmS5Sr3kiEpr34SvcD63k/gv8L3wY4bt
Y/lX7fU+miKYVKW+ekYFNy490je8Gs2ZgkB5pTgTKHoPGG/EgvGTQOGtGhXlHH/R
9S3sO2jcdJZmCVv+QeBtdsuZynqC4zWWwoJXWHfjM6WCcfkp8Xp3iCgiUWEjwAn2
cscwoiPD/Gohc6hFjaVUY7fG3IkqhMGWPGEbqB6HfXoa+FD/oOx0OsnovZGqloyF
aOKlEJmEjSqfR7Eo1WXu33OvJ/C6GaAm1rRBrPA1ab6vYyXmUpEySKVqi5fnbWY0
2+OWJdpYmRcJQeYdSEIhUc53YHTs+ls+Nx8PhR47zYz5FCVvfwip1KWoiLpNrC/5
FaCl/JUHcMJCLSw/SVQtY6uqwPVXT1hJBtcXHBY3ttjeTngUgdERqLjd1ibk+4GI
7YWiovE8o05T/PxPY5YBQyNfbxXjJKjCO4MnUguG7wd7lYPKHbS3d62+W2EymRC1
Xo4lNKOzJRDDmMKEmKU0vvYEKpJnYz9bquAIoUY+Sk63vZl8iN+LA4KJWe1H8dnV
qvmJ+p9w7QTwEqDszxf0dGRSbXZquOU3kwqGm+EeH4UZ6UpDlj3WfOkGwZ8shDTg
TVAJKpkf9C9oYeSO94Ut2SeJ3yxcIdWJcmx6PXSW2/0rLqxTdLw4eknyTSXqyE0O
/tvxUSKFTpvl3U1ZHuvKBNaFOKbaJzWNkDvFMW90kxKSxh19ZwjoTHXcYosqIp5S
yDXQPm3AYclA4tL36kMbPsl3F4dbzWRiFGQ0SNZQG7FykJMzvR8ApE88OAQyAeUQ
i8sgNVJmBK0AVFPACvvk1Gi/mYa6MsNUehtQci8C1/Bw4Hms2fKZSn6ETp+qs4C0
k6G/0G3fcEXbAjMAzZsUM1qWopQ7sPgeWMpXGY2T+TJbcBDqg2AIIVRFcG0Kxbp+
BaLsZNM478AvikqessF831GalFDrGqr/KDpENYHK1YIYNJ2gEZN0GUE41PVskpes
hTQq8LuTmyJ013eGYMUGMmWaVXRGi15KOr6LLiLz/VWrOobN3OvrdxIDKQ95u/d3
LMTnCkegwjSsLKoVy0EuU5kcnLewTftqtATzQVRJf0Fi9i7/ELdGZXAfl8iHmaKh
m8Pe6uJS3aPTjWxZRi4vgW1+Rc9prdlUH1xScWp5U9sYcXuojQf42Or4SgsEcxvB
dnDSikUIZi2wSJRp015BrGVQIT8iNaExG21udz6z1fyPlZed4jVWGFYN9pM0OPVO
QTbV5UiNkDZDMKlpjvLKZro+rTeXbwv+viGcOanz+8fTTq2VF7oN8WEkapU1Tfx2
cB6XTfP9bFxCbVHlVSvLj5ekhpoqphSjZsCrV6ysR6MsikSNSGMWrd/wsZFQO9Ao
+mZoByVh/Re82o9hT1NmNDx+5ucg9oOGnnjgDDFunITNyl/tfLvfPiGObyVm6+H9
jpamC4VzriFRV+bDXnTNr9kIyG54kXG+E1cDmWbVN0oSeoH7vHy5cPaDQKomogFg
2298tygCnHgMBHl9SFC1Yi86drBMS8tAZY9ahg7DJINkUYywEbjB2g3lDnjldSYD
nHZddwQpsOKDHDqz/w+7eU4MHxCcDiMvS4fINr5PWjtw7h68UUmEAgboNr23/Pm4
YMbv723DwFQHnPK3DJa5i07NzdskZkyM+bMuBDvAwqale33vLD3AUXe8qXClVgt9
kkd4WmLov0Bic1fXqy+HL8s9z3jiPEKlN3KP8C4jeYW1uSeyHN0Kioqr57fAVDMr
X/wpziZBxROXBOjwnR+MpAXUGlutpyPe9BLcaI/myCOTZL9Zf6MNU5i0qf9OHmg5
+RI1o284WhyOpJXWpbQn+V7GQOgmBPHCsdReh/0kfZG8cXgHMaAiq6vb2RZOZZ2V
NI9y8QBvQfKGJk+dpNDHMDAtd5vLWufq8Q7+I5DNXJEeRyWAKMWFE4olwHFSQhy9
gy99ztxNOvxXNW0hRSUovyTY+xsshE2v7cEgwYZqMwOmCmQSPHys1Kma1KMz8SIw
7CbysvCu8eQw81SG+ujkSMy9MbpWKm40aDu0Wwjq79kjL8B/SGnPIW1gNkcM2oaY
v4hGcUSa8xSyWvXT+ZH1WMf7ARBTl1GEhrfsPQOI0bVxnXeVLDkI0MbC3OqunSzQ
p79SFYY6xUEekuoAi9MiBaZAIJu0rcT5SIJMfj6Q0nLxo/ZmnD0AQHWy9hyFXqQI
5gkmJdtLL5CqfeFPy83ZBKnDyeiUGoKdDdjvug6mO6Vj1mqJIPIHD8k2ZA7Hy2Jo
0ANKQqvM4EKlFOesy73j+wUvujSIrueIlfAkLkBUc90PSxTbyUq0tFYCcw7PS8t/
B7cvDJCNtZvxq/EtHq7CVrTcijHGmwG8kikCGheX5IPnZ+1szdsFOetT80dnqfMx
FqlCYYdzIJ64jfyvFwFGcPgcdpKZ4wKMxpmMAL9/2JHNGGgO1nTOSEk3rxhmSLYM
wadavB4lixoOMi8JE6At/u7U3z3ijV1BFv70wqjIYCuWyHxPik+MITkdpEC1FP8z
RKKlWU89Xn95Lj9UDqvZC+AMiy1KBERkG87K/YDxFJcmuh3ornY2cJdtHJ9TjzI1
XcJVpQXFjzZUKuw9qN/mbTe53hGidD/FtNum9k43A4lE9zVh6c7Inz1aBxXb1Sn6
hSTf6wwK2Wv9ZEG6bM5p/+uBnrzW0JrNYz4V44No8Xe/8jyRIU55KW6fTkOvdX5p
uDH58kep0EMSCFSanVtDXnW7UQRozTPsPCSU1AYMV4vzEA2KGrARMUcq1DxGjcWX
oEMPtz8JWVKEdreNvk8jr4OaCfq+mgYXAdL6401LRtYPvqOdaE0WIOA1sThL6Rxy
xa/4cChzWhZPpAk4YuTmQ0usXAXK6mwBFf7emLIfkAHEiNaGjKNKeJfPiIQvAzB2
5D7FFGGnPnPzFNmVfSJ65Hn+GJBKcWKoNWQgngD39VGSSOO6R/67yEzIjRry5hR8
Ya5siJoLCfv40UorqkECSGaAeR+dh0YceDHZIc1uZ/hGGg/1mCxZOAp/qw6uKiK0
4NNVxHC/pZV1gStjwdfGge5AjFacZ6lvakQsQQfhOwZ06ls67mtiGOSLewcs3at0
8Ce7BchAO80+9yjsojyt8x1Oa/jBCl5TVEFFxCvVJsPRcd8Paak3kmd3cQVyBdo/
vrZopVcDqCCRUhE4IxIuikKMBcIZ56tG0rPGzg8I27rDXWbeOabc9PDKqfT8122k
58+d8eANEVtjs3W1pbWImy7JTN4Sgr1xfxobmgR8M1xjroVJ0EQGxqoKGe550UKr
xcs4ktaIcKbyR0ATz+A4cUOXAGLlf7qp5fd7y0+nUU4qSge03iRktArj0ilsTUYw
5soSaL4lvPmZ7uNDg16SJ+CqoTlh+kY1HosYJN6vhMKKkohKbkPKR83+ZMbkfMQd
EzMrqvPLPA3cFXfyse/Ysn5+/TGFT/oNwXP11NdEcS7CWbNVFmGUEqfUhm3/bjEH
UuPssROzSai+hme40DjKkw==
`pragma protect end_protected
