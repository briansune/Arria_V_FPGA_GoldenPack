// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:02:29 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bOAdQ9BdpnDRDxOleiQelfHR+ji0TwINczPpJmOjL5D0k32HAtY3h8DcCDkZmNWV
sZ2J2VSyYkZkBARbvzaSM7hoVT3nlrAtCIt1dAS7NOvLhTA1HHzZQeL+yR5pBLAO
cEkuJWl9Ail52Oo4391Ppj5lvLAXChZoAR7310mMLwA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3792)
4eA4+6AaOCfMtj6g70ciirkvb78LhgoCJpeJLOme8mt7qch/Zt59lVwgJKAq01Nz
Vy+kaUJgqt8RXFQsx6eU5tuOae06qk4W9WVjvvd0JcdssZsXviM5qe+uSsR++o4Z
lQe52f8Q01fiG/Ic6jVKLbPa9Ba4HKRAhePiheE5dZGCvWVhkcc1E3Ql9qU1a1KF
j4dNTnhIxO7L1J020Y6hNkGF6TBwoRTLurpsW5/zBaQ616z46JPsY7FHOyEjWqh+
fM6KVOQ8OWDYFSKAHYSONMgeh+SU6PMFsBMNs4Y2jfkMmzLGzonyrsebJoEFX0YQ
59qcJQzUT1W05bAWo/38nR4NW9k1KXhzy80EAhQ5pUyAMoOISCF6YR9njQNteVL/
QMRaljaGNk22OuAkdRpVEnWQ3c8pNbQYxz2blJgQBAF3tFoGDTFHJO/fgyzE3ajb
dh7zNjFtizJL3188eS6KekDaze6g7fpeFU5vDqvqzNCTG07eazF2Uon5SxE6VNax
VRjH7LyZS8ubHEyJMF5y7yMY3LnsR1J2qbi014UXWnLE191sBI6zokjpRpLXVLbh
zeLM3WzglRV5CkNm/dn8RLeG2ubXOPNJpnMZB9HMJ7gKNlrahrFBreUjL0pcQgtl
8HFtQYge0S0amrmwrdJ/iv5dUYdS74n0efagaBaVJUhBPFilSGeA8XBjGHPZnsQb
+k1hm0A7Ho9OwawZ1J7bkNEHcVnJeOB63l5c4hvD5vld+EZ0kaeeVr6PrJnS0HVr
9i89yhtIOVcWzXE6B0nfpLFfJXfsav/kmrz8cQs/A8cLqy+3h1/yonIDHP6yVgOr
PXS9niZ4VtpQ/2FhILoaRVe/NRac/R/94qWAeG+M2VTWu1qS1b4VAXi0kjmjccoh
0QC66AIZPRqWqw58ZOmC6FUQtUAYe12ckj++XjHDvJL8gW2Z1DWbnYAfgPGWlo2I
VKpqrWZVLK/xvAXztvVhU0fB9tmGiSzS80nGeLEXlFXdxlqofXo9ClhhoGDPym48
eI0ZYx/IvtBdh6YxA/6bs9Np1T8CqvZSpqnRJ7i0d8kT8+Ou4byRHNVDSL8zqp1p
NRSXe1w7God5R+thYlxQarFRupdw+oJIWlydZQn8slJa471KZCEJ3S9dZUKWACsO
MKtLtBm+baA6JZ5PTuBdVlzi3l8hDtMHi63F2NdRUGjC+JcfZ9lXLHmp62anQh6A
avVLR9s5StVoxcdjkEWp79r7E1q6Ti78DlvkL9q2YHltFgyWuvHIG1NgbjejQWIB
lFwmM1kQnSN/P8/66kZvF1msJolJUMlHnty4QpgpLq+Bud87IOx8rp3nmCeayXTq
3vk/qFtvYwZKyR/7nT7BvcFYMOgH+9HUtEBz4UlJTsudMu8BKBSQzwrzFn1ryubA
iQ9Ne6duNrPVRsoCG/IGbipNIvNoLSYW6foG+yeDbNKhA6zKOcctcb0n3dJIUn4C
e71HRlQ6Q/cOENygzVZp3JGqyb2GlxsgJUw/P4DxCMNpkPyulH+joLS0oYiJSWsK
cXmocMeIYA4ntt1n2qyKVDAheS0O9uxM2BAwVcYjFch0jRXkJPljVXBMBPIAdemX
rKLKNj2mKreUMU8sRcrPVkZ47SZGqXiQmOl44Q8DGmWZExHlva5TNYiL0qHsZmLQ
9n9yKvJOmsr1FC9jlOnTtcMtKP5LBM6IdFuM6ixAzx5QbjldQdbSltVCQ40EIMFu
2kMcX3pNSkp+PcnOYereFMRzqL7BOWY/QGH8rZSrWkvZLxOcY+qLWAZ3FhgU8rGw
d/DcC/c9Bzo/xVoOCjFotz43acp3OZ/fpoQySRY0BSC3WGEaP5w5voJOSoL9mkq3
wIBFlm9v7nz3zNGB7SmD1vMjtFq/cL5j5G0LrOABUdU58rats6CTcgBY7KF079u2
weF6UaMhA/JvJYuvp37XcFZeM3nnWMU3wnpSZ9d684CaepCqcstavyIiTeZHM7kw
RUsxULDz/qlv6O9podlwdNMyKP4sGFPSTf2Dd3PknGlrZZ6eBFvjUxZeqIrvXz3e
SOLtEVudcTD49/6x4NZPsgV5HFXhu6vLGuuUpKc1xP53w9wrSNhbYOkvaOILTGih
/tRq1qBUJrpNRww+QZWGojQkuMQwL9IFcUJKDG+yeCtiTYKJHjYqnze5h19ohlfo
7yynhZ5OIND3gm1ZUKsX2l3fBNlrbCj7mH1MxG/eT+rcQpUsBolA2vIgTHFeV9AO
3++qJawy+ywSHNAQ1uBOMCdqVXJQF2J2Za4WAbmltW4iKUTMOIN2sxFI4a1hpwc+
HDovtPJs8Dw2Z1v6/WoLNY/wQtvV3yvipxKWqdrHDEf/7npEwYP6/YNHFmrlySCw
J7YFCsCIGLmu1LiWgJwRPrJoGsQ5T/9K3n7SqAXRtpW8uXzNuexiEMyvOlfS9e0M
2KfwQ5kX4xspGVOnpfy7IaKMjBBXUaiTwuMim95YhogZFyn9Mr/MZKncJJZvaq/L
aTYRtp3mWJUkFpiPuMhzSX7G2DqWyRuSu1rf16x0T51NfR2yp5r/qGv3JvwR2VG0
xUK8S1NHgB43JaEupLlgk0sMso7aWOn0fefc8jclKkPBEyGJQb9lfBdlzKfYu2rd
g7mLH8hLKfhGLyOsae/JD8HRthmUHVPoMTiPdnTqf3CZ5Hqx16BPnZgNjiv0v7gG
ZT6D5IdX3fV850Z2NlCSNu8czEKNNOKgZuqr95JE0edyMQ868EzxOJhkgktocDNh
NMrxKcgZR/tLTS3wYqH6t2hH0vscdLa3uqFHB/+rIyK4mbOiVGsD8628eipDca4T
5M9EKwEi8WAXlx6k/S6q/HCiz9ax6CTdD6Ejq7+xTYGo0Ev4P0e0rqiqF4XNUrQB
oJ5iluhZVWVy07DRP/lUhFX3s4G0e0xx/9aG0fneN5cDOXDUnAAcK1adhjHvII5V
fluspfpKXwsn37nFIs2PWkfQUYIg/TDxJ2QMUObAKCtQ1R33YUL8NQY3Z3ngDHBd
JmfBv+Py+QugPv1YMWEFCIO/F/kQd5ayc1t0EyI908kQDnsSJcpiQQI2vQtnBN9s
Wx5lLUeWrbMbI2ibWQCRu87OqxLM1YcyLqvOi3NJYuySbxEL2y7rj5Fh5Q6Gnw87
KK2yfSogd2YOsLn2GYdDlUo7IoFJxxBQIMFQ9+TH3yDPvAwVk08XRjF6CIZOrw/h
++L+fxHYFj+MYJIKcBISbCl1hpQsTzY9yUzSoStEerAxd4DqMQlkTJrQKauOvJk9
ZHm7jdWLIdLJnqAFQy4UXa7hlQA3jnTI3H2JScvZx6lWIICuAO5vwPE+u/p0DyqP
5nacvznTfxnrPq+ahZ2ytFIW4p01WX6QpaGoCAFSflp8oGTUEUDZpgbjYQ0n6iSI
3Og9uxvIuAdqFJDoLXlH9Xng82kSTnX54iaVOC+J5nta4yN/rt0LixymZ0CqOQQM
mnyGU5+JidILnZJgRns0BoC25pPhJhfvc5IfDkDTAey1am9NNYPU6rH5kBiLyRju
2ab9Zqq3bI+7AXxD2sGmK+yg2K9V0yRkwnlwlNpp9elsdHJThFWZQs2GMcu7F+9b
kFEuPfZjr5YzR7A5gTUqxohV3AHHeiUmif9vFNjWpZjAayq1txP1gyJ3f0gHFEuY
0DKBYKr+tEt7Esx8Cl3VzFBZP7DC4MV25u1GSYAMeU9cJ3pesQrg0DxwZPRmhI/M
g2rW5mIe7h5rsOkiAdOJ/JJI2jyOQAxWg/nCSkak7ZP6azQ6EdC5mwtaQ5gamQQH
5mL4iJ6z7XrAbJOOXdN1y3CBGiI2hTwma4usd85I90MQBUq78bFxj+sJrPXPPZcZ
jlW9ETYAtW6fyeWWWhWJLscWwdEE41+FRCs3Pp/gSkAtC81BwN8OAVClpV/vDLMp
q7yv3fDWcqNVVg3xTxkQW2KWgfqOZ2XlQlNt6p+mD2ZTZpq2srbvN7Zy9dgpZQxo
7zE/6tGw3SKoKGVe666SejE+Z5WC6GObW/nt9RmRY67JZxbzl+59owTN6sPlNCeH
TyJJXJNfPLv71xEZ6C8VtqpVg+K9d0jcPdMErxWhkkAg6C+nbah0K1j0V6ZjjhcX
o+tuAKFJ3y+XenQ7B5WOJxHUrd6K9nYJbqaPlOPpbPu5dy6iymjtRb7VEUuWx6lM
vsfH5hQbpBs81ZhHz+0kOuV2Q/vlTxoDK3kD7EeNyzR5dGgCLdAmrwdLrYr1pv70
j00Vg0qzkZNVcGKRiobvhKXksPnRhYUH9+fdGhdpQffA8VB2MX7+RXbj3dL/cywH
sDT/yus+bNAAQkp0f4MGmBRmVzmBMRKSeJykbftZ+f6DaFH35IA0fnMPLAocCwwd
mGP+PLzqMZnhPCIj0qVVqpzry8Ny8P31kU5wlz0dOlnrR3p/VNzc4/BmtWSI58fJ
U+/GKJCQ7MzLv2nqNxvF7R+Vz99tXdnFezLG0cmghV+FRo5vCQw2NLiwbNkxPJUi
dwQ6GhjujSrxyytqPD0uxa3IgIi6FmAhLBy7icW34RqxmJ343lJQtQOCQVkD2TTJ
ldPyov1gAI2EXnsOeUBfsSmxhWQkbjGnZpMeLE+WbXYPYK0lX0dYmZV9tYTTplXj
ZxFmJ8KheUZZWmcd73U18OmAc+47IH8md8PQ8rs7jJqaXipZumQS7dMKyPsochAt
2P8thxMorjkm1iyYNJSflu+YhbRZH4FuoGn8C+vF/id+5rT6eWfwEcV3dtH4KfNI
GWif1uXFcnUM4agdgDVIg4IKHr77m0XexSIMaVuW/6tTlyhrOQeY8zLbBe+zVVjI
sO5p3nwZSAqWlWtBytSMYroI1nVKe+PzK5FaJ4obxdLsACabZocOlzOPxFH72zeC
CmwXvYHt1L7VI6+colB822BAk3FY1aSUjynfiv39mA0Op8U7QEVytBWE7xGMBrqD
p1SgzTccudPphwiJWwusd90g0nTirzLSKCFqdyAdNNyrYXuerK5V2zsA+Z7OG0kM
jXPXYL/91P44VQtUI3XQ6KM1cXEtgGkRgqct4RKJ+Q7W2ovuXfkd0U3q+7Yge4RR
`pragma protect end_protected
