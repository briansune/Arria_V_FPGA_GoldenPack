// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 03:25:16 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TkXlVqEG0vwujjBbXB83sJUboV1G1wwB5P1ecl+Ub+w3bXTQ3qrsG/rLbLmoLRod
s03yHpa1N+1FxjjCs/OIAscnTWpOC3wR0k+bLRBSFM1XgaMjmlGxieWLWpP2mS/D
TigFi2QEykWFGUcL3jnLIJ/ojIcNNVhWfySgs2Css1c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18192)
ceS3xM8j0+dW2y56+B553kzsFRUtMUzQNUMwcnMW6OVScegGeC7eUtDQ2+blUlSf
Qkgfjl8YYF5/OBf8ddqtEOiTXMw84QLcie38s/4T1vQp9N+8VcboC5Dl+sZ0gkCu
aW+SW/ybxrWFB7yMNK8xkkhAbmjd5BC5j56bhK8baAXqp6FbTFeOdjB+XSFAc7fJ
h5FDsy1Z7TtCJhLw9RjQJrAnsg2i6DQHSIPnRXRaDnd7TL3mEegCk52D0PUHyVo/
Orw3z0SEEUZah6V1vo9+bVVHF2bJl+Ee1OckNcDdPAHFefC3hQ+bc7JgkZc/DcCe
VUXNqrEXyvJF46ebICowqIQQ3jMl5lFzuXE2ijVLnpeen5xrsSMKjVB3k2uvqGAE
uLB1ijJxO9HSGUBsocZssVGj7eziTxSy+RY0CNB/wA5vK7yD4+lSAmeCFXkCR6vV
NVVPoEsOf2LUkMtD+S3RdnzFv3jvvigut4QBf1rRIO8eRrasp3GZ+J6wLhHX2rDI
5kWs9xxZ6LOyLwEfmLcpCq8TETbNKzQ4TkbgncUTs9BD9EfB5uMjbdah4KcK0G/I
n+EZfYJxHerx039NZTYcm/P+9wuE/OWvR7mlVmRlh5tzq09XkfD/hCDxdbBgD/Bh
CVBzVMWfXYhyXdHPvbtEuv9T6Xe0PA5ZeoAeJ0TLlY54pi2LoIFMpt8UELgk+zFO
35cQpRoIzmOnRPQ6yL+i85a/hWY7F+yngXPIaeHit+igKgPaRUpSfEdKFxTPPBjL
E4LibA5tXlbIEzaX4ynBQRCNX4nMhkmx2H3OZ+EpwgX+Sjz5gmrB6EIcMdQMpl0Y
GqSseTopYnUOfGi6MnUOUd8ZEvxDYOer201iE/CucgLmt3Jv89ZVEP95/5liTTTs
Sm3HvuFw6ePK1u6aa3oNrmcX4CsbSOpQ+xNpQlKC7S0vY2hIrqjvhVkbHdb9gVyH
eovgORCMcmjEnsw22rJkNaMDIZdaJAPJN/Hlvjb7m8RkA/sx/FgoZeqFmNfJa8dH
4G231o6EuoEHzquzXABU2D1xoazborYJMxN0x8DSIO+ZVcJonuDydcLCXSpx3eFI
vrUU3NatwW+s80HSvT1T5aPnOabc4eMrCmHnGOOd9c9Ri4i3X9hITBljItXiAxtT
hM6owF6vPe0ZKW+Qd1eWBU7l9b3Uv+74gdid3+vT1KOSS7V0vKvN3+9aMhHguzSt
GiE3SkqACPx9zkjmWGtJp3EpEybuAvK47mUH8BDkcRHDtunzsuDeQwjZy2DSFLBF
i78eJlQTmQTuYkRuvIQi0+MOi9Op2QZahJkpad4bjrLc2pmuA7BkqxKBxMLPDVOi
Ehg0YV753UkMl0VS/sGFJ7r+2+QYP0QZmHrN2PeskSQZqapmFNW+M0w+VANUmsqf
YVOn5yI0DBrhzDIZsjb2x9pJ7JXq8dJosRX8Adiw/gdlFWUguE69W5SRpqtnCGMg
tzXKhQ0owPdNpM9s/Nhtrbw4RJWVtLupLSzNBcDjszib1A8uCgEc7ZVsqGRfolBs
Y/oZ3d2p02FOBZTcy5mMRblCvu8oHWMVBvGGQE2eh9a7lubpPpvBi2y82V7q7Uau
I1k2reR+5swOt5XK6rwfOC113VywOamLnLmrlwMpvDKc5uhdWLgT5GqVjef2OKLX
VLuV7rYvMoQAtbHE4ibKYbkAv1r5Z0p8HuT+6AAUcSOPb1ztmtXW+xXwdlPpXEyG
mf3qZ716Nm5svUqsq59y76AZc3eLupy7d+QzaX5YBv9Btm+3GtnVxo2oDUdzM1qR
T1XHvZ1E16CvHsQFPNYJE/3lQ1FBpebGhVUuBPB9i7fhy8SxtU/FqzBGPwZ6ncI5
ek021AkrxjhHDXG/oQIf6RSM5lQKZwRED/mF9+B3Ev+GqLnOB5xH0oHW1TO/CcIS
tskY+aW2yVSnWiZjPMJpZ4qC4sXWp007WL6mB/02CHkr999tzsR22vdm0Qurh17c
YDXFLbjOvn0avkdxwe6sbQxCY4RDCSDnEXfqUsVrAZDCfOXNe7u2zjjcYdwALpdt
lDrTHe4uuUUUNIEGv1eaUahHtSlm6ubwYmzD/2G98Mt4Fu885Nllnq0rJ4hd5Cgc
BFObzMK0VZxnFOtuYMyT0P2ZKnsjobgDD+jT/xTH87IDzzE9itf9A5GO1SqBUe/m
JeADk3xWqDMq6rr/cvWuX3CYEu8Qzvt/6zWJl2f+5OxQk3tNr4OfzWFI3SREgPcd
40OoTDAsAF4TxDnhAF3115gDVnX9c9jCtvmeRH/8nOiK/pBdojJFYJTqcBFRWCuv
MJjV86y3TnElzGU9pkG93CAHPkMSdxzoL9vkJvKWM0N4F2fhvQI3Q0CAsyJPWt51
Sedaa6rxxzojbntaEgwW+XIlm6vFvHUl06OnstgXglk8OY6p4T6QbeMoZxOjOEdW
VoZzLyEcyDfdnZV8BaQ5LAxmG2Bp/j7Hw0km0v9Ai0UQ9rWe0lwRljyagxkbpQA/
wYt3L/Ca7aILVest7/1yTS3+Uwr3YORzP050hnHDbC7SiAh8v70eWll/8zGAJcfU
wkx030g4curQ0ozOeOpe9ujDJzsN8kRnFNAgJPvcMbd9hgf7sYAiOksLUEz3FtOw
mH1f2T72IkoVrLSe1dkdbZZC+s9ojkLb0OIaAYflHNx9WlJNnlaxmkLkoiXjwRkb
vk/xkNElW/nloqQV0do9Hp00WFZErAJoZH15nNuLNIdJCl59/Y+0/IWk9BnPF3lw
es+j6zZMWeeTQx/rlMRhZzImqVt2e4xmW6FydzSoRZUKHHMDzB4pJvOm7op7o4J0
qEAdq/sm8uP25GoSNUMfvJB3FBgB3Oc25zwD8Cy/zcUIpNR3znXE6XkNllKTLMUu
sbT6X+ma8PgIORBBfix2/y5U3DRitjGVW4KOKbu0nlizpAL2+D+V4YkZU47PA8z4
Hh0RTejlIQn3N4CuO1LwGSYy1THvND9sjxjuH/oYGeacZ23NcPF31rE5ttKPsDgo
mmo/xPMvLAixtpGNfxISoxpBqEmcB5QpqICXtX94O0hjirCcpYHuM95l9U9VKy+P
7KflSKUg2TbeY+THROQZ25KWMRpGo+pxbfxDY/BvGAXmS69h0GUEv5zOXqEqg+5r
PE7uMulk1APhqiYmKqzLb0vB2khGZEokCUGlbQ90Oiku3oXnx2papKI6PPsO6Abu
EjHk6atQoBiFgUAH5/9ievb1+ouskweUg2XBecIfU8On5GRXBzE9IJCTnuAl6HZ0
fPaFGNY3w70/FFxP7KEVIimdytG0t2HQeWflxIV9NpMRyEc/REbOt5p6fgR+NAkr
bccFGpgYRGMY+dLf9Zdk3H1oWjIKgnYYwAJnJZaKR7oBmLFhCgpxiKyvRD+bz78n
35F9qUl4LOqQwC17Y5eGYh1GslMd2u7T2LsB9hgR/TcZJdSj/u6ufhPQgT+U0pCR
HPJ5XKzVorzGHsR2GR2RC1EgXpEXUVa8G34IyTiBwTAh7U8ALK9gfb223QC67REb
FNwmWYRhJllIlQ23c6H+UXLuKgr97FXpP77UvHjDTInuIzJI3AqQSqayFPp3bagH
qT4K8YXdInAG93iVhkVNGy0ZNL54EpVQtlNYHHVwA+vNMq/aS2l2rr3jUkHtR8fK
rRj6jLBwIBsxpSA42vI6VAQg0yTnoeuTyKwn09ipmO8kdF0H/C35HDD+au4gV0qd
luMdQ1XCLdowNTGRbZok6KgIK2fcQz4RXKnAAqdAN3QBvmga3Yt+P1d8/y2XEKzP
EKZixh25vySnJ6TI1Pg9hYOKujqC8RwGBkvD9B17emRxplDWK7Cb1m98Dd7dka6z
r28CXK4Cm/70Qz02/tekUqV2uNQ7/MooG+Y/WqviJOIR6qLSkNf50iscg0Ga2qRl
m8fzHrJPuSnw6havY72To8Q09AnuRZxy0tMPeeK/E6gWMk4iiC3pRx1PqEpPytvA
TxnK+l9aTJgMJ2Jr+F1GB3AdORnqjoNYd0TPFNzZ98W8sfMky3V8UzetLj+EoLfz
5TLuYS+X7gr9WaBQV1ad7fW8bjrqbCyBTqH8Q4qVdL9idt3QPEzUYWI4fJ7lJIUl
5nht1RXs60Q3i5cI4F1JotI6Yo+68F6PBPcA79UjWYMCtcsfCj7TB3EkMBNBu9ee
WSWifsuibC5s1Yi2Re2JM05jqfePWwxytbNPNRbC8vtESxbIpERuMbTalUjSP7+Q
ToECJOI5HDvVBQWOvwIt5UKCLtaajjSSRDRLSVIhZfRFK1uIt+ioNnUdpYzQ1sVR
uba1cUUnPIsyQMnETw1n8qnqQHQfEAyO30HOe8A5S74h8r7dUDKxLhDh7tMCLjXH
q5gdXWgtKYKrWRlVI+ezHgF+9IBau3o1O2cnwy2b70Qn6et3/Qd3zyFbtQc/0m3G
UjUAebO1003Rte2Lkd4SKagCr+xn1FcdtEJud3zwLsNeEHRa9Sn+qNlKjM8T4Rc0
DuTxvMSDgP8qR3PkkbVI0XYLP1kZro1fwZugdZJLNA6g0np6mp9udKSP7fxPx2LX
GRCTeB8uhtndq7SH90W/PIw47puOy9nfXEWDYO+eJSyeiqmb0HlIc8j3ulHy0fhh
uOtVMbxUOkKXt50Aa4ele6PXFrhbEWJs405NR025W4Pqmah0pyEOXWiZ0FAPY565
0jz3KAIgDWny/animB6wBjO/Wrtl+ptOVG5n/G1KmV/oWXcKSFlAzVezvP1aIrAF
aAxWdy6B0SiYLpfb16O/3PG/T+MZVYnFpKxCs7q3awWKhIc8WpFpzA63EUi4bhw1
1/tfrBrd9ThRjE4IijL5AH0Jc3XfMS98huwSVXvw9vYHhFCAJksvazqRkOQODAxY
zlfQSE5a2ezkInwVPJhrxe1fI5/TTgVZDVez/k7ePiV1xE+7tx0BZWdwZRVGPfWo
vrxzHZJG27oHOi5LONOUADyrb/ZsC11nPfghaDXFhKzqdReg//MfwNvGLalUWpEJ
KChVBIew7kxIB4WG++pY1w3mojGCxSfuL0FOeKmHcrznDEc0Jm7nHCWwxTTd6M3G
qVpZOZ2UunREZsQfqAD5RqkT1H+0hm4yYjqBlVIktunOX3Dp9JGKHWEmRwloBE2O
n7wSqQNYmvbu1sMEnNVW8Uk4jHGFq/lH57dFXpYq9wlP7kNv9MVfuqQerSThbcod
XQAy8uNk4piJS2gHiJh906eNhCzsamaEmzMekytDpQ4mOxDbnFEQIK0t/lgLx2vQ
QsIgxmsvzVVlH1haiPP/npgghmfsKJZEDZdsAelFWqsbteGSLwL7GVIeq6O++QS+
WJyw0euveExaA4iUVOdLFhVJrBEKB52P3jG0XGAcSce3p16XynmwnkBI+fmwD7c0
6dtF+L3KQMSnwa2+8J0zWEhAerDYQQtlj5dGf7SKiKeYHzQ9KU7ctCAudHuMzWvT
7+8tPLJplKncHRCsqdGuIUGxa5nB0Le/qK8men1ts8pnLX8piNCOzsXf6zlGwG24
3Cqlt/Qc5QgwS+3F3xUcFSieluq9eqKh9FvN801yWncn0OoaqjZRryyYWPR+9trI
kzipXSFw1pxxqxGtPLDN2T6ELcilkKzynpbB97/+PeV9bn/rASucyYl28xlcUZEt
XWs0K+ezVfSSSZJTRf3Uhfu4WbiUEsNTxHPdSvOv2cp/SOCBSl1ijdwmMhmO8gYr
NE82GBcp3qctoQobQlprYb3tL5QPwlgFvwwGwA+GRz2Y745vZ+tb4NAUQLWB6cQP
SdSxwvk2u3W1Kqx0WnVmrXJLVA39R1cbpFpatPLsi9IccFNxgCGqUmk3mOFH0i0R
eKuNjE0xhGzMx4Wvl4RYRmFI6DLTfcfTY8psYckpmosJf3GTgMw6SaYaEfyYbMRl
OIc0rVNZKoK9C02+oaLRJ/YXW8ZpIWU1svec0rU7pfdsX3pzbPesdc+whQXosC9X
9lwaIQHu5Tx9W4I2nuR2TSBkKKUnQIvE3RQ4T00W/tgaUKUYz3by865Qm7WkCKgf
YpjkMBYuKxENXms0oq/ga3dKSIaPOELK67YYnsvoSoZ6/LIQaPL75A0HwevWJol1
/pfJcrpzLAPorodQzzbSK54q746i1NbLaLQwN50tgcx+ARkVuBAh7CylsJFgahuv
hhIYyscbWIXIY5Yjw56SGg9ukwuR4JfnR42l5/DVYFT9Y7FzlQtqLSFxq/WBbgig
Ia6K81fuOU8oTQ+VuMHLpqDMDxaduP63vxmvWXA5aoJI1AaH/+FqoCyGIQsIPJbp
7fuiKiiD8IB9RnQYjMpZIfuikhmcXYoBnYvg+fvWvUK2cmiXOTzYnj/wohnnZeRP
/YB3CcIpHv0YmgeKGcpmboBkn4VQBarCMBSohUcdi8q4m8rBQczj8a5mdt9u0NVq
KagYK8LRSffaA6CAXcxY/TPu3Nlryr4Us3R1fEsvvapDTyP8w//+ov/wKVN8Dt9i
FiN23i67kY6KiCRTZ/5vWnt4PYnbziqW0+vuYS9QbFhoqw2YKF0LIN77nZLi5tzk
R3VJBMn5VNTEn4k/aMRGi4Jy/q7iu8VX4VEW4DonDw69WkAD279j5UATYHKiYQIt
DgZ3pRttJwDzaVvCkwuoIT6SuGcwdB3R3M5gFugGtPPhkKRvmMwtey3JPNPmwya7
Vln/nkJbtUBU/mO5cIzOY/ouc3IhcrK5jtXNIQnCSjskkQtB/ymEYh1SRhJ/xkEm
lH5wFeaieMClTD4Uojh9tI/1hDzfGJUAdcIvis214kPfgrLYSbDPvl3taSccoyzA
1GOL1tpvLKb/QvvLlCzDtz2NngjwfhNz+URaF2l88RztjQ71sTdJw0O9VhxvpqaQ
CWDVGJkECe+gl4kApo2krtw4vN6TVno9T6Hu2cMspqKbQVY9ZCmpcmRul3r4A4ds
rvVKS/stHGggQVGho7mCBEQ9/4B51w/P28Fd58/xFnFK5SDaiSXDnhnsdIzVSi90
+FUN7PpTzx7dcAJyc5+kh91c8tlxYDi9HYK91kpgQRvX6sjWFruLdapw7xoRk9T9
JNIarvgqYRSCdaTyaGvOfBYIpB7+pVBcA9i3tG414uB8NSYEsAoLg5rAm8dCfA8a
zw2nTZNs92Y5Yr5S7HCH6HuypgeXXim7CLSfSZa9LZzriX9jc7WmJ50lvg/x7Vwu
E4vLkvIYUcpR37XikVdH2ZLCg4F0b0xY5+iYvdNIX6SdvjrDbksrKyepGHAU9dbI
WYS5hUnbXsORzLsyg+LBCPZxMsklCj4ESkuG2EKywJPbIH+PqhYXI/DmMVRBBquV
0AkTi0id56NNb02csHIw9ZU/17pwCblgdzjADL96ZxUHwml5fch/qh7nyGeHB1FU
fH9HN24jU978Miacj+WpGlMHAWZOYx51aWsLoKrEaN17FAvw60XyxiRR1TDkB166
33d5tIqvFrIUJIzdSSipr01MkBYyvtEa+qJbXYlPHupJs4He7XB0TWtDvkKkvaJ+
0vWMEJgXhZMHV4M7+7+eZcb+yk3VjAdAob52PXsbNiVyEKCZdT7a38X/feZVACPc
R2Cxz7OmLsfmoBgaUV6qqS/MksH4cYdg1cmgmYaJKYZJ5HhnRwYNZHiCBDmmGUcA
LrorVN3VMzb1z8xUOwdd/WPKBFJNFYkSJqMYkZ036WTylryKsQU+B1mlr0MLMhbX
xqiv8yXJNho8lIrUaKePbbDdTSDQxsDCEinOFhxE3gB9plRSs+gUiqmgcSxJNCxS
10iSM9MUStI8da00a6mtYUR9i3IqnrH/Z0ni4RFc/FyVtQk+s3LVIBXYrGFozGvx
vOrDSnwDbEY42Gbr1nwVA6Ra7Tbtlis51p4kRoN1NGs5fYtIDnQKIZbHWNdSunQr
v2Q/b8DAmEfrPaLreSzwOvjkd5B/djxo50NVtl0OZIU59D8YVZ3cpZziCe9+jAz0
htHHPySLtdgFq23YJ39Ba3fQEB4zQsdmyWM8w01i7SGLQUC2d17qTvBRhR1gkS+3
bCEIStkeWhAeI0HnXJQZqap03IgS8IU/rnPHE5VKQFp7rO8LO7NaV2G4DWEtuv2K
87nDpDOPrcz9KrpO6N1dE+yBFfgf34/cM0cVHRWaoFtqDeKn8eOYWCQc3HMjsrzi
vRxtwu/Q9fYLmjwXjvNhMZTKKFQfIJn5ttAnxJNl02A4/wfS6iNHwC+hy0FPzaG9
QeRGb89E4e1kyO4vb5QJmLu1BqaAqmjYFfq8NMNUFlbVBWcW7Cw3ejaCHrsl3Oud
wwv2eRWWfHkAzicj+iiK/HArgNhOhjpt7JLpnxDX4u/7UOCt2o6iab8kq91oliKu
nFF6xEYWHLRNQz42itqpc2uCndChkXd/DT06IUmm2HOtg87B7C4hB+kr9kawFjCb
5uODTjld/jLL9QzuUeEwrxmUJddAXrR+ebFnumuJ78n8uy7OCvZ44rWPe2eruFmN
HyaEtyvf/bdw3oogqSXuirKdGmCsMcd1buYl4RLONDFVHT8R4nj3yW2qmTqYixTi
xA+EewWhvW4yBW+ncqxOHAutTh0vvgPDN8RPvGU/AhwaCKF2xfTm4XTwEsQ0qanr
98t74Lw8ww+HSPbvmiKjp3PBY2jReLVWAHrZjUwIGQaTXuQ/nEHoWj7UCjHLx/gq
/wOUATpp6euFcHkmAOoUUXJfK/3+FEAZnl/xVoJKruPgLJbuGiXBk6At40sWqZe4
WDToyxowcHmQSVB/1CJE7qrI3B1FTRwKO6N+BAt9pJBuS+Xm62PNsNpihOcfwxy4
rQS+Zh7qW1FHoYKoHQo04tlvry5WIf7WPxUUlqL+ky25fN3N31cWxni+m8f0NfAb
PWSbCsuYALCMzTllYcBO7nm7hBy/TIpBBmB50pekmKIiuBx+F+x+Kxz7JfRx0uKf
9pIy/l20dto5Qjt22qcRfVq27Kwc/NDfKSDQ0HC50Eb3igUdmj8CySiaaH7O6+0Z
VtzPpHsHtEYyZx7uEBq8KrlDeDwd4njCBX8BncZQV64nEOgh1+Z7Qa32wUa7lDmd
Rbgykkqc7O2N6BJR7Vpufn1l8AGzgYa1C6qZ0GeXdW1IKfhv7bLEeK38KGJjLZwb
lGxBn3HvcClnHPCZjiKYH+VkpbCjqdzxVFRB/sOcjHg2uCftua/OsRqp/PvQ3uM+
vSsqkeOvogqUyKvSu6HQm8yjL4sCRDjqPqtAwIfDpVTJPcjp2PDDORxyeV/955Qv
jnc6LkBh2JPL/HVmfQwTgxKbdCDAedTQlP3VZAZftH60LpN26gO/6Xn61k9nTarX
+1aVdlTnwHHhizyw3h1hizcWrcftCl/4lH/mXEvsXerM2PxuaxbhAqKoJIKknQDk
YcLYItO1mXAccxXOJV3kl01GvXDHuZzg1dTHR74HJOeXUmaHKd3gOWx6vRNRM/Fb
NxFUBcmojJRpV6DedCqKD9e4kSEBgWs5deGYHbIroGVjwsFqXo4/zQvZVGuYjUq0
IeavehsLUopZmcqyCTv/EQ3mp04pwudGMR3aLqHOWvxMuORx4UVdTEhY+8Rfn9m3
uVbX/pOgI1RvawLXr6XcHCBOVIvuLdbya9x7vKmZMH+51TvSeYb6PI/BXEvUlVQ7
3EX4in6suaBmwYChDDlT+bylrFq7EcBIaHqYt+q+g3OaKuJKUVfYzZkEPa3Gcw9g
Iz3PdGcpK/PC6v2kIaH+I0/cSikcr5JhKuVhT3kLJrkCdEZLvv+Owa/9pR8k3ARy
VZVLbr/A2xRrl6rrdoWiap7Li7uupUz2p2yHOSjB4oViX2C0w9KzyhJcGeUkihxb
lAgezo1BZPfu4tlpoi5/KhATRLlmiZuAkIvwadk+CN32oGd4LtHVmieRWk69Tj4q
W4lcUrGoSbsrgd4fKrLzIQN589z4t/O0fUmmT2sPPnnP8pxWgBlUqXujyyX2grY5
nMDYM8qoitTe7kxz7OYc4Twn4qxdLKrvPm++eJzCNg/EcqVMMzHdh7UwB/bMT9kw
ybmCG+IFUAqFRNNpw/BpZ8pctrBN2dwldxXiOXA0+89McwSqwTZBLWstl7u4r+k1
nrWSDhx9zkFsXsJkDJJJrYFC+BE2klPByrsHGYsHZtShl1JKYN0lq1lzwxUInmxz
KIQ8HeywgM7NsBCQVOqiNBcYzCzqOK1nXoHib+21StnBy9cx5zhkTOPDnXyMzzjD
XUvWr9zhMZKZUXoB831Zxwx9aard6ufAp4AXqj9JpvVPgUK6cOL1rpR1yUA9Hn+M
d8cV+Pj0EIA9PHLKEjvk6ByrzK2jYOPIw8J8zj3dmc0naHBBj/29U2/Hz4CZPLM+
kXKHj8NXg+Tu8TOsXVdeRgpCCZHPpsWxIc3YfQpnnZ/WdGkl/kPR+NQykjU288ER
//Lfe6/dCfKM6+S9UFxaautSoT81GUJM8DB+5J3g8+jGIeLO3cflO121FF52sEkQ
W34CBO2OlnK7KmUXnWG7Zp0Ceev/gBvicSnKPzv13P8NqnIZQz/VStGlOKkeCrrk
hoaXm+yWCoFwj8xPFidEIT9ikNRPv+/O9TWx0wd4aX/uqWN/2H7Ef10yiPivAda/
9AARqyLcaIt2pVDBYKunfthMULqnJmuBRsFud677KySBLpBO4qUiSeMBhqkiTrQO
ACbpn98I3v+GnwN39xBcaFyVMB+52GJa9tZ/uABPnpEE+ycbhX711ZuDHxIw4Qtu
yCXVvQkTZv/EmErZXbi78XLkbpEFhSRVh1LGiiswP6xR/IZZy2Sv01LG2ocuPAX1
aogCEygDZrcBFWYxysk00Wl2BNlOBcBPtKDbba0PMp7OUx+4TldTpqeza395bXkf
84JedgspCQiLCHUoKUyxM0IiLyFORVbqdjcNlmBCopxf0Tnd3/dUTHGeFi3G+f5J
ihRco5mD5rKMGVClF2T6l8/dTW66azrGaaGY8VUns/YOjR0YRNZkFmrjlAT3zoc9
lbIUWXW7S6JRUsVJQEbNdnEgJydO0OMngj24XZU5aG7+IONXy7RaggrOwkB39joO
O95whrE3S3j2oAiwn30FD+WJQSjtVVWj/f/PTAD3TlDv+LY8it9IHzpn3jZMmzv2
tpAb0Z4teU0kFK4N55c/fZYuuiqP+edV3xBHYJOYNx73fg/RNonUxNTD9EPasehl
7ypUCBjtjO1cPk9s2HMDQKxkW9YtvBRVb4kZs2xiDCNdDs0TRz6C2z6V/BQYjlme
qhp5fdYD/Ixbp7mEgHJOw8eKo751b1UUuOkNvPTm7ICOUynquZ0OeDEGxsI1JiLc
IUy8iTi0MIjiOPtNrdorUNPvcZaC1YEFbg2K90AHaRKteP9Nll9FVtonnSN8F1FE
X8j+KVI+DPV8ugpnkqjSpM6h3IIY0RLPdcj4lfra0dC+8iwLRJQsvghnDhvgUhrK
LOFEafVarZ9bEmKau+OeTobFiUvjOM+k3GPzCmjyDQWzVcdEVgWcMVmu2stFS9Vf
K9+44LAuyqVe/bzTvF3+xZsfjxaJM55QsKRONuCrgDhjqspmrsOY2J5ckWqd/XI7
lH/I9FOfHWSK0PPddm1jC/JBRq3+lyYqVxnsoqDdpB711AR5+Ao6Ub1N1w6Oka+/
ij4xsKOvqaiFv3uJ8dD6pGxfFVmJwfq3SeE2aBto4iHfG6gzsNzdbfHtgz/hlviK
oySOjf+MB2R20u8RBxGC1mdqAKF4Jk+RCdgMaL1a7D2WonhRjyZAPWnC9l/Bq6JY
YgxrvscwuKFj7DHAgkAo0WtpzABmADYx83my9bc4/haZRh0sNzAt4s4wqrVuUOR3
z0kKLvKnCtYyO+aldUBSZu50tYvlnvfwDgciCh8LiuHT3YDTwItIlKNyWMmHqLVC
4x8vNbRxLxILgKP0ETrUIPz/73RRhaYO+/erAr0gMeyyj7UO3dWsTp96M+cdic3h
1f4Mt7TVF15GHPRWyKKiqVqIsEdDr2sgiBofK882RLb2nhdL8UqBdUVhF75XlfZ7
xVDM2QLBfyNIlrDJh0ZitrigpFu70mnWgkJ/FS0jFFF6L8TuV92fAG45x4GdErME
Wlvx60RhZt5oAm5aajL+2g0DCdvT/5EMh8eaNzK1MbV2A1xY0d/WZmM1ix3l4Y9c
ikiM4DS6HF55VI60SHzmlG8xYb7ski8A6oxG+MmFO+C+TYkIYiN2iSOzTmaUzSZg
WW3ckLsRJiFuuz5YQN+SZyzeKfh8XstQEwFQNi2rjPQtHgR20OlhmcvV5pF0fqqh
oM9wPoPWC5XqHnJwQ6x2jiwlJHBhbG/Lcn8eH18VJjVMs+2C4au31DdkMfX9YCIa
MJGXJT3eTV31yPn097hbpakLafyTv9xp6dJIWtiS631fuRMXsvlHNgkk0x8t0vy0
IoTu6BzzUeuo3q4EHCmcdQ5qIUDUIqsTU0i6vEAy/K2uogSU20BLVVc0qZ3viLp/
/f3xom6eUsmnb5JL+FEZq90l2kkakAt4hLConxfwULwYyf1wwBlryB5ann5JuBD/
9XoA2DrepC3Y+wR7MdmpicJNbVsfGmp2u/gfgZPj5urp4kIIOFqZyzOlVW+yelum
dQaSk15w61JBswftoGoAG9GUX7xNy17/RS1aHWUL5PocL8IoHvRpmckO14nmvk4P
nLvkWKxS6UuE+EM/4EHaWK12RFXdNExeSayW3wLPH15gUH301xEu4myujsRaaFty
P5sxzm4YIda8oXRNQ2gzVOm6o2kdVMq6Ca+cpA6SotX7GeSTwylEEYuLTFU592j7
YoV7nSVV8jpsLk/1g0ubqMRtTv2fSNDNDOv7EhXuDzdIrjob0vrDi92wCt1FqNEG
6SgH8j4yNS9ORS6xmVFngQtrAJ1K0EvhtgfeM6HFwuiNUEASBTTvcpfYTJsWhVDm
eq31nfhi7AqshcoE6Zbnv3qI5qD9y45Sr/7R+woaxdgGxE/Iw0a2z/pPEHNISNGR
HJxLE2YNm70t4EvImOIniHcgNRKm0DqrTpS9AZ2OnYEc4jwRVFQ2AZDeKbNKusg7
PodnpEmpGnDS9KaaRPK3g/xBXftWvbXVqaNczv4rlmuEKxxJruGG/jk0RNqEs6pF
GAvI7F98Xg1a58c4XjJcxBjzODBC7f/6sMz7BXvmQleNwj39Hr+YWIZscLHpiYPu
Hd61F2/JoY1GJoKPw6eQL2MhEavnTr8VdpJIzmpk3sqnqzI3IsmIA2DEtq0qk3ME
KukDp+I3k+KCDYLvLJrjku4IBiVrV868OjW+cBfvNNgcjaP5QemwqYXy+WYlgnCL
ghOOf64MF4lmqVwi3f2QQDbed1nxv0ZfK8lDu0qFx5wzEmY42mwENvC8vyiwCGRL
imrDNArePSR/n7ye2Y81KxdyEC+Pzilc8cqTPtbFn6i677hdalsP1AbPjYuN29hE
VbqMui0iZi1ELRDN5Zw8zoypdJ17qdbS8NrzuIdg1RnsMnn7WSJ+GWDrVBRYGQN+
Jy2b2Ha6bStRc0fcbC4ygkXOj2BpYuU8t5MWyWjq+wtiLz0zhpY6S0OEUUSGM1Hi
4UfC4/c5JY3sDF1T8w2ASWr8JX0bW0mKNFp1l+WWKqujNqvWeRK2fOuDqNwHrTri
JUAfV7xXtlcS5gzbmMTbs1e9hHnrD1njmzVMgEIgZNN4dGcs4Oa5B1G+XxNbYeqz
bt4SD+cSSNIsVqynXfbKN5aGxxT/257iCU/UkZAmw+xHvHq6m3SS3geHbNXNgeN9
vrox84Z3jrYbMH3y5Ci7TSLjT0DBNQWY7o6FBvk+9KNYvKzTqh6xt352hTc+w6pP
o7nELLUQSJStaEduei0aPD1WcXx4qCbAUXvrDen49kjQmJVspRkMfTl5UXR8a/xd
ODp704++ahBjgojIWcY6q+vk44VmBdcTd3cquY92h/vceHM7kOGnAvOGQhgxQPqR
uNklGznCG/Ekabgla0My6lLV7Fewt4CjTVMlvYkGpYhsIX5woYGIhmDDr6FoovV6
Ra8lqbn9zSrb+zYVtl+yr6SOCkQoyWmwkSrJ41oX1V0FRaJMz6oL/Lw7+V/6e1UC
SQWmxnWH8G5VnNbExQejOCXQsDZS4pzaTfl8HxLX/Uz1Xsu2N2Hl4uVWUNyvwVF6
d01AclHiMj3aCGX3mNGOohznC5o/j1mo4yYazH6L+LaBcAigWPQu5DC0LyRDFenI
Zyu2J9n/xz5JOMqMviXwBvI36fTbmYWw50enERwgZlXo+8/lfiQ1NE1xi2I/ANm3
qyI3mc6upYb8e3+xyvSFiD78XQG5OZhPY4E3zceziQv9chd7K8N4YkaNy/shLINL
t+9skIte2qMqDG97zX2X+lS44NjI4v8p06XVLbmFMeMKGMsnYXwcG4DZ9GxyVvE5
pP1Z5Qs2LsSZ0xPoZhO85zA0MnRyINuxe7f2LDfjPlpoX2x8rsUmgmmyhBxT3GaN
31qsQCmCgchbVqQ6inpskd43Hwp3QOWTY5/CWpvyhVAU0tLr6KjBGQcPDWPIMAx1
jS4C+K1DU9VfkysoRBuA5jMaTN2MKzMoiykIqyf67f6/CLEyZ1Ees3nWYjozYfKs
ir7WS4OmX6v0S6u5iLvuQw432MUUnlI699ffonist7Or1dafyWpm/WeGuBM1Y+ST
W+XmtzJVLK43FZyIKguscb/9kQ4YYOZqivWFkGBvf3U9SOc9yIpA7R1RLjv1lOvX
pthlXt4bXr1bdqrKtG0gwaO8TWAhX0GzpgAlxMPdT3i3LLyTHJ2ES71psl2h2yPS
OzeN2i/3RPQpYN3VT1t/mkfb97IaXWQ4VL4fiMg94FF34XqIK6OP6h8dYaOpN+tM
p4y1XBazFuXhGWOCiqkft3RrVrkpKsn28U0tt6O+XCSEryaGyFxU3Tx7FNqNTaLK
jHOgPt+xcLGtZal7E8SGpp2BczPETGUyFGvT7XE5eehvCDoQDEcBrYHRUXAADsez
jonrQs0UVY61yUWAifqCB+YFEMJqGeqbJ+RWxOHMVztHL1E6Nw6qrcC0VUhopXBk
JAWgiuZVxZG/OH/wA0WXn7fB0gIwYx28rDEyrApeMLZkXfeseIAhA/FGtbJ6Zk9R
oECYjTOaPryrCqi77Dxfxze3ZvyO2R0vUlh6JkWk/9BmSC5t3mam1PKbtZbAO3A+
VTbjrqf+Arpv+zgfTSc2GcIoGaavWpfsnysDlJ4rFxbzz0DG1GHy4OnkSyg46wFj
7bDbAK4SNAergx2TPX4Q+VTyfkZd5v7UyGEVLD5Rjl+lCQ28LP83nMzq+zMyzv9g
H2wwSnw9/gB3mKkF4RY2rGs5OeUfjfViuT2cZDlM7rffl+zcpfsIiTsaRsHH9Hs3
k0anTYPI7LGrR5FLzz59NFCEJjaeaaE+9RZqme10iAW5KlE2S5d2P8O/8UwrQyWP
JJQhEGHts60GYr0VHtmJLt89nZ1osNlwWxryy2FthxGi4FFnxuI9hjSGQfu5C0mj
DctVSvxx9IsFQl0Fvg4TApRcEqr9DxZEl6fdVD5WjjFTTC7F+hw45yQoXmR7CdaJ
pImtsmvvIwZJWF4IyF0Ei+RjmXPzC5PDSsZmM8l+Ldy05u1dyfG8cTr07HCF9RJr
9NhuyI0QGkkM93PWmpvi45hOwQDjWSJx8b+TPZEt8nbU1au7Y+Ao1WeLd414v0ge
ueLWqvGGsqPyKI7uG5AiCRQybBD/u+4SgAAiMTSBjCEottURKHf1RP8I/5JdU5qf
Jj7kxU9Z/bgPAX3OoCu2Eq9V7qIqiPicQR8DVgLwdoitBIlIWtc4ND1KPr3LsNKE
9awDRCeSj9OfVNtipn8SLuc9M8tC21ngoS0Kf04CgEUKZKTzvGn82hFieHKbInhE
duYSdHBAAPUvGGdGD6YeA8Dd/syZYJVTf0R7s6xpVUGbnc4ZDty7DauwZ/66E6Yu
22Vd0n0hPKBfbx71mSm08QDb9eQKLeOaGcSVrfh6TpIigBFpYolopy58/XFHr2l1
7D3MYoirHHABqyHPjiwx7O0rSRoBmiAYqswWqBxEW22SVm8uuRIsui9rS/TggQnl
J/ACdlDEm2F565BIroPvY3ALHDRdTTBF5rrbOq8/2K+vr6SZtmGEJizPdUsv2dIb
+RhR1VQTJJiYppyT/R/7IF08uTot8yMXqpaGccuwQ/YsDdnnuhgEd7N98+70iSfT
VtYV3blYk80oOPGB8bX1i7jUziMe1eq/AkaKFTC0pgXqV+4fWQogNmjX8+aIV/Fn
36M77dupgKtsetgJzHYRG5GH+D2Oyg/Y75x8vFcwq6f6jF8Po8qDsCwWvqLlHiE6
zuMMuZouqBAAZpKcGGMY5jfJWw9VS6Kz+M7Cqw2uTkJiKlpKEuGxvZ08XlyCpA+a
+n76OTMnhIcpxtD08SicYAMkRK9zAVWvPsO/acgy1LmqHwSrYLaZDWsKGW4tXtK4
jPX+YqJL3WEVoAEWuBk+NsR22edqlgwYfRhCx5z4ZDdUsS1qkz2ZqyCM+1MQkCPA
TJZToOfRoty6tv9URU4drDSr1BKEUwUHj10NhwdDlLoCx712VlEUN3GpMY8pDs7S
vheSg/q6pILIO78X5NjpJoV6gnqOoBu2r37ZiTfZfu+MMQVQzeL2nRAfm8H9O+Iz
rmhOgrBlSK54njhc3HH8rZWXA10xlw6/HsEUKpLO5Ne/eYhHrSuSkgytoG5A6+By
Kmn2rvrCXaqVWcWDlTg2AdnGkmaeNmQ7L1TNL3r6CNGRu8sKuNkXt9Lj25DojMqi
ut3s45JrNAwglfXOqd9W9WmLNxorj/U3AwnrjakFIfhw+rmY5cSvwoJCClFQp3gX
EsPm2t8+pVeux0iH/QcJrvmlh1VXZ6OReHzCI+eelvuEhYuM+kXsylrIaa2g70tB
otD1eVoI6TwCHDO9O8MrmVxcvxoCvUkcT21/xI3mO8n1/kmoh082uh45GaOoFaXI
Afy2QTOofGgnt94b3KBtwX6Uh1sNnAoyjboaXgrkCTZh7HfXX1rKWK87IMV9Semz
RBLL6KltdoUXaPIzR6Oa2BpISqPkfK1Vh/Ac5ueT3fUp+VqwGoqCglF72fKcNFWw
xY215ropPFcRqL8N4QrEejopIvu+GE8BW19qsIfhWpA247zQinSEiJdLWgeOg2qo
0LBRlMDI5a7r9qrbjL1c8dcPHzG9JfUfs/LDgaoKGDFOvMD07yV8Z+zlPsc7vuar
PO4b3Nh0gf5KobzY7VY6vqVNe+mWy6FKJLiNahZlTU1XvQIcPvcnYb3aXS+qWOBl
+0Ae9hDw8WKzm25gNwNZKADr8bMp9QvYHU8MT0A6lToj7EkgPJ9j+0Ds/VIWSiQp
gMmBxDfhCzSMPfKxQ/n8KVg9qMQORJRHvCIEYRAD01cPHL17QDo7TgIfxcRycotX
GIEmf/ZQvOa0iJHX0KxbrXITmuk8NSYvShHK9vJVc2VKoIJo8F9T4HhrhdDsKXuk
OD4V4GgArEIN6WmloCkJl4FOW8gaiLv6QEJqRTqjVr4k44L833dGXxp/nn3v7gJq
p/8wxQRRRX/vM895zKiw/iroonby+cc7PVkiLF8t00oKKf6x4xJwfeEx/symvhUq
kHQivi8JLDzC2bUERtiUF8GYfmLtChoYymHpjsQTUVhORtafDtafru3u8iwt+Zv0
eduJp4iAtPzNHMKMShMwlh4DNZQ/Qlbw5/tJgPp7ExHq59rTpyRi4VyoHBmXNmVX
yy8mz8Sh38ihCyEdy9FFXd7obCKG6AAkG0C++nE3WtP80MRu425ynyGbkzd7TeWG
w+zHp8sEfpi/BAU4ESyBaJTe7Eb0dbyWN25DMYfrOjt0hdvQbfNlCpJk2OrfnYfH
UJYO8DqyxxD+/KdTixoTnHY2NDoO0tLt1utNapGpFCQqxL2BivJdq5qHkPVNwkVf
xFTdKaTcicHfn0TmwTfZCRODvSoJ08eV6jkK1MvBJR/yQ9bQVKIZIamuqVQnaXZL
80cXZlKYEaA5G05wGae2XXHV75UKzjQjzZf2YMPt5jT5NIItp+hG+iPqmnYPwQ1z
Vg5egn8spVrkx/x2hDKf2ZfY4QA4Q/P3mznUpgVYF7PdzPd+lPCWF8n76r8+Z7mM
wV99y7VdScx3D81SVts3GN6RUaPWX4bQeRys4l6C/rfbC9+c8CSNsZcEZZvjHp0D
WZOzqs5Dx/do7eMccVSCsdPp3ZCrKqG4cv9bhYHGWRwpaXhm3ozHRQsdQWFRoeCg
ZrmpLxmgV+yYBaiyYyz9jgwfIPYmxFr5HbtgSdwVFGNWYkQLFe3LeFlxcN1dRHmn
nqREg1zwshLZxA7RPJHvWsnk9YAtM+Urhdw5UGt6kzCaVL7izoKzl6RpGBZPs+Oq
ldh5AcNjP8da479f5re5rbU8hokQ72X88IV8PO+KjNlfalfIfCiWMu/1CAd140Wl
yakbcaAg9GDxtLKbMTPf/sxwisvdIugNyWVa4058kzEJzxN1pQRvkdYj5H2IGPB5
RxOqYei6aE6QBq9sV55nj9CywnAWiSlDsDrhvAStfUxAll5jtREtj1dREKubY7Z2
nysF4K+uDqwgV4mrDvG3jch08nAj2z1ehKNSi4oS6LjOXp8NEtQQoZWqLmKbDNsy
GKvCq0SA4PuAlWHIjtyORgMFLspct0wsPREp1gl26kKJ2pNaMq21CSbKg4c97Za5
V64zcf+NNJ8JiXy12QHos4B2DLYLiMMSpRFOmdVN2terhj0yDFIYmaBUvvpA2ac8
9mWRdBy1rTgaNo0lhDdz7LKapAHR3PSJPDF2n3zW2sdLm3GoIgtBAm1hGxJ65YMG
/sdYcbihVld2OXvcf0zFIMrrU+dNfL8nnqK0yVLBcF4NT0iF6i1tE+LuJCHmjYMX
fTAwFxT2tLr+VjW0TGoDRe70zDrErRd3dRGtAFafRyBGqOeaZK5KWs1HLiGniCb2
AND5olw+hhnh3JZFC3HibY9C+o9PK3eagKqqFwnJ82npqc7isRQuarTIfSUstK89
5j5hqWsWBBcxmSmMtX2o9mnBuAEcOaBNGz/NpOP5xPrDgy1uqCFhS8zSifp3zOqX
cEVgI4mqQozNHCBMUoUplaplqDi+E9No71cvpSuuo0gk801LkZ7+s70VaeDhrJnY
VX0NTDLIKhaI9CTq1jAORGxtdPlKkvtKN3jD+USruwTXRcLdGqCo6Dr7TXpodXcH
vmWqu5ts8qYiCyxH5yGlgAkWtc18jCyEVXyIR9NVjlR4VbzSoqGC3et8biN/0PUr
7d6FjkIM7ZilK4VEhcwep1pvlW0pR92AgpZDFMaQDubxBm0JDUEfYE7ebTPhGHtM
3kBuqtF1HraN4k0jSTvW2tU9RzdmqrA9xBYCz3Ve+w6RuluLdyXGvDuMdlTzWTOM
vSKizzu7Ock7gz1tBJqZbVx5UDJRAlA40cs+3TQdB9yHZIwdFHG9LIVjI8XzUNZI
aW3f/sgOKoghvP8cxPcKrzh5T5K4oe5rhBB7yp3pPm1tmXDINrrun5VeGwm0f96c
Hs9fzi4AFQcMp4aGfho1BNZE4US2GMV4gJfk1ckqLP46WRrSh8nfk1DCci5+foxc
DozrYdHzdchWXMWOEzzgfxjRRu2mgA5xXW6kwl70yUrnFm9wOScxNTGbqGLcEtB+
S2Ewp9FbwFEYx8Ui5SFKaZSIYgXcsJIf0MnUcHCBvtbUiSjO6WL8zgtZlYyaSgAf
Mu0fYqfuwdFuDAVCDz1UfE7x+DNyACoMtIWCxS026zah+CN6xb8vLMoiE9Hiejze
mj1Nu/jwyS6dIft0IsE7/OI28iNyQ+Pjib4Vn9t7aEQMG+8y3RrxpEzKX12BXHMv
Bl769TOgi/iYghbig4/65qr831wu5IqJNMfdc4/4yKCtAbB+Un0uem0mkWuZxIUt
qAXWh4v9ASmKHpJAjsZ7bY4IHTm84qreddazheVpKUmxfMRLQxItjNUXTqg9Vxkz
1e4lalvy1fJkBul6UFJ+46MH3HTz1axnk2R8m6NucBGUTfC2eEN5U62TX4jJ2RZo
ygQ92XYcJ/QgrQB0XqqNTEMarO11I4yHaXw8eo5X53qrcx0tzMJh7AJHhQ3iSe7X
2NHLIZQFFa77+QsHIN8+v6ncXH45C5xpen0tsBU72KfOKKeTj2Yx0louTArocqag
C5ALLbPdQwm2Q9z7KkmVp400hgRmAm7lG5BWOYiGhDjpBNJDZRiyl/S5J4gF4IRM
O9nooopKMt80x0JQtP2USPWn2u8k9c/JTeFhWZt+wQ1AOKomCxz+5YQwgLt7jA56
fP//f6+HaOaNRPEag9uqcm2U+WtAN/OQ2unnH/98pFktMzIAGVdnSsNRlxPejq3i
R4R358XzfDLPI4V3K3R4rPFN67d4fY26E/PyGQ6n2TjjDRrJ2KzzaBGqbMkWG9DG
ZrwF7stqKXKhil21plys3DEwn3OXgoYgu93cmDB3TytxiEQ4HTf1R1zbylaTI0NM
fV868osOimO54W/slK/EObXbZZW3oYlXq51lkeO8mEA4rUTPsnuTiQySfAHuFAKB
82g9XSTNzw8aPbMPOeHoxEg5vELNkrfvWr54cum1Oo24jzCdzUqhb1dEVatd4Z5/
e90FHBpTyf1WeZ6mHO8JYcEivpqHGCf/QVmqPhXbi27INfDgBVg+Om5V8UyhmWcF
bqbMLREmgCw+CDZT2m5VodaQzk9aQ6uxYMYUt/jSM18B4ZPqIeq4IS8GejjJdn1Y
Q481JTTUWZSfpLp1rDsh8t31OEdXzaUFVYVvBFCCaoBQ277kWErqewCokV5sX8Fb
JwsmbsgEazmA0rlfJ+fgwBMONO9dGmKhmd9QZF3j9CuShzdwTLFrcCmMfTbUs3Qm
X7ZOnyjbIAz4OS3J8mFOvbTTEsN/nfhCE9J14le41h7bit1Y5kQqmHUKIPSgGE14
N8mGSpNq5SrjVPqPgdrJ7ezg/88Alj0AV2oJ1wRRX79Ye8c/Zrq8WdLjDa72TQTX
zVhbZkmzRlZ62BmaFiH3IBX6ytbOlnLDlNMQMqrkWr1XZKuvqzP+9wWmuxvte82I
L2WOdHqXWZOl7ZxZ9kXCRwG3bJBannnqzqBmHwDItijEAnmdU2M0QW2CVpGAHqWE
LXcCmrqmSAn0to++gxxnEjxqJvsKRQzs/vb40Sr1eAbh/5KCizhLUZzW5hyHLSQ7
PwsIaRwuS9C0idGITvqroCOgkx+rfeInj2VGS0bfYM6dk15a/naRdRiHINuzyw4A
WAycMjS5m/6rL99PLVFWsUBdlmc8DHAvYFV5aH45hanBe8/2GwkFWaeXV+r7EhhR
Pjs7wvyd7A9iH2whv5Hl7Td4XxTgVzElBOMfRbiZl0kT7UMXk6TrS17R7VTeZ/j7
XL42KAoBpKDnfZ0shjmjihGMkyOt3gIsGT0ZKeDrx6jXFYmognwZ+vpAAjAfw10R
ZuVh5wW5wm5NJ6Y6CSeafpaIeuUsxDlAq0kk41P//n01l4gFG9WLXUtiW8BiAwVq
EGoDpCOztAeFnlZ3Jg+xD2qnrNi2zPYOy/sYcyyPpwU4mL7Z9VF9AAbU2Y9Lx4lN
eLMeDQsp77zqxXe4m4xJPgaLHsNR/1jwdVyPXj+K8I7b9kCfCzBm4yv+b4hY4bxd
iBKe7wq9L0F/bE6vcQUc+Z1gTSwzOfwksWUey9Kfpw3vD2TIEyuWbV2Vt1E1ngBT
ewOifN6YUTFt7u6/Q169aVmKhIpFhyY4k5szOkzudwp0N0vmktZ9alE73NDVM4CS
YFLXws1/Epz6x4/G54kCw3QG1pllFRbJcqS4S5og6UHKBjFZTL+Fd8Tim9sVRBXL
hRrbDx7JAFXG1TVDlinJ5S2KQAemXnRkTvrATsujabP3MDo1YtfCh3ojGiksWEWI
bCDrZr9YlFCfc38NJNC1+Alg1b24qp5xddeDhOBIXTq2gTT3HjgDj+VDFHfk2ag8
jP7YKWe75p3rL7g7MnISu2Y7+6hWm5WEi8Qzx9+nI5NNhfuzvuX/lKnkrq8hH1Ic
IMtpHCUpugDZsSSCtocS286qqDbzJkRk4IYjxVRPGsYwiqU83Tt+Fr7poqYDroBP
mvZniduJU8MiKJQFuiGZJC9zSzWCh/O0R7rpT+D8KZ4Oh2Qh7IhUdDG37L8Ig21/
YzLbpjqqWQMmTRv98+ra1dm+xaDhAg28LyP3Ox3Ct+tuefkHs2btGdIP67REKaJi
a5+hdtztpxwRo01uHng/AshFQJ0cJjzd4M6KGgKWVyF4OBUf4iTGuXVh+0cHqehD
Iy/wUDatKELWEL+K1R3jIWsk1LCc+MarSdnuUC3G3L1ktdpqaZKe7N21jo/iQWMz
fpIuYPhtWccSBhUvSZqVKWLzJ6q0Q/3n9/2XYw3B9O5yRBYZMGqQvGUKcgecfhFX
BsanvV3GmcPFvz2o3LuixYaD4OOpgT6WuQQpLYUnIMnvT+db/iFPwSvexde68ANs
ERukLBfAnIcSIb3VXd1bcZpIOzLq/4ijEuQc7caPD001IpkQo2T3X7vF3HLsJbzV
PPZsn2V5PiiV7aDKGGEm/3/G/L5ck2+4byrIefCFmSzU/4eqli2WdUD7RFEl6VRJ
v3RxMIs93EmchqYVKOrqHio7sKUxTC5hW9xloo2WJ534HN98Eh3oiyV6tyaNAlN6
Cxuue5jkK3GOH4cmKBdrFRCznlKzE3YfteinI9v6/o2i43f2+Z6w/8rWgyVo0992
Uuh0f/5XMI9+9masVmzGq7ATihOcdzF5y03mSLL6dOOMQRK+sdA6NgRrXVgy1pQb
Hf8q9dWUJTl+Xt441WGG/UCpvmPzUrNGS+mXRt+C03Qndk17WZoUf6KdMtIbQap0
E5bmCgl7jDNf9uQ9GZeWSGcLGeI1Rz0R9eVTqi+g1lTgwncQQMoelrTXmWqYPuPp
X3NTXEL5It5kdXWM685EnHNj39UltgVM5xEWx7uBMuu7h9xSs81FphALXCcVUE48
WC5PwBGYJVoaJDM5Bdo89MenCFsIcgvXorG3eOnw4Oq5rx9+IpXnScdrVyTy10AJ
wCq7garBr/nZGnduypm/gGK88gZnY1AsK8bkwbefZIjYSXGkvYTmX61FuVXa5ywL
Q2xM69ZJVOpeDJlIwqUnkXrVaKXSz/P4hARZh6vLw2Ir7zRYx5HQTWM4J/STPqfB
dSzZEzfCtbhiKJXpI6l2GoviBj4ItSYAuRZfM7bWn9Vspj/zZen0/0luyUCGB7Ty
8+JN+11O3sKsX/Yz5kwoUqkJ8XjiPjfLV94q2CcI0WFBxdK2fK0uxkFgYVJ97jfQ
7kje3o/DU3P6vVBTGBfrUH/D+hSOCRMXt8s3WZNIGnIf0j95gR7CrA2N+C4rQLsK
uKNZvhIlT0xWFsZs8ttnvviu1l/FIU78hLMjKF3QmQyDqvoh2o7lWiChSNQRbUti
lOfyxb6At+BlIrKnK5AKdpHwuFeC/NNPMGlaqdX096QFNLQU0FhyV0Q2/vUxDjM7
EMCCTIrxXsFRim4iKFDb0xI1hh2ie6lw4rJoHlow25q8HQCyhzHGW3VdvtstLMTb
fcInC5LBqNAZvAswDgLr1b/DhDf2OWaYyCgoWOQoi/6TjGQX3JRq5urDaH75FeD6
3InrsIkEiKSwdbe7UjwR6k+zXI1qEsHTVUNyxRSwL57zSYL6Mc52QtRG2kmIr/qz
EdXSQI4EItjeL3jpV21lD9jHyjQVSOcXj1TSwXihUR4EcriHinc8zGKf2y8N7nEj
Cic+Q9ielc0Y0/wklCNXnPLMOpnaMIGRLKdqLgWwV8es/pZQ8g+ws6TVxAYlvjcm
Bj8k16ZSGcJ0iRmJQPGapHekIkEJbFGtcheNFycHsGPCzG2jw7tPSIyTeYBGV2LH
GjXzerFiBFdZfuFyoulgfXAZAhj3tG1hYWivcqN9IBXgRO7LyCO7sUT5TNhlMT59
yPlRL35kA7PfJdLrIwxr6w1269QGalkzLN94Mm/LkhZkQyqE1wZhVVIP9JSQHpZL
0NDt0dYZVTkeknjFcyDjQM1Aj3xGVu9h4GZ1VxkHweYWJ1KyOvFoAjBWM8YJ0hXz
O9YEY2WgEeMPR8gmwcXFLdaaUcyz1G+ZS2O3tR52R0b13df7zN2ugAP4a4swpwvI
jqe4U0Y2jUejSmxVqZYDrHebXd5kzdnRyCk5w/BbsJay7qApY75E/DLxqNWQcZ9v
BSG6P02jPlIefkwSA6UAAP1/a+xB/QKaW+2RtfrdUms9HJ7bL8VSe+co1zuHHDw6
3reLiadxsjX5IK8P8zfC7COGezze5kVCuxXVaiUV0PTznvG9xUxx+QfFy1ZEM1CF
`pragma protect end_protected
