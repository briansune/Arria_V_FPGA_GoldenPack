// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
dirpIjc0cWuACT0zSGyy50Fm9nmx5PooWqI81VzctdW5hHynXcILeau2SgPSoU+ezoJOIGwhO5gO
5RHUdcH0qTVKN5UtYJRgMU0Kzk7g4h/skOPqcebpE6yH8+BGEV9DtgWXG95kqBZ4tM3fzHVJRKow
l42cqgAmuQY46hVOEomZTrsTDPiKOOfaRGjElPqNiQCVC5uk8oZkXhnJ6z5wFIvmPKckTnhC3vQi
nyGc4cXASI/7quO0X9QMkMt7tVd3rgnU6PQs5170AEcAsapz3Y+Nr6U/CMPxFe0zoavZ1zZjNvI2
WXCjWk+2qXCK13ekysm3us/Bu+G3YckkOv+InQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5440)
aJtlgm7Pv7R5K/Xf00X9N0asj0InnEHQPybDXAbq/AtBbL4rXcFIu3CMMzqPSU9I/5bJnkCW/6IX
jjsZJiSt/Dp5npFbBcfRQDy8hqOaGs0okkhk7aWc2P0KYpMXNr7MGj3VAh4Dz9rHDPsXrcQYK5m/
mxy3q79+Vh6KQsIx33L9QaOgWjIwOJyABDxZHvpIKZILBF84VkZ3XoNB73NKJyW1FiHo/aoFsXZN
WJi6OwAD9KO5BSWJ/FFbFPf1V0M+9Ip4uu8MS6W/y/TMF1qD5jR5cZh0P8/dQOoj+tuAznK9Rggs
b0HNR4qM3yRYPnqA/PrPIFMyC4C+7Z6hwBIAaJF8THL6U0DUebtIfn2LH9w2GppcezOY03e6mGWy
PYYB//nTsUJTzGXOEusL40vBgKOK/pKsvpSgva20rFZXGJlBRgh17BvmDkbbb+hN+mu15EaL6ZmJ
DIzpjlTSnnksW3P4ndCVpvdfqv4PeF4jWxwPJybayhoGfPymZbVKdbbSeMNaCCuq90FfUo/l35H8
qsxeRULeK/Umpvd1rIC1Nh5HFaxlIKbH3bVvc5+DFzfzyA+3kEi41B2/LxPp2sOlzza+tGIb7alJ
inRhAi5k8wLFGKRvdK3+E0O9SxEdqWvlJ4CjN2PvfYmZcsILBV5OwsTiwiR7N5GGKwd+1pQEKFnR
WEHybCvZJ2i8X27ItTmZInSjaMbLdYWLgn/WmJgPZVSZnN41hScXlgU7/cpZrACAYFHkVAS4P0D5
e3OoeE8EuDeufolEcxR8T38CTO7Y3P7MtO+8wX3kSYnWqENDOCuJWZ+Ws8BnbqmeH/BDFnBs4W3c
zeTyhT7r+iGhhJnrnH7M+Z64SUWF8rIDAcOpaV+TbhUteC6LM/gdAsSfT8pR9RRqyk9D1H9R2fPX
qqWlDvjD3tDTs0zDjaFyOZoIm0j8T6Igj0S2NDQzhjAJ6/H6Sk1+qV6Fo/JaEtbX46prXv8Cxew9
D9ZA6ZF/N76LkcbL+/QpzXxaamjmFpOKemgx3hJNAUSB3Udqrd1CsbWircMgcRVo0OD3lVQxhwQu
GBK1SZSy6esRNRYuojPeeHdklX226RGxhV4zqSnLmB+Zb3BnZpg7q8mWurLgysDwVzqxO+0Rhu15
1wmFNM0jQXpw8QwpCD9k/E7DmyIFyIF0DjbyAwMqn6lQ5Fp1lJl7bufXNs8ABxHzz/egN3NwBlJ1
6Ojai4m094qpKgz9Ugv6Le8ICjltguTwwi2aSmkosADnTsVh0ZCfiQgzNq3/uWHVURhKTW4hKNCE
CS7LZunTEEKJdG92ltNkGoYaBZOlXleVf6hbFw8l8/i5atvOJ1pUylNMbLYJyG8/OFp8CP9B5wyB
t9rcAYpaBHcKrGCN84h1YcqVdh/fRrFnADII4P98zjTA975p4urBJqELqAg52W0mTl5SndaTo3o1
epaOaww6eCzR5Vl0EwocLjTemO8uT+//wlV8/Ondf6iNbFqFjtLr6ndUtTQXYXHN8JM6JXermq/S
VzFPeiSrYz7gWD1EFeedPwi8vbckZnhFMrmRP5um/CKmwAE0cO9oSmE+i05lSVkH4M9OlXdGpS9G
PwlC/5CVDhwriJd9Xaz+txAhFzn82d8whQ6krPRiA5ldUMbwyT6wjJ81MfC4yGSMgdAyQT/rdmlG
3evkEl55vGhvt65CRmqMBOzF5dj0FmYs11jNTqXG9192+sc3L2kQ/6ae2RljNSVL9494qHZavoVz
abjITHe0x0rS8AD3qTJ0oRWGqYyf1faaV6Hjh5uKqGhxtxKitdYwecWbOZ8xRqycGvwXOKquA2A2
U0QjKdrfBeocxn5lBK1Wr+oZPGiReUyggDK9b0lc1EQBeAxmgmDONktddTr/lvI+DtkLAmOcJjkf
iI+PODKq8NbnYiGsZBAe788+rT0jvPhkt6ZJsE54vmfGLWNK5BZ+EEPS4oE9VBpAsVix1V2QxYpY
oa/8/e528AFRQbsx2t14Pf4BDZt1+4pEdXiiMq/d0rqzcSiL7EpKfmAdSdYO8HG4XU4e9zegAnye
NcsY7FhjeQs2sdO66qC8ZVH/6ECHE9PSu97MnqobP68ofkyBBuFYTh/QWWXV9dsbQ7OqHPSp/7ev
j38xYtGI7ZYeqFgm/6WdbQy7Hx9Z5Gt8kODQzFCt/YMMMhn/8gocACpYAjZ7aRtB1Id6BqzcCWvd
fVSGnRTY5xvd9Vv4Sg/wyE4TArNwnqXI+7s3vljfZW204FrYDEh/STi7RNkqz4U/q6DJTGBnApkO
i2IUjUAb8YqvDLD3bsyfiW9dGRARqDC5PNxbZAwR4UitDzenk4ROxMJAAbQcc7p58dhq/VdlqOlA
Lfkp99WnpMz8GUQrpkiClr2woK7mHqMkOlkhpaGSnK9Qk6J5XgddJQtoGs1cg0ZW7yigEMPCNZFz
DKUbmpwNIcIrWgaxkDb4npxgEVDIMMclqelTXhYxAQEN1Cgy+PQTVioqnv/tsSGQiXL8iSCJwxJb
aC7TwROlyeThj6Ra+pErUTvv7moeNdiPKV/cnnmfyl7xpMcOqkrBFOrKK8vMm55p93ymhlD7revH
Ie0RPxBfXvZHCKMD0qH0enIcclQj+5/VcCiQbVymnClZQjXgggr/bMoY9u83JYW6UYaXO2xCFlPm
kTm4qMTUppNWHTd4LrAYIQyUEU+TFmFjPahdG61bGOiNkvqBsSUKgGziyZUdoOqHVV1Cq3SjAljg
TDFFhcGCgCdkIwsVlVa+YD0ezghRbEqrMxLF5GH5HpVrlxzH2ny5tku4KHcL7IFF6mdTT4HSidzQ
HdFbnBixpbE+2Mv8CmFS4QFsOVVKJq6hbXCP/tr+OVlnJO+GXM/7tZ3LYIZ+ktl0edKjP5bjgRRc
oZqbEMflBEHCNtb6iCconx3pCvgZLZkn3puGVlu/vfip/uk+vLmSsnvNnyHhTNOYPat4eWxuN6kB
lnD9ZQK+eiilqvoxPNlANwy35RsPVrgY21wFo7OmSliYRON2b2rPhHZRJVyFKAs6Gdm6F4B7EkGt
Z9QOoXPmriD1nPnuP0AXNGT4sEjpLOctdLestbnpwONoV+zAvZRCS3kvoNW6H/nxELcZ6qbfhjDa
3czslzjrIdafCuFnL85BCFrbRSbzGudb0LzMzZHyeTNnw9U0z3RiBuM3/Ygygi+1ZcuVnKL/WlG7
E7JyIwF33fSYN1QqvlAHZah/f+ZsFW91PYuFBW9jlQRF1PA2hRU5/POpIy+dCcH5Qic0wJytlR/n
MQlblVtXttyCYJ8tqtXiXB9DhAWlnoyQ6w628yqivVRjTOpPjdUTpauLp6b4zyxK37rVWsAFN5mV
2n1NzOZzqhvVu3Si2Bv0Htrh/iUC6I9+CVb3jIuN6E0VoDSftOnCuy7y6K5HPnUPYpVU7avvTlkk
0dY6mHShBMgX9A8cH7y1OF/Y9RC58rrlo6Lf7DU6G0O3xtk2kX3JICxjRYuVy5u4VIuLs1JWJRBT
pRqs4fphmYZLGqnwVNd2Jqy52XdtMxRehXihv5tWcsOT9YcPGFKR5YmMVdmlEnawUylY0Iz0s5ZZ
gX2xQ4Ym5q6v4sD+CVmdM1ZdAcpsqGaxbu37J2LqSxwr2lmINn+TWqsKQQFkXny6raa7jGjtIug3
25P5L5ZieAfpbJAVS3bdTHEJhBQw2RtnSnM1fa4LeORT/vcarEhxKofT6YtQoP5PcQnH7NJ7Yxn1
06aiaRHeqNsJn6DySa8cmizGTrIGtTkJGbQwTyZOhM5dRJO9+KifRwmiBD6Ya4soZaEwV1k04Pr3
auB9f7UsHq13DhhBDchP86T/BoU61KoCfefD1ww14vK0WGUD03OWf8iClFhiHxCFCGeDe/pN2F3U
MHaomJzdThvDzGzyCPvQ7z6PlHxFJOYyJrndRFd8IapbKZ2Jj0UjE6mq51JJZL2u8LhpPPcmfzTu
sh2woKOdxDN6uMPfcAdHr7tHBTYQOFeek/rWjJ+68VSv0bhOdm6DpNuXBFtWgLcR0Se8InvxCVfv
MT60+22cEWUI/A1A4y8kSBjelG/n8bnktMHLP7k0e80EqATN3XBXUDE659kbqbo/vhTCXY0QKqF9
wIU1Zn6FZWn35mVGHRHyoOdg+xS2nCQ6nXtCq09cWHp2qyOn4jPTRMDqJbuzAKLfjzcWRTNbq4DS
htLBx5jONjKOuJ1a31V3NKCQ5g7mSWYnZbtGHDTEr9C6grfR/fVRWjpzWh7gPtcMLeR3dlvo1NsN
ohzifWuh+2XWEkR1G2jq/w6s78fdzHSVLggB66Gd7Wz+M4oMdDu9qPzccE/XDk+hgpC3Q0T8bvdx
Mq5rNYMHnxpDaU0JwOmMW857J/Rr8JC0KEEJOWcAVDjOWb5zS25zYllCToG4QgMQG3BOmVtLPteo
KMbERl0V+LFn2Q3sJsiHwFXaxwymfKY2zg4TeEadsXmEG86/aZYivW9qdsHKHkmq69ukPix/gukM
UHYv6wESZLkkoNsb7R4LqVpQKtjk5MMsWIcbPSUcM/PpsgB/nQ0LjzsrBtFzG4LqcJ3HUovlMBI8
TWRGsyjNjnaTOFZ7lyRoKdvYtpwiM5sLuJ0Dw9JepRg7tZra9RcEgSULJKDCzldseJUojc5GROOQ
Ja1zwzdf0+3v3nfSBO9bUzPivErOb3S6BFNAzAaTtn+rZSXC/qnAsC9GGJfCj/03pqxdE1V3LKYY
7JNPsY0FSKTWLd83RnRaknsFmeID/Q5hkngxFBQUOOUq1eaEdiToqmJSXpZgiUh8yaOEwSeBEWgb
01j+mhUrQ7j8hBw1hUeFgvUL+V2pdzHmU8ordOJkZ6WC7b6fTuvY9y7UBPz6ELk1Y80EG/5pd4sI
GjHlUvXtwKu++nAo2KD2j1hzB1WEy33E98R0ixx6PhpS7lHJkwUYp8wDbOMJKZP4aXnvZRDDp/bz
K/kzgm2JbfQ1dnaHNpVn7fphVarXUHP7e9Z16mkBHttcLtXIIrElQooWWYDqbXtepUE1JkreAZ2o
ASNPO5lqhDE2LPPSZmBMU/K6hg8m1RoTYNE4pJ9Lp+vzqMJYTMJsV/dgqpNqgAZK3Eb7AjZaFhcM
VzMNuZcFhg6tyDK1kVFqOuS/cjEcxcmK+lES08h79UY84nP6r7SCnDAmDQo3cg0l/WOCq9A2aNGX
Doe+w9ZbzJ1gjw091IimlhJNVw61pcJENrKJb6B/ryVXAO8lkeI0xvBjRvQJQzBX2j+myGILpQXn
SSkbz6wyiumLshBM1bL3bewrcaLazMuS2ePeGSx8R4N8CvbFyDLoWVOqfdjJV5uaT+bUDlFFevzg
s6ujYSWwx6cl6FHyZtBM077c1msIhUuB7arbm3JMUYOe1k5G9MsqjieBaQ/PrcpLWkK6RkADdHHN
aUprGNi+L6gD8p+LthMgi3I2ol5Kt8tzE1ZviwRrL+UitBpzDdXMVsGM2r9oPyiN2m1SlMcptneK
y+gQ6HvSpN/Zansh9pIk8HVdOeknLEUyI8ALvYxB4Dbe58McpNtE3mBTweERRcCfvYyCm5a4eEGI
p0mVFIp7j39pnIuJCNUVj4F1rt5M3Bte2qRtOap6e7bWApGTRjNZtQacqn+x5LkDO6jmYLxPPBON
k38m/MTJtMOW1fDoRnUVlAMcvw/kYUqmBlufXxzspr2UgAPta58GkB1odixAkytdwpS4iiCF1elF
hSCVs1nve/sfRVaOUdKxhpNRFlc2uCjvooRcWjbraI3lOFR1ydm0Y05nhRVmchoCzvt8qkwmPPkS
PD28oQqXG7rgpjMt3EwDMINF9Oy+b2s2CshD22+TnCEKe97u/ZJK+FRwNHOogegw67RDc06uBQbn
THFuUEynQhrS7ZrORmzGge07xdwgo9FOMMM6r8YhirGnoQaxzGgjSytiK+/rdlL4/BVSjq1kMtVQ
d92iO3WRsayCVK0IL+0PwNjGNWP4Xe4YdBsWk7s8vH2lSMMVii4rgvCNDYDWYcrUiduGtW4O7XG6
qon6BxP1ZlndXNbZQ7iqhj0C0U4Aga+mcyhYbVYb5RuqYCO4Ue8F+S4KSqR2eP6P+BcFpNEjeUfi
VaMWE2Sv2Q4uWQavecqACtMhBTQA5WGNcjC7rr1d7etQ48hQR4qeEAbbQC5pVAX/ckQ9y0N3mAu+
5avN9bC73EjbYkO4cAN3W1gfsUT0VIoUGhuf06LVwUTGyHRYP6yiKz5U0Oqq0sGcvBwT5yRaVlFe
/y2K3bfTvTp99hRU2EwYEQ42dTn6MDxqcQlstqHZ9B2MXcYjrAIUiWuRC0g1YLHP3MCVxeowgGsm
wEQqwSEifUUGB6hcMk3H4Kr32DzOKxROhHhWLa/jh9oj315K5+j2+ubhRu5y1EZ3qWKF6I9V60ME
K57ngZm0onmo2BnvgiIUJBvDcFK51Tb1LNeBJojkHSg7cWsetZOPpmphif7uNxVIHLhoi8J0nTkW
1RxJmTo9AsMdMGaxO7LCkjCcUP8o0Wv5KPTlBHmqzDNHPHlil9ZKeRl9rDrCSUxEt6v3LQ4UZ4fw
drjm16N1P334Og5XvYonSSM3bd2kc1CmOJzoOK7SCTNHYGU4iaThqlhgmKbvA3TrpymT6MOfJAuD
H3FIcz6VXAf5aGJuVcHzS9JcrJg3ZCN971ljjafQ4BcEnCG80LSZEbKc9jZK3XGcCfYb/6sC0uoy
Su1UhZGK4XFPLkediA5HrIAi7BSAH8W4LkjoAHHGOZlzVjptGNmR80zQ0aJiXbxxMFuZY+gmmqFI
flftk1s92Ni3Bt2OUrf7RCy7vX0iA8XM1RdpPlQ2NCltvI7AuKgcTrkkmF8Typ0Q6EDobwVUmz5W
/Qm08FSX+0PFxJKE60i/J7iegKjOhvgbFIJAHcx5bWPMiiBW5i8d0t8BtCXSjBTANt0RyxkgZ+uK
RJbyo6K9qS+Cvp2HVRdQCaE/KzOwn9pH5FC97xHNVBHtE2n2aXwAVfz0mePcd11CRQpsZpoK7lX+
/fFDc1wjYvxR7mmkN027rXf6iBp4luKDVjCYf5puerWkV/CjNhYKU0Hun0JDb4cR+dvPoUjlNqgS
BsOAtQ7KEhhGn2UNzjfdB5zF9iSEgtRPaqVF9gq0ZHvcfOCE8Ppas7XGJ2ffS3HbN08NCRvnRFKj
4Z1uCclNJ7MOzl7VvQ9gwnHPDuHjh15f4f84mZXlwgP9ci/0c7MMh/hYNDsRRjz+sX51D3GVcUcz
zCHsSskNcMSwGgXqjcezJ7hKmaPZu5Utnw==
`pragma protect end_protected
