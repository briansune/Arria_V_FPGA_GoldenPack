��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t�6$��}�e�Ra�<q������(2ߐuoR� ~���1d���e�|��|�oI=E�={c�Z�)b*ȧ���DD"&�8�T�u(��L�!���V%@�c i[z�W�g��n�,TI�|����f�_�-')8hj�Y���	AbB�NH�.�$H�cU�xL�A��wA�>]���}l��>�����^�8�w�Z?�!��"4�vx`guw�w_��-�mU��0�R�7�ڨ7�1F��\#�W��3��n7�s�ʞʛ׈��5scWB�
��m�Ɩ��I����B^k��q3���AfH�c� �gE�d3���[��.t�=�	2���>Bɯ���YS��3Frx#���خ�Q'�-߫8�ϥ�Щ�	9�|�U)�z�Q�����#>�߈�w��=x�� 7;
�o��!94Fbg�d�(oGt�M��y���@�lIn��6�U��7�
.�J��X�<��j�� A�5�}b���F]��ו���N���D.���M]�UO�Q����v
�#E�S�u#�Yp�X=�薉RΙ��lD�X'�Y.<"~�;�'g�BM�/}Ͼ���s����\�/IR3!�y��lD��N�wM� ����-�ϪO�	_��¦���;��8��a#���Iqo��`��~(y����0�3ŏk��eP^��Awȍ��u��I|���%�ҕJ�-u��?�k�eDި�`_)����
�vg��v�ՄD��/!/kr����k�(�¤:��,>����!"RU��\�/=������t�J�����xm��i�j&l��l7�s���AY4���թQ熺���؉^DGŎ�<�2Ӭ����za4���&Vw�t�Ln�7 pmEVY�5����O[�r�v-p�{筅,�䆷��LhV�j�<#@��+2+t�_y���~ D����f˛?���7-��3�J�	��K��C�J�	*�Rv(glgnA&�e�D,�u�/c��w�ɠƵ�D�m��X�*��H�FK��"�'Q�~g���N������èf�#w�U�� ����~��:wWo�Y��Y�!����Қx����@X9x�.<�R퉦=�����UE�9�_V8����siX�BG=ĵ!�����.�;6��4�Y�V���OK>��| K���G���C��z���Zb����%��Hy�N`R66Oک�J��C{��np����1�\�ʗ�zUJN��۾��߄H��@�@<�3���p>�<ɱcB~;m)��*�N~c�_R!������
�y`�,s��pj�����Wd���Ŕ�^´�=ۻg���cW0�B�X	I"f5���V9�;h�dO���^F��A�]r�<���5����O�y�Z��Uv����@���{�M+$���6��Y��|�Ҫ����}��vbŮ���"y�ߵv\=�2�v��d�E����ֻM��o��1�;����,�`�ޢµ���0Q��mb���-�̑��,�|rE�n@禇���w�S'�,��-_�&K|�-k�=cY0?�	R�|D�J&�O�z5�0��v��y�9^�Ua澓Q���g�@v�*{��f\���S��{�p�P7@�^g�Æ�$x���~/���x�{�Dl����}��4X�-�%�O��{� (�L�\GV��m*��(r�8��?S��c@���Q��LV:��� !�}r�N,
\4��at��U�SH&N6�5���~p��cZ��]�IW�)��k��+d�*"(���=Z���х�'ȴ`+F�)?����K���9@S����O�]ϕ��DO��ʟOD^#���u�pꬣ�#4�����B���ϯ=�������՛��^$3�^��٪��;8~	���('����4����O���c�7�� f[˥����)�Zd��)�GPkRIʪ b�K�g�InCk�F(* XmMǚ��Aݙy��<�6��Щ~6��M�Z_��#6%�SN�A��Q8ѻm{�΁���8%h��X��@��ax���|�?�z\4��̍�,�����5hb*26zO�0��^#�/����Z�F/Q���Ժ��RL��u�F��RGю(���0�ק��~���� �*a�@���>ER��Z{߿�[�:[��A��ː��'D�EB:�T���-�{�`4�b���V�Ps��>���ټH��V
٦X��V	5A�)��4[��;�$�"/��0�|ލ�hx�s<����"���}b��$�D��C�)��L^ذ���9�-vI+��6�
o����5�����o^�u�T�{�#���Fw��\H *y��ۭӧR�<L��s���{o\���<���k�n �j�V��{�L���u����X~��:xϪJ��I�bHЬ.nv��huغ+Z
6��r��Y����$�gS�~@����tQ��37�����n�H�2jͅx.C�[���Du29l4K(��IH������(�;�ڦ��4&ۖ�d�h��h9}����i���i=)�S��|$�����N�D���v���l�e�4 ��׵J���M9p$����AEA� &u�����NYޠ`+i�A.�s�2vu�~2��@Ni곜sSRj x�n����zq#3;�Fk�"F�E���Y�C�O'7���� b��kC��T���_��� � Hd��jS�ק���,9������ P��]D��7f��7�/-�:b+���Jf���Ѕ�y)UQl�����r��l����͙�]�z�;����"��t2�ߙ�'���M����EFЍ�3�Î�K�C!EfQ�L�t�j�qlY��˚E}�w�c�A�Җ�
��\�m�a%(B���\/U}�10���J�\O����=eE|6:��C��N=�@�ݰ��S��S
����&x3~ɟ}1��|o]�k��׳��35��u�o�� �e�Z4-�t�F���)b�����/i!�@JT,	�!6�m���^�2��2䧞�g@sX���J^*���X$���]��:�1C�_��x�b�X������d[]�M��v꓍Qɬ�!�]�GV�������m�N8�<�m!д|RY���$�:��øv�H���d ����6�O���&�5<CM�!?�����^��.u^�������
�EY�����S�]Zm���gH��m��󛑸�}c8׸�1<�s\y�#�վ�/�TL��LY�XU����[as�nn���V��}2��9Q����{����(H��(����U�o/����zZ�� ��Gg�2�*Y��h|+%�s̈����ͅ�F|�\�������kz�b��k���|��k�3���f�@�
�ngE+�f1��2�	�I�X�ͥ����eC��f�@��n��~�JJ�Hw���G5�8uQHoP0D/��s���<�,�$�� "Q���
R�`�'�����}e���`�Qpo�؟D\z�~�K��W4x2���U�mh����~EQ���� ��Fe�ݲ�u��9H�E������s���̪� �	��8��x.&�-��q�H���	�eW���#xF� h�MXH[���<��ʩ��si}������Q��QT�\��r虘Mg�K;8��U�[�+ү������o�O.��*�ӯdyעrc�K Ax�W�fҗN[�:,b��\H��2�	/{�3(�����������|~1&��^8�ŋ.NpJ��t��o��	�@�b������o�T��5�2��(���W~gO���b�,���`NoL��v�^�TBh���c`a*����ҍ^O�m�:�cUU_#s��Z2��[�48Z��Bh�[��d �v��#�F����������P�7DDK��t��E@�^�����.P>N)�E�*Y�P�ZF{�T=`#��zhF!�r��>��y%�V.�������밀[j�z������� ](�A5��g�*i
�����*�h9��њwH-n�y�n�����/�d�]
�ƴ�G� ��P�w$�P�ӈ�����;�Ͳq��_x��6d���Gw\��� V��؍��Yk%�>�wx�~A�F����0�4�âi��1���;\�`֑C1�
��.��IR0Y�^p�>�Ԅ݇j�;Z��z%7��N:|r����ϼ�	�pW�.��T9���n� ��+la�e�@2�,2$g`�A�/6���U鮰�}$��J�y�L�u�ː�i�P�x6�upB^IXJ���]ۘIr�^:W,�uY�w&��{Y(��ݸT˄�\��l��|dRs��ʐksv��1�C����r�Y����K:�t#�q���v��*cn���s.�[�b/N�_�ɝ�'��s,�p�#�Ug��bW�ɑ<e����<��1N���Ȃ�a����46*J��RٮN�:;F�(�Gf�22���֍��B�X�PbM裓���	9{��"�lfѯB�{�ֈT�6���Up�XTgܓbw�Th�Hَ*r&fG����ǭ냛b9�X�c�ftJ�W_g�W�;*�)vğ;���6s������͸j�i��=����)�����n8-�����F�b�H���r{���z��%��
��� �*���&�M�2z�k.tsP�)�O�h:Dޫ�n��)
�"�-�p��� ���'�t���8�f���2��F��_�D�ƗI�ʏ��%p�3T�Q[�~T�&�(��yYJ��ip���R��/H�mp��U���.�� ���0���|�:�ϩB��^� �.��˨�s�)lL��h���L������2����C�YȺ��4���?X�y��#�@����k}mB��T��Δ��t�6��qz��jb5�SJ��S��E����+1�
��t�蓊̿-�u������B,�69���;��N'
��lH��Q�7�=��n��t�5��#%�u&9��L*�~�	U����C"R�ԉ��CS�Q���%�(�%wޞڀ_m���d��m���f�u�sY�C<�q����@�q���
1��
��p��S3�#(���kC���`����%���L)~����e�1�V+�Q��;�@]�G�p q*m	{���L�_�x����3�K{o�%�/b2�����cm|خa���L}�=��m\̃7W]�e3�TV��g�-wi�Cћ}�̬�d'���	Ut��y������y���
t��C���`]���zo�mslN���A#Q\N,���NP�#~�m��p1�.�=ӌ.��m���"~S�hC����2��s�/��'�Ύٸ}��-k�'�������O�r!���\B��d�B/wI+��9z��͊@Z���ԁ@~�^��7�.*J�@�Ah�w�f<�*�>pѿx�=���z�y�I��.#�F}�!��ԋ��p���xSP��>�������I�;���֖(�k���
CI�ة�+!�b����+Q��	���ڴ;G!�N} %�ݔ�Lom��lp��[ɷ��ju6�:�#�f�������rqt�g�}�B�����a�N�*>R� u����#��4cK(w�S�'�p��W�K�/��V]a��0�J�������+�ia�ſ�����ݿeJN��j�~���N޿�?��l9J�d� ;�R�$�~����|��m��D�s�c��è @G��䭈���S�E�r��鄄b�&x����H?���|�\��D�$d�C&��Ɛ�����̨&
���!�=�w����-u7�"���>�\��������ѥ��D6U�h�Y1�\��y���$H���3���q��� p�(���K�� �K;
>g��s 1���p/�{��'B����.J�0��E1����?q�a���(��`���g��\�p��&n��b�J��`�T[y9w�;�\?�.���oa- x3�}�ҵ�RU�ƚz��7=[��#���e4f�9qw�+�-���Gs]U�O��>��|W�Խ�M��f�	����&<W�q�@x��v�+��6;~e\N�Y����w������� j���J�<�~m�[��*��<���t�_�+�iLagF
 �^0�Y^�aB����{��(��r�L���OԜ��\�� �U�Al�*>f�aF���R#�M�K]��Ȏ."����~4�&R�.��|5���7�r2\�K[U�g�Hһ0��`�w��C'�lXu���)"��-$�u���Z����\NNX�~`� j;�$�N��^���ѻ�KN��:N��T"i.2A�
��Dxb8�-�-�H싁�ߦ��z�@t���k���˸�b�%�Rt�L9!��sol���KL]�Ǖi��m��1����ꏣ�D��î���^i�.U4s�������9��?��Y3!��3<"f鬼����;�X6���t��"�?��@a��F�#m=b���z��	�?�Ol�G��!�0KS�	�~���Z��fߡ����u(@���h)f2Cq��K���3�&CşK���?�ZfD��d���%-d�_��U����zH��l��@:4���O�F��� $�yiz�����=l7x ��w�`n������+��!9�e�
gz�9�τZJ�C��DD̯��$6[�!L"1�Vxd����6�	\A,���~���`A�4�.�02�~grM��Cnʆ÷������j��?�<QW̺��lu�}M�m���t38��<��Su�n�Ȑ�	M#b�/R9�9K��d]�1�C���S�L�*B�@���|ߔ���?�WN�Ir-��bF�h���#@���tq@=�'���JOD2V��Bw�B����iu5�NUU�$�t��)�Z5�bè�f}��j1�wq���i;������ն�u���<e�p��~I�Z�UL'�I����l�1��q���?��p��EP���*�ub�ˀ�.�<'[��-��d��6M��Zy/�q%�[RLXr�ij���dQ�N��������l8m#/;g�����'���󟰉�?������tLg��L~Oo47��ƒ9UUQ:J[�w�ՕL1��TǸ��l�&��{��r���X���F/h_M��<�9r��gn��C@���x�����5S�ms"���QQM�����J��Yn�����㖃���G�m*�
�z@p�~ĸS1���}�Q��DdP,�1)���:1��b�ѱa��`<��q�в�+�ᶭ�X��
(2�uYF�ծ|c��
jk�6���^%�%-@\�%�Lu3/	I����h�;C�;���S=iD�EJ�~i��U	;H5~s��ֱ��w�C�9E�P�r%Lײ%9A���B��)�q��q�e�+"b��#��"c�m̳u%��U���x~����8���_skV9�cHs�{������X��~���R$��a�c��0�X#(��<��f��[+��ݭ�<ǵ����(��8�D	c[h/��|�T�}���Wu���j�A�����y�@v}"}/�cO�-/qy�	4�g�W�N͟�/z�
FB��`�uDu��{5-��~���&��+�?��0Ww�#�J!`G��.$o�� k��IQ�'l��}q�{v�v*�s�O���WZ�nU�������1� ��?�<��h#��o5�:��Mm�dl�s�Z;FɞC�t�X|D�P�j҇G�[��*ȟ�ǋ�X��./颚-�;����J.�_`q~�Y�K�x�z/N�,����Q&�x���/c�;u�0�Z�y{�H��m����G�P%BFܽث�$����}�}�B;!Ts�M�.pBEH9�qC���=��հ'�@��t�:��w�Y��Nh�#*A��:�@�hG��ցr/d���F�a����	B>~�h!��?l�'O��1<�r��R��*�GVj�-#�2q��Fr'�N��ra#
N_�9����=�,p_��2%�������N�s��V7)��,.��j�d�� �~���LHI�_�nw\��?�Z]ʇE��&H�o-�\� �Qt:��۳
<��;w6]�c�X]2V{�ԼB�j�f ��p���h�<au�t@�*��*���ݳyGYy����&6Ǉz�BU%;o�յF�x���)BVm�(b�u��hV��
A���<���W��4�k�-*;�M��H���*a�B�d6�x�>�zg�?��H\�I��
� G��-Q|Z�ៗ�@�&&��J�������
֎K"�^�^��^;��A�|p��=�"/���k�΅+�M��?�f	v���7��O���E�O�R&bJ4kF�>�B$�L��5���í�/YX?����[�]e"�����:p�NN�y�~(��[�,{�C{�9;��٬�	E���w+)��C���6J57>��l�V�4��)nt����'$<�7ǘ;n7_�a�^:ԛ���r��%i��H�uan�>��^�u<�h �ð�&��`4�5�1�?<�g׍
��K���2�y�R���
��^��	�ߊԍ*Zjj�m��X�"�^���6cs�(�'�,�O�Z�N�⎊2�+^v����QX�%Jp�hJ�T��w���0�UY��n�#�sy�D��I�#�}>VS��
AV�T'�R�����~$������8��lK�Q0n��}m�J��9Q/śP�d�=�Y�@K���i�"A�]���������f3�Ѵgl�(�l��Z|XUl~<Y*XN,�OE������(�!C�SeQ_*l�H�
��TF- ��Z�:~HQn|ك�ed���s���]�sk.�{�fCx��S�f��\갔��&�k�pg<GTY�wVw��H]
�b��%�ebC���!�<���S��qF~�x���,�݋~[��$��N�eR����n�7��u{�Tם4k�}|�����i�I�=I\���U���Ɂ�`���0��QX=4x ���[0l�g=��v�@_����n�~PF����Hz�#��������Q��ה��5�����q���l��OJ��������?P�j$���p���ϑN��ˠox`�*\l�	@[�A�d�Q�2ƥ'��2�j 4`WnS��Us���� Ce��*|�s=�\!����g)����j���^���r>��^��?vvT�O)��Sk�^%�a/�
��Ʈq/VF�Sj=y{R���Be� [#�&�m^��۲�I5K���籵��v_���?�pWKάA���j���������	���rU��qq��K����֎C��藊��OK�a�����7fg��1m�Bǿ���E�4]%����3?ń{<m�����ܩ��֨���H�7%�#���-�I��ᇄ�Z@��A��>���#��g��c1-	�O�[ ���pR�,E��z4�F �檬�Q�U�x����{�x���&�̘��k����S����4��ƽ�{��Se�Xzv측�� ����xѻAN�8�GJ��*b��B�S����[��������Ǔ�D��'�H�'����ET *�ӯ��4�p���*�OlC4��b�*�'�;��p!�BLl���t���ߜ�5ѶNY��(%���>ˮ�Y����#��)z+տC@��)�j�ʒ]ub�
;+l�L�~��d��&s��Ga!���9�ДHxQ���tܼ�w%�;��~� F���G��m�B�T�<�~+a���ڱL�����x�~��0�b�H+#���RN��y*��B|B�F��*$t�o՗3h�x�ʽ�y�\�{�sq�:	�l���qڞ(���_�OX�TYi]*Բ�Y֠���/��Mc��"�37��m�����H؂�M����22\"��)��^qA8э�0��0x�W=/�JE�!��1��}�Qw�)W�cYK\�,��QR���l�qc1�����ۈ��du44�"=��3#?�Yn�+쑼���ە�����gT��R!a�lp��wIݡC��5�R5��s�@�-5�o���5�&R8�W�~P1�x~�t���jȷ���P���p���;���OpF3T�fv"y�*)�w��2&������"sq��{TtT�9�'�I'�	���ڇ|ڂ�98�6�%hy杫������u�Q��O KJk+�����:��a;��EN��U� w���e�aW��D��ёq��ݧmC�/�U�{�O7c�o_�@�{� �f�S69��.Kb]�M�[;p���.����@p|�	��+e�r��0����V�|�l����NyL&>�;'��-�~����tt�g.z���Bx'�6�a�.�$ �����gS�<�Մ��Qx�G��-a]%�b��L�Z]JO��ؿ��T�Q��5�b|���Y��@
W�� qvf��x_T�!RU�)C�k(���7�"�{����!E������U��s�C��uLn����G-����cF}V���y�J�H$?~�3��ގ�d;A�k�J(�a�D�}�|�B��5�Q5$���1,q3Ȓu�x!0Ԗс?�.�jm�sL�/�7�YHR�r�˔�bi�=��=��&y���|^�"�� oW��R�-J��.`�6����z�G��?���j����Rr~u8�,��V$����O�Ԗ��>s�ɪ���ߌ�"%ʹ��EA-��:X���f�t�U���^O�b<R�+:�����/R�b������5�͑�Y'Z�@�������	���+�p�e�e4�e��=F���g��K��f$��4A��w��`.�#���YN������s�F�\����H�Gp��>a�oF^�Fkr��q����̣���n���j��}m�\��bf}���$t��7L*�לּ��W�G��������ǉU�6�B1x�!p[O�3ؐ�i �~�LI�%GfͿQ���������,�ț�g%B?�<���\�'VI���!�fP����	�������V�uDE�ԡ�/��`Z�wGa�yFκP������ێ
@�rzVD�%f��Ek�H���;i�&�����sv'�)9��&�"q�����7)�E����U;� Sk�q�F�&�!���3��0��ܿ#w���̐�J$R_Y����=/ER�9Y}�o�;Y�@���ܐ������Nd�"w0��.g\D}V;�s)�j��}&!<m	�Q��-:�"��2AE��.���!~�O�>��+�~�c���T��9��lM��A�2���3��N鰤�f�u�o�fv�%o��e��%b����s��C�_ؚ̓齀%��!CI3�+��6��������Z/)t�*�
��'�/��Ƚu��G:$�5��9i��倅}���|[b,�D�(���+4䩂6Ot�S`��2�0&���*�DS�5�bY��oz���U�1ӌô���!�>��f�&����j��y�k�3�Ͽe�D�����׆�c�J�Z�U"]��hf��v#x�0�&}/�*�Bۯ=��	����E���r���O�0���*�����v)��f;�_!���wn9��&��1��_X׋��8�W����y�Ώ�2)�;�ĺ��s���F=E�V�#g��G�S!B;c�{�`?@3� ��@9(�O��G.�t�+Z�4Շn��j�Ϩ��ܕ�0u��.{|X���w+�0ZMz�,ׂ����͎�T����f�P=G���UH+~�ֹG!߈g 2�8(%��V����M��A���+�P��/hiW�Wͥ�Ņ��ݾ�x�P:�����,,�W�&̬CQu�;���^�/����8"�Zd���h����X@f��jmi�{1j�d�^y��1��d������*�� �heO���c�F��@/�q��v_�q�V i���|�$WF�����<�\7{yN?�H��F%��p~�S��L5!���@Z��4-����|i6_���2�:�T��V�B�Wa�#"�hԺ���̱�o�2uI�D�E(�ĸר7��_:�%p�u��Hj�-.�N�'K��E���h�����W^����%Al�/�ۇ&a����9[�����cAU���%�P������tWL]�����#���	Tw���8�k?�w����;��1&�@��Xg� �
���I��B�[�ߡ���w�'�}0��	ZIya�2G^��%Re`c'��]eԻ�_N�~nZ4���u���V�3"�����A��}1xn彦\+mL��.HVIx9ZVew�[�|#�
qVs�ˢ��;�l^=Md��}CG���t�<���qҠ�M��<�t�QŽ��UJ�&X^Dk��#�$3+|T(ia�/v?e���m��2���H����`%���T�[]��qe����d`֨\�qq�Z�?���v��E��Z�$�yI����6j$������E"�군�3�q�ăs4[hb��yޜ�	d�yX���է[H�.�^�����͊(=���fS��>��Kcĭ�����쫊c�0D���9T�	��Z�_���L�!n�F-��ʆz �5���9Fz� &�W=�HY@�~NC��NV]��o��6^s�,D*(�TDu�1��Ĩ�����ZB�7��E�9{T��9�Zw	�ɼ� ��\�H��V#�y��Y����p�M�Y�j��t�&|@3΄� �]$�j7��@���6��(圧7K̄�v� ��z��*F��L�vi9�V�A���(.i�"8�����#��unޠ�_������Y�qx��U�D�]e�q7p��`,z�2��eMq]I�(�3c�\�*�l�ҒB�9X�>c��70���?���i��C�^gBuN9S��RѺe<&��@�b��!�Q���<�W��Y��=�X:S�q����vb��6����op�]ʓ��J��{&�N
Ho�q�^z��<|��X9����
� �!m�1Wt��B���4��Ν+�+}�q智a�6�؞AKp�M�� ��4[
�ĵ������Q��j��<�S�h��s$t���#�:+Ae.�-���➁a�s=J�
�h֬�U������R��`9����6�at1�C�=3������?W����ef���/qjһ��经�i��\\��$�ج���%�%z�O�9�1�!��ZQ2��:@A����Ŷ���In1�ie�*�y2}	:c�w ����7�5�T���̦�J�ѝ*	����[7*!\��a職�g^�>ǝ� 	}i��B� 9|�U��a7�0d���jF0�C˔���X�d�$�B"���5.�7�;M�^�: I�,*�Q��B�I���j���K��t��(��}BY d��tćPa�ܑ �˄�W��Zg��cκ�����qNB;�ާ���N�$Y�:�^������L'���4o�̌
 ���*��;)���q.8��aJl � x_��"�G�r;�� �t���.6���*��ݛ~���Waө��*P#�b���z�">�*�J��܏����A|wc���p�}q����R���q����9&�����{����d�cx%[�.�tMY��rv<P[`�pN׳�{��T�+�9!���U{�-I��h�R�G�+��#���Q���r�$T��BL��r�+(��Sav�z�AN��e>���Y&�aͪR�M�G{��ҽd�����<A��^$��.$�|U��cG��d�d���֎�loAx���AOqW���j^��c�/���^X����DO�l��uPz޿\fd��H-�� R@=C����2���f]n\�f�Dɢ`�m�~G �	Ǝ �u�L��q khF@/������$̤�&�3�+0ƴ�	�Y���Ndm����(��w5� M{���l��=�c�wU���1A:0���5�w�v���w��`Xᘠ��� $��f���e��9�		��z��r|��"���ɵ��S��GΦX�o�gQ�k�|H�I����z��R��x`j\��}���4�U����:d�'5?�wC;Xt ���A�PK����/������v�u�}���*�ؽQ�co�E��ܜ�Jx���E�j���K���q:�<�أ��C��a�k��rR7 �z���wȧJ�	�2�B��3u�x2���6��/�7���5�b:b$�vQ�x�.�)2D�4<��iY����#���-jN/Z{A�W�-Ar�aU?���n��Ky�Zoh�y�4Q�T����aZ}�~(�� $��:������o��C�l��տ!�i����-���kT�:�h�31D�tC�|��1����+l��#��"��	�������\1����
|�j���F����Xp..8�ԗ"�˿�+��joW��i���[̕xw�#0�Q*g�ΰ���?e<�U�#�<�sQ�Α[��7�r.2�1��ќ�(��� X]K��)�!�!��gJ��?�=����f�-��A�Dk�Ƅ=�R�?��G��;)bﰹ-}=������t��;���ZP[av���2@�7S���S��3|�me�e�f˛��!ت�t�d���7cgM���
�z��
\���#XL�?"KW	B��5I�N�c��I���Z�i�l���ҡgfr�w�H쮑���y[8xg��;>b.X��l�>{7�35OsW?�o{�8�_�Z���`�Rq��N
2v���-_�墙��&��[������Z��Ҽ����ٱհX�{���m��5r�yxaЭ���no��̜�,U"ckl��
]~�º$l4~��kA����y뽧��jŠ�]���6fmK��GΓ���dGz뢓bￆo"�����z��S��mmf� ^�"�_E��w�c(c\�L�����S�_ӓ���q�t�� �}u5T�f��z7X�yW�Bn�!W͂�1w�Eb�|w\�Liy�wtuS6�� /8���>�f�^�Z��H'�{��c�����_��������Q�L��bhAq�����-�D)Q�l�w �T/�]`O�;����' y{i�P��~�_�QŞXs�$`��۝s{�p��l��A�F.��Ek���
|Hq�b��K�J��Sɮeh+�j>c��1
���R��f8 �y���G���p��)ԣ�7Ҵ�:���M&��:�i1�%ؼ͆p�:��p�KN�r���\��PڳyW���bά*�R��%��B(��b8�� rݦW�kR[�����:�mԧ�:�ño����c�[�9:%heBx9�����,��:�M:��׼� Il��x�1i��Ű�F����[�Y)��U��xͺ-%�����,f����j���!������Y}��������I��K wG�������)׽�#J�%;��7e<����R��<|��iK(#!OYKuk	S��qT��@*.�-�j0m�1t�i��oJ�T::����&�����@�٬Ĳ�l �x��<n����
��6a���D@-��R��<�|�����Ti�[2M����C˵&�j��O0�N{[���(��*m���k?�h�x��K�����˟9�~	K��n�Я�q��­��xH�8[�m����h� �i	�A�}W�\�?4�˄�R��Z��-�ҽ]g�E�'��L�/y�m��W�a:!��4F|�a<[�t; '�?�ƶ�#�ʚJd�ɢ�;��ҹ�%��@�/Z:lLU��\��B$�םSV<�����<�I�0��4d�������pP*����d��ζ �SY=�8ժ�o�e��e5�gI��k�� *�=F�tF��(�pLw�I�`��.u��|b;�~��TYEۄ��z����?���0�ͣ�� �|��Ek���@�'w0���ib7�}�����B�#8K��܎��(����Uc��⯤�R��r�%MD9w���K�3b��d�H���]��XI�O�eȎX^3ſ?�ډ&�7@jHKQH2��q�u��J�>��=1Ii����;�]����^�e@"jJ��,���*Y�qXH#W��XYS�k���LG3���st9v(i`5��1�%w#���OX�ږ����oF�J	����F��*oo�U�H~������a��vj/ĵy�J9�F�t6%�����>����yj�y!���j������^ӄ�HyQ�;���>��!U����66	��L��퀒�r��LO����`R{(�2��|IB��Y�O��p��/�)L$h+��]LSD:�ݐ�PH�=EI!6�(W������\�|֍c���l�Q�:nϔ D�s�ER�i���u���yUJN�Pt���T�q��կV�+��Yĕ�'A���m�L�dR�a�]���n&
�-�ƈ&P���u���4�"�j���Yb�~�Bи���E�U47��:9�X������)��d���6n���~�Y=��(D�q�u��Iҩ ���^*~��6gj�]�8���(+�ŵna����v���\�H���&�d2�k>< Oh8����<��]���)z�)��E������c�����7�Z�yҲ2
�C���نޫ�C��y�؏8��@�9أ����S�LE��&��vә{�Hu{�.���=1��Xc��6.�3f���d����'#��w��}�{G�x��{�WÐ-WK#�1D���x�r��(I��O�M�<�������B�mo�1<dJ�iW�d���c�)~V�
������"�8s_���ҧm/�&3Y2K�r$Ţ|��%c%o����Oގ�
p���g	:3 ���2��,̴�]�=�:!�u�c��*��!d�_������
�����I���_g��M�l$�����^����p��>r�QU�_i=Ȩ{�0>ͺ�M��mA�JI��n� A�@F[)ӕ�EÔ	�zi˘1Z
u����;(&�S��K�J����t|���ƹ���h+2�aO��q|������ʪP���xJ����{Y�7�_N�5+W>T�#odg�v�Vg��C�U��瀽��j�]�4g�)y�]�e�ʺ��C��}oV(,@�}�KZ��o�c��㎇A�Ǔ�&���6��Ƣ�/N�+8�����<����چ����pH���i�?Y���Y��
��d�t�st6�a"�"��@)!�������e�A��i_ |!�<�uN��L�g�*�:�%�Q���S����Ā}���~6����,�Kg�=`^��\w��X3!��9p�V��^�C�b�_�rdc�ҽ�<�&�	�U�����0?�[M归ϧ��g8���dl�O$����p@a��ک���LOi	��MIF�A_J��X��ӥz�B�Fݢ��W��ZO2��I��V+9i�����FC9�ZX�w���Ϟ���ʬ����=�&��Q�u�����AGr��]�	ݚ��l�/C�{"-��^āew�8˲�-���2X�m�Lݙg �ޔ�yq��&���&P�Xoe�.��A4�m`�g�O�!��1�od$J�mE�D�G�8y�l�� ʢ��\&��� ��Z�ڎ)̉��2z��o�f6��)�q���:Ρ�_L.���>0xX�H����4;v�Gi~�4�L���l���:�u�f̗('"y.�;e�A��X�>�ug\D����Y RG�_a����յi���t��Bap�(�gSP���D�λr^U����M{�7�Y���ߩ�	�V	�(=!�aa�;)��w�t����b<��nN�/������{�a�i��3<�Ix�n��"A���#� �ڕ��<�*O�NB�#�T��*U�"�Ě�T�û�E9{�7̅0�!�o��\'I�6a�:���TX���hn��ɯ$���z:���L���ﯴ��A��՝��(f;2�}WA'�&�����pj�B!��kO�l* OF����y�5�ǧ�1É�CX�Z�[l��K�)�-� �<H�f��{g/��kg�,�dT��Qp�N��%�F�r�B`m��
N��`��s4Kn�}]7U�M�� ar�+��i�6c��alPg���o(K�ᓲ��3�YbY�/fL��(<�ġ#�����Q�F�8��
Z�bd���KC��_��������韅f�l�W�۹,��"�)Ɨ��������j^]����ʘ�^��0��aP^��o����$v�B��V��y!���<; ^��3�/3썛z��0%�Y��Ү6�D���1�Y��W
�HX��H`��7��I���_S�b3�2�?^���Gឨ���x�Ɵ�&Y��3��3(����e]}��-���t��;�HSd�Q����'8�$�C:��Xb1�$�
�4�*�	V�b���j�\�Hl
�E���'�HD���ߴ	@C0%�-���~�o���RD���b�]B,ܧư'+��N��v���+�5^NQ{��L8cv..8w�!��Zt~Ɠ^]��I�y�#S�.����`����ͮu�wq=�W�_�w����ޱ�xfVu2����:Wɰv�0����Ū錭��^Q0���8���w`�ݢ7Op.xLt���O,���x~�h�50����}�ʁ�ڕ	9=ft�U�F$!�@{�����ۑ��Jھ����YWe��e�!�O�*���I��`�H�g����9-��V��7����C;:�@A	`��;"ݾ���s/�?�.��i�ng� r�ުT�j"�!?���RS�=����s�[e	z$�\�'`����}��B��E��f���d��i�0�������%`���C.s�r�y{�уN�>k������^d��{�f�,�A��@�Vo��Ϲ��Q��U���s^��M� Č�p��ʧ��ȑ:��U���Q�мn �b�1�L��&ů~>��=o��(�7s9�okg�z��]T)v��E�P�d̕���`�c��q�W��AC�/O�d���u�^x�z?	g����k���"q��ܖ"��N �83�Z�έ��8�F��7��YY����?���f��YNcfn�6�Ž$�4���P7�[(����.0J&��j!��Q#�zs$����ڑY(���lh��\ى�F�%\�r�F�����G|G�ݨ�F)�����t�`3��5>e�P&{⥈Z�j��D[]n_ ,X#73,IA����aDA��!�Z�l-Aмg\��y�e]��,���X|�LG+�����{J�3a����4s�d���5���
�Sv�,�nCG^ŀA�G�D��(��dĿD���ve�g�P�[ ��Q 3�3��_���:l	3S�R�Wp���R�,��7�S��Ix,��Ή�b|bUޟ�5IiT]	<�t�Is�M*�'�F�z��Ϲh(��3����I�l��m�i�)i`+b���-�ۗ���i�����U���L�7[��
��>��L���X�j����w���	q�K�)�N�0g��9X�<�m^���l��I{$��|�q������x�x� �x9����ke�7��zz��,�['h+YM���d!k�H�\WPZ,�K�|�w��b��[tVR �N��D�S7�uarIEItMӧ�g*R��'	��`@������,#�3�����zs�p�Ѿ$S��ns=�(���O�G���*�g�_g�!�"f�˦�5h������[�p4��"�h\q�q���[�I!C�{Иc[�'���]��<��JE�?WU�p�s�:5_���!�-'�д)F�E��V�Ao�F����N �B��q�[t�
���2j��0��'r�
`d����ZML�7���	���
u��$�g�
e5/��7����)*"�s�d���{���@y��:��;��b��b��|P}5��h��|˔��n�C]������[�U��$V�P�츐�#h�2�žΟ,�[~uL��"s{����A���;V�\�Oi���_������"5C�+2i�~�s���Kc4<�\C�W��#x�X�:������I|{4�j�g\AԷݱ��F�@~���`�sR~A�x�?i.?�|p�MH5��� ����Jt�`Op��ҽ3�,��EEgE��Ǖ[�=8�����^��3sJ��h� �K�f}��7���@t#�v�����.�'G|�����˸��Cđ�E9p�D��G����!��=����]�UKpL�D�<�'LHm!�C��RCޑ0/C�^*[���s�~��7_�՛S
�_�M�(]R�%u��{��km\���"F/]��W�䗒Q����ӶTj�I���0QiD�Tu1q�ŭ���z��P5FB�;�����Te7�R��w�t��e�R�=m<�^t�b����ZG,��q8��K�B0Ww�B$"�ثZ�&�N7By0��!���	D��dŅtt,e�fUv��)�����Q~���w����F�0�.]Z^*tn+���bJ��(�´A�h��c�:��e�>�f��d���ԷT=�f��}�!4�������["��b1������т��K����p�s6T���dz�2��>im�Ѓyz�l��Q���'����$}�" 8'�W�/��S[�3]�/*^vf�l�n'��cL_L�!>zk	.����f7�{���l�w_<��ɲ������P����	�Ҳr�d���c�c��N��j�<��+�6���*���\L�dN5 ��
5���N����J�>03Ũ�Q�W�"�k��ICu��$�<`)�$�WeI9C�̲eb&��O@hU�~t���瀥a��fSkC�{R���g�&0W6�Z��ʴ�$��g՞5�!�o�%ݎ9���#�2wF
B<q�G��6���Y�I#�(�![�V�Y�ճ��Pb�i��P���9�%�����
�ȋ�
	앴E�heΉ��purVgʏEso��I>�Ԍ��f�~��}ި
�d���{(I�8���T���]��i���
ɲjk�~φ#�C�l�P�OQ_l��N [MBJ������,�5��Bn���m�uZm��b>�n�V�Jo��N)�n��o���b!)���	w 3X��-�2��kG�>���)�"(�}��s�)$?X��zB��1!����|im�q6'���C��)�C߽�X�tI�ZP^��`�Tҋ#�P�,2!�J�8�d�3Y�nQ+v,,��Vz;%�?ޔ����(:?`�cL'7��Ƴ�h�c-Xn\q7W���8�������м�1߀m�w���e�-��	t�+J��i����_{'Y��C>�Oy|UÛ~��X��!��B�U�����8�d�i�׆!�	��~�p_r4�XT��jq7C�Q������T�����c.��M�!q/<z?�D�1�yic����#�ֳ��MIUޘ?�U;�:P�)���G�Z+�7i�e[��ꤻ	�߶8â!� {�٦�EmٰXW�+�c�Ş�ӕ�?�)�2�L�(.Z��\#h�J��8#e��7Aߚ|�j� �Ʃ���1%�� (�L�l��'�1^�2KNl��b�����~&�z!��
z3eV����nXN|a����o��Yql��gKW�?��4�o�/��t���Oa�2(�:�sK�έra�hn%��}�kW��b0U�3EΉA���iո(��dv
$_��v��:w���EV��z�UNo ]�)��^��`��w���hH��`�Բ�D�V��[ߪQ�gb<l5�q���(Ux:���)�u�
�
�%8����CiJ����O��+��o*��|E��2�t*�SG��99Z�9��@C��J:�����Wwꮲ-�Av}l=jR��uz���!3������_:ߊ���O�H�̪�8�8grc������i�T?��xV�x���,	���s��XP���W`�Iy�i�]��ia]�R�e�C/��'�:���$D�}ܴ�Z̹"$Kp�ZΧ�\�˧<3�߉Z���wʾ<F_>���4��F�`�,�Դ AHE�JY`Q��ZI��<�- .�E*��)��J:�z���D�)ـ:�CNR�.�-1;��<D]C�t=�����  ��.��7��ňC'�����IA!l�,Gj&�jw(ʎ(+��Hs�?c!��+�J�������)�z���!�t�	�$�C�xv���KlL8��p�ɭ��)�4�����g��x�I'��wz�K�粷O��%K�����;��=�S�zFD	g�Ht��|�D�'_[q�MA��R��> B���Elx\�@>n�y�'��SC���>H�/v} 5|y`��/<��d���R	���].�P<3�N�-(L�QjY�y��ȡp�9�{���B���]��N�i����&n#���FZ�|3Y3a2�Ak��a�?�TPއ�nWT4�P��(Tp@