��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����՗߽��F&����B�?��'����n'�۶�a�P����� ?�*]�)A�llCϮ���F��r��t &B�X��I��� <Z���uI��g��zr	�I�<��cX_�������u w���?�(і5V{�+V���(ą�n���J�7C ][c��>@G)����$���o&.�L�W޻�^�	�Š��Y���P��r�F��+*���ّ.�^M��~|׏e<3q4�M��lFb<V%"gn���H*�[CP�C"���Sn���w�E�1�N}Xu/�j��}�?��L@e^E�n�LE)�N�t�aq �R  �ag�"3K����ep{08x.%mJ�z2��o��3�0OwGS+�8j�?+������z	�s���?ܠ'�z��ğ���K��ڎ��dp[�S�76P�85�B�-ҵ%~���Wj���4w��,J����/Y��Bk<*u�:�`&����y�?Тn���D��L�2��ԻvC��KR��� �aF�Y*CP��$�����Q�%�G���H�I�վz�↝vO��(�D����s�	�*	�>�.����h\��e��!Ϊj�rF����X�CF}�L��5w�f!�
�)��k;��U���m�3��(FֲZ���Zʾ���הwP��g�;���aL����2`#�ت����������DL�1.L n!%�g��2H9��eZp{ј�_�($mͷ��h�����p����K�?#�fn,c;��B։�*RP��:��&��|�;������v�*Մj*�����	�%�(#j��U<�V[*4?`e(�YGY��p%��/;���*Vp� ܤ���o&���g��km<��	X<:�KY�7�Z��t�H�}�B�����,p�a7p��X ulw���S���ϼw͂d���P����#j��-�Ppw�K����0w+���/0���r�}�?�Ĥ�q���wjύ���t%m*p����~�(d���+v'+a+s�Hˬ�b�����M_�f����K�F�hlv-���#��Q=�@�'�L��l�#�iv녁e	>����w���9w�n-}�b�D��k�3p��>��>��ItHX���L6��� ��M��.L��\8ǿ�.�*%\^~��x�PZң���Z�s�IY�G��Y��2N$Y %{�	ڙ��9O��Y,��YC��2����@�_�ƍ��ݹ�#�K|��x�Q���]I��� g���ܠ��o�d�����&����9dn�-�#�G�Z(Qn�G���Po��4������G��7܃�y�Q	�x=�� ���g�:r��R�J�» �v� B1�Ff�Dd�`I~X1e�e�қ�6ÖQ����Y��q�u#᪶�V���x�Դ޸�*ʇ(/qɶV�ʭ@R;��0��挮��� ,���B[9�l�6���,��en���s��z�z�K�����D�;Ip)��[�[R����҃o7�h�q���.�DFZ�Pj���_�&
����}Zf�H/�f����Ry�PeR�M�\����.����0�jJ��-d�e��.��Y�:�W�W_܉ 1��򨭛C2�w#m��pM�E��V�y��@���'�9a��bt����y�2�-IrE��`L8��-#K 3������$Ӡӳ���䕏����4�ު�.=*��U�.���Gi?rq�L�lȇi�X��>�6P�S��&�l�s����&�ʊ5�b�)��8�Ҽ.�X�X~(����d_My���8���D����>�G
y ���v����ZC��R3q�c@���ڨv�9���PNj�����R�(��G����p��[�}��W\�E+���X���ߪ�(���X��ڶ����"�3��"X,���ě���q�\�c����h�}�A)�U{�PWRސ�\F��3~Y%$�#c���A�-�/$�P섌!�ߏ��Ɔ����D7ޅ�Zm�9�RT��p̟m"�1��+���a��տ�L�'|�h��Y������YL��:�����J��!�io�������0�o� �#�Ut�AY3�Ǻ�X���%�ks��:k3\���}�;Q��g�|J�Mq{����m�)L��;4��� ����|JV ~t�z��M��7�f��,"6{�0?T���֔�q��Tb�f7@�->���Ȇ=Mx0�������T�}�J���ED�^�T���NG-�.$O懨&�G�0�vdS��29�m��0[�d3ȿu�9ϛ%�R�u��$��W��J����N�^1'3f`�>%�w���p�ͤ��-L�v5���qoPYe@�֑��LI`\���bnI	%��NR��%csY�1��[^[Q՞�#D/,QN��(\.����}&/_h0�+7����|�Evj�'ZC0C�_6�N�DъF����ɥQ���;O�G��)�Ԅ�� ��.$&��s�ꚦR�&�����7W��Ĉ���U���\�'�bF�e�PЇ�U��㉨�7q��(�ZP|֍��]���yz7?yZ+J�j�|P�[�$��z�'.A4.?��<��q6l���fP�齶��,5M�2ޏ�:6���H��A���r�/��/U�Q$������~��un��P��%|_�N֗8�M����
,L��cr�]�a6-oY&�3��c�B��5qu	�ɒ[i��X�;b��^@e�i�:�x[n{�i%8N�.�棷x�1��%�IR���j��iW�����<�D��j�M��t7��ϑ)j�{g*Kձ�b�#�3Ƈ��W�4�4�4s��lG�̜É�"��3qI2/j'O�`J^~Ye�0��_u�ۯm���}��5�#&�e[V�R��-h�z)M鋬��\<���Y��9�-$y�V,o�*8̠157��{+`���B�ew�5E�T\�։^L�b��0��5��
/��-՚�i�3|�s}��{�o��+�E%F�rt6O��5���[˳�ә�J�I��Y@��k��?�I����ef0�w�G�J�?�� ��ʒ��u0��x�6���Mcщc��0�@�\��b���n[��V	���:xa5�8(�`���fz/p��������RgCەq�	�i���.R<8m��:�߲2�<9]���[��.�!��o��r	��,D5���[�pΣ��ƪ=`�i��		浱W]�1�CРP��|w?��(�A�]a=fЂP�;�7ኳ���Be`��9��J���a�(,iH�=�C�L�.��&�`d&������w���Z%24h��8vh�4g��;C����i���տ3�E���8E�'�c��l�>o#��"=�-�����_[��K��Ɣ*�>%�õ��J�z�2P��W��c�[5�&��a>��F��M�����e{�]��c�%ހ0Ƅ�c!�0cʋ9Qb,�]οM	3!�I�=��@�c��6���p�_o�eh�KZ����=�ص�~M0�8�g�&*KW�٢����J(�m�Td�Vmt�nyoXPZ.׆�PMG����*/j�t���d {ZԌQ���hQr��J����L��~iO��VxC�	l�Ӱ0�(r�_������'��/+�^�4��+Fyo �cґ��N����H+�<:؎�r���2���=�E���O%fۿ�Ӻ��I_����F:O���?P�K @�hK&7ԟ�l�=XS�=���w�V$�9S��0F'
H�R����A@�0֗��1i�y�^����ݱ�:�>�BI��ԃ��Y\%T�.M,)XJ�����>9v
��򞡳K������l��l�/�S�&�S$�<���!�4;�s=w[�����0�B���Y2}��o�Ɗ*�����O
����
D\����mY�<��if8��çpn��u1���؋�ݲ�in�iw��<qA��@�����A�v�Pc�ң���ፇ���w�t�M�o��P9,�8,�Q�R,BUk���j�-���m�[�qϒ�~�炄X�x�}���1s�l�I����^��i�Ar�3�V%�q�W�S_0?�kQ墅�����d}�k����ڋ~��������2>�6�r�ÿ?����;��%͊3((@`B"V���%�ʒÿ��G�n�6n���C-|�+�GJ_��A�� �3�������+͈�Aki���-�2���fа��������-���IK ���@�����{W���*y9��{�$r����N�t_ ��G����>�؝AF'�T��ޡI���&��s�='�< 6Q�W���ܢ�_�6��T�z�[����%� �N��K���~4��)��-�6O㟔��Ʌ��V�3&�g4��	�W�J��u�� ��i�.���js��1��^�FLY��Q�N��$C�G�aכ[,|+�Y�8d����fVR����q���gM+��t�>�:������x�ꅙ~�i4�>���%k�(IQEv1�"�Ti�2 Ey��{�ɔ����������R֫��mWГ֨�
A��F�
��Yc��*3��v��]����e�<��0*to�ַ������ ���%�ta0�����'�*�5��d�,�l���	��hQ���S�`�n��+����`�� S{!� #
��oAcV��L5Uz��a��ݣ(�Z����y�*rSh�5��y[�6C��L�93����n��� �!u�52��n(�O�\�삻�q���o������>�C�'&�*Ϻ���OR�H�S�vɴ��!<w'e�=��8��O�%c� Jf[��t���3P�����:��(j��%��6�3a*�#L3u�DxpĸY�L.�^�%�}٢ 1^���d�S��~�����:��'�� ��򛨝yI2�ڱ�a˚5:�K�D�������Wg�&95�k9k�dW�u�b�.�a���v&����Q\�H@�{y�Hsg�|�	�F���(�:��s"�!��≞��H�1�g��!Nn>43�r̞����P��&v4����Co�Ԭ�֍�_f��J��Q���T7U�מj�Ǔ��/Ln����P .�h�(�7Í_l���ӘS���/�E	��W�%ezڋ�Y_�H��-]�H��mj}DLf�whyH�oꨳe`������Z����|.xX~<��nu?f\
t�b���dh����������q'�Y�/��E[V['_����X ���i�+egB�U�%�U�?)����o>
��������\w��]c�{�1FZ�Q�s�2�sW�E'(
H�}�|u�ePB���_���*��(�S�s�$�g3���'79�_���&�b�zǵ^{bğl0�&�<��<ߢ��T�.t����Xh���P�2�i;{_����z�0�̔��ݍ�f�L�2(��g<��V�yPͯ\�d<n,����6��l�u4}U��6�i��^&�B��c:�9I���h�b����X�B���5R�$S�M�冀�7a�㛧��	���Oq����J$�>-�Yk�Y�Ef��M��E�x����ސ2f|�����[~s�,L$�2_�x�(�X9��d��y��������.�V�;���Op��)V�?#���P������l�Z~�"gr�@!�u������¥��P��R�t��q�[�����Њ
t�>��K�K��mO>9z�p��ͺ���@�6��B�!�M���8�=ۺ�k��%f�a{��z��1�����T�wS����;���S Wm3�m��fm꾵��%����h�&S��<�Smi��⟈+�4f�n8��,��`TrH�e]��ok��q�8ct��[g	��!phɌ�������'�q! \3B:�_,&>�(���^��R��\�I`�z�s�>O��w�Y�5Ѵ��!f���U>�Ƙt�N�)B��G)��M�Ac:�g-��P�(�	u K�D׺E>���	���e�v�E�_��=�ی.\p	AI��x�{��T
B5��
�`���^�~�B�B�<�T�����|�hQ�M�t��ڥ�l�H�z0��:z6��7���o�ڲi��6���\/���E�[]5G`z���L�h���l��:�>P����Q	��3ҧ�:>N������̣�Cz�z��u`��*����]�^��kd��;t2Y�9]Ŋz�h�(���~��"#�,�c�uJ�[�����{9=l�0GO�\�A��& ~%�U]�����:�&�P87�++�W[Ls��1)���.��؈,��l���Q����}(*i��z���W�7n�� ��L�.+4!��!nZuT^�m�yP��<M���}���s��(��b˖o����� P3+��<%
���pmAS�������0����A������^ �Fk����yMbV����z
@�%ê-i�?7.H�3���V���fa?x���$_66�fj]wı�+��|�PA��B+U� -�}#!h+o(���ʯȫ�4���^Cqm.�$��,!Yv7� k4lZ1#{Ap�@��������)�Fa���)
D�����B(Z�B��x��r/VE �̫�)�>i�?̄P�wP�o�^oL��ܓ@�}&;*�����IQ�m��"��zn�8�vbQ�Ha���G�^�׺g�lѪhe)��A1 �"hl�*���z�"9p{DX���$�����"����yj��'�Q��;�\��2�3��祂�F���RI;�ׇ��YP*	�͏W��|Q�3��u$��L��ٞk<T�;�,3��H�;Lͣ�M�z�j�a�6ܳ(|�ls����A��������;BgG��q�D�gJ�{_>�5��y���.�����z��^Q#�j���oĝpǓ����x{4s�0�e��u|�GJ�|��U[�!�9��:�ᔴ����[X"��Y4*޼L8�[�4�[�u�"b%Bؐi�H�~K�@+�:ffHzk�y����Wv��`�X~�뉝E�����9�|���k~�n?�i[0�J����"���i���G�M����ٰ�R�h!���m�Df/C�OP~F";Ԑ�S�DU���'>b�]E��5ϐ,�0չu;���[X~&\$2��L�o�-e)�L�hSm���@��]3�~R���;�I�����j#	�c יr�7��K\�����׹�">�d��Vx�N��_�&�+�m,��.B<@�J�e�mW[���R����ŰM3�<I�+ g���Q8u,�8��Q�9�����t���~�:�g�BI\���ۆb*l�����q�R=�Iߵ_J�+H�J>i��ʒ8�(��[�b:���Q�C"K��&s����E��K[��������>�8ڽ�?[?s�F:6jt�v���Ysϑ�"l?��mB�o�r�!-7�F_�[��5�������]\���L-{�N[r�R���1-�P�wP��C&���K<`���g3W�g��>�Q�å2m�e���1n4��r��
U�)t��BZ6�"�R.�0�&��828�4�惆��^(p��i©S��������~��j��c�]'V��
R"k�Gv��#T����kդ!Gn���r�KGG]A_%I�E�C�x�L�G�����������Tï����qe)o�#؃E>�Z(������D��rb��%�2d��X�����-��D�dk}�oe�o.^{ݦ˳@oB1Zv��z����|�:��-H+m��^nv�*w% 2�=]A��QE=�Y&#��D�[���煔��uI�Z��圧�|�����"���=���43X<�B�H\=��A�b�O�nǛo�-iv���U�袺��O!J%�W�{L���Jܝ6�5>�
"'� �E��\@���ZS�.Ͽcؚddr	��G^_�7�CdCm�T����#�*D��;�M���#n�͎�Ӽ|�V�����'��d�eh��fM-�Q`R�re���}�5F`�N__s���V��!��ytb����'�L��Σ˾�l�v��*"����#��6��ʴ^�d2��, �xw���
5���Q��*`� X��jI�;@;�گd�h�ﱬJ������P7Bδ�,�����]����,��s1q��F��d�>���4��L��<2e4�q��Y��#Aі��\���G��XY}�݌K���v\��.j���()z�)u��CpO@OI�_L!��9c\I���V�@��;��;I�^4������Ǆ���ЯJ��5M�΅;�}�����w�+j�J�;���h��t�]���A�j�p�w����IY$}�|� �7�G��f��E�O�&s�=r5�O��;�kj'$���g�n͚��ݐ�s�v�P����e8���L>�߈��I�����+m�U�R3�J�[5:FHZ���a��Նe52��J��+�H�� 泶kn�bwx�.����a�Y����X<�գ���g� �p�Ib6���������N	L��ɂ4��QY�
l�;7&�'h�1"���R�TFq7(����.��T�d}���9�K���o�v.�h�M���sIp���R��M����FT�*�@;م!�&�4O"Ɨ�����%�[���"�pd��6�H��*	���6�H��-1L���O�������@�J�JѺ���H,��~��9�zk��k�!���H�.gʑ?������C��D��mw�I�����<����M2HZ�sF�Y3뜸��1��}�Z�H�o���M��M���4X�6����{��?���B�E��qkX�o-~��wR�O!��ԓb���d��g��V!(�-��Mҍ��d�O��}s�/ː(�Aץg����mLV�Z��ꁗ$֛k��ĻgM�O ʏ���4�MM4�N}+�-����#��|!�M.���,?��%Ҭ�K�}?80��o��r���AA�˙�z������j�g	c�_N{G���<���R�φp��Z����|\��Q%�_����p.�o��[+lDe s�F���,K�|��$�'����D��!� K~GӦo��[J�p��D�Z6�BJO��v�ܝX�
�v��J�iE�j��X�M�8y�$f�^����XaVņd������\3�XI��W A�!P�����>��NL���Wp�S��(�z�j��f��U�S{*���af�R.���?^������#;�>ƙw������[�C�+�Y�>��ǳ��{h����O�9*1��Zl<�C#�K���q�ϢDw)J���p"���|h��m��~�db����L��j���B%'���}��sۦ����ҟw�h�S[ieOq,�Rֶ���_�&&���9F�na"��3�(�Ft�+Ep7�[��i����Ԇ�̭�%Cs�Hx���I�Bqo�?�NK�:��!�G�!�<^��jZ��lW�̸YV`�,�� _%�孏���H�V|2�E r���^"m�#J_ W3,l�i�����T޼p�fwN��J-��g�K��P�ic�� k��L����ԑ1Bh/�k�oO�x�M©�v^���$>:�W_.�ג���N)Iu����΂���wsգ��2؛�n:h�"G�hX4ɂ���a�lZ�OsI�G�m����v9{߶�>����dP��5�� '�����J�t��](�A�M�ʇ#��"��{�ԓ3?@\�On��&?;K��8�b��q��~��0,i��N =�M*��d�~��'6��e� 	��$Y���^�����%��{���f��䠅m.�%r�P1�b�~t;��|K��:񎀽�0:'o.�k�jd���1�[������D$qs.%*q�y7������x��e�a��mV�l���'"R��<���Ͷ]��t���1�~�52����#�rk�C�{؁�C��B�X*�ax7�@V2$<lFj&F���E�|���w�E���TLlkH��̘Z�%���[�fu=���X�k'~��G����=ƟC���:�IQG3	3e_:������-���;��Q�BXZ~ʭ���pkM�ZDw��ka���1��Ǣv�������p<�D������ϲ|�d	�AN����b� Eo��i�s|�C�u��h������>������g��C⅓�m�45�����N\���HLS�&�I�Hޮo�-[������C�M�ȹ�-�/��x�_�0��#�����@�x���C�4=�)��
0䏜��p�!����V��j��c���u�I�:��&�p��;2���'z:'�G�n���E�^�7�$����]`���n�Q�Xu��}ݭ�t�O�o���af/�VE7H!l�&&����F����b?�)�������i��`�=HN9�?��G��-��U]d��1��p˓;{���MJK!��� �ќA�.^L����}5B��.n��{��c���@6"�-�+�AK���r&\���ڃoS�`Q�Ncw<�3�<1e^�]���y�Ki�$�G��s���cJ*ג���c�-m?��*
�5��Q?���Ri��!(�S��"��x����z���DL��-4��G�P?�[EY�)@���������,�Ap4���v 0g�4�I��N×w�Ѱ�Ng�ʎq�!j�G�^�:z��T�������������Ri�p����~&�/�nM�iG	�3���<8+y�$k@���9�u�����?���g1�[4ՙ5�>�!j�Kg<�J�R�r�'����g�Q�����@�
I��*���P����Ua�`��0�����8�hV��I�R��;/�%��}�yY<aa�>S��p^P��gP� ��<�p�w)k���|�� �g@,G}�l��(J�"�x%��۞�*�(,=<��[TN��P���z�6sg�dξ��;<�Xm� Fr�����,�j�Zdխ��wc/��M7���*�Nz��^��[�m�<+y��q-ڐn�`�v�$�{l]/�t�Pf����ڮ��`r�}�Gu69���e�͝(�6ጺ�pLg n>��m�F��־�Υr`>hvO�n�С�t�i'1�����Zz��)ӯ�X�.�Q�Q{�ї��Շ[�}�6��k�7���rÑB1�)��S��j84׀�Ȗ�$^1�)v��	�e\~�^��c��x��m�{tJӾ�����K5��3��}
X��a��Mvu`�˷߄�­�t��%_'��Z8QhL�{\�z�XtE���0�a��Ԑ�}��na@8�/=gt~���/h�-b�0�a8U�9j	w���5�k�������į����c���w�X��:&B�3"����3)�%x��.���y6�z��5�M�n�ϼ�o/�$S0��cH,[�\��:�7�؜]��I�+%?ra�<�u�8�OY1N<3El�(~ͤD��������1 Rd�=e���d�Pq�RD�x��m�HJꤷ�¹=Z�9;�3<�����}CK�-��DX_�A`�Z��Q	��ٿh�M� �g��j�c@dej��L��l	`���҉�}�M�3#�Mg�L��˼��r�O�����lDz�,d�H`E�;�k�"tпLIG�s�N�Ƕ#��\�T�X��XA _��9]!N���s���=�wL�,_���i��;?�K{��f���Q��?k����.!��#p� q�0Ъ��@OJtq�4�� ��p�6�Bm�h�b�F54��o��(�����}�FB�R�U�`���T��摒ߝ��X�d��d�����S$��,���=�`�������P1&k�#��,�M[eV?>	��]�C���_��U��ꄎ��c����3�н���D�K�� ƽ�k�/H7���aTt���B>.(H����ܷ��W����� lƗ�]dP+�AML��\'��g�x�d����R1��7&Mg�Lˮ�X� N��EU�M�W�� Wbg� bY�����"��Yݧe5�T��)#p������X�|]�J+AU`h��A/���=�X��z��=���|�d�K��K"�g��v�
�v�wQ��n�w-�E�G!ۖ�TQ���?�0����]>L���'W�#(Ф�b ExH���\�m�y-�����~����Ʃ�I=�m	�X�WZ.U<�}�`�9W�+���l�3��ю홒NXKQa"�On�o�Ŭ�Q���8ԝ]Q��Xl>vC�>I)D�Q
��{a��˃&�'Mx|_˻�xdv�=�&/� s�։����� m0w��|2~�X;�Vڌ<�a[o�`���:�lö�Sj��]��ϩ�r!֍q�k�.a*N���5�Q���g�=㸾�:;�������N���*(5F�U8S����{�_d~�
�7M���",b6���f��+���Eȣ�]ե���
��7Td�����?�/��yiɾgۑkB��u)	��+��q��3A��b.�X�����
�C��K�����aXq����"�Jߥ�/|,R�[q�C·Ya����Mf減�q��1��#dQ����y�a�1�Ƈ��$��+�?�f�P�조���J ���z/�d{�u�d)�<��{Ͱl�[�KՑ^�ݫ�Z#������n��9�5��?���
��
�]��#*e���%J�<K�p=Y���s_������)�Aѳ��(#O[�F�����2�G��4��_(>
pm��YRV�Nq�9��ު�"� �[!o?��)�˽�o	��6Ini�aZO�J�RUXzUaU~ߛ���{ #��-Ʀj�A�~�\	��}L��Y)-������3�M�Na�=�eǄ"�੏5���O3��g��� �Ń���N/�pZ���\w�P+ݿ�,R7f(4���w�;aE��Ĝ"���a)�Ń3����!�
S�J�DQ�h�^#���Zۓ��1@��K����_����^���r��+Ӌs���m����H����-?Iֺ��O&�{�AOC��1�@@ҳ�PLu�3S�^=�g-id0���X�_ kZ���j�A52�?��
�����|��]¼�Y!R��
]�;��<�w9��DbZ��/f�� �S=,��t�XJ��{M�dJ�̨Ҋ�-w]ĪO�:b�Q�d+��L+E��C�ҕ~���2��Ӓ	��Z�Z�p�$���S���[���Nq�fpns�+KT�O�u��$.�><�_�M�
��Q�m��KA�1X�%�h}6���v��](��%*S#2���˾�l0u���ص�����R����N�[�󫆰�pL�[�'W��>¾�mL�:5tN�@<���vC���U�"���3�ʖ��PPs�޴���I����aX�*��]�pn��g
��GU�h�D@�"�;�=���ty	�{6���*�Q�Ei�/A�5Z&�0�A]�LP�Uʷ`�`�˭��I��?��ԋ-Ұ~!`��&)z��~�2��n�8<�l���p���(���4ϗ�څOr,8�	w�� U������h�ǽZ���<WH�K�Hޓ\9?�`���+^�c��늨-���'4�!���{X��O(
z�(�}��O]��I�A�q�@>��7�#bظ����\H8�X�C)rԂ�?C<�\k}�Ҧ�d��5Fx��h���;�Fm�H��/Uo�%qJN�M�i �-�u�F�\���H���&5!>��RᲝé4�6���M�ւ��0�u�ћmb�GmE�Y�]�<{�A�b�E�
D��Y[�n�&v����.�l��#��ɿ=c��*z$|X?�
���O�)�_,P$*³���ҍcm�;0>¤�-�l-{#�;��k鷖޷��!�0�B��bj��-}���!�Ǡ��ߙ:{bN|��k�i�=����N�2T��V�f��Yr`�̺/��Ș9"���|v�Ȕ§w���n�x��o:r���;�V �Ώ˹3���FU{
ρ�]�Z�뎐�iۅ��ba�__��L�ND����Ga��,׮��-9aȱ�c�S	{�%�D��[��cF�C�%�Y�|���v��^�G&I��l�I���1�R�i	'�W��.�t��	=/ێx�H��5 |��lq
VȌ/}(���W$1�5��@؏���I�q5��D�ӟ�k�ß��g�]h��V�Q~�|�3{�fD��)L̷��ڧM������0lmn�O�8����(d���²�(�}��e��3� ��� y�K���^+y=�� 67b�-�dO���]�"�g�V�.����c��A�C�Zݷ_#Oe�p����	g��[�Id�����j�h���y���K��Qy���� ����ҙ}���O]+qvYA�~�\�%Ea������eR'��oƳ�SxM�.jhLa
"�-H6g�ey��JAB
�k8k����v3
�����W��MyT���pUiG�\�����HWz��U'KY�P"�7KJݤV?S}L7��(@]� g���A�Kd\�`�4O(�ݙG� �
y�_��`����ḡPՙ����f�|�z/U���6�e���el�e'мt�/Z�/c:+ؘ���_/ռ����t�a���&R��[��=�z�xf��IH�&�4�'7�>�rP�#�pOyp�P!�J������������Sď'P�͙�'��o��=3��Z!��1��r[o�t�_���I,c!�TDK:+�:վ�Y�}Ǐ��M�h6�(Mx%��W~�ak7N�ja�<?�$X��Jh9%
x���V?�:òh�U3��t�c�`�`��H�������Ԕ�}/�rÈe:u���G������$��d��Z[,W&� ̔Q��.�JKdc8���j^�U�K��U�-/�N�#=���~����<%���a�U�i@ CB]|��e�a�/w�C�ӕ�py&C��+{t6�NbmX`:z{q��כĨW��5��їE���o��XK@�o�ă�(Y�7��j��"
Sj�e
�avo��O�� %V��t��u�����&�F}WC�5y	�� �je@��uP	gs�Qta��Gb.�m	������t�����D���s�Q�FQ^�!zH	ǝ�,�ڏM0Eh��{*>�C�q]#~i��p������kd��g6�+��?�G�;��#��^�w�����C�,�]���O��v8�;���|����)U�;�8S�_-m������r-�H'����Ǉ�
j�c9����  i�H���J�轉5��!���4�r�h�B��D������Y�鱆�1X�&�5�nm�J�B>4�	:����K������u���YKNk�5��<���x٤r]�Ւ��wV��I��p<�G�8��@��+��xe�~����(�w�ǝ�].����&PNڼ�X{x�z��Lc�C<��s6w�\�qucRz*��<O�?�?kU��1��|�H+�ױ:dbJv�\��@H,H6!�`�8H�����I�k�|��Ѕ�'�H�����ϧ�����]V����%�^`��R������B��@�֙ǈ�=�P����؇C��L$2�FGY�HTu%~Og���� Ts�w�濪��fG����E`�U�P��G�|��sMv�B9�R�.�i�W�*E�g��	�x"��m�*_�kɅ��Y�����.�QxqCNx���z�(���b�'��T)�R#Z�̡�(m	�+W���-Dn'����#˔���	���=���J7'�y�y��W�4ޠ��q���5�OĻ�	�V%e�T�pT.�s����C���R�3k��m��v��>c�*�t�|�Z&9��R�܋��H�L�'��P�y�^����Bw�?Ev�~�c���k�T�u'��|'v�L��ױL���~N�Y�;���&��l�k�څ�].������n�����=ו8�F�7}�~�ާ�A]���
NŌܙ5��_ŀ��?v��]�vi�щ�`]7Y�����E���#�}h8G4���V��j�}��B��~Nn�nD��WT?kWm`?����*�h�l8�j2}�e�엿�z��;���8 �8��^������%i-��%sn��- ��0���ѐ�(�g�?ώ��Rp�}���&����D�l↔��E�A0:�gH�4;��ݘ�����Q��/��Y����Pč!�y%v����fvb����n�{A�)w5k@d�[����H�r�%:|Qu�e�.��`��M��X�7�]���W�Oa
k��L|V
�;�z������z]ԯ�wt��cM�d�����~���u���{�A�2��oi�z����[o�7�״�x�zϟ{��R���r��]��:xv�&uag.�������3<��L[]�k��q�.}ã�!��ʊ��M
��j �>���2�����C�N��xd��l�/o�'�,�u���q�P�"��>v3�����X��-L���dL@-�y��e�� S���Ԅ08��9�^����-��F.V���Y���g>7�`�`7}_8}�z����ZW�就;`�4(�UOmhn�7�d6�h���gW���-��մ�LӕO�Z�����wI,	�AJ*c���ii��K/��H�U/p�ZOeu�K�6A��sV7��b硗�pk�Ч�Kơ�>���L� �*]�j�;-6A�ہ��Q6pX6��x'���1��